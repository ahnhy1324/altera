// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Bsr/FVcymsHK+rgUxX5U6J4vnNv81Ki84cfCX2A/Dky5S0qbDt4aY8D58jn3GI45
Q9VwXVz86/S2qyRhTbpDxpVDUWX2ZUxTACCVkBiykYuKkxKZdLWOOlx+vdKrw5t3
6rveKfSI7Tmuu28fNHX8a6xT1rbt0Vp9LHzb3XP5//U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24528)
4azSiplZtMfgAqp+lTzjymzzOEQvbAdXN1xiw7prv6u6IHv8UDxIigtU7KyhpJmY
554DX988jilipRYiN8UzVzA+pRSabaRPRof/HWh/IN7Kh/nE6CLZzGC+j4n8Slkq
AIdMWMHtheKmLl6sJUWBK+hsdDPIkFpOU7/WtwqUxZXED8U2usl3VjQMqM+RJlIf
d5PrXpX9KoDRrQMZiIWrjzKk+AOX+YzveMoSegh5hJpYIwdzKnonA7wHSBMXNZxT
mcZdGcGYpyzsDvQBGLgOz6mt1w6Qwoi6j/3SSQnofg1zp9KRQKacpB7Nf9arS6Zn
eBXMVqhx7eo61g1qnrKBwuEaIQOmQq5a0pJX3xbzJP6YIcXo4Fo9teKpFl1sDJSh
xBsDEATtESVcwLEWHboxX15oYzyD2tw6CBe5mldsoL2XJdCqRVXOcEk/QFxkIiHt
OiHG1+2mRY+NeM5vfGe9r1tL3RBdXuPeRjmZ9Di4pSGW3hcrkpgwzwDzFBIw2GUW
pm0vkRrBlq0n3nAOhTogSwFYoH1S/+e2+fW5xU0hB79BCwLRBvi2NUnBJ4tLDWfv
R3DvaVYf67O9tUSlhiDdMvkwq8Vx86H2Bn3j/cgMDlyC0+rcNKTZ5VUQX4DOQlYM
Fznja1K8DepvmuTYMycMc9lKo2CYvFSt3iy2uVxuDZJdKyd4heUBngCa+z4GSyjQ
pyPpkrPeLgaT9WuOGSX5ykjepvzlrz9ZOTlKgzbgWfG918fj9pz1Tuyy+OOLIu12
+Avc+E2JIEkwoKJPbUBsAn6I+S4FPpN6Jn5z6ypNUVIpWVOz58TqM04o81pTgOoZ
F/xeUtM5pi87/r+x4kfL/GLT8A98I+vKkyzr9tCfmMjJbl/a7Ej9LuxAOvt5hEyn
SUPWjO2hTuj2I92n+ZKhJUS1lTMPZL8XSMyyO+2//+LlSIWmcFb8W97j6SCGziW7
Luzm5Cggi3sTw0evZYQrmu9HVF7BRwlDvDi6C+Hb8awxM4/XY4Wu2mJu6j2NHvb6
7YjEd/URP16wgxIqG8hmmIw0eZZlSUO2gzNUbAGSAUYaOvZy4dkr7Qblpwe+Rw2K
Wubew4gF2VxE6Cx5OYGgOPmekGw4fy6ynky37Z+RD6tkBomroo2BxAX6rLtb7ZJN
rYrUoLwRb1JZcPSvbzhe3BCzXrHHF4D0HBp4wkAXsctdkKy9rTuXsqZvYgnHm3+K
rsugmhFcqKugLQ5zjYtmckR6U1P6ljXmnL+QT6i1gA2C/ziaUlIUN8n9TmF77C9r
ZaDzCUlTCGgYJzyBw/75nJ8Kx8tW2LHcfqzJb84yl88fdFfGrpbkIrzn8IpKfVho
QtR1g25616QWVHhganAKQiGMk5PtQuMCnXATfsMfqG3kdzJhNfhgA8wrM2tkTV0/
1No+PhROCkcOf4NiWw+0eIFMA2mEqkK2k9jJr1STh1x2+JvVyETKCteRQ8CLU1J7
MKmG6Qw0A7aI5kL5UzloNMNOiSnc7FmZKVDXOHkPnBjQvS8HzBswROCF9WWuylzc
jbUg5wdZa1Pa0WNPfjispatJynmg+2Y30xSiRvezyoHBIQ7eG8ZiH1rpr65depX3
JCLCMmoBJDZTHF+LDBGBT1Q40QazrFqRNbYpIl9T7oO87nNBdM9f+6ReFvZ4VH0I
xgoIYqYgFcMIR2GP1w5JHDF6unZ45hxcZ3/6Mh8+Pgy0aDeKc0lROrwqUpp6QCWB
BzoNZV/Vbt6neV2U9FoD4jEFKtCqroCzXTtwcnKMNXlZXrBRoedJMMOoHwUTAgbP
krGK4f22dioVf1W2KA5KsgkxNhmbTzCgP1mZ6znsfnDAKkTy5GlaHEcFIKTYLc+l
4+wb16C2+jFyoxNX7cnW+LLZImfFo0PBuc1JjbEfrA+y8PPqaTu3hQtDAXd49Z8M
NopyTs/CFmoSXsqYiO2MguovMw/J2aRiranWMdu31dvZl0Hbfzs3CW2NOck8CaC9
blY7QDelA1SOZyWHA3bGx7k3Gq5pWdJ0fI9DiPNkGxnpTyeHjidPaM7H6TaWQyX7
PHfdVHLuzbzDp2jN5tfRFDxIYnnGuic92x2nr+Q6TIV40IS7lupOilPPvRfKilEl
9y2fhZ2gG9shCPBfI2PCOupz6+4tlyDSrVrnPOA3Wv4k62XEfeZSv+YbBHaQQc9e
QYN9BdI55YVRP0Git8BlsmMauYHBXiaJ1JaZ/RzXyQOfYWaDLScwHPGRvLStolyC
OUw6AmK60Qxl0DU1fA5mnDQUkBJL0xCo8Of1NT/zNLyfNItV1KDr9/LrLiSwdIvx
S1BegY7i6HliWs4+9TjTHt0ozgtZBxl8EiJ0aFrHVkHCqrdDM8jqTeeaz6RvoH3l
iTFzw6xGFgvoHKS7CfLecP+twFpSgyqXjD7mwz7sM3wchZSOJNmPzXYOWn0+MLis
p0HOlc0GrgamFUJCI5fS1KbbBSm6pKfwX3Ny+K0eR4PdWZaovgwLyFWhsEqMYL4k
gSYPpv2fzPvQfn8NRCNvl2FuSYa66iZ8UEh7xwrDcMcvYTDTet9bz2+7L8eS2G1j
Obnn8CNuYKYJipm4S+7Gfbpc5Dl5tT3sqwmbjVir+ukYCVh5ocbpzXoI41O8BSWm
EjAEn7kc8K7r937gMlIFpczuq2mJPnqTjKYp6mG7YhFzaXHBWPmM/xZ2sAYoOXbl
jlKGxR05N3tLh4q0ZdlzdbaPqtO5652jQso/ruBZ8aZK96c1dYOI5qPTbxw9fKp9
mx5BBSaP+Jt5mrJ/y67LnX0foGtZ50rBZ1TMYVLK0OECo4nqrL+W8nnNPkka/M3H
eVenBeFiZ8HQQyjeh733GRWtq8rnudz80KJXuyLGvTXETzYx5INrsxRK2/nipSlW
x3CzDjlKpRF43MS09LaXps3HcAqWUahlQsYWwmnlOHh2YR6sCB0bv4VgHPEHgLXn
NCWTC80OUVkktlYEus6CK9Jx7QcGNzpqlEOFWsXtka7IP9lRMbphZT7TqER9vUks
PqupQoEURrjJZjm4FUmg5YwSU7LHcKlNH6QcpXFCl0v65WYa5eYR49mus6CDwW3Q
42d8rlvlT1ceCz7sPekLskFta067rwluu3WmFefBHOu+d0nS8O+e0YUzmqKhYCyp
YCMgVVZfCrmYVto1gYA5f8l04vYsUaQ0iFyWBFuAeIuvCLqmFduaaVWZF75KpzH7
VGzMvh4GwwXaWt+B3EndxF3eFfxv+DvN0zcdimXGBKlcfqV8P4yuY56Nn2wv9T4x
6nNoVFxaVQONQVqIFKV/qIYStrrLALYrwsBUtV7NnRIaHXAEFLH+HHsbrqB5B8pZ
QNdjssN881mHfQtBy1yY93V72tP5EYU31+2A+YaLINjREbQ7qdRbA97+O41d8XgN
GXCMOMel+4yu6MpPI926AHGaIoTHCvd98Oh2Mi2DOJDDQJFAH/JkRwIjwGGu6Fqn
hJkmsJi/eDbqAeKGRbkeZQialtnGPB2WGzIU46JvwLigHEa74HiL1jxhobfkzpNg
XPq07UY9cOz1ZRQAWosCfB9QCD2NKUA1KuwtNw2XVAFCw+M/QpGuHBMgIdjI1XS0
mi71aNiTO5kdhKGy01nxgcOrYhwFiCfRirVwQ9sgQrv8Sk8EnVBCQlOOKWNwF20e
aGgCmg9Ah/B0fQjBtvJ6dJFoT998aorYeFsr68P9bvjDonyx9A5Q0r2Q1C+plRJ/
BRg+SgFwckAlPgJAeEeyKHqyjNBx4KRVaY41E/v6bywBKZl5Jp1MuIsolbMrkOU4
Rb9PZZPbBJatZmy5/p8COyWPNQxQI7XauW1X4gq7sbEXmNLpOyAQHgwU6mQcGFyx
R3ZTnXG4vmde0XSrEW/peOyB3yasTnsA1Q/K+cuCY+gyzQzLlqj9j0nPS+oklKEX
+VtqiJ8MwW1R4Rragw5obZget584HWR0UsMtNcmT1IQfD8+FJlXtbYOxQy+0a41Y
sWwtyht3s1XqX+ibWttIDBWDWEKu7H8eD9yZgzfSZca5zW3jKSG2uNvHDxz+Qi1g
xYj/xzH64Gm8R6YsNUcUWofXxSCsn/KPwYNzXx8YJ1O+hU+bnZ45xC4HvuVHXk4A
gzVBYekKoxwvSP/Qi9qcCUllciKs6Tn3uvI5foF5Ea8X+euPuMVfsEukwdIV3+gW
0ZqQ5VxVXCAtVh3YlmKw37JJE7yrcDu7TUoeeO8jFmMha2AN7zt9vB9bDRhGYVbM
6LWsWP2cNqE5UuLuTFN6CjDstn5Vi7btb5wIObtl0K7TC040GjufDiBLvA0vAk2t
yBTQol3yDp3FlmJlBvoiElNNkId9ecN/3MeZU+7JNGmWW0DJ3WsgLG+J506SXYD+
mipA7sxNK2Uu2ELuFLj1wwy3J8YkD9KQepA8q0Et0A6/r5MLEXkjgnecHikuQdDC
/KoU1XeXtKYljmd8niVQQaFsc5R5VMQS21o/2sEioejJqxBDY0gS6m2rfhP1cMWi
OVLIcWX7X1WdtpPRYVab2jsQaV4Gcrn3KHfQwdkX6foxs/kpHOW71SNOrS/JoBot
msQLhaM1uVbvHAT0Fjcsl80cLlOI9FhdRwBj7+N1nQhXjKHtDAFSEuR2Cb1/L179
Vh/erDmwPoPKN10405DWjBdwIamAJYb3v6q8y9xqX4Gc0r4H6Sesu5bJtDTNw0Aj
bFMt8AWED9Ot5AIb3vvMB7FNfYZLHSVmR8iXS8/PXM0tdKjmRsgDSYSvSV+iIANS
crFxWKpEXxy4P5QmqkRGFJG0BLYcBOTRWtQn/yu75xJRTaqcydpkJ3arZYiJGFf4
srzXvXtT3ta0kG9HXeYvYkTjcWY197ZH03EM6mzDWaPC7aDCy+8+W0kWT0tuOS1i
v0jEO9l1+aL4nDiqc/Uayskx5Gx+jOCBavNlU2TYmBp9G22XO8Q63MsbTxT0oLat
/gr9rKk55168qX1BEwH2DrGA548BAnYPuUEfkucGdcFDQ8SfH9ZMsoA2mOFKUBRh
9ecAtepMnt1fW3VLzTIKHpZTcrvQ7XOwA7oe5SYM+7WFA4qBovNiAGraLQEHscA2
6ijljz49Mhp2Hd9z3WhIWHdf9GX7t8t3x+4DYaNE4dj6yjwGQcBeH+p385r5dNNH
rObOxJB1aq+crOvepQw7jXVrx4IorX/J4Jf4rN5pEJnp9mIFWoshuwlItibhOs4T
8xSxtJ0bxtvROz7e+Y1cew//0mFgnPeGrIhdCpF6+bvqDXW4lwOhZTUY0stoOC3u
S2gh3jTnyPT0gB2fcK2lXaH2zOLy7lsbaZYJqDG5YtNpHhPdem6wxXVdsxNuLicX
FduE+MJ+AqvzFMn4chj/iNCyBtBJACfrvQcQW5S1AbrZ1iVkF3Zy+uSOQDsHuqfR
NRVRQhNS4xxST5hbSjb4C6ZMRx++cQDKO/7E//93MhF8P6Ob1EBiQ9o+oiToImSA
IMdec31AJV2RAt2OOgPrwgisZP7MWSo/YdZGTjj45bduy1xWU8VtNoaIZv3b/Grr
hVBqnBPtkOCkrxZf186O5H++nkBK5bXpcLrPMrhE4lOcYw+bnNsOECqrpKM2dm8X
6gEpmJnDi2vv1liQFMqMBL1PqGhsQsloysYcGrv1f1CHwvrcEkqid7hrgPmPS6mX
KXEsAJkFafoWml5gYX4y8/i429E8qzGpt1EuMry7YdAO0HMecys81V1n1UXd+0q+
sNdrIv7PRvKYjzMzWLoGStH4tYeCc+mU0kVktFLCrJe10NK9kewigO12t1VYMVDD
ITQe5HPuxnVUqW6IOtkah65nFDtsJYasti8MDPoMOUUSQyxbUYqB1gLICl2ejHtv
QHRWLpAfFRptoehLTwGqW5IfMjRK4Z2jvdmjDbvGtSNh+GXxgr+q1zijMkSj4Zio
peReDYiSg/37qsJHxZ6juiw6uFbs2s5oaMK/1ge+BA9n6G5N8GdxkGTek3U95+1I
KMVCRB8zGMVHUlopjuv8piv5MLmlINEbOboPX6NKbWh2MINW4EyiTY1HaXbtLles
JG/xRZqLLeG36XEdDi7oGPda4TTv+aPgY+DHQoenRPdGCRObDb0FTDfzpp/s7bE4
oGLBvYW0HZsAgRgG1zWiVdKm9wSIUv2dJt4kw01AwXy43o0+Y2qkhZm5TEPqgBV1
b9iULvnhDSErrVlFXMIegGzmYa2QLKi41D/FNK2p6AEAfAltkoMmTy5nDa4qnL7O
6eyC9Qaec9K66UxK/SH4xJZx2qwYvqIreoDjNH18xCWp6N9eKonixXjr+J/7qmqQ
JDh6c0gjqEA+Dxz5B0X2iYi3OhEvSI2ZLAtgfapWLp0eVIryGjIeiGc1h1lwQpbu
5gRQDKruVu+K87xj4NCQCXwfUPA0qc96tk1fjUP8V4Cy9C8L9utnrim5IaTXmGtm
IHumIx+mJ7CW7DkLnAgxqnRiJqZOP7yayKa6PFMkQbUToKjMnusmcic9J5Ns9bXk
IFdZ5wXhTu/LJ0z7FF+gubYdEqARObAMNiEyhsZszb789IRghRlmnxendA2nBTdV
NgXi8U0W4U4e/77gxavo+VymAvIrAdYzCmrO+2CQ5flR/D66+UGQvC1XReqEfp23
vLrOeEFWqqUDagHkHCCqEXreMA3VRzBQjC21eekTNV0dKQMl5y2UpeWn/FSTTH4y
Dz/RdqSi40OftQPTEddezLwQs9Jj50aVbHESQ0/WgL9WlsqwIzO5gsB9LEIRSq+m
O84eb4TsUqKJgPNc7VSZ3NjBAWAy8sJ65npJESi9JVik9j68eFg64Bf2dGq5iOUy
+xwK04GqC9i9g0CZ3s1+h/F0sfEbaZL8vzBmDY3qd3ksdKb9MrMD5YVQ0zG8WI3e
8wGhhBcBXlaHjefsY3u0Es6a1A1WX9sNRaeT1/kthr3BgIZTPYhJ6rh86OJkTwZO
tr5ldReLIthZ2xu5SFEYw8Ty6rDv/lwGddxYLfFtacXb1tNJmNhHkER9QZS0vizf
1F+E3u6ZX6dPiq8WuzFxhth4jgAsTdF/hgyb6IYapxATYF+NHMTrZNohampA3FB0
/iTVE/sGfIdJQ7GfLdOOwoYQ8h5omKlN3MJLoN7p/xjj7Onm+I6TsRwPGXjFa54r
v3RpRQLzuNLBvJlrtC8X9UkpV/0TuBbpvPbUxTfppkqv/qquKOcXzd/iOEJFAwKn
4TMrUQ1+9Rp6GGLFAFV+VwcUyVNXcLBdmLMNGk9r9jfbhpdyF+iszmtduhM/ML+Y
ZBbcASsI7LneZrzsizkvrJxqwUpOURn1u1KMjc/pufiBkpLSmiB4Zmh7MguP4WQ3
mWuPkFwJvVmNgN44z268swzL8lzdg2swKNfK9D1JRj5X+Qe4bxELoyS6vLesIOuO
wWLjJmHMNz3XAKZwKXuv4X9Wy5IBqq061WUUQW/t5oD44ixBZeG7UDzthkWO/mQv
8UGkKMSIF2hQc5uxM3gAii49Grv8o0f2oIx0YGsabDikAMQJKSuS6w/kdBrkAmSW
O7H4/iKXUvwCsvBoBluJOjcKef20aDZAo+uFDbwYi+rui4kk8zAoF3mkc7yVYgHa
4AijIKUXlS4FYWi1JsAkSc+Uh+9tbB9JNFlNChv2dNjNp1pCRfj1khQhA0FJ24Me
zVMDFLE2J8yFl4DxeVj1kK3+u/oTFEvMQA5mFsEnIfyDxR1EiBO9Y6+SsFukU4MP
Wpqo9iVaVon7ivsGwVq58g4e1CccIKk6mg1xbpdincMBjTIKUbh1UoRFxHPqJrPV
efrnsuwKMv14ENsuRoZBooyWt616NWIEr7nhmi1WEBRChdLML8vS85bp1xfS4DTF
fNZN+DIiYoAr3x3wMvNil26qAOTdTNU5AjiVkmRC7SvTZ23ayk7fjq+Km35nV1Uw
z1aODede2MfjvkNaiwV6vV5PUXBSEtJH+b6jBvoeiKjzWL38edjf8h29EFz8102N
WOvkhza5e9xYgLRWAe2U/SD/zgnoNjvkQaSEavTo0WNkGlBtHt+5fIFKg5+Ygeow
h3mVKc62X0cGk35cKa2+uZnTJtEIJ3mQ9YuKlbuZzzEk142IHcE8uF7snAf5NDzb
fJ8SbQJGX9PtxpLftZUgANToZJWggN+g+c8ctFnA7X9rB4CucD1cGniddgzQZPIU
UYWVzQ/Mxep57yAGlRJRMSNzuah18CcwJNwZzox/Qriuxz8QVfYLro7i7o2u6RMg
S2eqgJbezJPlC1MpnaEfwbeq64kde2zYgPXGYOTCKBT7BxU8K3OjwtA7idV4jW43
qGpvk/F17yBEKYedknBO9h7P9qNLbKgoEvzNq2NYi1sUyXpoh2PxKVEcHAylODQd
sieGV/PmqK77FnfplL0ZqQlVPro3BXfVYKeuuD3v33DrfvJrXcvk/aUIRbPc46pX
CxEvEfnV+iwJeBMjeSw2RNTTrHon+YzsDUQIj3m5UwgcekGwL0glmVE/w4g6D8jf
LgrDyqqQoktDHlvBSu209LtYwGd3yAIGJXe+lk/PLwTWvBbWyB9ro/0nZQVuTCg6
hANVKfXlUUXqhBXm8C3hjZmYdYWEsce0JjkefUEn8YrptH0CELOhUE8m50BY3WR3
WiCFwIYtN9Zaf8IgvXmJQ1zvUFbofCP7DNM983SzszCrihvsRhUyiahGQMfzC5Iv
pB0puc+HqPcn1Qpm/R6P8NOcD75k3RXdxR9tGgXnVYjYPRrEDDZ+iOvY7RkwSVLg
HErhu/+tGTFJygRrodj9fBO4qyzdSfx40LtE+d3wPIrYKkGt1D+/9zwWHeDbP5lt
/75bdCw7R8z8bsAXe3xxq5rfU+y0sjrHr0V16TTZxyISPbPjmasZ6xj2zBm/VpBN
CmbDdC1UBDGIT1Y5m+V+EcIHiP9L9br1o214O075bXoOTA72RAJUwqmKXYnUX3GA
c6FalxvFSCa36thlVyokv4c+/2JdJ54/4ZJBhaiXvb3K1rtl2HVMtSnRu6jaGYUD
27VTfcNVU+9yLkhgC5d6UYWn886ZNYTU2THFx9BnDRe2nGlJMowoXS1PBSmfFW36
g7S0TlW8uZTXbPZMvrhRE5riX4QCAlHaps4TUgLjchDn7Y8LW+lEwdftE1Ruf8s3
vnzV9/0hp+Y7gxGq4Xo+DGyxOn2dnhWi8FZaIMH7OmExnMeglAWDIQEWZJPmC5gB
mCyMng4u7ZAheC2Ux4aVuUBG5Wl2pWyt/TqSblfypXlbc4mzHnxU5U8CPGWSfe5t
tX3XcDeRbDdzyQFSXG0uoXMSYVmtye11C5RS36d5rAPnh9ugzP++jJRBh8o9YHnP
hkWKOaUFxYFfHcSCy6NwlXC9C8qhzPh4uHL0gb3J4S6vhu2MV1ufJlpvNEB9Hgl7
32qXfmldPkZ8Acs45R3XWzwPsB7f0bHjg6jMhZXDliGUJzXY4t4ldN0vcaEjyMv4
oPU4MjIccck6MVAC1edckhnYfiM/05TQly9xrd/3mafzIM6qEkcLqO2p/Urq0Z4K
/22NVNUw2E6xiOgeNvTvnpfrxWQO/eupynlz9Di3alyBhUjg8/7011E2HxmUuzLx
ad7vcgrfUeXkhU4jLr7YY8PA0767fofyFqAKBeyGml3+tpRv3GDonPl+iuYaS0LN
xZVnoMdtM2/kw52mtpRZ7s0kK79VY6Jz2t0eLAql3VizJw6CJHHGWSm25pWaDoMj
yxot0pp9Tmxs+k0d82X1IPGpke+6mU5de0U8J6xlnd0qIds8od3i2nW8ZNCza/Ij
0Lo9fWs2137pN3m95MRQhAeNclIfjc22LYBV8q8+Pakih0MwKnur+bQnXr6VjBeB
yefKPMKSQuJmqMrnEPXqvcFtws6ALfHqQctiVEBwanzbfyeS+KHAU/maRv0/kLf/
foc6Hnabj/RGwO1IO+s7eZUbuScHWnC22nNLwmuqcWhn5957S6/kQjCB/GfRbaU5
k/CqAgofrXUVcCLVv8ZVOoU8a96crgtKvNj+sziphAO5OEuRO9lcjXF1v95/NclH
/NaBCn0YTJNlCJLnnvV+MVbpo5eAt2zSNfy6KBEYbR5alpGrfko5cRcPpXrVlt7n
DPO3KPJmbYnMyOkVPOAKFXBuV5aIY03+BKN9gLnb/oqCspFa6ls530gPXaiyGBeU
OgwHzhVKEB7LV8Wt/QVRm6pQkBCetfjpAD5+kFApsWb2evEvFbX6hWGem22FeyMf
lE6vEknDAWNFdI8GoCO+Kb6BRoYzFDBgL7PogOPMhgOsTO9e0GYjaEaqBXoxIYQY
ZJwCtsXZkgCu4r26PgMA+vubQyd0h8X85axQAz3L3Z4qZUXitSk+lzfX6IF58Wnt
jN8W1hF6CAsyJtmtUa5X7rmfn126Zm9Qzeri0JE/japeBfXlsBSfvXLSsKwmrlWC
gBfgEt/H5j3AAgOvXouGX7t7roWeNxN4gQWi6OlTtvXstU0h+wsbi/tRhkQB+PIQ
fG9ZRfsENrlkzbY/uRDMkpun5MkcGVmSUEPdvPkihP7JaztAL35jIMyvmPx2xtQI
SQ6r4lJFvmZ+UK2W5As/sNPniPj0XQYrVpTVDm9MyIIWOskpbEco4w5ae9TQmC+J
CAWlBHL6d22UafA+CSok89gpo/W6/JOFmC43ESHqKYbHBCRRrs7Ww/OJaxdebE6T
49mc+xBZ3H7y3el5esfgcAtLBAfq1o23NL+ko8bFWcHoQJuJTraN/DD/0X8jIK1K
E2Qasv2FPHMuM2nF1VsUyGPb+8fWSyshu7e1fMcpv3bkhIG57vESMbwLACzHY5u0
N/AplGI9peQe5ajIb8XwWqE+Fn2lgOC183bUqd41gNuqYfZXPr/zfA0M61iGWiEJ
KOnE9iijzMJ7BtP9SGOODo2ypYgRp9D5lsXAgGinulaJwFCoojss+syNtQA0kOX+
QZVjyusYz9LLCMnitOn+WuYQaYv/tQO4oJTAMeRQCOpKr9S1kolFr8/13MXPzi2T
CZffXtf8eNdbHRRsfw43xmZsL3kFNw8oe6Nfo4VpUfXjdT/0y2GFieqA0YWh2M5w
GJjjYSR09wmO/bUhaxBOx4Xj4QGCHVlZqmgGWRBj8XCEw72k/2I4cCZdIdYl47nv
gcxXMik7y3gznNU63roWdSpf08mbIjHO+Sw9VLZz0/38LDKDcGHbp8wm6GsbEVy+
ToQzgRsxPZ7zw5J0TypXlWgD4p6VxUbPYyCcNQDs8R78HdTG7Edm41qTh6aw+Emj
T4Fm6jt6791JCyc1mL2XcYIcxc7sozl59qNUN2IeL217l5b2cq0tGQBM2uI7mlzc
DDO207rsSl5mm44+IEjYgrLkXI+MXy+8J9GupI6soaROBA4p98B/SY/kEVMVgQ9g
h/0dLVc6vZG/wDBKJfc3AlmyCZHWwmc3to4+G4xWkFGOiLV/bRo4mUFIHT+wX5U1
NOqAZCgcFL3OknxnN7c9ggE6JYVouFsfXCAZoUcmQF9+nqb/20ZNVxdlg5gBgaZA
DK+3Y8mG5I2GmAsazv8nTN7nZBJsNBlMIpXU7EzmSoujjEbs6u8KMH5+fxwK05GM
/nJhFdSy02JA4oXJtYLc4FYaB8GPoPRfkJJ2ofHlTt34hn8+25maBbSCljpBOf1F
F6CHDXuByIh9ByJZhOfuEaZLXUZGyO7UGNfvC2heN12X3QRa3TRkPK5zC+jyMIxu
O6tBrf9z4UCyiwn+LYzUZWIEOW2fRj6cnXfzOiN4EVGp/LZG9ItkmkxyvbjGmZlS
UbfwjCsZB5stM6iIaXXUYIZ7xIeQHc9KZLMH1dLG7/yEFvNMJrVRoCwzbpfaX3Sh
mPlzMJoiwoDEDk0DImfu1iv7bNXCJ3i0sKzNINxKCpkGJoCLL9K0ELG3uwd4B7vY
X68ExUgI1oMDLBMgS+4sfrgyNNXTIGqzhNSVlmNIsBNAngF7jfJFs/D8NOg+Orin
dxuwTFsHik/S2Ruu01vZosmq0Xee5iQefrUT4swz3mXy0ZGP53kAnLQRU2r4fnD9
qwHQLfdCTs7m8q+YsFilmGfSvhsoLkUv2nHQdN8h5R5JKT0GKHtKBvJjaW/J7B0/
+5ugC7ugbPmqD+xO7Fi560suh7UgI2II2816ks0AprlCYLLEBPSnRXaSDGVwIfn+
pDsPAnqUs7mVo0KhPCJ2MZLBrhOFubtrIbgJFS61lhUKRpTJ633Rlr1ZOtSh33+D
ziGaUrXAbXtGeV+PloibV/qVh0ukgf4lwv10kXhVtS38NbMi31H4zqRe6fn2TfaI
1zbPvVbB3IntdX/U+2U3vFjXQrBPKvM8tVMLD+U1s1oAVSO9sP3ES9NvEA3UKy67
PD0WYJeTqSg1uc1T6LBkftc4T1D6uSsseKH8lPLlTb3sXDCdo3Zurlq3uqjpLOly
Sq/nzZOmo412hT4rKx5ByhBMr/6w4NGqtox4sEXd1wN/WEdQWhDcQHeBps8xxNju
4gOkXFP/rzTX3q1FwQk5vOVm410+PqBm+JeeGy3IqwPB0j+PJgxx1bef7uVJn8Dl
iRgpqsfobiXWqOJY3ZRpzl6NmM6AAtpRofVeuC9uj7OzP0mVgYV7iIlrThGsepMx
0BzfUHiTiPR/+QW72iSXrdMqq+8eFl4+sWOMU/QumFZLjc0FMoIJhIF1yvyII73l
8RSu7yHXmeRI/WI1WaZdretNcEwJbeOdlModwcElxLPAzh4wFov9H84yVp76L+55
GwnStaIZbqbbeAmXGYOqToUAaQto4Eg9/O/vYBhZKEkvnoCQwGZ+4LrXfoLNrXHX
vMlYHSowSmFcGPB6mzCgosbeujJLkAZ8Bfzv9S/HfPiLgN/gGmk6kxDqIzLEkP0Z
JoPQGZRV8vv9uM22NRwLOzaT33ScIyMywIMCYvWivNzwpjnZdBAIL3kCeMm3e5Pe
2dafjpcahW8oKhE5M2/ZKKg4myRIwLcwwKaH58G2ovUh6oBgBQZ6V7y57YAtcCen
iPiw9URC3JLL5gHVH6Ox/HI8xGwA8iWKabuK0TgBNM1PSffH8cj8VsZFYWt20APs
OT92wjqWBkXMkJo5nayR6kq2kML8OipNU2ZABMbnjrLhacgfZg1ezshvXEYIMmKj
di7Ef0lchYxs85PbZaP1+jfqgHaoVliCHgys9h0QIaNGeZVVf+sefE/Z95JlBSqV
rdcfHtfTQmgZLy57EUeTFMaodmBFlFsFeMKdg9EJsmDde4qBYBb2qaqt0MUD2+oZ
dPdmysBu9DvaLyWgEehnm3Rbg8eZcKWu6W9gyO2aehLTa9DIaHqRgS0lN+wO9w66
lUb0aeWUtEZ+b8r0PYZOdmiFvo85ituUQKkRwyV6S1s8//HrKUHx9XHUOV/0+Sf2
A53Z1Hzj4oDrZY8NrVY0T1N7U8ATwA4lFPRXsTewzLVKfIHK6aOsdjjIOaoAiJW7
g6Ie5a7dYyKkaCJdsr6eVd/LCiM4AKK/vbXcTte5zw1GG16MWShDlwOQQABjFRwK
i7Kiu2cHX1k5bu1JlWTbYRimRcgYarodNwL9RH8Pi+JRLLeQ0ux8M0obnes9KqHf
NCtveiFPpuzLpLSAZpyrq4hLj+/lqSX5XAXorA1tcZt/UsAM9jCk66nQ1kXjsP5s
49O/+yZPWsfcT8LBdIsqcPYjQG9tkHUwmbjmdRzDuIMnlxIKyeBdqAiFY2ghee/3
JhZiW4S1R3pbROvGfjF5SC/4CrHqh/M0cQWQ+49jecRXQYOHuQT+HXHP7PyHOru5
E5z2YczAqsrifTU7pxHsUb+dI8U1qWRsIeO1W8auY44UrbmCKSDnD8qwl/kG++HV
EgtZyCrYtKs3KdBOsp1ED82Hiaiyl3n9tAw99SMKxYwRFn1/trf5yABYqr+91SRA
WkkRsZu7O58dC9y9RUAjv4hY1xJEM84U1JquRLIZzybT4iR6KsPpL97D1jTTNdZP
Qf3HeILMOONf3wqVv8BT/vDnivULuDG8miXq2b1C5L8YzzK1fFFdU3jKBikh1gNg
ypNz6YACpCOi2xhoBldqwXiwhuBCLwmK2PLW3ZWfAezIdUH5dMv08oA5O73MJZ2L
yZN15zW0kMNFv1L+v3OhRFU81iMgjrbJGYd+3a3VD7jqyF9j8MlBD9XmcFKD6QWO
y2ViiJZbCuJQbCXfOGh5g1b1+s4QP7WUZVpX2MmmeIZeXqT1uNjoVCfSPREqVGPu
OgrqzMQx/4GZBaloTODxeKoEi+IhaC2Zz9zgpWxfP7xhCwBJc2Odqe8bC7zWt8Co
Js4ouUFsWFvNiMynP/xXTzf8KYxEfu8iiZ/JmJao0tb3yk1AR71SFFW2var63zeF
zv2Js7yvTrajoiXpWwNIKc5kYTIfkIwfNSN3V9AEge/Xs+tlgtT/OLggI5kNjo9X
h5VpS2DCTx9BXXGxJ/gCTR3DALGneTu23WWVcVf5cn6dazIRKoNd8q+CUGxj5Ni6
EkcW9P2+ii4LN9tot1Y4lG72lsFJfkgOgc9GJxzkakscYnUiGk3Ev6ww7Lu7YBuK
rP5p4FLPKtOYxJFwSrvtGgXqzAKSrzRiGJ2HD7HPY7zLFC0kS8KlP+WR791VSNGz
CwKOUoMcHnu570zfRQmT/M2laFbiuUN5iqqv2WW20E6Kc0Aj4vbM9Tp06GrooX75
aIsFac0g+mEaL1l1H99LspzqglyFBdPApJhYY19oenqtmgqlYKxfEtxtH1Gjg/wC
SPHMT8he0TsdceUCHRl0uppCD91sGweOlQ3adLKy0Y4cz+ahKeb+gBKcFPLVUwG/
tZUniKZngMif2jNLgsWKWMMhNi+bhR77RrdV7F3lhd8AxarPWdvjp+AmEvPuPAZN
Nrd54106oCGsYA49YvLx0DdbowYXLB34fyIJTsbF/Pvnb0aHf7mBIAX6ak3BYjRd
miAOvpDOTDxVCq2vpTyu7j4tNtyut8OzoGxYU/rwmMDQ490+JoN4SHTEfnB40oLj
upcbyjI7XmXkLynPkhni2VF1KZirV1i7GKUc7YHnzCgUlKVd6UN4iVZQfSyKkuWR
tNABwzamGG8ROR3d93xroUTU0HGzGQUTaSy8frc5lr2XCbiZHG9hUwPHuWacU1c+
TfGT4dHih+6/KL6dD1HVTRNhEZMZJUtzkkY9qY1EYP0sGLg6T/8qitfYpoWEsDKn
CRW6/HF+5QiFHLe4XwfRa96Xe75Jjc5w3UK0TeeykA1C0y94ngcn/TrAFkHYrImu
9awfAMNH8Sx0FIYDTtw5jBf+QIN8p2uKzbfLWv8qYqKI5qAcqhA3IvQU2uozcYCh
GLNT9m6trkD2LoSLcqfUha8Sh7Tr4MJxFHa0bk8pBLKaq82tShPE/71b3VfYfDdG
VJO85X7AfZ6S9tNwMBKqFlT74LjKcwUeq+kWLH+Wy92GZIDQafSL8cIk9X6sZ+RA
Q9a1LjVambR4pandpJMz3wkryRglEdB/NiRTt58jcJ9Tu4WM92L12hOHb1000Oh3
LtvbSaC2dZTYmCLPjh8c/gQMJlS6KAFPJFYc3Nr907F5ob99d6YGcdD/qK0XNenc
Qk/COT06kGiBreOGdxkb6ffMGg+NVpoWkPV31pJQyhoBJ6CeoKxjau53f5d58JRA
Hr31hAlnk74dfDByl7HREiG8f5jvNED7uuR593Xw0nvlfuKqB0lfI0ucC/lnVFAa
EInr7BZ+b01gGmbtEQJgBn9/zw0LcebIhuivqHKWBrCMQs8q7ckFzHKEqf2h5fYo
/SELgLPMqnIAX7V09jlJQjaUNozSGJAUsyO0uR/Xr0fnKntFaWcJtdFG6RWh/miU
4+UO29qSocH/+CaPM1Ge5KpDBMg8ELUAIW0N3EcR76I7D/CH/BDmT5WSSJkLKLs+
N62IoqZBTNDjRpTKTWb40u9TvOA1vQVGChfktqkFJGD4jdgLv5SVJfbaJYPBau/R
F3JkLi9HIExLbd938j8FsSu/oiQsXX6fcW6CETX5uSeY0K/EarezbewhtFSu/1yA
j1xB9Qo561sF0QxLEiXu4YjyYkhMJDYDr8NM+ULhCdsM994Jp4BYmZOFVTGSGpHy
IOAoSb7/MRG2Yr52L5K+Rqso0VmAl/ewIzJvEhbisWUDrkKR/1f/k2evX9eIxAfR
NQkc5hkm8xKyCrA8sLDjDNn5k67cFfUB4/zGZC3pRjUiWhadFgEVLOfZLMRGiKfb
JO9ou93F7fdVu30yCXVdLd9lrB/WuS5T4DOcBHE0+l8pM/KiZF93TDiAFtJkdzqe
bkJntdQZiKRlWZ3pOABNqmJs/0MoeC9XCDnviAf572rs3SYewycazwWUt5p9spX6
g6D3scA/a4UsqS8Iw7TDhvQ6BS2gmEIeYmQ0BLzXdueNLRikzioGjhKZBqE1k7hg
JHCH0xkwd2GqmnPm7uKKcaG/Tz5f+ORXAlTSZvgP1bY3Cj9LC0PUExGvXRjxfTW/
P7YHmE9rV7X720/w7cj4vVs/OPgIZ/RcfWZ10+rJrgCltAinpQPiUiW+9T4xK4jy
EBLuA8rLGQSaeOIzvI4gwnBui/q6Vm8ywmTyagy0642k89mBtiJL0k20Y93uwAzJ
RQ3v0d6JJqSGPEZjegc7c02kJF6C0ejZXOVmWWhPGwkLnWulc6jWuX/Y3+pgvCd3
vwWew+cMKGlz9ROIiVe5rWsBP6LYTGs7fWza2SHBu2bseZzPR+weod00QkdQhf+L
Ny4R9kytMleHPxQhmIw3sy8ccmuXbB/zfah72Uoa9FEX+YduVwUI66L5qEThZxuy
6Eayxg7zaEZcCko8b+v+TzEB8toIJU1zHYLokBfQm7UvRQySA5E3CoPtnbHJ0zXT
obNi1R9zXLCdNX/ntIjTQIYfqVX6FtxEL9fasGlVXy4y9266Kh+YX2E5jBzWe6uU
IxORi0VcAshk0jGthEnRY/sCO2fKkFD+C4GhNdFXYwoxF/IloLYvak1S6QUW1JkV
aseunsQ1/gAdwB0jrcXdbcbcAEHJI0Mi2RhEUrLm/qZ3pgBjejSO/CFXDAW34xml
QW8/5xTQknQx+yNaSm17QMoaNlO8zJJVoAtee9NFhJ1inKpSPJ7U7YEXC9+RW1NA
+vNIKgAKwNDf7k3iKt7fN4Ux5G8FSQN7TN4g49Ct6rW/ener50cDapEyUnUs5dB3
snIqqR5cYJyIjInvsDpoyXoitGN6CEOXhsn3Mu7rOPKEt/3xlIJLX+/BXcTHaeyf
HSl3/cZ+vwx/UgiD3R10/t1wMd4p2+z7xClCphGZ3MZ524zFPQghfFcrOqLvxbP4
UPXTupsLzRrAMd/peSJY/i6GjW0uDz7UGBChIJ1wOtbTk4sV2y/ps13nAhJEhdCX
7qAFF4GyIowN8PTXZBP1fuOeuoETQyHGoEnxfFmIIecp2RlB+hmfl6ev1sDDS1Aq
X70Vz9jEUegl5SOW9w30JOSkDvd6NtHkwiaMBGf6/XjcCyCFyhwtEJwfxX+TVCkp
oThd2hEercn/49FtXoM/eHzaMmUn8fKvmMsxFp0bKU7ePSIWbTDCiZWRuRjTsQTc
LnChA/GgsmrPYgTgYPWnWmfR6hVMHhjE6yFXuf0Hu6XsPa08dSwXpOkI3un06eNA
FkYK3HVTXN+4Kjd8hrXsb35djE3zSgQ4v//L2jaPcck+Zw8wwAiS7Gz/2Xt7G4LH
KOVyLXxFsoPEvNYorBpLPC5xLF/fVmHW7Y7Mzz5VbwO1wNVFoxf5ZFyLO73ZQ6e+
vUs5NeCrkGv6mCma8CqNybLhtG2wKNbk0xqLj9InxN7bFXU/e7NH/tgBq9avkmI7
5656YIIuB+ZGAmCyd+hpBwBZRZI3OsCfteWZFAyZi/pUWTFlW3AFa2HuLx/nGMTp
cBUbI4KQilVCIMGssqLisaJmycpZuP1dpF8BSSVMeGVWw8L2kINRhFcjbZz95z+1
7ZXlSdaCHmdje/Bypt8+patzljts3ZfKorht4f5jOEXycSIXfrAVJ++o+BpbJ2z3
XOVwKjJGhj04va9XCyGHMOnLTQSgBnzKwDuxl4wl4tHR9JN1YYFu3HfdfTldY7lj
sxf+rZzWmWHkxpQHwkYxSUxYoQS78A6U+6oMLV80VID8dAuJRH3sIFRXSASBAY9M
jWft3MyQy5IFpyKZ+O4UsGkDEyuxU/UCKuQwHavbqGaGiLbXlgyilwFpQFMRVcOK
fjc405ydiuF8mj7UN3e6x3MiZgDn3BAF2dxlXChonNo9o9aPFYQqUojHLSrFyp6Q
t1mMIvfIMVIITmMRELYdDNpmT05aMUpX1hT5vYZqE/p+QC4ZiFIvi67darMug06d
6acCrgOvR5rzWLsQNeluGPffwV93ld6ajMljID9uPfhlJQFIOcqB96LXrwG/JHgC
yh1b+TCuLv4lgYmKN0fyvvOSSnDKsuW/EvhqoEcyPJzfoZSwQutL4q4HoXlFxULO
sBVwkPyV0WNjw2xouvTsGKuiy1Azu/TGPerINan4E9ATxlQK9AT+ooSSRa0HY5hf
vSsxvCStODaQZsysnoprN+dvqpPx/Ry1shTI/uiGOn2E2wyxwPzA8hLSVN45eJzu
wZCzI/KAnr82wLW93VVQpSZ7M6+e43UD+DG91B66rQYfvt45b46q1MuWNMvSGeoT
Ufon5DEC6a/xp1BE+sBCthRkbyMNA8hu6vzg7Im4yusK51kauY6ELAPLkFDBAOIs
bo9/+3fmIlPqKs9ijITvKCJhe956UPD/11LmYuqwtAkwucsZr4UJGtZ92xFVv32p
uHtH67rGqLJo5fe+POjQ5UUAGZe446AS1IVRP4z6nNIMokZzWzZmMvzISvVBgWr+
RMsw6xrT6gSkzCGL4rmzWgenMQG+Kaz0NT5jM3ZCsqiRt2B0gMqJhih3U4Nn39+U
NNolpP4zpbyocyvPUNjU04ZqRupuWhYplLjNLnMvCO5MzIdQ9f2EnTeuaY7dfFCr
z29BFkorIR2eIbjj7XXztfK9eUB4v2b+No7j4c73wsb80BF9dZDyG6LPKjP3WC0e
UkVk8kbL6kKAqYuYclfaiGkSo/EERalUHnmxHU91M7Gf6AgKX6bCVagfIV9r6p/x
+UuBbTGoKxA/EN8OkdmQBWjOf1jYHrcqTLFArfiYzalT1CSotDsZEiY/HkzSkkxx
igXsb648+piHzNveWQ05oWjC5RshMtRhBcCbN+M78HBoDXP7714p3JrBR+eWgBLp
Q9E4F2V3Z6pXBMXiq9ndJ8hnoh15WIbwNAAFUm8npmnSp5VzWycWT4N/a/7yXxlp
IrZ47ke8XM7EcUPoAAF5LCvvEMyzMt6Wgg7wKdEKtpXXSyw90VzINCsbZtZ6Ei+T
7iCGR2GF3W6bLkho99j2qwu9dHs/PqPi/2K5/D9IO++5s2fYb5owyx2kvjQ1WpJt
lJreGKp6YmYIMjgaUPfqFhTOdxP9p1Fxk0huUfRT3R3cHs/hVfk/walBnVqitlPw
h1BlY9yNsrTRLsH2hV7HQuuNhLNLqls6Nd07anRWMjpqT6+Afh8EYHH4793485Wb
hd5lkxAJfXUGpqxagNTfh0e9Y/Qe0GLJxpPrlNntvyy0TalQwpQUl8Sp0mf4OE6Z
OM1Hv500vUobCRuX9RKFXTuvWtvC5gX9LZvXFhRJPtukpK5mDbIoENyJ2LfIk4Ek
paxGhNaS+hAQkDlF8pYY7y6h6KfwHZvAQAq/1knkjZ6IpGV+iJbEmXig5YNGrSpH
8mLnQ8noSYvwmfpd/VlqRJgsKYZgre5B4k1lXrT2SypicRCguLzIShZwUPBcglwE
0r3Oh5fvZKY3yIG/3/b/w2IUOVa4b9mlNPMU+AwDcws65rLrskYMcrKBlNM0F3nw
ruqeUYwHC5rkJ9MXDDjWLJDw0wu9cQrfz6ArQU42XUntLT2LqZooAsO2PKPWW7SR
/dI76SyHS+P3BH1x6fqAddbhg0U4EIcW02gAA1YDCLYDJdoAz60Kog+1aMftV+k2
wiMqGa/0VeAt7tMLUq9N1HrwTBGJGVX4kgZuyshzi6zUIUNAV73Q6rFCv7/k7pLZ
nIKaFaOaAXRYYD1B/MDtUyKasu3VR+xDJFJ0iCxzOUmNhOk3Si2l+6hfK7MjWyCb
Er3Dze2Boo+0/alCtZ6DJR0+Q/roaRXfHgq3pPfIKT0btvAZ6GyK4equaqYmbZg9
J3A2q7d+WOHm3C3xs1RUcWhgoF6caGEUvjBtBVvHyNrcjt/vji3V66flUv2aBZpS
068IlAxEmh0qDwklaSqxUrLziBeSsZCUNu3RQpDCjTHjhYp4s8MAYW7lB+rlrrUS
ijGkteoqlc02+opgMzNHqNkcTAqswTGLMkkZPGGYqxTeV6F3y7JCn53YmXJ3QNLw
T8nfjc/Z0WZmWhEIiRwbwI0KM3loprI3rNBA705d4qthX8IzM4iafBQOrTMQxasV
OCdaYu18eP4eab4vdUmwSVAA5Scswq37mRTvw/hqPaAL8RvPJ6xMNuLC1pjorNbD
RnL7qgvp6g1/XuuyD8wRaRc1f7kIkbxVGDC3kLofThln2QlRVOu2lmUxes2yeKRS
3mONgVI2sjE6l9KQE6RunlXELudVS2mSnxX6T3L33K5raHWcWNCtewBA+xK8juH0
w76k0MrVUik795jGxIffO+DjwSG4IuiVLGlDLOLPxM1ypc42Z8pUwelcpel5WYFe
Cl0zriHQloQf7OSlDT3IFfjy3M6EFK9EbXM4Drg7KJU4LG1oRRacZ1cf1QwiDkSH
etZj4xJMiuFrYjr/cXC1Am9knkoJhkX9PB1IhSZXY7qL0hiM3sEpF1YOCQKCGAD4
zsml+o/oxg6EABhrEPDJ9ui9wIY2XapYL8ZniCDpKqOt5xct9Kq8qRsofiXzO/9e
FrHlJcqmVZ1HzbTFbSyphQUs7tOgAaHQutLd03BXxIbtOgSWmv50HarvOQTjcjYO
932yTTd/GH3Y1IidIgNV5Pbw0ddEhJa97p2AiN9L8PHPzrzDL3j7ZezhxZAANz4v
vOjoKYRs7vjetkcHVceO5GBM027H7eEKHJ3S76tjguTXuZFiQMi36rtarkO/gdzK
4ol0Q14oBpp2tESeYcsIKor0/7VHKJys+xcpqeF98VikIpXdU/XM4Nv/DFXWPfuH
hdSZdon5KoZxRkqGpuBOt9fpQfPUOddmZSzZ0zG315KmbdcXyXTP8HFy04Smb6iC
nwAnY6sCGfcYX9cGn23uz9Nmj3Lr2F5Zyq8uLCp55pUA74Q3FpuLrpG0zT7GIt96
jrhuAcYGaMWIEAIXJn6nIZTs1yAJMfhn1/cbk3ftRIBd0ojvjdrCE8Es/IZ8HLfv
kXsfGp3TypBPHGxlVYRFGM+tJde4KDDwt++wVgyUMsU4aZjn8iZbwkt4KGH813Yr
272Wlrv+y8SH5+qLgNs26DymG8VdJ4+HW2j4Trrd4ziyE+2etLiyYHj8bz3HrhKK
0Ya0LXjzRPToZf9GgebUi5+9X65GhNkCzDe4s5xnPyRav3IcivYBcxBKsS6y0s7/
bfdGnMjRGE7oK3nx48TbjqD8WKX3M0Q7OfdsZiiaUcXKFcpXAZH5j2OoXnABNDn7
k62DnvpcQGXAmi66V1SqdPtxcHHu83dXhLBQ2/lJm8CfxObbGWKGbv9seWSQvwpn
7RfW9ypZfEjLgyEeMpLdpKFyZ6wZfvhs4cTWNJU+pJPuWyR2hEc+59/yW1s/cqkA
sSOadLJc8DXD2lzh8YzOdHs6cdLCqEdWBH1mwCwAyQz4gRZnQ5cC+ZibRwEBjpZS
D87864d8bSzCA5LFeYM1gkeCPR4kYzI1zhX0FmGOCFriUs+eB7B1xsjWBodeIQgw
P1/8MRRG4ErPrMHmUjXsH/Ehp/9VXFK2cO9lVahkqcuVziCgWmma5xar8g1a05dB
sew1f+NrIAsiqG/8m/nUPCm+UGrsek/C+H88M6J0vYAkJSKLcOCCo3cEnTPvDK0Q
CgC2DUvsPYU0hmyDzYAS0urv8jBh8jFOy/XXM/fwYtqh6GBnHyEBP1g/39bSFqJt
b5k9/hGO+gVPp/ESmQkT8SdbrFgJuHF66v/yxce4MX2kuAlFKVh0z+r7oCj1V2hw
uLJnu5XVkZiX984AmPsM7s0k2cQwncDgQc+UR8vj/2k4s3a9br4IqDIG+QYcZkEk
NpwNRCOGLs1L03kjNWskpJd9jfYz6dgB/OHX3IaUP2YSxoN4fGfjQiamxw3aDCdv
p9v7aQceMMT5rhu0mWoujxxhMXgnfCLcjVYQBkxqDh2BXjZujg+tah8Z7Pk8M148
ZST42xrXPXpot2qc2nUg2oTTD6+rmX8KrXGdjLFndmzrbb8PsFEvlrKco+YzZCXn
ZYMlJkB/AFbfazD7klWL4q/aQy8MyRujms18bdGJ3ArbxmCNQwVx6bGm7CeX6c0a
nchaxbpDUqNFy/GgJ1EoeKCTnD/nRgkX9wdMXPuJnGV+GZi+W6RVw25/pB9XsX1E
yFRaIZOmq9DomIsB958p0+km2PpfFl4qklGGTHfZq8GkbFI14NjI4ndaSY5b3XLy
GdismuqPsYb6z4ZJei+gfu6k7jKCQFUtAR/JKrfOoT/b77huQmZVUPMPo0rLwIoV
eU2OfpWF3uOKefdeucS5Fq4Y0FGvmjXvO/Xa1IUF05qmVHXYR5pkF7ohQBVe3GS9
T+0DUQQdYWOtYTrXY/x4g4e69dBjrAY1nLVkJoqFnBhpQcT3LjV3r1V6Y9EfYWtU
HsGK8KvMeNvKxBYnQlaD/Y1xs6sTcpZWH0+G34RyDuW+Po74uH05HgeAyC4pUt9/
LbiMnL1a0/DfDhhx7taskVVotpvvhXCsC1xOxnvJ8gmFvozpPZCAwLc2oZ94qGOz
L60bX01aLSG5n840kbQUaEHH/27K6p2jZWgiYsAUFq07ZMrC5lsytWx4vsBIJed1
tuFxHZ708+hVs3DymbsoCWBHpZwWUFfvI5Za44ZLyboDV5qROgUUAYUZqsZ37GLm
mvSfddfzCa+g/Gh42uwSph+2P9x457J22HN/KySPLToZg8Zd9nkA0vwyd3sIB/9F
kvK7DZc1TuNCgivwMq8mwrkBeyzs1NaCCqMs0qVC7pda92pAkvR+zirnSV/Hsoi8
DZE6RPpFZIaytFKs+S3BoRAdsJG+cz2wO+ASN8q9NvhiDePPZuj5XnPTWHnFY0NN
O98lXMQ4R2nemWQX+ChI/Yc0/Oce6rZX+NEj3H1Vb0D83MtHS6HeFToK9zT8v4R5
gftbpxv6kxEil/s944jqulyJaus2qCF5LulaO3jGTf+6v0HCrP8txwNk7SGAeyrA
OoPaqrtCyKUz6HHIGZ+PqRd9Y74D8DSV0voIOqC9YiadsNsxcDWetrFIyimgGcFZ
7JiIRSAkhJpbMBFRCWyFWBPQGzNfI3E71/DqX2JsMUBx10rp4Y/LtaEQISN2fEay
ezbpC9Rf2KQpU0NMFZD/h2w0SnzEdUW9JowAwPZ3OTvJ0Z0y2HiGskNh1ZHxOC8o
Sxd2tR8Nyh3DrtY87C/GfHKVpR9+5RFWPkoezqVWwauiepUvQf9ofz6ZGdgQ02S1
pOB2wI6It+TGMQwsFPAkjKUOFnAoVlBysoD8FnJjP4IbHUyg50LKpy0Y67VAsSYu
xIMG4rKUBE/cIokDEBKo0fSrlIVcPZt20I/S0KREsRHm6mwVIgFMp4ozrOH8b3CB
blmuT38jInZQdqIeW13YYvwEtwuK942XSMi49Xj9VBWZlLigp2ijkRs1CqOx/Cdt
qSZfpVVZ37DMEnhTV1VZhb0uqxwocm9yAf6wzcU+Wqy9G2L/WhFVh9KTQMvID0TE
0XOgApSW30V3g76Z/FPjtfePHI6AhnQI3A+nhdotsQrDjqATWM/BSgiuZtG2Cif9
rn51G/aEVd8iXuIqJou1zSyaCfsmaTMVEEQuAdQHXglmx02M61yvlKqszqJTgyeo
RAw8P6VqX3GJETlv+8vgKMDR5QOOtZzMN5tP0bbHCekLLeH4mgN1L2DxiX5AgO82
onoGiDZQE0lGOyOKYwRMp5xf4KZ90TrH0xO/h/ZZsyEuxa0NlOO5TE3WYxZICNde
BQIqettAU+THKrqE7NTmONdI/RVDQzj3EWT2y9E9vyeA68jjtwd5HbsQ2g+V2o7P
9X8QZrPSk2mX9VF8cSwBhENV27aoZZNtAXyqAwExJZzWuDSFBf3jqEL8UPuhKOI0
K8M6ZVLsHcOkQdV7ENgYIWwlANPOtjP6dc5k5Mk9h2heGTMSJV+7bibTZW9cYLUR
1Fpguq5fBpKTgGl1qVv1sqe4XckABaWZppAlidJFyRBGH6JVGrq2ZzXrWLTcX9Ep
KnXVPG+OzIPpWO/FuG7KYLQy5y4LoX8P6ah6X420QohqPg5rDLPGHUq4qYbbDP2w
vAR5FnZygMyi7scZFGoj3pReKnlFJbcOcptYn2flauzmMzRG9am/yY8HtiuzXAca
BFGbGyKwxAcq8P23y2g1KYY2SxtZBl29UDjkfiqLTLUhYSxit7f4JMXWFS4Qvu8P
LPKJLIv4eNRq9MvtoDpkHBsHj9+XunS+LsxjmqVqn0K05WpoHx2bEG4K3ZIDfzkk
fuwJSkcLQQq2q0LzbAB4O2Z79kFSkoWkTz11Y4c3dvXHkMBVqdib4CEdMKulzpWl
VKkd3GVbKWwpdlHZ7NyNGzzh+EzsuKKfJusitOEqG6I8O5JUlrxi2an6wNeBYUWL
pEDBRGRG63touKlBRP69y/+bABFn1GJ854Toyvp9JqT/AJXEffdmipojpYE0mpv7
WaJf3raJ1+h/1c+sEPMXD2GkYhMWLzJcZOibtnm8pI2jqo6CbochOrTr2piE9mUX
5bbHN/Ckmt/5wJoYMuA+bxOJfwsw65WrUy3uyZPCTNZw5EieBO/YuwGhqdtZzaPx
4U7hX2QbH3eqBc94rRX506h8FyIJvOxopf4UzFmuY08eazWUm49MSNnT0HwQobSx
sjsvzSX8XMRBkTeOGc1lcKcy8vvUF1CF1knD9HhPK9+AOqsvfoLZ10Gbx1JXim51
8eogqQtL0YpTvo18W8v517/hqK6nBdpRiAt49gvsKafqmYXLF6xncjQT4WCbjPOp
iFQ1oj6MeKu8nhToRgLLs2R1tWKfNI6433DBfbGQRO/Dy21WSbqF+SUT3dpEeiu5
pe+yi+B1Z4MRShy4lvOif1Im6Zfe13jN86Ss+IT1klZlWjcMbAxDzM+zmm/jPKON
p1tH4+e9R8o0VQ5K7XAcvLXTHZoqtAkHRJAgUPNk4Y0Ad/pjr29V7yPBm+v3uS0t
F806MzBz30lsJnTmjb3ZXeYj3DzEw8h2NQMSKCRXDQ8FGeVx3PKBJXxmicr8ShLc
P//7CAGocV67O1Hp+XLlDwTbI38QBUJJZzmYs9fe0uWR7SH8UYBYceb8rKEyZzUB
FirXs4zQP2cRZm3OMpyHubcbacvXkY5JrsRTHtGy1IpCVeGICKfOI0RywExogB3J
5q/2v6Dp84pm+vXba8KFO5DPExtZschWREEJPHvEyF2IE+EPEl/2hstBXmfYp7yV
QiKfS0iwMnGHcK0Pbxk3ZBNsEB1RR7EYmm7scehtSDom2U4ydDxMpqaj7z+TE2gG
kG7SX7O9hXliOjFNHt0vgHLXjItNrfu78MkWcx4IgUfI1sIo4XbRiU9sz/pKIQuX
HqrLVbGIkYO4CUlWy3v6DWcjJLOADHFcGmvdTRr4wRnnuuArZ4KBt3BXTeVgEtyl
ZNyYJLd6Q1CHh/NZlLEU/I/xkEOxgfPwHwB/n4NXzbGJlE7ceXc47awpqtzVD8w7
BPeWJS1e3Dxh+J0ggZ/5Oo/d+OJVyNT+t0sO144D1VKxrgJB/NzXpxERcodO8zcB
BOkJyYwJTulI0093RRKePKKWmtUTx2AC4VlloNk+wF94oEDgQnQ2c/B/XOVM4uZR
6xK07N+ydljVjdc5atjC/ynywg8ueCXO3hpYQUVtHN0rpa4YpD/s4oulOQ2Jq+6C
brvCaLH8PLpHoVnALZnKQDGOki8jE0Imfgmv2Xeu8anJjUWA30qyZH+wPw1y0sRx
0JtC04XqQn/iVnCToRI1UBIujmHzSoroQXDC6i25o5zEiNkaT7guO2gFO4up5ShG
0Dfocx6Wtk3motDlwVozQ0kLJyRn6YxuKyxZTjDRX/Fv5KpsTzRcY2Wb+B8at5Kw
ofDHtSCWIq9elAU+VhomyflZdR7o/b412GzbRvVbWIgFmtg6uq3AXGz2dgsDC/Lm
H1tNRT+T+XuujhFnijt3IOTmD+cY684ZJi19/NPlU+MOrjex0EGIGjDFuRMcR2Ce
saTolKmzWhqNEpd77NY+pIBYZ/pgZFYkKftnanaDCicDuBT4cwJ7FfK6u/KW43TZ
m8yi5lBigBHF06M5P39NS2dR1EBSFvhJMCy7/Uvs1BA1UT3Tm/spWVkjPFQjUlow
bMLhTKZeqTq5hKVutEYezIgpKdtBVv3vAkoSUuvVtW3xtbMfus1DrqrfaBI5WpWD
v9udaJe9u1mGhG7Xr889cC0BMdBS2JG6spO/pajgHy3o1a1r+gDH2x9ErrLOc/af
gWrlJGRUYLLeI5b4dGS1bEPTvLJqHUbRouoAznBq45ylWdqz5Em3ZLE6zIAeA0nW
rUAMnyx9Gq1Mv0RwR9PCx1hBbN4Vj15IA9UvGM+10a0ZtJEGSkdQMpkfeoSrj1zz
E+bmrVYRwBma0/5xdotku8Sj1/s4t4Fq8fDykQSLOJ4YbO6oUa5YfO6G7Fp9nnMt
XEgTbJBQENZ0REqIXrNzknzf/MGFVeD5F2fsOio/PEdJO5zSvUOYIPoXAxE9kCVG
RYI5rhRDWNSw+I1v5qacrKRSA6CDTY+TBda5C+i+gTPM8+4CCoHwl7j3+bkqCPTe
97UorlAfzCYjcCZDeggfbxdf/hl9SGGSj/T7tO3Xjh7aBu6lIs/mbyg7IXSyaXlV
QNceRr1/rXpT+4cahNAV9TxlAVq9moqIZ4FmtNyOpA874PL3E30tLBZZWZYRmGix
hsmKMJVQSS2gXDcMkHdoEtz1Ym0CWAGl1PsDTVpUKgeiRne3mYhQy2PgP3z7FKYN
5Rx4/YT3YwCezci5PS7lDMSNf+A/U/xkxCy0vTXeu33+V4gMh1TFdTqxjIllXnoJ
rYiM2ql2FSHyAwKs/RlB2NwyUHG15Tf4jkjAjIIwvBZrwOkhHhKayLrP8SalsLB6
qtBaQIZD/9F9TbfhXsZs+0lHI7vW9+avcmxxLrkn+zLyhpFYuR+sp2U3noJO+A9S
CuWRhaVGrVGTw4YgGNzMlcDufb0+st5yI8cQvUnspuwnMGlSAwO+kOVCT62egQpl
/PnDxpV3PADm0YDQrERndw8bmc3IjNH+rkncDWOB0yK/Y+ksRoVpVKDB9H+s5m3E
go9w0h6Ug8EMwcRWkzfqdjlsxsmFeL9hLP9+lvVQ9/OFfpF6LKioZSywzKDSXSRv
Ia2udaf652LijyQhFnBjp9epXSaCH5VcfMASZS60cD/Tpc+Me4ZXi1eA/eDLeq7R
cJdCaHiGXlhS4LPROo8ucvX5x1q+N1BZPEDrq8PzZprpQ9JMywwLC1lTxOmXQepL
8f+n9hzj3i1c66znW24kjCqY+8mgyUrM+E9j6JF91cSrrdKVePJrQ0yVXTZc5h77
R/hpcs8jf8vRShW9ZfdPn92ITzTxzF0VrIybQrFTxlK43QjJ7SlDuqowvTCtB9ZR
hdDPcg4b+rFlqd1mvlYoKnytKjZiWsOQ3M1D9OvyEoE8WNTGZ3nTKc6+FIMsKPEf
/aBmkCmeODU0e/gIsFp4gSBD+S1IyK87QxLzCMsjLi6Bz6DnFvVSzEzLPsE+n5xN
XO5LLaG5dpnKd6Twf0/boSONZV6XG0Cq1cNVzEu7m5xGBTHjR5dNxhtetXu8rFtk
ykkXHG94TFssU9TY9KjHeyoeALjw4xIlsIshTMRWSnlTJbyJjLggigNNmeEqmnQ6
3zt5x98dJ16Sr61/To98LFL9kf/hkwcJt0mISk0Q6JqbhAbirwSpt+YUEvu7mfdk
z7PAnpno+eJgvZt1ygHsMSdsiinwD1T5+bR/vcKWm9qu4ZYF8TfTcoPdkke/0e6X
5cxG/wcmkERd4LJ/zlM4J1N3R5O1psQMLODPBOLsCSTp0J/yFjuKa6VvC9kMwSUZ
GJdLSV6YNP3vJttX+TxP5CbsWy9Ef2I9e8wnOypxK4QB3MdSbtcBMZeefVLESW8C
HY7U2kdYdTrgplRAVAtR//pOOOAgRdpdcbV3VtRJwucN56hQqWvT82ovSJbJi0Ku
+eYcUY/gezoVLcwDRgW6vzYib0AOg93QDsR9qRvAgjhmIuHmFF6LI+INP52B7PRq
smMWwj1f5O6GLyVInS5ATBk5+qo4hRsSF7Lgn0FpnRnztBzmNh7LjFYar2JYUNbk
/tbPnjAN9+WNvpodDefHUByJMlpkmAdeMPoR/6o9I96drF19zvJPl9T2xFiSf9SV
A1opFFNSw4OMPXnh693rKn0UafqqIZO+oZ96JF9k0DqoEcaxSjoorpO0GifA4JnR
pHGiLKWVEUMTzHYgPbT3fR4G0VbnObJeU2L1gZDZPpkR21tXt0qkb9ZJC9bJrRr0
AxKG17Zg20EqlKskNGYyBgPUZ3C0SYzfYPnn4egqLLlh6ScQ4b0CO4Ga/yeTb8NJ
eh7jEaDmGZzHlX+3Il1wlNsL+NRp2x0knu1iSlXdABwirf5aGizfujOXGnrHFYpK
dWs31BTN4aLfj/iszZBflukyGLTnZOdc8tL42ZU0Hxv3g+OlQ5KFXYE1OYLbiAaQ
qcwU1/bFpIEN9oCVp7gQQ9sg3d4Z7rYPtiE8EDsrjrh+exmWqugwIzeE1farn/OW
qvgbn0jDesWYSh4H5J/NxnmU3vY2InDDZ8A1S5nHDSfWWu+ijv26IeiUSVa4sq7w
O3acsRaB1ojMGOjS2ufUD3sVRult1d7oQGdoqb6AD6yvKfXiovvHp7dGicylNDNU
nJsCf/vJ7x5Znj8huhI7hyxS4oCGvulRJSCxB5XnrIAI68Bdl8mv9pc13cUert9p
PY0oMSfdVFqROPVYHtsgRpR+vwotYxGfAI1ihQiEn9xIae4VIPJUzcu+zGemm4Yv
7PJZKOK7xKvujww57p2rgaG5aoEmtJw54x6GqUFE0qdzvz7uZagSxTYZBarcouGf
KUiOTy1Jm/gGZanMrsQV8+HD7D0Q7i9SFUooYMjjzVOzYTRWqlZVRarKuKYNVi7e
HtGLDUjTvUJJFbMJbToj5dLg19pnmVEcQjTB3YqTDB+ss5m7848apnLWOzqvLosP
Hr9VxdhapACa1CDSLgNHlw+0KAbQp3zktUn77q2j2l8rWhZrwJ9BeZY1jjMGAnZo
Pz7a8dk3iKigPpixIud7xoa/rCzesgnQINxctEfl8Vwg27HZRW/zvi8vUtQI6vq0
5nVWWLw7t/pPhJhHinbCFGKO+rZEB/1v22yiLmeLa6df+gayuoZgKTLWz78DwHmf
Q5m/3sw6LzM6w7jeuwYwQwTozMDOs1r2AhLTIbmpjfHZe9lJDthUCHLLQvOMG/Lo
1v1rodhHNA1YucZhOGB5BpDLiTOpvD9x1qhtx6Fi50QZE8h2kmprjJEkL2qTimkE
SMQ0Uv680JCx6NcQNSVEnrOeYxxd0wtlEdNk1V2go1OxJPWHyIupqXUgNZ8STai7
TC3JjoacqOIJOh1V9wa1AFVpweFZTEt/ef2sRw0fkElDtBLGkIytbU0BmjbT+PzS
kZk/EAsow9YvKeKm6F/r/xoJpgrNdukdFr/R1ZfGqfiWB5ISBryes8WQpmqtLAlc
LUCiT/+lztdE6l9/kn590/NpxIKs6EweROaDxaCNBXmc12eQznrJrN8J0WKDP/Zq
C2DwWIWnwK2F3Ub1iVg1eMoFZnTjHn+cEI1p3Di0EcLmwG+3CIsDBnz6mRobZ8Rd
hOcWgeCCMnr8vdfwtmdBDk53zeyXZU3E3cVvhwqblK19L74Q1Fw+eF2mJXCyYo4X
5eHCErUHbDja4KGTL3syD6bYLqpAWWad2fJ9dSeUiwaNWOTUB2LRT+pIgE9pxPd1
p+4FT2VBRChDl1wIqi2POPXYmQtE0UIU426gQtR4bR51I/Sym2LMMftxd6mnLA7Y
XDsqEzXQ5WEaQCajA8SuRkkqAYiEHJ5RCIiJyu+kuqliGeBlJJqz53WOTU1fC3Ms
RaCC4/0Ic/mQ7OeDnGmcm0yHMhUkLUjcAXuVe8eWbNgsYXTQrFtVAH5oFv8uta+X
frD56rl0i4D6HzV6da2iylYmH33gp2JTmq4EJguRQ7A04gIzrkbo1jSSlCtMC/5C
Ack8uIrDcF+0/X5+MPC1wxrWKxJlIQumkPS78ZizeQMkBWzob1kIpW8fh/3Dj/qn
rOGT9KRVwESKTHJYAXqqq85qpqhlaAHvjmJDtaS7209/FZYaJg8LQWF+aEpJwsFJ
JbJ/Igg7HQlEASqGxD7xySWOnAFzkz8aOtEeCZQfI3OPWmcgpGFU8i0/So0zwKjQ
6kxovf1jRDQh4w8gfat6OGwktui+aWNb+4EF1lJmFhwZMJR6DAkDyOC88RB9wFCJ
OIzL7UGkut7mkspi7R/NwmMPkT7liL3Ek2YgVQIv2wV6vltkBwucSYAvZswhIT7l
oLLRtsODTsGW8OY4PmxHRw3XuuCbl6YoHDHKzqWPIk+hBjBTE+KRZKq9YPZNTad+
FvAErl2Rjf7JcWo4jSGfbtMgHXcrqXWs/JT9q8ZqjoJjqZhdHRkxMDAD+CE4QZBx
3PvX7OXhXT2KbAQtWsRFjLb3JW/KHzx6JeownNMATDhaanZXHjGZ107NxDbqxudT
uFfvQVCtnnqgAAPaS5xZjS2U65Ifr+8zv8dZBVyT4MlVlXTakz99cz3XdhB/Ov2a
yT+UV9yMRJwGIa8+bb7fAt7B8mqdmFduIEc/YqkYQdTK/w0H00hlln8INoeQUsue
exhlpmSE6bw7Mi9rZ3ImfE513tZUXOddy0nqVml7eJLWU60Hjzb4HKQwZTvw7ulh
DjOnWiI0moGWuE66dXQWlhDNBWOk59YgTnxl7yaUO6e8gWuli3kmLHTFbtRa4WJn
EMaa38iIaSSk+5mnwt1jPN0b0tIa1UYBpaxA5b3M4kRsSDcbFC2bzlB2guc4uGll
eHJaZn1IN6XK5i1uY0e5MYBkj5+Uqftm7N3oHh0i8Ib4LjpxEqmk7a5N2sOTARho
rc4wheG8XdNmEPTAUzLXKzXQdMTOadI9J0uKvR1wV2YGt1I8dEBRHnBn1cF2Lvhu
R/Dx/JuII1WF/5RHy+biMm4z4RFoxkRMW2aNGgwLVIr4WbBcsCgh8zWIcdz9Mgol
TUGjrhNaTzZaS3njyCD4FSAOqSiSoNR8g75xvJVEkxNT+jTKOEhH3DcnTSp9MyBN
MUEgbCA7yXoLp6HWXxIy3wPB4nfpe6hjyEskzruBNxs8MJQfspZd516kBHww0wFb
TuZ52D57IidmtvQaMy7beCWsmTYsRKND77ZRO77hYpYFBnXo3qSo2uReJ2ALnJJ8
xn5k6L06QqGmNkhyDAwGH0wDXZR3My0+IzR44H00TPUqAiK5GmyGnh3Am0Eo8rlM
hVlVqo99b2pic8CT5iZ2vY8ZepJstv3lbrveixbn8Agbpj5NT+N/uIqtW2QoXPjz
5K6TiVKTZOoQLQQOSWj1sn8qZGogFWmFakvGbvBQ9oCdwxQq98VEyjH8pismkuYg
kSdLAXoXTtJaUpRuCE6Go92Cv+awk6/tuWZyYif8FrzgD36hnC2M9zrGZqnZ6qdh
53LI9ig8YWhGMVSkW3r+5Vp/vcOE0q0tcVEIjLNI1a0+Ut7FxtjdO8Cnjraxcat9
v1D3r4NB9YcP2b8zq6XcRctrNamCpC3JdQQBJhgtxLgIFGF8gMJyxXk/oG84zDux
zfA/R120O09ReTpTMhclLUATqILSeWrflbkVuQPoBg2Wft3bQ7vNqvlVP8GEPkaW
icEayxrRS8nC75eVm8VUyZmK3yIVd3Wt0KfL2M9/e6Lc9/vYCcqP0NRZWC7oa32S
JwWjAzgWBj0aP+GJnP0UitmcFAkLVm8bZuJ4LWFScV8rDO7hWEs7KTgUvH9l2oE8
aQ0rgkLlYs7PAP8o/cqr1oKhkBGRzANuEzimTdglSZIZWVdeyp+C3WfFjh3ZmsuS
PBhGAm7m+g7nDQ32g/evIzsLB8JBdihhLeGja/TQK796A7LJnWn+ATF4vRgxDoBB
gdCo7GbwDbRJQaOTM3YAYohzVtRXsvnwb5du4DwkW2n8+5zfL7M9plD4RU9uA6iF
GQiHgSxxC1c9GWPd/2YA+7AmlJLAXywvsiZywnMIkUDXzSmisPVblnidObTorC3J
xfy/L/KgnFs9Au3cp01h2xjruhqR6lqjTIDJSBcFRoHD2b6mXD925pQHxE1TFH0k
+deAyyhEQHB20j8GlnlIUjAmBx4zXpRMCFWE6MN99fnVqsipyHYXMcmzf/4SII/n
h23EjfLFANr4vcBtvaPav7SJvMTXMc6ll9FKg46fILsKdrdti43r/3LUzJQxSZEE
jt5Vs3QGOJy78yvsTfobpDS0BlLajvRiwniwqu/0K8qVODu7ZNWOCs4VPM3yy9Lu
EJ+uvcCaXdJmyBbp+HedBCXkRAVKy8cnII0IskzyKxQJsQJImGK/WUXx4lB66HR9
iqxywlv3pjKw1yLcwbUZi3C2sGTIR+hxe7Um8iZ8OUt9G6lIIOwaT/2a+ZbG8Kf1
`pragma protect end_protected
