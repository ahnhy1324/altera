// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tKtg1/zqsxlg+waaihBHqtykAHyq2vyeLVlepMw4hUbu6By8ZY38dBPbDUUnjbZm
rdfXbl4w2FbGsOzfwW9ig+TXtCBWSNKpGTAQIUE/hUb0E/cPReWg0gzVwSpNTAmr
+wWTJHH+fWfl2jSyJjHVejlizTMWVnnNblyxhef6GAo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 85936)
RUfXmAMe7Ho+iEWSQEw+10He14oRIhKvUYZIjNP1m2SKkzgxD2tVT8EpaZPiHW4W
sf1M0TXdT984wHjV7EJbnazHwLTjjrfai2aHXjAfXgRcPMoq8bxk0NnHGQSc6Brg
VQHcZSkc7JKx0Ll75Rn+pYXwJEG6zqWRaYLgJ54vU9jbj5RW3nho+AjfCzf4EGjl
So1GD+VG09qSR8Oj0crWm1yfZvOEy26jZDy3MXGrHLTGwyJvlVLeal4zH7ikrKeC
YUqVqueFRXil1NGyVBKmZCSb5ivBm/ev3fjoTkon3Cs96nDNY04tdAisms+akpd9
BdeJN6RT7Nd7FsF3nKOQZ29uvEC+5GFTME9Cvhy9GNvGAwnBbqldboixka1xEYEn
muAplB4LUFOHINvDqp6diPA6RxpUfEJa91hCeFAAWCvXpwOmNbwmgYMbG77Xwom5
BD+qyKaaAzfDi8Ug0mZBoIa9Sbv0krGx1aRM7KtzKugjXQF7qtlm1+Bg+q3TloCp
adroRXQhXdHPGEBKLlSslfngIFplmfB8i2zXqmpqFQksKPl7BozthiM2vAmMfwfZ
HLI+IeH2NV9SQHU8P+JiS0hlWPT31gyCiNbah0fK3iZncuInNSoLVaav+NiCIXFZ
lDZmpGTDiVbt3FSWA4RKf56aEliAYJJRW/jo5fVPeuR8pl+152KOxfzgnMMV9xl9
nOaawldZ1LGnAHw+ps8SBWcKF3Tp03FWPGYGfmeDzpw8x3to0fxsV83eY2s0zOda
t7ruRjRhELTLC3wHEknzkdCdzLxja8oX4OrNmfkv1rPRQ0HPkce7TFPOuHgOT4Lf
5geVmBF5pcH7kmkOjyw7f0FriVDQFbnSEYL8TbgZjuh3VlCBC1lQdKhxiqFH70N8
OI+lRGdC8/fB63K08g8rI7cWwbo9wQIof9Njw1LCpqWQPtByREAqkFXjSQBh09lb
l2V5AkUXO0qr7y0PsRDrU3zeLhNZ0K6YtbP7zhLOT6ClI/cXmQQVnvSkmTzU3Ti1
9zpyrVMTMQZ/M07TIghSRs1e5IFBHnER5VEwPO95frvsjfb/V1ZX/8P/3zBls08s
EFCPZ9YfX3Qt4H7ZTIbxkwrJB2ETBeWq3zVeTMC90KYR1OdfjkY06LRXOris8ole
eIxJMOtbWVABdmhvvk1Mni7AAKzEUV3v3etOrSOhbRYN6MBZN8iX1m6bwZ8/OOgj
sWhzMiIrAQlfTa5/X/BXNh4tFl/OpteeS+JLEt5PSLBS0U90cMVfkwh8Gl74GG7T
SGEKFvtKf0eYCHLadrpoWAndbIubhPo4RPSQB4D8tulyEDkmbOM/YKoRBk38VXmN
EGg9PR3Mt1de66o0D2z6/R3DLAPJspOU7cI80SIJiO2fVVSzLLPH3Qz28HRvQpcR
Mmv5WHleoRyY3gTbuZOz8XavM7T5JpnIw30efNaE2uQ/vbXt4NraFcQATcrIGek1
KhZ80lAQtf+Qgy952MMD+ay0x4WaOz85YFt+wL7KgSIuPitauMCIZryDC6PZ2pbQ
rGNd+6qU3VTh2dKLFoklfyL/pL/4wt0rPdPxmHDLcthmLI49qAVT36mcDvQ6qPtF
hk5QbtMS4g7MjGuXgaTBlfi7mKE7X92vM0237kEiHpwHFscZ/9FmRjAZjABqV1Qn
7ALvGtR8DlZalgjMAXWrwCPrXOL02jKeI9JlDHeXIKrHYy+TMciwxc87pkm7Ncni
rN6jN6yalSoIi/hw4ADBrGCe3VmW8LCL/W9KbHJdXWm7tdegxRcyvfVyJg5q9SG3
bnDgwUDJ4CIy+Mmh5MXd1+y7F+TfjzREbCt8pglhJi+TZJ81qF8M8Frzspg7i0XK
Y8wK++58LgNeGBg5Lvfsh5ntmP/fFLEU2S6zkdZ/LpR2eyPpPaIELYgMpKUIr30v
PqltHHYhtr6B1y1MCrfUi/FFz+rSZ7f+RmEuUw7AC1LpnukbDN7RyaDlLtDrpHaJ
laMZVK7Zq0oJdw1VR/3+yc/UyFMrvCOcw/dQXcsXplVHMjCO0EXJmMWcdcXf6GSn
4dLF1B/xjo2UWmnj8y3SD7VZHczGyksie5Ry++k/lz960KRJMvnisOMr51bIiqKO
tPQbFiGRyrr163oEM27wP8A0cdGHW79V4j33YErTyOHaJsW9gA3c7Cw04zBVxnxT
QEzBaSP1T0W7a2tGUUqQkAhM7Qc+7zhM/BlAAh5BlbuEeTU28AkZOKNkVmuKHf4F
fvb9hAlf44RosamOVtU9e1aVCPVrmzWGJhKYaUPqMjT6ecLMWMxdkHIn2dOMhJA3
wO0p6ry6XbK3FRgzHadtfUwS5qaFDh6KfmKqiCnk/WmAu0Xb7s8BJgdAa9puGK2/
cXyfesxuVib9R/EeYcdlpTYnOrVGQfZdjr0SmLHVcEndxQJnEDBNwUAlfHAWbsVk
YeJq/TQw0c9TXeI2oCqjb/7E137YkvAK5r0BJfxGUhUD5/5ETcSsyD0tq0+iZ9O4
OFQqJQ0b8ZQ9j3HQ6lwQ0i8Px5b44Q8XKAkT8VovQRxRDEa45B45ghaQYXzYdB7o
hlnMSdYRdWVhE7C2Vu6hiSpKfsv6v8SWIA9+b6kM1/PHd/T46eCztBmYCc2F2JYM
nl/6RfYwpDotj5s58J1iisI6Eq2AcesIrIzCDHL5kEuXlPNujAuQiWxLHnoxtBuh
2AX3i3Y4eAl7Ykaa24g6zqSpIhidz6TkFdmmJ3GBAbFctoPPM7bs2qAUaB1qxlhQ
QjxRJ/+bolrD889wXxwO7Z1td6LDNenykpaCbfkZNZjFfr46uBTMVKxnPrNqBVmW
WoiT+MXVT/ktBHkzvGv7jaamR8MmJcpz0mk9Jbj7ddZ5DNMoJ8154X3E3lSBGv82
8036qqfAB9FW91AzwQkTPk9g8R0DhXvtQfFghfkjkf86XwML14D4Lz0EjWUnYD0n
gmJheMkiUL1ENUxCDIQZ98BzPlWjFk+Qs9lteB80zgBkTCbOWapWoJeZQpa5MLHj
gJ3SKx23ht86yXA13k0cZ3RaANx5OHEy5jj07juFZ5CTJoQ1GKZhHiLVR8TJRTPn
apTvVZ4YJ7r78uRBUmG7hJRjc8iOg5XrY84Bo6ZrA/oInqy2Jzot7udnrbsbR6Uc
BENNwhd3cgvSHgzvk0kcENqeTVQ4t3uq4ZywlkG3C5kN/2qKxoT106tv6PTc82Z2
xFvZQUyLMxKsMeF32mSnyfF+PJhRjqE9nv7JHgL64D1zRHwU7p5BZuofGQnGkDHP
3DZ0dRg7NmtGM4TTjgnz3/b7UOBGDz6fhn8prHzRxiK1o2JOkE2nUT3mIKAyhJar
nLXO1ogUgOh3L6xLR1PjHpB2QAumNSnjegkPMS/TD8vVI+1ko3Cv7whqfGTvWzfq
gCMXj/uYuu5yQzuKVulBt/Ws/pIpBWtqnKtDdfb+sFReWsbngBkdjcujBbIR5Qq2
HVWydWQrjnZRLxUvgo2KglY+sa97NXyamS7RHjcl/CcEvSDfIaSHAk+nFVa9XWlH
fW2tMtRvisvRgjUxZELZABDUzsIRYcb1fasdAI7P7GhvBQQa1Dug09R3Ki6XUBPY
HrRoGCXaX5L2eh6Fb021mZeTBIZ27iX1Y7SapWNvV9pFECTKa4wt73xJYe//c3JC
4tXcQYA31KCdow9Ztu2JDuMx3b3PYTP/1CiHJ3xkBzOiS5vZ37BHqGuR1rAqkDec
Xjf8xLBeHeiSlXPvSLcSAHZSXkaiNxgD3ql+YiDWdRa3FX7lCscck1ctDERdxTdS
KRZ7BoDMcKASnwEFzpAfhwwBHeNV388Ntgq1sgTq/65iOh07JoSu/NlUqZyuiART
hQzzqaSIZZReRcMQI3CT7xGEhA590AJuM2vGL7pp/4acclEUSjwA6Kou2hQBTzer
JXZyC/AQS1ZZk41Mv4PUo+d7LDTdv8S78hAiwRGMeJB215oYVlWV/WLBm0X/R9wu
xE1s0g34bBvW1weafTSJ7DjPtY5zQHMN9M2QlxmeD6woNh3ClrJVZeGRg7y3BUdf
ZqpodSTxT+P9ZePRdT3BTpopdzdM7UZIgQrCH2U5Ja/VIyOzNDQZMooYNjoE/x+y
JgV1W96tEJMq4p81+p0tz3HJM7vYz7cr7L9yDWAkgCj0X3s9Qg/ARgzT3sg5Ajkb
yYZDSGbkq96axJoEXsMC3iiwPm/YblGuGr5O48fKb9+GBaBvAyBkLNpleLyy+GIp
QT5nUF6rc0rmm25fBLVV0YsCHuXRqtiTeLVZsslE7GreZLZIxmJKmnxR8bCSf+Pz
ik1cE8vQyO6jgV4yrg8+YCh5J0/JIqyYk3ptUXtjMMXtqX0Zi9Q6axvdbWJ/xzIq
TQZHh6l4yC87jTk7G3cziW3V7jVBbzZu01js40pOPWeAIBvjp9tRmmftVTxLeWFc
/gNGy04mwoD22IVqRuEi2IhBbJmGjx162JxwMiqErFQoybA6FHeRvNRLJ3HPvoR1
RU23C5YlW5eDCnvt8ca/KAxBVDBY/Hym8dyzoLHS9wOPDvPTWAcMQtqtvFbxzGz+
8LE53ckZSGmmwUEcZV/SwnafdrdTwNAqKH5XEZyBZulj8GYvbPetvAXXL06Jx6kp
ZsG9DXXIczbjJhs9Uv65s3h+eB63LpRw5B+Nnhw7ClgtOpcIuHryZx+iquih5ulD
hsoRwUMzXeJDQbHx8TdHRaE+vcT9CdGuqWA13Ki4rJypmmFv7VGu7XUhYls6JHj1
wHeXXu7twdiLNAw+6wZEZObmOhCxjDZteH++OSIIs91SrKxUsIYxGcipg3fz31r6
BTgMFuarbMj3cH7v8IXVMKNvYZNLWIMbj/UaHQ3nXqcMmhemE0o1j7a1/XFtDtQM
Hexek3ra3X160u0fw9GIVfkz1YUC/hMyvV8nemFX5VbJnImPDx3lgDG7w62SKtwQ
kkgOeECIZiZBI8LpAXfkY9iFMJ2rjybuEOgqUUIgto49TL5W2rt+N7XEQBsrsx39
FzC1HGflJYca5K6mdVFs3/f3/lmRSydTVNiF+esgunXy4RNYH+NrUw0gJvCzE7Iy
GKcCtiPXE3dEROqxV4kNBZ8dZuVxe20jcZxHjEnpbYJVmWKyCkZLy3DCxqnqvRPa
oXBoe/F+P8JWCyUCAviGFTmFUehDKPwCzOm006agILOQrycrXbNf7RuhwjRXyg5v
E9D1zHTchCTa1ZDjj9YpFXbKSTciispFk8Ekq7nLQgMxnLm+kxep3nrBizHS9TbZ
8uTt75Tm47ZgrC27Zk8v98oIf3GpacB4GAGUlfJp2gh4JcVTAf7DfrH6UZwS3lGx
iL85cT3x5ltligcELNWUpMgBIV4p/WO51C6E4vWqV19NBEl7BmD2L7N+Ddrp9vXo
1G3AVB64ypWR2l0xdVJN0qkAf4jYLzKEXavCRa5o2+R1dtsoskQOzEqzJo6biezY
3Ruyr4hiRMZiuHsxWr1I/x66zDqM4BLakOnjL/XkrIl1P0TKJF49+AsGI9cH6vHw
QFlJBKrmE5b9+g2FJWbuovw+W6gDWmFMIGhM/OS7JzwPM0R/all1Ihf6I0NFYCn2
2UjoC/47YfyWe6F+bylf62VJIujDLfCTz3LR9Gt9gw680rPL3LnuzUqsDk49xMV5
je523KetARJGhGC2OEanDAi69FyAkWZdE8ALeiEGAUvqUnaG45E3TQSQTSbkLAOV
rvx/NIfVZk/Rjet6IACXoEb3kvBIzOOBBZ334v/8Cn1CKk94gZRrjeD4f3uZE2mN
ihPLRXuwwypuNr3sJwKWX68hN9fU8mOxQKyIzJwo9mUfbsHKfyn8SAZG4SeIVtKx
m8KYwVxRwur7/S3xAb9JKbb4v3oGCr4AMq1iRR7GmEpVnYw8vn9jUCGogDjcMltu
GWoJhKVggwIZubt3qQji7jGKp/AfD1HKApgGS5GPmeHlvQwwo6q8wvpgW+DoklL6
P5EtuLS3mYAqzW7APioG8cE/sz3xca0SsZ8zjej6yUaS/SY2+lsCsg8HwABegLMr
+g2mZKw8/+qGIKh72NaYBilygKjFYWfVYLNxSamiDlNBIiqCh6sngr5hPMslwAxB
35o1q22Zzm8JPNIiSs57x3T+Sw7Kd7Zk9+Ra3cl+qxhuCmI78oRHWihNM2SbQbWj
IA1jJy6TFuhtiUBrqVjajMDSiAPtfpnEwee2XRvTtEvnbyKP12ORkw5KUW/SzYmU
OOAXlqE2iFIfxzdzl7XwWWG5rIZka8littTIbzrfGUfhqbl9tJI3h9s7Mq28wdud
pZ/OXYklQIuA7yeUtBEld/S/6kUixNAIGxQisa1l3tDERfIRkl/Mu6VzPrqL0ugz
ek+Cj/QjYDSK2/1C89pvnVe3s7URx+eyrWdR3ztRD/uATJJCi9M6f1DZvvV6pDWm
SEY4ZeyM3RCDD52cBJ3kaTi4ylQQgsRvBunvteCyRHn9iATmDl7nwRlQBAdoRsdV
sKOkpTJ7/YvL1ofGjp6AKJGiXj89Pxs+/dgYhEi3sLT9ldBNA5NuoK0rAqPlgDa9
j4+OinkpK42DXBT8JQmkE6KksfYAv/Mlw7X5YGMtNAAILHgBdnxZs6suYEJPC6qw
aM0e5iuCASiFtO1vPSa3vOW/Vxk55x/D3FT2lKnSrZ+xUkFx8hEdYKA0rwhJd8+O
78EbhW2SzP35QNYhZMOn+zSjEm6khd8JJsRlhVfP1kY+C04BFVIQ/6U/tu/ftyK9
/p4XvxCKtgAUtWEMNqE1vg4gRDD49G31J4c+7lTKTXKtCF+ksjgHO0mOfY9B+mh1
sQpxvV55p+OCF9HsZYTIKhkQH+/NnBlKox7K09rgMrXbPFv/FAueWPlP2FOsktUu
tsIsiEGmWtqCsD/4zAkddkBzSfEoLip7z6io79b4TJlmvPu98dL0rAUsboDKgHM0
fujatdzrNbgs0WTrLcw52ZcToelCiFEhwPo6ZxvN2TSVey85FBbhUzuSXd1QkBth
p2ikQ5Ah5tcVvSsns7IrD9/D11aYC15y7Dnr+gAbReMYhQAx4nif6Y6rDZsCKUeg
JRrRqEpFXrfO+rtl6wUcavquHWT2drH7Mgp37PSRXol8QFZQ9MssEjbC3lFEUR1d
UqtUCKnqvSDfkMWfi7/SUSEjsCmhMrUcQr6+lcD4/8SjtLVz2DAMKDtEiXG3o+HA
EaPYz5xBahCWmeF8LkCmgKHqB2jit8I5NSajZyzMZall5n3V+UfEuieBdyquqEbd
zpYWzh35bFLzHNGdHEeY4qJOWPiF1Zqh6C/F7soF2SyCQUjB7nUuFI6ybqBA0RL+
JizgctRYoTJvmHApT6J3hkzj5iQ/c0wmcc85vJrPzDnhlqY1kitNcFhVXH5XxLde
FClikFtQ9jIx9CSH9Yun6Xm4lW/kVN5FqULa1lAZA3ArgEIypC6zQJJ0FTurL3GH
W+UwNqQXNO2P7bbVbsZS0KWO+Rez07+WWy3PoOySX0hSDE4Zbv+VWSjLdGafwntq
hYwpc17VtKSxt5gxV7ZSBNA88R1dxFZggNRqEVOvJS8IYE92WKXID8cS27lKShoE
LVwqCwpWs3rFgiQzi0KSjdbfbk2gBQ0Vp/4Syxl1YvlHwMzv2KXfix3ghq0cvCZO
fxJnrwQ9/dl6NsBOvpJ9Ushc2RC+Ea6aDwnQhuwgWF0ZY/dSrE7eApUO9/2KK5gO
TnQ0rkuNNDJiTz/X9ySRGvZne7YvJ6sE8RcA8i0fO8iMdMxpWyBV/2pevT7QGIK5
qg874NUrRQdBY4KqDqPEjFpjvQh2dFLsKr2AAehiz5pFOwcyizFYNv/Cz6KUTMiW
zEUfZ8BaEpntr0avSoqoayvtxg2+Y13Y0NkzgiFqAZP3wAyboXpAz0yUYU2jT87r
ay1pQwoOwA5l8J3Lw8B9HfrzhWMhe3R6ARnp+hu5rwNmyFoNmDB/HW1MdvrpUmR1
Aw6DFNeneG2fBbevQZdVoisCTTA7Nk+WATpoc3+19vIAyjJNnV2QN8FSIehtP1VQ
tH7M1hxa/Pbe4FdN58Xu/1FMxLgkbUqmz02c2hXS2X91U1vK5W5H9MExe/3RYHxr
HpExxDLTN7aYYltNhuijFCY4mNB/Cx7VxaNeyJ3O2kroJkUmi9UtOcOKMGDv40pH
iyMOa/TgkCoeUmCxy3tp+JvIYuALC8EAkaLv6Ym2NrxHb8aTW5AWOSV/H2C8UcxI
zdt5aMySjbhGMdH56tV6ym4OrSudw5N2QPwiKir+ykE86QFPdafW/vzS1fBLxjdk
5m3B3eSM2vUH8CKAYEzFxRYWCyP1uQKXjkkav8NvJY4+MLPrcmOEwNYKm40L/F0t
pegCoVCrWI6wto6pSjpME9OSa49Hpp5zPFeiY7Vlw/J8A8Xtzp4O4gCtS9z2c5Ub
mZhq85fxmAA91OzPpF5MC9Dh0wVV5uomSaaNyxQeoaWXSkuq3HY0RSvrJ7FXt+sB
Sst50xHeTu1IA2Earq2EgWkcCppFJgaAfFaLB1RE4SIzUNVnaRHVlTs1wJ01hqCU
PBpD9XY03F2oDfoEBif90nizstFAbd6QXzqSexD4wiBrId4jgF6LxaNlGuiMf4bO
phNRTm15gE2jbYlgMQG6+AVrMuXVnQeenjYAJrMZT4jFgml3QVJlJhepYlRbbiHr
z9fiLiLfdqP47BrrXVqc6Y9W7Svv167JXvRpunAnlQf5X1Wui1Q+Zsk7wKgJWRhE
kKfoIk9RK0bIY8s0NSL+PVLzUPs9oMZwLPbXJirKdP6dY4o6exhQlVyRDI0QNFH6
knlazMAmmTLi/spvOqVL+9ND8kWXHpR73ZeGsY9TnwzhKQ7MsVY20q2vDJUtwPbD
oQ15XiVP3OszIFE6fT/GCSVvEmuSvMDATaOMLeVNYY6+U7qNROR5Qev3xZVJU6qF
mlWGfYrO99P/en9YJQgsJ5zrCQPlWgKv/jHMWjhbKZ2T0/BXN1wfQ1gqhhyskdpe
1OdZ4fFIPNoQbwtSb3OVBAfQxlJlWPVUBUrp+dY4aWk9TfBN34k4m85ngom1Mrkf
ZcKPen3UBDSWNxWV4DgGCZWW4mrajF2G4ow7rKkZdwXXWWCzBY13AKMxK03Z/QOo
GeQ111RyL4C/4DKeCH33DIQ1yj0IIQx9UT/EI1CsJ5mTEQtzNeIfj3wCCvY2+mSn
K/nWjjQj7gcQiXmU3BxobNATmYV2O3PbFDLG//7sSTmPWt4LdHjozDlbIjHYNlYW
+zyrr72oyo/BalCnLAuT1HEDfyjJAgIR4Fi4R705AsN4lRGCLp1B6g0uZMg37SpB
Hu6WT4FoOdnVj3c0AiWilyR54scUQ1Ly7f3MiOhoVoxve6HHoIB9XbsZctaZS1yg
7U8NvPr4RxCwMg3B+hrpAMrH0FBrU2+8L+7avsWM98KxETmWeg2nIefWXKez/7i0
LyrJO46SZMeMOA375CuaDZxroFn+e0v0tee0rjD5IvNdll5iRg3UkyMpJk06xYvO
+8haryUofWzl1F85c2n0xSNQg9RQpcuJzISRJmU3RKwBDHZf+rblCjejddnu1e60
MckuNA0eXxMCAZAEoX9DcqiF7iv364cdYRKN4mfdC0iXzzRme42+ye35lO/HQx5a
+/ztUN/rgjuWsTjqZMpnT+ejsmqzAOIeJVvNZozeYL9wrK0sjDxrS+H5Nj9w7l/m
b5/0XSzGxU7Q5JSHPzRO1B+RWX3MOCyfLCHvo2mOD7js1b29kXqRDExKjMqaxU6w
4liDmW2Bb7PUSzykZlR6l4h5mshaU/2ld/WSCHjK/q12FgICqpYtJgZrkXdS6z0g
u6uY5s6uCa83KFV7ElquKYaA/NThQ1SgMgghADIpz12nvyrmF3asUMEjrrdWW39Z
hg6Z4wxfuBQtnw0VQvGaogLUR0L9b0/x7WCg4c2r/zA7CigQMa5T005P0YOJQBgS
yKIwL/prddqQZG6DmRUhMKlL9/c3CEuqI1TDSHQgnSSyPLL6f1A5L/55Hi4kxZTL
KYz8ZFL+gi/6x2x5L5dKkoo4YAifjQAojWh6G6W+7TPi+8YL9wdn3E8Eby7NK/Cw
+rBTxuy3AWNMzgKust899nNcGbd9NPOZ6t7mO3twUFjqyR5FANV+GUs6tb9Eis2i
7r3IogoLLEP3Ck1yY/IkgpwcHu6nK38ZDRKp7iQ0KutBu3wahahN112N8BRvrn3W
6r9ygWGvvreVy3bvPZTBiDgwkZ4kbRJ/OvLqeTkpM8cKBlDe5JrVNfDGoGeOdSXq
U2MR3L5tRz6MUAj+YpYYEFEhcOS5L13Zs9uhIa3EDhoRUgAqdn3BWWX42mq4kPlb
7OimC6YIMzoLh3TCM+OUk544ZNk1XQtrU0XHvlo/C2Bor/oc/vOdGlVv2aQgtfgE
Qvvh7JqNa+2g7y3LUaZu/wou0mbvxk8fOTIiyR4SepsVQvzItnA3zAk4MGZFT1FL
N2bBFAOeemkGbMfCcO7FLcc0QVRPQdl7RQAeE0Bac5DvVhh19pztQw0sBTNbqwh1
tnJqTspo/53GH1ljoxVRo0lCSQAKcj/5l2q5CVWH4GtDNWVsbbvw+gEH6lijuG5N
XKE84mkETBJuSqtAvFfc07Ivbt1BRBmIHK+V8Btt1vUwH037ohWPKVgdgGaw+6O9
SVS9M/NVWiUJp6tpM1YCmfi97tiqPQRhsrd49sAxnnGywRK2arSUfGdaOiRCk/ei
/QG3ermZLBzdHKNZt6aFWGIlQ9OVWnsgRDOgNSplLey+amEMPpMG6nu/uwz2QgQu
Sj+0MuazN0eSXxK+rXVLsRK3VySpgDOCMEhhxna6HjIkeftnzB3qJZ6YPWOB/n2z
142nWkBIyEztiNJ2uNokf244GdOt9j6KIYscnvQNhvnaBUq1/5044Ns+2pA0xzyi
016bvW9Utgj0sLAK92v/Raz0p5za5Tmc9dy0r1lv9v/YvxzB9n16Vykgbyp7SFIQ
RnsbA6QHRhrFnYctY6a3uRyyNZEcNR9x3u7BUtWaBDDM7RUNfULPMa99jkaEz9Ib
KZbjzPM7muFniLFcnRj8Er8zNYeFCRJXGe9YFzF9LZPxlek7EbXgyZ1Db4Xniggh
tT8Gx5HJUKnzTCux3saZKJhIr677rEnw0lw8AztgcD/HoYP6TO8Un8RgF6akkoAY
izKZznXnrOYPTm8HNhft4OTN6dDEPDkJ3/PI8ljlqKQFBbyArQ1O0nAB1pzOGGu9
kBuriBh97wcLYN2XbNKhqS/b9EEq+NvsHJH+uLtrwr1XiRhkKbZ2F1x5r2xkWQRg
GGExDFy9V/tD1HAb9u5q47mRV4L9MvpEUrZ3+j8/IDgwHT9NN8cMcBkITqh7L9B9
yP8srPk+UgguqeOPjq7UtCDBGV6VUu1fpdtC5UhAN2QdLbdctznSpK4+UquniVtG
7/ORWO4FfkOYvErrLKYFP99X4j9qXl48bPNm36+FfF6a9jiwU4gtwn/6qz0v34jD
LK/rQOOCMSrNXQ/f8LazBgunZAanqJL5A3EOGowY38CHzrYv1khqlCzQwyWmb/BT
aV0jqGdAe2dNhtoa6rFrN/ofvJ7yMW0jPJYOUXEMM3TgUIoF4xsOQ3HLSOwsjQ99
V7f2u3y8uedQpaFIulmYboDjWiNHkDyIgbNZLYK4Hawx25+PeiBZg+m7C35fbSKh
MGYJrF7UWnw0wug1g7oN5PM9MmaZdN68kSC3aYPsjxYDFFSza3l2xiYYjthiIR5F
lu/h+M8W1gxKEJuW8FFx22RvKwkBhLrVEpLR95wNV+SUlA4OiVW1TLssvPKrQ77Y
BdSf9hhq2M/IyKle+tF7zwSV02jdWLqek8X14S+57b2Ddworqv6v9BBZA0/LaVxr
Zx3iyPv/OptvPe36dQZYcXTIie2MdyVmzRSBB+nl5kfSIRKQL4LuxKm4oSLRaHmT
GsSNinj63WlTYKTsOmML1YMDN6xyng0BfvKbsume8dBL25KuKsxqTPLQJo2GVEYy
5nuekszvCr3RWKHlvjuVkUwKq4UI9lJ03RvcNdX4DO9SpR81v5FQNOKBpe5P9Frk
VopIUlI2wFKrQzMiYoPWwDPzIP1E01/gx6Iafpgjsm45CgraEw+hAKJS7YX93IV0
eaAOFF0Fxx15EjGp8d1Bbq35m2fxOgYcuU18iD3z5+FoAgG5nuLlIbtq/BOCcxXF
gMMlDaz6RpZ2YrXlc9IFh7IDuHV//nbCufAgxYG8SH39mYmxmOECplEBr+WEa1BJ
PWMmuzOMbVFfh/uEoHBFKsNleYNSCeIoV7ar/9SA7sg1r2J5MIY93+HbLHT96kuA
tyMXSYjiLNuwZdnBWhpglCOcU/ElbF3P93vBK9DBl8+q+aT+RjSHrE6wy/c7qb+G
Jk8ql6SOu7hRHNhS0evg93BetnZptAWNBNlTRsmdPmy24BMBUJY/F9/+Zg2FqT1U
pHkkwK1cs2xIY/qKaARlQzNLdP8x8tyjOZkcOgErZupwfSWsZxTIFRe8S5OvykAu
LwK+LJihJA7DCU4g1zVHI5ICWaJ2CA9HAlEwebkGwyjXKTPfaJDNYljybzBZlakR
vhwLs8wb4v/G02gVMame2qrcsFTFZZemV18QxZrO6IdhiEso82Kl0ie/MCcmSi5a
kM1aWnxMFUjzL1JYlnXCcP5G1AK3eP/pRJPM9wkAF1UNfXgPn4qnxheUNk8B821F
cHphA7+jaFfWk634p9EWP/vzEj1NkMI+Ij8aGqgztM6LslpdpZyHbfXkfJtkzV+I
L+heL2a1R/Do3vggYo/AVYkS7Eloep9LfVCvzx98LSifGqJcDmOLYNc6N0OsDGPh
zlfUOWaESStbv4mL4Wav0JFN9ENtOxdpNe1cEsVTjCxXqArGdLSGsZb8ZLtzie8k
JfYRwh5MHnMeWFOoP/0QAlVX4Q7sDK1jBBKCj4Ox1D8CUPrOcWaf+xy75wZAmjFI
JCUVfUl+D9/BLrLq0wCUHGlhnXZj2Xc8InQTsGn6mYVeAyJXKRZCe2Kle1cRYXaU
v0kHbE8wWdxIu8Eqarg+3nbJM1qdfLIRfX5tvhnj205fQv92QFMJ0FyJpeQd7SJE
rI67irYXei/fIwU4gUT2Duw0Ssm7yl9poHfi3aLu2+26wtjqG1F3IZdd7/4yNU7i
LWetONi/jkW2i2gpfIVq4j5wiL8l1HobhaGB6kV8tRFt1JPS658koXeTW3ehWxY4
HA5/blnsOZNAe77r+Na5rolgBYiD0SOY1WFlJFDZxewBIF360yVgbTAH8o5sABs0
pgfSE1/cWL0/6Ow536T53YwjjCNT4QWqYsk8/flg+aeelyko6FL50k7qZxpeDXLM
n4Qw4FK6o1WgyKOaEfn24M4ApQkNE44mOYX3tFbrktwHLONVi6sWpwdQooONNL7f
oQ0iZ7+Co+PbkMsSKPymXKhik+82h2Uno4rZQ6r5FPqvoBl4HknFrwvL0mxUnYEK
GyNJQ73/uAcrBCCfiQj1gu2P0LBZXkmZCB6yR8fKn/6Y15wLoTVjTDNNrtH8dSSc
YHDEW4dq4iS9hYc7RDeI8U2E5W0B96nLAtjFsm+F6mlP2KQ0Ow7qPGjwK9jR7XHQ
GkkTpovJvdVAvjzqPflR9UicGZiI/szLhI4KArLhxSXXlgDmKagah9/PGc8yrfYb
4Ws73fabu/QqCqfODQIA9bBdCczDMmlZ+wxk4FC/+rqRxtEj8wkeKsG9bIE9yEHi
+VnUGjkhIp7NjeFmKqqnjO4LBj9+Wa7DT8o5v01XegzRSdjcy83Y32W1rcl5sxZY
K/ON2Aq6fq2NtUQh9xXFoEnAeR7XblKXQetJU5a5Xfef8PY9unu/sQMhBJ2bYZxn
Zamt/R+euNnnAkP5IrjneWjfyn/+NNaeHOj7l5c374+zH0QTlFe+1oIuAiwR+bI/
lThN5mJ3OHN6FghGIx3SZOl8Vk20zHdPza6iVEA35wV0H5Ewk0GsqJ3gw4sQb2zj
Q4WWuzpCZ1ROuU5nylh1/0t86Nfs9BePT8T+8UdXz0zeVf7CzkOA6tARVp7d4pXE
LfWrCXvxLPtpS4nX1wYFvz6JaNEFCC8xNECzaaA5XSFXt9e3WiiQ3r3mw1Ef0LCf
2oplhVzxtEruXUdu1+xqS0rJJviBmlu4YEG1qhKpMF4UPe5ufgveMwWntGBnwRmJ
UGXmyIVQ+UmRY4/mLJ8CVhjnmrKz9laIwdm8C7hW2xshE8aKhQ/YaD0S7JRUApll
R7vuXbsojSzs7rloBnNWZ1kGxuvWY5cPwKQwiu9hyn7UVr3WVZbdY8BGWineqzWy
bdRzYgRAezeL8yHZqc9c+omisWRVW8gmF06a+h6BmKDVvOTsX216CR7f5IzQx/12
y82w4uIu7j2xSgU71fc/Z3Fo9TCOilgWJou46/9pnPUk9pHHY9eliCqhCdZdqmrS
H74BVMa0deQ1GdUcpFYQH5NI1r/og0oMqwo/MmM0W7beMrO2v610LQv19+SPgXQ3
9d9u5x7ndNcHcEhG/mrGps8mYMRCvJJsJUY3n3asEtBZliQCC/b+EnwjqyAF5Sfl
1UACt7NBm3gLLvWzI6tuEFbP8fI8p2nGNuGhy1xRSU3FL26goFBiE0LQN0l0mVUw
UOZqpmMm9JD0MhT1D9IesSFbnqrF6DZYe1OaihBIABhj7pykrj4O4iOvK6WEkXR6
QccHlJ3ndqWCgThahNtU5toSMSIRZCj5i2qBzIM3ge9OVnzk6AhDDeravN81iJaw
zwZK0Jp0HB0Q3RWL77QuIzTm8RhsEyKhGrlUs5OKV2xeswNr64BW2HDBpyogL1ip
JrZfehLeMTsBwLJVlX7rvJXFKZvrTdnUK+VydYFGeSKfU6gOTUed9DJd0f/l/Ms7
+6IMlDoALGvdJ3A7VjCvySxkhgvD7gCnwXKu9d+EMi2Qnk/Qj5WFoNSTK65AENym
6J4YCM60D36s/UxsshsXHPgRkjPnfJsA54zu8f8ajwoUauPc/MisxUHKDCFzotIt
E7puSRtUH6+oroAvKF5y4ppi/XaPaf+z2EyZ9vrwglDOToWUSvhDuVqTS/g3q+Z/
yiV/IzDp7khkH/78pYYrbT9DvU8MEjKepDfqLkdYbgauVNnOMB4m9AcmvCkW6anW
JnEHqKTZxGIEck5AFsUfk4xOIZ/5sW9R6w7Nn1WDHLoRPNlM/tgLZ/Tuv7m9WQ8u
AMeksqJCRjfuaTlXSpsoMn0DG2gK/zPMgKb5MCRx82sedyWFTpiliNXCCpTTBWsw
/WLHkOsQ+6ekc/oV08L+naoUWqZoqYnjHhfuK/9IqhArvmXlhraUh3Penv1tfDid
1lSx4gxVZ1KJLEHEikAVXzX6OHqI7Ldcry8+IqO8rHuJFz1wEQhp9uYXeQcP/JD1
v/iBxRXS6S2kpMMjffDnX09ksD/BvC77SddTh7I2SAiqvS2lYTFTGQ7RQfKfbZcY
6RZGXuzTEDfN2XZT+eM9XIiQo+l878m/tHpLmtPpEAbcgU/l3QXrrkwe6YV6ZaYn
I4k1Mp8/vhGSbRuO0qalQAzCckP+AvlQI2PfZy0qmzix7UMlGHbjPFcKN+YKymxV
+cPAXCk1sFU50Nhgau2c47TmGWWg6DwYH+CtZlJuwzmx/heDiesVesOaSPPlpW/I
NTgUPhXT0N7GpfwFywNGp66XphklGy4kf6PTexL6nJeJvya3+Jz8EH+OrAwLgSbT
R/5aRper3i+RjpTc7/KB3bAi+8b0rkL6gyBqqdscM5ndSQyvA2ILYWccu8C3VIwc
GcW/U1o0uFEB+rxUUmzxn8yLGeJuuc4gNnBiv7u/bMOjqGNDIBgcuGQtXgNc6CLK
KNUW8VGXWb5PmD48Yku0X/H0t1FUtOsgF9/AhVvtOOPIjKT6NA+6/A2AitcqtJFu
YNqIA+uAU8/qnSEWEwvrnV6qtdSN4VF5i4/KJhrVhsYTaOqoi/hIU1GVo9Q7iJ4x
lyHeUNsBVAVNUjqGurLTEdVwrCh+lkbZrsnjUO1DjgMilgsLCptApiOZ9TA4cVkX
tsHcpcgoJN50ZhJ46nSrJUG/AvcfqQilgScnX1coPG7jJEWNoNCSVqKvVHfdtKID
zIuigezMMN+eGRYCX/6b34mrvC3sZ6n7WGH7OBVoz7KlE4RZ7r5C2I5DonFmfK/K
uwNmpVi6YvqCjkGwiJ4tOYOL0DP23UoWhurhj616t76l7gmrf8mjIvA2+q0QHtLM
eN+qBqi0fzbDJTEJQM3GXKKd315L1ib2Qq7rfy7rueLTeNL5pKp4sUnZk5OeKSjf
AeMQHUV7Tc93BMJcZYKX+2Zf1OaZwf4zythF0lKW3ClneZ+HEJ+gCE1IBeLOJB1n
ka8cGHioU7xTzKuSpt6ip1BSSpcq8KcMUKegQZi6FWVnU3aDuAHS7xFdGJCkvWeH
pXvsqRyIPrwbLBOZVdC5GpZi+S71NJoKnIIxTKbyMJb4Zvk1LnAwytFp178xk3sM
mszROKfwHSp40/s6G5F4gFJHpK4pSUZotTLZYDrAV4T+LbxNUtidrVHfBZoacXfx
5FmYQbhYaK1qNUw5FU3lFdE0ykQJFSG7ZdeW4nBkAsLGwe3WJdEL0fY3O9W0BcZS
TPqx7uOB78RlL8zWdALhJfrVQCtq7lbnP06l+O4FWVp1N59WfO6vvLpFpMJCW8OT
RvE3lYr5gj5QoLSicAvLrfqe6Fsp0oGHadr8ksGjJwcnnHhyD6cij8Nnq9rffx0S
WUwidPJGeF6jJ7UjTlJvnchkSmKZAKa7q2GiDwC3fDugLD3IfautvMwDSI7g66/s
I9P41t8RID+bf/bCDPHnA9cg8ND/cQo8WikXKZ9y2A43yMibIgEsLV/bWmTuls4+
5Lp+ablpDyYIf1WnDvQVzd7/tr2rzCJ6sHDXcAC3pffMZAjIzJXjOCjPjEbQvHIn
qYF3chhcbs6/2iEMOK+iMwfP6Y2tnc9rs2RTBUK1PYXNcZh86i7EqFGTTCUxEzjk
vflnRqRH8AuR5a62fYLno9K1CTsBMN520+TUgv50xYkUoHBpww7a86qMnPT5jB90
O7f1YnkXGafFkuEwNIgM5/M+e1V7H5CyoV6OP3sX13lXjUnZK+JWKZ+Oj9yQvK/M
q4u41Sz+TX23gp19KKeVLRKfU8VAkgNs01cLnZq+kVO1j2DShwrkyBJvvAYEIVJl
BqEwGoYug+4IuPMKgq21NchI8HcMQoMxK5spwfUK/ajIAMnhfoVxB7Y3a72m9+8Y
PEZShLLGM1usfTNQK1I+Cv7+fxkhoFosVhLUl3Gd3FnD0LbdRA+5frWICrCLeh9e
kYU+46HNZ8A9i3IhIxAoS2Kat7cuWTIMb1DSvuLRQ0TgKF1LSTZLX2E1AwbxHF0/
ix3pe62w5YD1fO3gY6Iiprb5mX0RGxUFog1LUBdSxYPPvLqTZrnBs4YmoQU1h0AC
OsJg6VCMD7DmTX4/3zueMIJFb9wvK4BXaNmsafEhabAwgAqTxzLx1GjsLArmZw8H
wb1nwDej2914lsxJB7XAt0tL7g2IEPyI1mMN1VOzINZI9tho8EosDw7uW9RO74ns
DqasdexsGdT+m1SXtSZnrwymnvMCtwLVTt3g8wRv6QKF7ExmC9y9f4Sa9nm9dnae
EaLhnKSeLc5GOL5syB+0Qg0lChGA9aOMVKXejHxwcFf5AomN9d7IDIjGeCM0RADR
0F8pdiFWcJWJ3f+39tQ29+oj14SvYm5Y9PIlnZ7ASiOWggBWcTttUKPQRc2CT70c
1fY2uJdwI5QotLs9K6tuPkvFEK9rOsAzWQnai7S4w8w92+JeW32fWLMYd0oSjxki
HQZbSX+AAxlA2PA8MR6rrfqUdJ+QAl78t1adJCuM4+18QUh6VCQpy9qbmT0Pmes/
4SUwIa3lmvhc7L/fpq37ql/OZGqVF4E0myM2ND6E+e1U8O5Q53m1+Vgv1PMcdi9N
fQRdmlHymAH8wB6bL3qwjt5nCMpzWF4TFyovARZo0rtxmKSC05q6ZHSoegWcR9B6
4XGy6DFfZ1nS4fLJ6BKEt8S1qBZK8fRyyrdEMQeR/KwWHo2hv4mwDElJEQ0G1b/p
hrh2Rw7osMkJ0iPPP/gEnrx/dORitrkFoaW/9gHzS6W8EnEN9cEOvQcdyNIoacl6
k4yvFBy2iXghOuqMEWSIbLYS66cVNkBPWVjCJyMqWbS5IBjRUiCEkdYsAUl0ATvJ
VNcIwwyavO01rgQNw3E8Vme+jN4PnbtskvHEkW18yUpCurYqpknRj7PHe4EYUoga
dDZ+cC3cwCZTxyK7c6Dxup8OI9vPODg87MxTvT5KZClWbDfIuD1oYLX3p8+vkj8d
6FXHt+Fwiump3D2TTEAK3H03PLd2oQoe125y2KwSm2Hnt/AUtYX/b7jBvwPxRiN9
nAejSl9QC5qpMtDDQecAeMXfLyyhCr8PNXdlwH9RaMiwGcRyNjS0Zs2n500LBwMU
lLRNUqS2daYFD3mDgI/h4YW2hraHcp+i4rLCuTcY4J6u7oB6lQboGTJJmzCrogTM
YnWYvPeBszHz+EhF4+PTI9y/TBL3wEr/nrkkWgEq16hg9T1MmYv9pM5EC1wh+yux
zAA5hDhgWO76+J4+MIArk49jc0ztfFOAj+LluqcO+QNN7PT12tREeTk8nH26cyJe
j53XpohKRuYy9ys0imbO2WYQ0LM6IpcTkfLt8lu7E7BQkri35KvSNH6P+ZmNUDjH
rWfh8yFPa+uLIx34XugXRtvRcdARnl93FQU+8KulskkSWFySR7+RcGJu+bxGJl5c
zKJjDjApm5YIChWsXVkT5X545PSH2mEukjGueFYLmZRCIByjya3qF6vByOD5pfr4
lNnFto2G/IWH2CypHimxiJ0/56TL7NaDIkDrOudoP7A2zyrwa//oblDskr/YImCm
gvN71Ji6a+pB97CrKPqSSz024zC30KsVPC3CbLv/dNAXdyVEpMiiDN9NCMtTpqNt
DY2g5P8l97c+vxKZ9i9026EX5jzCY2udhtKg7uA1GrxW2QYEVTg/+ORGmDJAE/F+
ZWt40WqUFlLXXOzLoyJp7wIslfPPNqpwAzmGlLHEqqBUoVHfozX3Oq14nI23bYMw
tVsd/sDutRsgLHmyDLXUGq1z+frW6l2tbntDGd6opZdJ1rZthrvBBvANEfXDN++y
LXSr9woWZn4dQLIdSc3AjCuRYS9W5snihOs2Y6sbjLwaVry8YCgksHnqYX1/Dj1O
1HXWS+iUALy5Ol/gycgD+gPhQlqB/PsbfVUf7Ww0vWRmpLP0zd9il7cfq1DXCf23
mdjXJRZUBz3dfBUSJA4sXwcwqvz4/Z2T0c6N6TLNLLK9khbufvaKkvwqwC2yZHzk
u9A6P2Yg7nMPSkJo/MkTqwiPwo6gOlZYRpTWBOZHU5f9AgQjS759vtt72e6rJ0sV
zxykUIAzAmdOjlVp/3JrvzyPIExFnnFB3WfO3zwGmBLYR1UCegAhhwy22z3ubm5S
YZXaLzoDsYsdjFdc8UNnAqzKfuP2f0U3Gjb25x97Bs0A6oMIPHSWpzo+o7NWCWmP
lydjWfOcZAqkK9ILwH4tn7qEcgxdlwgs9uZURRea0pZdpC4WGISq+0o3NuAUfIYf
Ui6HEJXmLxAmCMZJV9SWEnP8XVP0eP+VcFXuzETnVX2fKj+1h1CeoZKssbY0KxbZ
0P2mW6toEXt20LICzq/C7C0ZSSig1zRvif9/XBsxzoMrzLb1SB3Xgglg4EL/4cWv
sFwIXZwgbO7skFXOsLJs9hM2o0WBCup+nLtucxDqrvR6QJ0X4c0qrwZ/+689t2iU
0WUVYmZ0w48OWakaC2VGge8CZBCONQm9bgJmhWyJYco/7sQmQj1Hilocdqqo2tVu
Yu/yvVVO0lPPQZCPyh7o7FfYMfuAJFpaBVFnf/+Q9ZuNCWzMt1Xr9naG4EJ48TJo
nTbBvaNQj6HNlCXj8dlK5PV0c69z6BOzW19rXFVtyH7eSlESQpEj75GA+F1P8Cqv
89DMxsjLDa1M+Ao0pYntbyvVeihx6Dx3sNpAbK5H5iaiDyeSiATU/UpxSu2tURNB
yv790YXUJ1W2l+vprAN/LLeem4oj9ToDUum0V75roOAq76e8p1CA5slJZIjzbAA8
URVAXXDGQjQ2tX/xCXA1kR1XhY8QSIJPynaUcDuQnZKbvg1Kwn18GYEeSFGHmQc4
RRlxv9/poXQpLBCFQBa83hXNSX+KIx1zpMgrsUSJtH+xHmRkLvkMlYcEB6WmU9He
nBvarGTaW0enIhVmzDQMICu8MANS7XHFa/JeCf6no0MTTzSCoVA1DKZ+NSRSGiNS
ALHpcfR3/L8hQxMUmGiQxcBw/7Qww7DTZm9ABOc11HxokD4KI7G+3bfTYGyHTDfO
LV1VSOYm01Wr94GUeCgxUpTOCttsEJQo0C4NUhFTu+NOlsiy3mvQY8YPYhfSuS1E
UdXF9xIE7pXY+ufPHs92E3BGqN5LAFtP0L8Oxh1NNm5J7BfP/QdPdqKHQFkhY9HE
OtJaXOJCkwFQbauqLRbdqjUjHc6K1CmOqIOl4pfnoSXUJi7XtKpTAPu0aS46I1rm
e1lx67ZcEn7/vcs4mqXMPACRe3O2ginc/zMKs/ZV1QaThnkcZafEIjwgoWFjvFwy
q5MiBfej3frdiJACJg/7aZY3uRylYC8pKg3KmuoRVGqpTY1x0Ai+d6UItQI6dArS
TpK+5oMVpXhL7Yh7TnEdKb3Xc0Usqu5KXSoVYICYEmOwHn72I2NxyBcGqzSxFqkN
+XbrjrgBnDv02NpVu9mnSRm8YEnMMTqyGPdhvXV5ngFTH9Kocl3Xx3DroGwEkIVn
UDVWV8HNCCitjwm4FAyPE5mcStAO8Tu39Rm67mxMUEV3LGzs4TNXNY0eA9MmlBjG
ohQM7n3eiWALhxDPA2BcqVp/4cuDWUm5hv9rRMD8NeH6Pz8H6EX0AKuBS7kbw3zc
GVj5V54w6nCAxzE2wx0HNTUiOgWG3FcIYy99cjD3UglXeOWLDmLz0EZ94gBs17y7
hqBtBBbzSnBKOp1+/VSZCWlYuHldPjoe/QdaaNrS9MQe8ypeEF9Y0pcQsqEuRhSe
6TnngsfeiMA/bUJDxXsvY5loVvLqoEw3ML6v+fq0PTEGnxoXFce5ncXWdpt3bw0B
GfcAUKrdy3e7gQia0F0Yrgx/lUlVWkhzFoJVC3M0/5PFuE9WdXoJTBvIkStg/6tI
D6tffnhSsFUo7ce3xyGNDU+FT5xPf8rye6sqExF/1kycHpOPYmHEBG77CPKpe0OF
j6x6DXLF5jpq5TZLwRPh1vbq/6dqGCoPVMwJ/HGcm7c4Z6FvdrRfC7rM+/e533B9
2gfSz6sJQvCJZ218nDMzsbOxZN+RnkRgnmkE3kt8e78bFDO3FY/SrX55Ag5ZAfBG
pOIDYRd0yL3KV3Yv88fL6tuYHIPUW+ozrPl/xP7ehPE8OQN4vz0KAk82viGUWaDT
aYl3iGlXxahvywKJOzwVofW1pwQbnlonpaQ/OLDL3shT7udlwiyGfAlEmuwP1viV
G1vNuECTYXfDkYUQeH3uxmrbz/zChPwvlgp54v/pVU5KoiIft39MtyUcX4XCM2yn
9/Z13Uyj5ByXavywntAuO9YLFAvoVHXtiTzQQhbVhXO17koBA02Q0NsIO1rQFxUh
ev2fE0rFMBEsfDBzkup3pD9RalF9yLNeKzj4lWJuUd7ApWuI8tbQ9vjqNldfMnsZ
ga+4SfA4Hs35OLVLFX3JDEzwr7OlBNOEdxvoR4pU0qqYtndTiMziPYXpaD3lNgtx
xd8ZaxD1cZsrILtTDP1hQNyv0UXNk/vWVNn7AWMIK8n8NnNToYKXCw+kXeCBv8iZ
ZrQgoOGyYEqRYjhIoOWOtyqzRyzLe2f1HAkSMHkYsjog765oWnlgLjNp9ofKLdwm
jPrS39gB84J9DQV1hcSzCCJFeFiJ7jl171F/Zvhjjahuakqy1Wp07mrhEUnkalfy
eKaQGdTyRitNH/oqTAa6DQD2doNJLPEFBbQPZ1xAOlX/uEE2xa7SJsLGXnn4q4Nu
Jvx0yQO4S6b6cTq7ZEElQgadHa7y3ZgOXZgrfRkf0CRm64s9zyDzqcT9geCapka7
NFxmGVdRiByGABS5m7829cK2Se6X1jzfHrhaWTuGlxyhgF12Qe+djkTPkVQbguaj
7sMQbnadtOhv6n07TydC1nKAgib28OsSNG/1PsLv0dnl8KXYrTlmZR04NkUb2mnR
aWtuHMBMLaB6Hgspxh2KXh4B+xOP5a7dm9S4WRUMSCm/9dDwlKDIOGZEgw1eJZC7
ufJxck+YO3Ob3A+8gcvd3v31aiXWpcGgX/L14Int1X2ekFIlBxYJwS7QQJ/MKoNw
OVdFvDhZK6ehrXGqb2ybyNNIztAC8vrjL47LFlpwXYD6B0c4tTzu4KK3ykRWJwdm
Wy1616JtmeY7VGU7oqEIsnGoBiZc0PZMwmPmXra6Hg48ZY9Vf3+xvN/WVK0ZaGRK
fAe7Nis2ZzsZvoHU66htfCH/TpaceKxc3FjURwMKUcTPv+zTlBBVjBpMqgcDj884
JjYr8VmGw+r58y5kxiEM00Wc7+LmWK+ijcDn1SQsxWRL/+9grD5ZswTB8AggkvWp
MRaGCnM80jWZ3BRjiK/p8rgZQARgSE8jNLzXn0d0pQU+5h2F3l94SC4IW6J7B93o
kHP3zi6x5yWC1nMb/jijXuAGT/lhdDHLxthomxJYKVDnOV2Zz/X4ZP/pew2PbbbU
HFj0/8swfzQRX7+ox+KXyEAabyNxcY54nHauepgsv1+6aayQD+HeUfkjhzP3EPFf
/FOrreCLCmkBtbjERSKcpxbDsJ27/8/gScTJZ4QsBV5Za9w+SP/6vXjwSiiv9glU
aO8Xv4cdV0NSUF0ZRnxAVZByPpDZJchr52RDkQ712ddP2hf7NRkPgNxlN2TfrIH7
B6q4a8JLWCPzxfKAUqghjBPdPZYH9M5DQ7MobHjEsiWo9VuqjO8Q/SWx9oHKAuOB
2tdgjnJF66Jbss/9RbTXo036Zsf9ffYpIP/l1zKhD5+GouLrumRnIrGK6D3u8Kt5
SryLc16Pka04Hy9DYY3N5QzIOyH/0qLXVV9HwL0Q0N7yq00Q8cDwWhqyk/M3jU8+
58LwEI7gLRIAfoGumJ5jXwk7s4gYAmcL/STrLDtlkCv8MPeZJEkZj+X/xjQqNiQ8
A+xgDcB9fFn4nD50UYiX0m3tSg7P0Jbgw1jEt/U7vzdrA08E4696/AoPEqv1ocvm
WiF6URPr0c6b9UyVzjm00DpHszj8XUL80bnqbkR0KFTppSf1nnZ62f6xg6OnRK0y
AFKXMdm2cpwRwef8EZVrlcTasgV6p8pBAdtu+KFMW3v2xCUczsGHvO3Vt1JUdthQ
RZyswQhE8+Nh1wa8Ka3ENfGCLAvwgq+nC5yXZz1N2DKTth7F/JISi9ArU8iWzRGR
NVqLSs1eeodzPBrYUBe9aqIgHK2AjdGbXYtLFnJI8j/qYzfbYCD1x7HLcYI6vqX3
cd47SCDxR1XAjsAGVzRnKrb4G8oJ3cDDHaRpH6V36Wm6z5Iy5fdj1KFV/sUGwE1T
QmhOkG11Hy+RNFaI5RHXPlsDlSjVLfsiza9/mv1Q1tGo2sk1Y30dq97g2C+DumqV
pJljqG5uB5exJK2VSzKiefMIPM2B3V8wGXi7wRVqhe0z0cLpuLUJfk+vIqgD3CHi
kzfCrsPQa+1VT159KKKkrLsJ+NbatZXxzq32MOoSSFhWa2v23pqdfhJ+a02IYztZ
cZh9HDYdnT7tyqR4eR9ATdCdv6hjgDN0uBrrjlI9CAwmLNmYMjdNsp6r0MfgeFUb
xJW7RvFTxbBoHcd1yA+aOPgMTMhczoRg9A0+j3L0zaatqWKQd+sTiyrwgESaPJ54
NIl5NErOpjQlI5nRmtuQmutaztlLCpL7UM24QIscKn6SiLNfkHv/lQwgywQ/TQzl
h56rUvCNv0OVqj42kPKo4gbTDC9odKwkqMAGHZ/xiOmpZbDoE0C0ksgIV0qZCrBn
3mBX/eL3sWG5rPRIUZqxXLkGBV3RCzqC8dq5him9e3t6Cx7Uq45stJsV1CSAEFeW
PuVnqcJYAqrg++03y+5sl4EI0Gu52l9r0WdDzp3Laaz/afIjLC3xTRvUt0ZONJWV
qsKqiXPQnCDbaNBGddN2gx7nmRTPp/zFx+iHMtGQtWDu5ZWIFAMWnKzXLym/p4hM
9D0LCBZ4HbHUerubNxIB62xbeUmnP6Ijfyr3sssZkj+ZP7Ts9V2uDRQuANkrzcsD
xTBa4Q5Be/mOwkP5GmhI+s8Hd4if+GzujNzyea3zPeef8yjty9ZoQA78rpqqhZXb
0UL96I7CwF04t1rUBOXeLvcFiGdXluiXG0WaYoiH+2R0xqAiOCMo99VfQtR13rKs
bCVxsh2+cM1+MUk5bk3Ofiiacd9TsoAv09Or8fqbmmFCi1CzUbpUpXnsGhSxiT5r
MOhtYxC3fcFGzhtWo/XpfyJWoWilbPnaBoRwyMftUXhMDhmT0/n51Jai2wXjuwMb
CBypfjmivNM9ycX/MlXCnzI1zdUIz8HJdbaAlTLHds2hI4szq68MyFWVHkc+V6D9
4dX2KuAxDLFipgoROCUbHyOVvtYO0lVBJIzRyr2Aq5seLVFzENdlT6DchK99QP1y
OKmpsYurZ2lcZMkcrC1rpPBlhVurpYeRdKM2GvzfiwPoWtqN0+rEgO0cnSa/3mkZ
+ZRvJ7mQmrWl7WZRET3MQ5YS5FsfaMU97TUfN0RuPKVYgxF+xjpqFx8Bnbpgf2qe
ETtMlrhAZQZ9szBm/rXOO5olvhL7sRHCfWf9ilNBLP1zfo6S+iNZ909kOuuV8RX6
7Fq9kCiBdrqpFO4agrng4bQO8R4d/5JRm1Jwm6ffS8R42y8pfqmLY4D72vtuNQ1u
ECQbccHvhQnXKkjWm+VyjNZErTHyZ8WN3oh++A2CAePWBBfvygza44xA9Jv9JvzR
TzgpMkTWdP+PU4TyWOCHnbugjmZFL5RBGX50r7oadu0qOGfEDEmp+QnDhKHv/nOX
48VFtWjaZoDpUaKkO0f0iRrNLesCzSqcboqFu6w/zpNFfYAYJ+1RWywadKCuMtTG
R8/3vO4xq44WUuxXBr7eT+CvHNH+jNuUB0wuAbENjO8CCu+7t/a1LjDfs3CkbrlK
q9mzILHwEOQ5DnJqFzPxXraAFfH1Ax2rT82cL8NbAa191Lkf9buFgTai0lWTXnNe
3UA/2eeWRFZhqAMmu4eHO/psXEN7Mm07ycxeBv5rF/Hiwvru1I5hkNT4IW1teDmH
2gxYykOOSTeaBU6xoAxLv8fLoBlZPhmC3KB42PFNOKbiSX3032C0RNx54MX7Un6i
gNcyD5ZiE6eTTuc4tI5jkbKAG3oTqpr5DNsHF9TYTH27SRnjkmAVp9602L1pYCeL
+Ku/hzCcrwAZSf2wg7ahR8w31iVAyPT4+RLfosDTub7rd5StNQolG7geBWRyVWyp
qdAO+Qyi27YQFWZC7O61ThO9QS3VgGPCNYYZT0mLR/rVjuDgerctaM9rIkvALKwQ
foFP0T/YEnxMtE8FPvdRD0fwqOelZIwo3N90XX5j/SSiHJHlM79Tk1fbwKa46IG9
6M2vWIbbkmeV1fdP0/KeR9ZE/0ZGPDXldMqeRL2az9xXTmhMPbSwP54pjTIqF+yG
YTMFW7Q1scOnwmWtZLmYjB96I0BsOfnXAdv4LQIeLjHvgGOe4MjP+I18ArgAyf2x
aNsC4AfWqk9yoUdfhDNFzrNxfcdubSslofFh6y/5VnvF2BMw+JwhVoFYQiz5d3ht
91UEGSYfe8oHDnSJhbNxg4KlAXHGZvXxqD1slL53aY50sA+nwnALThrJONh0auWc
GilyUE33yUbLRTxbeR8zEqqXqwgOvK2WPjlOAo3yGvfqgSoHexSd78ysCgSJ8pHw
j4zom7ycSg2rCKJde3JUp/WUFVL8wMklAcE1ZjSp90n8w7jU4kpw8ukmybmdd1xR
Vhm0MeebnEv5D6j875ahg/C/IU4VRm4yyapdNUWIuKJkHS8foTYMMKp3c3CixS9V
OoC3iTkaWaD1Jd7QPujfpLyFKE0TAhBVRLYySpA0iydGNBQwvrNL8gZQCzGH6OlX
tRYGRqwaE/JgLOiMAgjSIk8uBjnI+felCVG42xNJ/P892M3lv/hE0fbv/n1wZSRh
JFpeLPe2Es5R4HCgCdNV5JeILbzK8nq0Ou8YFYoTDR6Jley7j79iT/OBtDxaT92y
1yk26vrIrdjOIR6ipQX3hGk2lRut1Zipva7w74Wm1GYnyGY9x7LeUabJkXQ+cuWh
DLk5xl5ab3tv3Ch8V3T7vgwZVEE9PZexkteBQPQl8wjvdNSn3rnuD2YZ5U6VUamv
e3aTg6PsfPG7MAqHmP2Q5Rg5AfjWKp6ag55RTLphlZYnsB2GAzdyvYLHx7eM/Lk5
cjz7nkQvBRzthjYzCN48K2G3oCzoKvLa8at+3Nd1tpmddmNEtrKfGwH++f5rQPRb
4en0k2faIhV2aYemYWuu67/Y5j1WXLZh4EHMDYXLc4W6jNLG/hOnXlOGLWmlIzVg
mBULsewmF9OtdDup9XYPze94F0iVPWJgXc8FhqzsdL4m5ZMtMss7spafaQBGNpnN
oIXN1spkqXOySe8kotS1S+5OTk6aWlC8ZJ/YoFM3Dtil769dAooUwCjENhg+3/SR
/Ezqsj1PxvyPOn+hcoR9OuABw5M4h9IHHTKiykUruU1OHjOUOkgkLicODxfH24zm
a/d/IWxhISLuHngczsKhyiBacTtChYWkP4bsXvp1G5GVlIRrXrNn0BG9aMTj6JIC
MpRy2eJtf5qUB211TwdvnBdFaThdsepqtWchWGyc9IO3AgED2xuIdYM9HOWV+8pr
005GaejDFRRvlfnuDQ9qcyj+Y7WrICsHk3BGfa8JrllfU1CIjZ7XRruGMZHnkp4k
WK8H2V1t56wU4lofx1OlRfmva5VdUmBPuMe69nXtceMZIcNbM79KtSHHf2WF9pDK
+RDJlZU/6/iQpm/M81+uQ9OiSLm+AMB5KIRiNONMKM4o888G91TnvjVzF/QJi1Uw
9zD50cnW2rK8ymRTeUKPefW0ocKE/Yzd0GE+0Q897VazM1+le5uWT5NTuhicaKxS
xsHX8eAJPZY5mwG5Z3g5l3mPc1w2h27TQRWHU9KhUflVBADk4U9vsYUWLSLV/Ksf
u8Wa/QG3elaQX+t+YNzGo3kKgVPzb7Co/YCtI6pGJ/N0Y5CzPlDglNSP8WYtQQgX
D3Dl8S8v/csyun0HBZ6TsY3uU69Wrkf3bTRST9HuCwwuI2XIXTpdqeGa4NupCO6N
XWNzcRy3j5RvhN6CKpqmW71znMjWl0m+JsBjb1uZ7e0+eD5FzexGp6k6Lqz3Av2v
zOilAnRDBXIpe1JPRz6FAhjd/3d+LuWulKuCbXGU/BfRv8HtQXBnA31aTgq57ijs
CkSFkGoHu3MsgYOFYlE3gFtpEAcKvnd6VQT+sha4ekdtIcZSdxQJrXD7ELUgR8/K
fYxiNdFXRhnGjiWjPhjmENgLso74Xz3CFRCwLkCUUYNIAdrrXJ5O3QCPlX9oaaPA
TkQWs+VV2WCWwu+raKgbZBNOAai8nQlQvj5GN9lJQLCXFO2NaXWc/QZVG4scD9Or
at0yqie92v9XIK5Wfwj6uFdABLAOZh0dFQ4AnDwLILXbzZqQ/+iNhRVWXGT03OZZ
QIX2FrU/SHnnFTy0oX+ES4bqngtl60DvExn72yzCe4QBU8Ps7voc1gVEsAKJY+7e
xzIM+ocKnTTnJs8cDKdHuRTEGkNWhh2Oz9tpg5fh+wxZXiuG4qg2Pp7SuvJOLBHL
bzGFKwr+P1N9qIQPXwfqgwI/Ge5zIo5Wvc0t8sfm9b4LQMsdvLWDR1KZtVjXg8BY
AesL9IOnBJ5sqhvZKYoRsOmyLJdGCEk7kN1fEx5luTouhtt0MhUKdohG+c9ruI0L
hYDvvzUHfCm/CqZR0/7mHY+yjQ1S3+vgUJHH7ELvaFQv6hZ5NZJ9CmXpLu0y+5ei
LDWkTpqP5X5onMBCkFpzmgBytGID3pyEuSHptYkla4+uVdmXPnYuDSqw1quWmv9F
yzJwN0mKdjxfCK8FkUGULJh5KheFTalq4KNs/X6essJsqNsdTSlfX98qlADNwZpl
vcx+hZJDzmVDsylSCpbnXMbEEttdl9yeV+/n5s4hM9WnTnDT/NSnmBdYNrbkOQa8
2dI34jFkg+8lFZ2mPYtHoCEmT+LhgfmbEfnK58rrGQWkG0vMYM0iQJeog8k5Cj0H
LNwKw6yVFOeg6Udggrtwv9qJxAQwROgzj/U0WwLcuSEXm4ij6+HbcYeQVUY3I03x
S6w2x83H+Wze7zppTos6sIT+Cq7BIkmK3faR4O9geKrFC81sx/eP96k440C343KH
rqJx72wRGwPCnDt6SoleeB+j96rHKDz0Dp0VLhOJ3Yj/mX4veEWB/BoUBewOds+O
mFjsS8himSJVahceREZ/KcyOmjw7vCCsBz4vPOtCLATFS3XKo3Cfop9CpQu4yX7e
a5I0dmMIsSCQK1QAGLBkOoKTUEoblXRxWFSq+6zmrbiBIn0bxPWz+VSrRPwAaQSy
DK9fAecrpUvqYrzuzUDhw8lS4EAebVseptkEFO/B0qjo282KptZix4eOH2a7EDlh
EXThPaSaBQOGGCwPC0nivsKX4zfWkf+3tB5+s+fPTGwD/Z0JnXaXS/EvkmMgcN8Y
iIDB0VSYYVRSR0z0PkVeulMkkPZgJXq0jqn1v+h1WBp5e2Mck629gzNoxBiXJYx1
BGiwicqFSYFrLiKuo22Nmk7b8DUpJnw7ppGjzRGk6sX+ZJ/OGPO9Fi83EtRsNANY
bQ4TWuYiAFO7TtxbFrx57Plb5lq8WeriMmfYTEEnwVwDqam+aYJLOrxX5KlQqpUU
dHebxOJ7H2fJWAkU/+s/fyfcUamJgoAmg1Rn1WRMxmrStso07CmbgxG8x8hcL2DX
hnflMIfFPPT8oE628vQcqNMwLscwYMizty7xsvndtMpXuIQ65KJatVX0RCP3rNGS
/i9elH97Qc2+D7BREHqaJryf800+0svKn+vXF4z/W1E5VXvoI37xVuohQUYfwBGk
q5AJxpSby3bP+Y6FY3ngP1okttha8CvUMT0UAFO+23v1JXhqsibO2/+eePsOENSi
j2LIjUKYW3ap+Dd1bupAk+TUB8764oQqA/pHblUWK2+7oQAskixxWorbw/Rmov3r
df5horijWK111MKbkJ53SH34LJg8OB0H+9Q8fNXhMJy+qXF9a802qIzMHAhpFCTu
rWtQSTt0rSh5rDR/Is8sJhf4T9t7gLcxSqMzGp/39jBIAYv8StDBAFaJ5YlIPvFd
zwaCKy0BzmqmgHk49I3IlMs99I+nJnIfRQAYwtN2GpPzGUTQkIRxEn8iahojBnND
NPYHzULr8bDpWzvXmK5DHSkmbadEa/avzQa4yW3LYQrY3GRhoA50UYGfyTpj5/0E
u/tD9xoI+/TAlAIrC6YV3vkzp5nGkHonmnT3h4GLPg1y8rKLoVNswTDh2ZCtTfxZ
6blD3edoryU9NAFJgpB3NB3aWZHbKj/YbKHeWgqPF/AKR9oQ0FM3bX10BHeKe1mW
u47WXCjRm8Yk/s8SNRF9Fn6BLHJJHCjaaOzYnpVUjldja716CLtix8DWtqBa7hlE
8jeHHlDWplsbOiVvfVwk3tVHApN1xuwuIhXlVWBh9uhdsgkbrVOjcQK2iF8vAOZ6
1IFD8dIHygeck2gTEIMiKiJ+WndruFmF5Y1qkZfgbeqn+5jX51G76SWrK6aZBqaU
QahdB+nlhSclZ791fMZatk1fQHR9ENjcpUrl0i4vfZ5DJRZj6dLN8p2eG7wcFsD2
sD39RTHGxvkKs7VobE58vOO2PNRri9ybh1PCAyuxR7qRRpynsVU8PaYNNbBu6Ybr
nttU3DR5Io3sYn7HbO+7CKxLU+PgojYSR1lrVpxJyDRw+MncfECglj/cLwlgMrsu
ArSc2Rhf+mMEPWTgGsh3AOfnGNTGujIZuRcUS+QEzXXofOeof1TbAbgDSwEV50zj
xU1Bg0/yOmXQiDx+cA+DZqhKxA9nccXhERSNdYQ7zTL5i1oDYzILfWx2URfJeJ2O
ofyFx8ucyBGvEwYsRnst5uEZP9OLVgVhqhAC+hFMP9miaOKUE4nEh76qIuXwdE7f
ZH0OAI6Dv1uPvwg3sjLxVHIRR/xaiABKYvuE8ee9kmsjz1/wvoV19V1sNj7hwdkO
GOBpT+yutIyCXXSsCQYVuwgH+oRVKZqR5nVmlLMtulp7vAKcQTjX6yQ+8WKDWSlu
E3mC36jdj9uanjkUGj/hADZ8l0DqDe/JM5fpaLX8hLEeLKMQRitFjV0/8FQIxF1H
Gceysaol+J+fBYo90+GQEDPbvdrx8UBlHYSLWWK9RQQL3JrnGUh7Y8upytSNxYxC
sCLo2/p0X5skaW1RRyRtlwkIeRRSaUZUAoMFTfVvRKQ8KZAucHnpX3Jj7vkM2gLV
aJnbvi808X9bHnLY24K5cUGcb8Uxd5kqnMS91LpmyTagFE/T14Sn8eJFRBl3yWuh
vYzHxaW6lmJuYpPxIBOOI2eiZyOhgzrIcJqJEWjYc7/l6PIVPu0lo7UirtEE3fq2
XDUepKJE8GEyw5rV83suuvvzBuD5ew2/qTf2OAAbKdg4U8kHgZYPgm3+qzMMSba4
s6C9rje1Qz0WQNC++C4/zxvTfkvZ8z4XGuu/gIMu0x8dqXUVnpU13mXWPQOXC13j
2+ZxYHgyvSfh4vhgaOKfOY7n+OnIiEilUFvq4yzeq3tz5bw4wZBdVkC8jFqcUMLh
wHTNcCNnJL6qFUd7hkmIzhoehPSqktTnYczSlDVKk8wsw1/oj2jG2V0vRAOuKx+u
efCO7l5fTlv0Bx0KA6KEmG5wUhhA3TmAOwejGoYn9NJ+4Rh52qIOcyqlUoRhJmpx
QXAYzwC7jeaiG48yIV+fLOL/vUNFjdIneLF4J8SyLv2BVlYbOoBppvr/fwQEEILS
f8tJzBOxGs7LvUvfOoICG4gVhTmyAnM+QlHmop5OpxtjDMLpvejOXZ0f1wJGcFeR
j/Q9Nk7T6tWsX08OVZQy8WHD2/4TFdyJkv0wvzGg8gBszkEVcu6AQUqojfHW9dMF
o+R74aR0OZ1pUo3YA22/gGUHgfwp+A7nrU+JV/ZQMDcHvdD/aoY6E1JNAieIhztY
x2N98McqN7ZfCaULviAau1jue9iNlyE9yCT43NGVaSrXENC3y8t5gsPUmIhrtaEd
vSHlw7ZG3ODMzDV8dNtA+9E/7s3NPtEZDPZd47QLSSWZJpjPaF/zssCybh6Wk3x9
3UMo9G1og2S7q+67LTACOVffKaM5dINvt7oPTH/Ydp9iokpYLzkGJRjQZVluaBdv
pGp1jUvknbYC087OVBbNaUTgKefIfqRREDW+P54E0KE6BIDavrt4I9QnGhhmM0h1
HfoL9M1mCSDWsRi1ZzS0SYr/V06MVTJ0hUSeSIpZobcf3hj+TtyuPRQbb2KSgvgT
wKFt2kYIyOZrpeAZ/aVUQmkYmx2MX5k9nzl5cM6SaTASgWjmnwqeYZdfxHPUpJcd
i0Lw479y79XfPZOBeoYO838fecuWmZXfTAq6skcDLs58AG+7qohNI1qt8VI4/ewy
j/7/ilkYKihE1j/eratKrokFl4hz8c2Dq02jMy3io04yWglsSZYL0E9PqaO8aana
fwagKw4tQpIzK3XCq8JkR3PtVPzlXV0FtEblai166EYhBZGfcSMp9ZQA4Je2KmUY
8eoQqnJlIJ3LTwpIn4xMikvqQBqQJJpwgHPE+hN+re++aKeBnC0GlFYfg3w8cESA
9zXgMcJEffIOPe2QviyOhnhucC4CdPY7rmUENP4UrapIaE+1UhGdPtnedVATxU7t
Mxd3rHJ3tGH4I5TeaJ4Mb0SVNoAsLbpAPNpN2nfUX1GVRrbi+vW4nZzdWeE2o8MD
/wvxejSQeR6qq6DhtXvtnwBDZPOOtC/iPWRBUNr0zpvj+0WXCz6gjn0D5UpDQpP6
pwe2XhKj2U6un+68NtPDLt8zBIf6eqrBhwFj8svUJgDYNEYy8kvRttqOhy3W2/u0
HKvWMr6+ySJo0y9ZKXNc2Vf1aEX1QsNCBPFHkkLE/tf3AOM9A5JpLiq5uQQFQxsI
vrSX8qDKHjOlWrEmkOaLZIMHhXVK6Pm43GeDYrkLGgm+fG0c9wGBdc0iYVd8Ro0T
f95uDTW7jG3jqw5OWm3WZNs4fNlqX2byRtpByg2NcQlpmUaEtf4LVSjJCb+IFqty
jiY0dIFLLYqcb4UW04M2S9G6NjLC6MXR3ufFEKa6lLjD4/22uySJ55mJU1GwX7ji
Mdh7EEKijGIj8caQOHYXOUWodhPs370xiLzvuQaXpeTnwN4jHa+RptymLsc06sg4
biKaWqUsJ5nY0r/srjEeHyTKf7cH4vH3b4ynh61q9swnK/fhll0+ITMg1LZfIy7p
chP2iQCQpSDSHVD/ucJ3HKxEhfRsPBOlxq7e8MNUBipmICg/G8Gm3/0R1zk6s5KJ
RLVgG1ZHGgfaYh60xGxCvQ2Sw18GBjD+MwT+h8+lheJcCNkYx+GWIGysi4/PNoh5
kPeaPcds3j2PW9j/TBuh6IAMGrZEdWt8PP6BIAil4EKWrEkb6XwQAAjdEc4ilvyZ
5b+Fb8DnnBRtUsvVxbKLdoKozjMCqNxlkbIxNaNDERd4isl29duv8tGdG7ZVP8N5
U4bYd9FqlRONWS4xqUvg0K5093zLKztvAtiqKC//wo9CAi6G6DAiWv8PCizyvWQg
+0+L2vRfiQAETSWCpIWZGWsRqpe2dCe915XSoE6avYxQbw9/bT0K7h+qlAUYlLCy
2phAIJhVs3SEnhmpZSIK+gkSGitvi3BMIR6T07l9Mi+lSxAjZwJbX25NA1f0vk8W
OAfhc31Ba8CKTQYCRgYI5pZ+H+TF8lTcBTx8k08l1CLKLWOiY2R3/EglLKQdNL5p
tS2gfrNbX+SThjy4+cVPUogPZ0HjNRguEOEBSoDIi2SPM1CsMpQVwFey4CXhy0L7
4WBbgwlmpIl8Y4lhcUzRgjEv99DQkRa7C7yXgrGidPkhb+40CBmynKcZlT0WdWq5
I7IwrUu/sWPrCKcrvvfLRTwuKy1fKy180bWsC4fsUN7aTHGzRwgS82edXcnBOUTn
In9oWMraR0mX11reTUKMNOwfH3rhRxACfsIMWCe264uHIXn7vX4p8y4tyxl/NT8s
wKu23o+QNHViqC7Vqjf4NugO95EP+l8iBKdZpSDsRW8Mctf2iaPoQlFgwEOUCpYD
IlK7qJxn5TIW7DsL8FCEBur+Rzn0+BFcqsXdoJY6Py+8KNIT3k3i34vVBKkrhrg/
tK5E+Y+iU8GUQtYH170G7DrbuozO1YFs0AgfF2FD2cc10Ne9t1R2bgsoYeux2bU0
VQz3ueC6B4pm2kRmKnFGsYmmSzEDPmTl0tR5PxKFTeUF0G8EaM7I6v6+CQhEreua
N+7cdh9snuU1CJk0WwTmE5TnuAYL0pf2420dwrJ7UMaLCVol0oaiyojGeZFIiLkU
twnF4d4vsIpiBkzKklQeT3cQVd6hKC8WHt2LKBMGoJ0DXI3B35U7M70wKdtlmANr
XajIs0Ul2HmuSxhwMMCyUQ3P0VS4U7a4HVlBSpyG+/3/1E0Zmk4Fd85VopVKmSE6
qHH2XlTRSOToNt4mg+e0DCsiogVHMFHBWJgBMJxRfkO4WUP9teLgTKe72yFtNfOt
2R/VEleObUk/vuAJxYNhl6BSTy68UsIhxORVqNztffTZdqEkbNQTFkFsayHIJuWF
T+C183TnE/WFyXbxiYQCs4Vw5NQd0bR2LM+sDgFgkX8PzBIpfgkxR2uO7DnLJxK5
56NoDr6B9dgUWZwh0Ce6AanOnPzEt2RWA3lSNrlwes0Bftv1RNlo7qtlMKEvP9Ia
TOr+O9HuV6WTywdMJuGUDf0SRto9L+WQhEXBG5JFoUFHo37Fmwf1BcRJxaQGtgwb
k05WrEPiWHzfRbAN63WnOf0pAT0Ko7SUCJw1DNCImOlELLuDK+VeMyDaEeRlJAuA
CKq0An+jE1ex3ix7w5rUglovsIs8W+0X6PUiKmzfQ2lrq+TZwtomT9EuDftphctx
DvMihJz0Xe6lFz7+68CGc3dW2bcplBvIw/z8xSErgTwaeIJHRQMnEYzqw0S1Gg5t
tY3mmYjfFkIpKfdATsKFv1QoIubkm7Rv0tyo4YuTiyvl81JmKBVoaGj68a40Mda1
MjyuEVW9HwLFm8q5LiBMLZ6mGUzLm9wy7x5Mz01F+rsNgqlxv/fIQXAt3SEigOLP
mNDxu7C2LW3xZqKuMrUC4U6Gxy/tf2Vsk2ZN+x0wHKwd0R5wW67TAkbUEZapS/H5
77G8W6IlL9SmECZs26uqLNMYo2xSpIGz7OC/FFOxq0s1hZHat2k0y21QQpbQfo2z
dT6o43mAyvTf3N9U10Xs7hyiAopo5myGZsQ0CrhSKyrWI7ia3JOOVgZ5pYAEF56T
tI8eSFUSKWmEr7riv3JvTJLTwYlWe8gsLdjYhrCpwDAd70lwqR1gyPiWNejY2wYQ
7Ynv4lK5QQFmrZR/3jf4n+CCklaINZ+CdnEPwg4LNOwpXpyiKwfM6mq3XibMP//2
qJLc0LpecmXBgCIaV7o62C7Wky5y7Y+OTbBv7pIh/nxj3J2l/PDyzzDN8/ibXphy
RqjQK3c1ItlUEF95asJUnRUyej+ji1DUwoq00Q9T4qTOO4OTKK8L+QuattPr/zt/
43RUbMzpu8Pt/EWnAWVP7Nd0MOfjNYuNePXZpgxkGeohXDxPGxur54Lnzxq5JzF5
DQALMnaKn2L0wbNrwP2doMhTddyejgwl57uF9Zsg1OhNW6pGEJ3srTZ4NzmQa7I1
D72RakLFzEuU6f8ZZNzoy576QtKHNd4ZXUxemoQPYEpM6iCEn9XPMnMnnexOzmPZ
eoYKISi0YWCekqtoj+ElH22qVjMOIYIUFNeAPYnNu46mU1mr9qAUtAGoxRbQR/IM
0ngBcTSv2iwWTxxbUARxkmA2W1PagkwFWRVu7ZAb+Y0IdcE0zjI2ic5MgatrMNei
kI/V7NlQvccJiW3fiKXJLNkSqgeplYUU97hCp5+gg0brXaVNNLak783VDv10Q4dy
Zq043rMdgmq5NwN/4xG6sqq2I6bJ3bKIDhBDSaDgo97UX2jsWfG46czItd88Z2Ra
/Zs5M6SnddwZF2bBJumFa+IeUa4wJdUrHBhXLMNtfWr2BwHd7b7/khgs/ilYTKjY
cwbrYdE1V4ZJyP+25iwirCeV5rsQ0arOLEiDhAuwV+RB4V5aYnQG8fheakbDNO7b
04OLUDWKRzJGa7nMWIzcCuPLa1tJhzoI/81tspQBAx6B5gYxVRj9vxCH8QxxYZ0j
qpnPN5wmaeW+dXoKAaNs1oW4m5pcyzkGvdT5FmocjxFDLvUIXHvB+gZkQBOjjwPq
jz7pUfqavx878FImy3mHpylYDn+0FusZL7+1oKJDMiGd9fDKUF9u/zV0RLvIQuRR
TxKZzrN9Cc5J43NC4MCj9g7Y+z3tkqESn+1r/BgOQSgALxWRh252nbPsK4YClHQ2
A6Fd2XIAxYbaBXKosqfHDtZZyCQXt4I6Fz0yZsMZecfkZs1O+YlP6bx9F4/EqmBb
EyIIA8VAEM9UUP3nifJSzTrv3kUnSOAI0ZU3ymk4m/k8xb5bE+9Euyo8uVp2AwVU
gcn+fY22y/UMqLn5wSwbLsrPhNpLH+aLfsEmZ5L5Z8HieH+L9Rx4OgseiC+TiG0Q
NVuYgQuPbq4USTx9QMx8wipEoWXcYFg+R8Puj9iEyD869bBFZFS8eLGjbccR3IlH
Bin/kCc7GvQzaE+BUaHGKlwOpVv5OPsJUwwhg7ChUDnye8FiWyP3kWePARLbaRCS
GZZdlHI5hRYcwD8ZbjpT1JEBQHKAZlxPvWsul3GNB/K5QaQPHQNpN/Il2Jh17s9e
n4ySrAwUB1S4o4avaTRhrFfbGmK5ewDRzkdXwf3cPuWQny39m9Vj0uVgsn197Mwi
0Ge+hXpsFpMrBtlXomV8f6/u2qXyMXo2xZYvimhZpb/SOhIMUEnlXgfKHAxwGeL/
2ta6fbvA4EC76eLA/Rc5mjrb8LkxjUmzgvDrzPs4gsebW0EXFxnjTcD38Dqp+plR
yGQOFt381RSqMn6GoS9IZ+G0zrPcKRF1/wDxXQ8I2NSW55lR9sGB356PwQIn2nWd
YX4Tk/kOQRmTUlhmFgel97p1YSMgYxv5jeJXGfWXuPBAOkI2E5JvvkVSg10dr19H
p92/oTiaJkl73xog/zndb/dzczN/bFtwR0a+IIw/RsQItj8GlTW8X0N6D7tEC+c0
j/TMW+EJ8MBOprNRG+TccyCwF1nKAmjTx6DdLcnaQut4srfyWB8MbJ/WctVtXWob
djsMHlQBqfxebUCWcSODPIlKnI/Nw8a2EA/ljvVe4YcoItYCs8UdP3USdwM9q6hg
ITEVZJkw0xtxF0GqWoHFHn3HwbFo2X+TbG1Pph46YlXV0j7N7/SN/QA5z3wCSDY4
gcZv/qRut59us1RghyXex6CZ1ZVDha4adSbyAm8FMtOYZ8+ZwnwpmyAbvmgrgGBe
3VHP3jfiu2E9/Zn1EOpWIQmZNXCpJmMRzT6Yj+DdUItCzjvHj0ora6crU2MsPZQa
x23YMGK98JyEocDSAt4lxakBt+5gRdxnslTGixciV5eYy+D3ri2e6xQW22dSW6AE
N6v1RQWhnp6YhMFqj9HAQZzU8X/MRis47NRDmwIja7kUVPs0qmOAFF/r8cN8st2d
pXB+32V5xVOwNAciCTsFOLOndPEEeaKEYr+DxtwjTkkqnzesU233pQFkIFSu7oIr
cj1xpcwYlFgu/aNlyAvUO0SaS0ZLBycNvAqEkh2FNiQIfp+vOYzMTi6niulyjZMz
bvM3ctX0sFTj2HLszIGi2qJyDcQix1hhnpcbBX1mCTanRZtcLRejjior3Zm9Jko7
nacA6QFNMgX+AXM57kZtn1EB+BRbh6Mj7FYuFqvL++DvlWyIwdR7pJuY5Fl3AyV3
jRoNIpkqO2XD3N4E253GwBQrcKllrdhxrJxa2PO1kdC5XUirwg/6ahjzSD0xnMm2
ub0qKGEPsi+ohNTgEMYq61vzsqJNKy37MFu+7yqicruqU5bmyvXMdD/f8m5F0tvt
5LA+AFwHs4qzxL1w79U4nsjNrjEXMVE5bQkrnqlPfZTcxXjvwEZcNFchtsFoalcm
8XT0d7dwi6gbk+Lr2AIP3kYqoh5sdh2rYzWIxrMp8un7RMnkS1/Q+96p77kw9EKK
jRLd0LKmUt5s1ttaYj0UCLgiTEzxZ/twLQwgXxQVaYUc1Hk+RBwq+38gv6CBpzVB
Xidg+9OqHvuRqjkk9F/dgHJDV2hI+6+8FkFcUUTgW2N7IgnuC3y7MLoaoEoKkx4u
ocwfisojj2JkPomsylbPIWthhY9pWB+O9bUCkPuvR/98mwdmbMPYQcalg89Ni6Gw
Ff2wk2l5GC1XUodqj04McCJA8xLxDxgh3MnOZfuZOh62kj7NEZAY8UHgb5mi+ckE
E8HstrJURGoBtgyiUyU7biAZLjTa4rBm/7iCA1C102vQfUHdzAyj3WqMM5kSToYd
Wvl6aEtl5DPSkR/WrZAfYVyOzEBhrEIFgx+A80V6ZMDegcpVReHZt2mLjfs+VLNZ
jkXMflXL2E4UuaD2G+DQSZMoTuYEfjbvbcwLrbCbggfFwjwgku5yZL7yUNKz/Yq9
tKE7wXtPz1Xzwx6p8fIEuId2AEwd4x3CCwaLeqSFmGFIT8e3me0kJ7GIwb2FAKQV
BQmV5QM/iRx528i4vpELfOl/o2ZSe7zrFQEiHN2K7hFShaylYost5B0IZby5lmWm
gVekRJp214FdbgQpvxhE1M9NArcqv5QUUoD0cAOCzPDZY6AS4LkZ4TfOr8AJtbmE
hgh9Yjlt/lyw7DD+KB75x2r2OsNYNCAtyohDHyyU1ymluvYTjdOTzsnhyKv1yJ0T
OXW1zrKwLu6S03konAyYPSNp95hzfZytw5mKUBONr3Q8f2/qixqYAK4zsz2enayj
SMM6MuTHwzgyKOheZd6nc9BZemdFFa67mzD1yz2zCL5uWPMv0WLyzzQbAeXCqQQU
Ify3rAjBeTY2m9w2nNrZrzZee8zRh181umrqfSJ7UwGgOvxDAaeaQ4LDGJZ+uMGJ
OyXEeC4C2vK6pM2fgPFPQhJIpUzsqiZ3M+Z2+BIFGf8XKy89SdZlwNlimfZ+/O9Y
NkW63QXiUH0C466eJ1ZsVxUykZRbEhTjluP9Pwa8+rz/X+ml9ZQJrhYXPTD95l2U
B4Jy9XSZT/JsTONpSTIvOFcAz/edmpUSp6oTwykK7nx0gVGl6nqEwX8V1QAVIFl8
UZhN4HFcdDjldA2qe7kLS0UCJ0ZhfqaAsfiDdDYsNQf/oXa7TCeg1rZNUxp0dMby
YHWRrGxKRFeDSmN5bEaFmyfCKcziBhizLLBhbFGDOlFE4FEA6L1MAx2U8RHQVNUz
W/4KAZLtMQggp4XixTLAVjxIjeW/Y+SwD3xFHUsIdoPD/nW/3sJBh1MtShnRM5I8
HcFXLzt5m3h36K/RnW18nrr96QJWhfCJgWdm5k/r85414OVWGYTn13UYnYD4/fbs
y2zZBiXlGDDj7LOtiKtvgAkSESJQk8bZvl7+Z02yzKxuzEAS5+QCqRD5bBaFNl8y
0AByQBRRJvlo+pjKH+gXLRZ8UqdbLSRnCpKo72tjW79+OQ8wPKNh6YkM15zHFMAW
SLBMitQ53HdTTw8ln0dU/A/Z5OHuuLMXCKAD+XdBTGquqICirLd2LHAXfQ5y4N6Z
qpcBkSeK1bBPUim5jpi9i+Z5Of131c/9cq0rISHNtSvuGZrugljlRdotL4N+7U9U
6WThz4DU6xkUlqgL1YUHgSvANXAhGsStu4XMipYCtvzuDF8VEpU6ZW7SzmYm96vb
gjGE/GYI/kWH3ih85plMaujywyRN0B7//q6DUJ9dKIvQpGDIDoYqtHOZHGMhJ0iJ
+WC2lXB88c07nA5vIT6USlqBB6jq0wmId+gFFnbHwzRUg8z2vf6YcCq2QhPRB4YB
bRfFjjtotlOlPnu8seo/ZK/GZvr2E0b+6nwKRJ7EY/SyV2wP//JSFzfDHhYvYPs7
i2WysTydknXHXIdvXK3u2yiAgNoPSyExmtanBcpaybay615E6lBHyUtkK+4wgP03
fABVEsktuXx1dcx/guhGG3QemfEISuDNpAD98CGSU0v+fHTQc0P7rXWsc+TyayUW
HmbdRr5G3dRy8lpnNKWIEORTilGXEz5hil8KOn5EjMmPeEVVnd24BB6MGkT/jvuY
ClTlJDLhP//q2kBM+PtPFvOBlNgPyOryQacT0CHBFlTb+8xkW6mIKC6alq5i0yYJ
ez5LmbVTq4grEBbmv2MUtK8URv1WaAQaJAbkPbQK+V73YEsok4MAIhT4HpcHnYd6
S1bkTgIIh9RTGBdou/lyGxUZPbXs18xO2gJ9cXSo8LcbGEV+HKpp4N1Ck5iMNSi6
gG5b3DfBH02/ZsOeVjNwXCPb39DzooQy6LuW8pc9fqpYQ2/Qki7BRU3Ar3m7VFs/
ySKI4Ba1408HZsLXaVu/Op4ZCTJZItwqNZa/t8qNoxcUKyir/igNlcpjOm5f1VJT
WrVeVgpJnqJOnlFRJ794OWzTC6yU6lK4SRcsTuVkVRSftItiJgYKpJWc8MRKMbav
Nik1T4wC8t/P/v1wEbnwo7eG5LcOGPzynb6SJmUi+dVQAo45qCgAxcxRfnNKZjZX
zUqHxQ2lLKprZutGbWD6N325jXlw8a7LopyyH5vMPDa1ozXnlsJhQQYMu0DM2V/y
110RCuZebdwvgSfoNAEO5bcWU7tf3ibFtYjhuvibzIPWUxyuHNSKgw+9iq/ouPxJ
ufr9RxBYXBFYcN6SztqYxFS3/0tUnlPSuE+caS87M8eXObNLXnpk270YwfMimEDj
GQJgaDcYLH5NcPvUvvfTO8p5+MLijFE/HdWCD1MLhLLmitVHON6OjDyl47gUyPNB
nyxCrKeOrZGMcIbpKWTd4Zvn34hwDxLmcp29T+kvJVzrPy8YEU0/7kdcVcO9WC/1
ctgidvg+MZ6F1Pwl2NTe/AbxsnAK1D1FlUYZJ1izW6LHq8ZfA3wkAWQkHKML9LYA
56sbGMHjvgEkz6St7dO3B2YEtl/cMMMnufD0/EPUSHqz2G0oaASg6z3vOseYTVOa
9QsKLurSXMkOWAH7fzHCdDXnnMm7XUz89ti781enXa2ItFo19dQEET0fFf8MzCe6
sTyIzV2NKxtvdXBN3ib6hJ+fSV0+CFEQWV7lc8JeRBljDIgpcoQIQD940SnyCZ1j
ycpVYR/oHrkHYNf6GJ/EHg+Meb0W9EjPC9MCTP5G/dKI92XtEa0DPIRq/M8GEgHW
LtEhxL8vvikRn8Nt7pBFzzlotDKqdsDRCrDlak4CDW5CJrzbE/5x1fE8uP+p8s6V
n7tMci7fSZ2iKFwOsJVU2XQJ7AE8LGdV/5/oqBjQXZ96ixSiHQcWS9I/VCG/BZmh
M2eiibTnMx+cCSJ3mJ7KvILIMrJ5RhQh6vnjsZ2xJN/zqzRLFGUpksAFFZWE6OAR
KJEfNJnbXPCuqNUuqsCbaYx8ip8eI/LeI5QizWAHHAaXDpM8FAFfcApPgsriartl
3V8BRpaWF6X7DAr4j85s/FE6sK+S941uJESlxdkCMyRQI9UV7G+4md2Pj3Ym2UMK
ImXcEmwbQpxpF87dW7X8vkmzMgVGS+hGvDPJFozPRxn/sR0YsXnwhOeEyXYXjP/7
U1vWPuHJbnaS3M19VeCVcRxtDUJzZtIh0Xfts4if0LEqT+eHgo9sGPSzEk3yZTAK
ZSF/Z3W4abz7WwEGwP5hdITTNDX4KNdltarfzh1AOUaNKxrTSMNLE64ix4OWCqbB
uVVBJdotxkyCu/q1poZzW5aO4vUd5M3ifxBtuz4DAkDQoYqDC1EVWCRUBYQCXbow
qXUkfIcKpo6sZjU7RTuMfuu2MtFuXEnMxOaAylrlFTW9SKJ2xib9hNVjr2VCyTuI
rkHj3cXAz2zGTDboN90Lz5ldWGuOwzLnj5C4vOUmhdJC1tE3R/sCkHS+kTrnjhPp
WzA5F5IqNa6Ty/YJXpyfir5QYXtilIHz5J1am2BQyCUll7cuSv+d36upFPGrsER4
mBLyBiQO4eYe3Erbt9gdrvgJSuju1gkMTlm4E4ahU7yx46MOsvofTfpGtX7gG0Kd
bHQ6P/bPDU51ey8Zz2QZQVB2LPkE/qyQlhuAL8HXK1Z1m2dI5elDJsWPYgBLbmux
zoDxns8oOc1aiSH/75uADtHMNXePR1YiIf+LqmJFTLhk/dbRf06g0MZCnd0Pooem
qnjiegeAQ0vxRXidS1IxlkOA4/w5PnAxCMft8oQ5dreWkeaR8OnKJWPloNEA4SyS
+m3ZEdgA7OTpoOMmFGmBPQunxxbohRJzhGhhRwJ+TeCvTSAL8D9N5F2EhcVG406q
VwUCCEnVTmIqBj6E8TcxrW6M0L/MChjHrR9DUZ4LusvJqevujsfEnNOMU4qwZj8g
185KUf8zzYjNhSM48JbVhpa6Q1/SsVScmhq2tUYtBVQXm+HieuTYCAfPXaJFls5q
v0oyq9hnHl9+j3VOwSqTWkxaWQVRsfzbkZsPb+ie3QuLNGyuO62ZsN7/DY9dT3fc
PU84VV+ne9be2vVhK6uR3SGH47m5pnMOpP8dUWysLfZdmzSk5279wWPm7YCbmaha
mifBKInIBxaZNkEWPKhyzMRPekcsADmmKz+Q0RO8oBaV8Q3NphRzHaKlCoZOV31x
2nRedD9OOaD4Zl84tzgdqlsBHupBH6W3RkVvmEgIXYCmLJQMNVXNAZxPNes+DyW+
hlKGCmeYvdFvqg7NZ1LzbRwnbxn4pcDDe8vM6eHhg4OHRC+lwahucuHMj2CVkX9p
Kl1FAaQrryPrLJjLMlyuLsl43RMiIqc38IhJwdJ+5duALMwnvDKz8uXYsNW0vocC
9HYDBvv9Kn+17dVDAiYsG5rFq9bNbywvLuCllmDn3rc5vSlEhFJQFCfzz25u+02m
Fzkln5K6rHmSeIrofsJNss/y+cZqloh0nqQ0EDrfmpUS9LouiFFrfO5kDpIG8ceM
BkCrOO9b1Tr7/rmFOOFbzfkU+ENfcWNe3l8bF6xMQqldtyjg7q8zUN2FGWtCWEEV
AszetSkJxOjPYNv12KxynhbQT8H0NZdMmJniA9K5cZctG65+cZcOVNq4vPnt1ENQ
8jIRPNFOGhZU/J8pCkvzd6XRoW7uWXm/x/DnMm4Sh4DH05Syn6DfSdikgVAkZom/
qYigZBZ71MeVHq++i0EL7ap1NB7vqGPhLtmkfwha9ev37PX29WE+SAuHiW9ghHV3
Uhh9zBrZ40kg0NkA3MNntPrxpZxQu9O/Uz+RQerZtM+N0PHVh1tKTstHX5CMgjL+
3Hq3qaIfYo37K/pS5ubIFFJN8lG++ZQa2UscP2tLBX5gxF9eJatuTvjQ9SC+JAkJ
A8Lyh/7Kuva/FV9hmooUfc9W5Hjpf39axj4yRDSOGmT/3MQryz4DDuydp4iSn4hd
FDIXhVtq/QU6n7ak/tDLD2lAZ0UFQ3+L/OCfxBLlJmLoD9pDbPec4vqMuA84zYpK
4g7+YJ9bFVjiQjnrz5hc65E5J+qS+hm7fN3JJcxt1n6XmP2XwB0qDpqiyKMoIKoZ
u7U5gA22wy8ZK1xy27tKM3FAXR5oEr4jozfCjWH5AzIklvW03q+T0fNp5IKuIM29
lLJ1qDQVNLR/DFTBQfHYXSWXAGjhmdpGT2OfxAa9r/C2dCSCuEPT5v87ZLurr5Ln
mcEQCSdM89rVSEFJgdoZdcwTuOsmSYOD8qMMzj5YTtk01UuGC1Rhu2UKbwz6jclN
C1pZCRayj58VyPqDU295Vzc2nAgqML/GLsxiQRUypjEaq8JZQiVBDkxdh2r7BCWR
IaJAbeWK6OpQHjSJUbEiBajdjKw3ol2ECoNIh+iJkRmCvQt2CxqAxlr9VOq1a3F8
etlkrAjxXNSWyBdrMb/dENIzPuRFv7OrqkXWN6YDoAOPE1GdpXe71PEoDyJknd54
Hx7MUWcahACFx4GF2Cd0mZSiyV+LOuVbmgfU36nZjACdwjtP3LfJFgp/ngbTSRWS
BA0aQ8t0FNi9GHwOmXBxT+P796pwkQQox+89DJPg/tVmFmrU+HJs6eK00MALMz3r
IlF9AehfSj9LMkYr/1AY19MzDw0j+hTydaAPTCpsST4xCRvdod/QbNZjyRZoDYpY
ZjJKGNM2fKevvCIkOPnC9BDTZtWXytM+eqt2w252q2WHbRkH4SzKSQjLF2NKtRGb
XO600Nqt4eRJ8/DCxYvsxEInEBBCr0lRJmNai0QcZcU/XRP8Nq9it5dk9r1ZTsqM
3JiC1UtHB8Xk6ySAj5a7i6mhNbt8ZasDwJ4ik+0SfCPv1pH4i+WjHwzibmx3QTnA
K1zn5/eu8XBijWFOtLi7do8kNqgxRlvB2eReNxoBTfeiQMcd2LJHUOMUWi/xsRX1
DwqyS5wiF60AXdj+K8/GK/HmzqkmF28005JLI3cxRNzkXSjbbodijnGchEQYe4AU
fmXpHa0RVpDbf/0Mwp/+KXVfZ9PiNo0FZjZpEMHiC3dM6TT4+q2SYRoyPGOJQiuf
Ne4CWW2HMC50gBSfi3CHOGgvdx+3oZoVjBNmyzA1xJVknMx4g77rKQ8RcLWjAJ+y
a4MgU8kjPJ6tlf3heXTxaBVSlh2XMrxynd4qjdlQGJElrevgEJAE99mmG7Yk/dF0
x09pkIi+gZRcSQhgLbjThdF4GxwVilZLw4Kza2jHAwYnpcGKKzhysUarBz9SXRnE
GEUOVheDaAR/zEJSMZ2gHsddK/hnTqMdcdH0SVg3zv1AhG12uPfzQDq2o4zJkoZb
N4o0A5y+vnwtZaDEOLJyXsy9s1TNM6rvZFHidHq3rd9kRdDt65+avz02QS48YRR2
sPdyEvmPzOtrbNYLMStoMXKE+FQDKA66uKAltyJK2A/hw2mRzAR+iuFKF9HfNNmK
vryGG7X7TfMpO6YseHwoRdsZ112xSk33OEs1DcCMAmcp8qJ75spTjqB7GtKJ/IbY
bFB1TzdLiaTFZapNzHKIS+VB17NqsktyhYIoidMb/AfZByhjDVHu2N0WSzpVL5vg
pazAmhd7utMEngO+3bhtr8ncMf7fVNrh1DJ7XrfHK99iPHLeaekV/9mCT8i58UBL
FE16+j4+jQArRw2DFxf5Y/gKp8oWd5Bt8MOChSYoLHuE6I5Cq+hrpHmMUoUfKgow
HPy6Eh1FGhXpczpyxSGc/hRs3e6u+WB2g9yFl+6xzW2+KMP5Gj5SHtO0QOhvb1Wx
QudCMGZdRgPaTaQuN8ASqwF0paiJP/8IV+igghN8EphI6Dj1mmBLdlbnSBABtgaC
6ZwSkbyTBg4YP17RFZ3aChfhWo8TO56CPfgqyrqGlfZOazaKweJLVS8Tefzojlzh
+mdeESl+2nCHgx86hTK860lo7rTTepztTaLqZuDNSq5iq8cIJT+ksZI3IKZ/KEhj
vFugrmp79l0QVJetOZ9BUcUkpENut5txHoC0EJINVyoqggh9i35LL+BBeBiEPPka
f7xLlzXtP3NIAmYyF0JV06a8RuEPmdFMglOpxit8dMFXhdmz7ne66FiOXa8tu/Db
R+4ClnJvcc5bMwUXDyuR9mL9VSUV4921L407oKItlSoA0prj2f8HCX8WEk+SLbPz
JxJa2QNlUrt2ZeMaatUu/B/kQGQGOTNlSX+zq1p7aCkbcrXVQeuneqoA6aLY+FMI
LMm0zW2PVPWjma7WQ3sNTpsqfiyOS31xcRzVxP+sV5+t+LjdYdkQ7NLhCGHrDQkE
j0EOOEUzX6I5L4Snxt+g5Q6070xI9tw+Sypfnvyw2xOu47na9KGYwSDK3FHDtDwa
Jr0ch+VyYlUJY6VBwqyCQYTyKX9EvubREn3WrZsUMRvoWOzQ+/HRtQDDC2OdwqIV
YhG1VCUquOuykaGU9PXDKlwwC7v68fj1rvj+b7eR3kDR8XJuCLMMbZy9OKhpXcBt
RKkv76xOs/0m9MMIYgV4Q3ZMQt1Wo+MdoUx62kIw1Qtct1pljA22A6tvzQIp9t7y
Mvhb2BPj3Yjmi4UJqNy5sRlMn+IV+FoJZIGb70ajPCRRIDneTPFTvoTBqq03aw9Y
Ahi4N54At9+2YYTk/36xIGCDFFPHU+5WiAA1Vbw9XXkhReIhhHAb5cM2xDmROBF5
uOmrkHQHGUHjkWsgX8R0El6fTNMOlLCddSzUEoZiGacfy1uRKEYCFHOz39hAjtR2
CYvKLTyfTWMPwFJDtET1UJSY+K6UsfbTNY9ko8jBdfu1TCbTbzR+wIzvt31TMshV
H4kYK+JFTfnwU6GPQmJdqPuwYtf0rD/PBqFdr4RYiEIwc9u+E1Ay7/4JrkIbKydM
MjMy/THtSc37daSUAg1WIm4qhIEMDrBybhJ8Q8uvxOzv157dqf0KxNCGyAahz/x3
AQsXe+pcF6+XavvCXOFktJikCOY3WIXi1gitwrgV0YdOpkVJDSjqUJAg17hksIHV
+AALCPdOhVY3A08xfXe8roUm4aPL93L9I4CVyiLniMGed6FUElsuOoGVfmwnnkSb
T+ASlRycW49vvfwYgfp0QTiIg8KOfgV/1HWOMSOSj5OMlOD5dvWTZQsdVSisV3ZX
ZorKh+86UOuYLvEKYI2fAkK5kiISKtblEpwaEFTKFZk6TprZPlHlO76q/rnRB1q5
IENizL5awLAqjfllLS5SCyx40VRHGVtE9olAvFuslMfKHLkyCwbiqZValOxxekNW
8/o+HV53qmPQfuEcdHwG232gzoMaW39rO05/ZKGBLeJSWkS3w5yV63NQvGR6Ey+E
4CPyxDD9jgaKt3pekT7A1lgs8dkD2Ni8LN2bo0Xx30lTitRmNl2UUM9OgZ1APImy
8bUWJjnsj9I/XCDwrbZbWCtHZut3F5B0+8u5USWmDBxb1AgktCwPTdNIQa6JaF9J
THzO/TfWuuWA1ip7OA0rp+brXxi4o166MBW9rgPXicwz0jy7NR2TJkrwh+E9r83i
NoqMyIfkLBU+mPtj8gptEImb/ZlNg3ww8l6OXpHomHKWEYGMtVbLPZkAe9irJhTs
QjNoSqQxvbIaAlry/09z0NIGzZ6lgSV2ZyVBfOqUfqKR4Q3VxA/utyDBoeSOi7CI
NyVKa+yTGJJZaJxOud3tzuhYwmHHyfdonwFhnsa2tjiAwZjlq2WvVhnUBPBOk+IM
ax5Oz3LtjZFnHo3VL79NSNH831Cuj42rLZBVt4Y1Slz4MlmVCk8BNxkDosDGGxZ/
mbOkqZug7vrRRqz6qndRUlszA1xbCB1C9b++ODvqLO64ZiohSuA9MFIzhJSDrYhs
O+iSmhb9JrwG5DCz+ZM2WbfkMCt3pm1Hefh5BUgHH/lQAejOwInvb/hWBOGB9Buw
PDXNZdnQ5UwndOUkDO2grguaNwH0M9vOwhZ3YAyrTMTqgmHFs3SdnvGxFCSDxRYo
L0JReCkGqERFL1+6vpab7DdPxi4kmNhE7vs7iGoL+KAKsE3CwG7zOovPA6yiCwYF
oXX8ADXYglD/xBW6eW9XDvMZv6HOTb8jBzi6qYusWfIra52Pp73OsWe45R/XJbWL
GOgkYiPQABAOqVttml+cU5rDskNCxwil3KudPFM3QhJ1z7E7vlb884MTpWVYWaIY
O8gdccFCpDvE4gfn6C0McixovpRF7OL4hcRUUTM7rTKJG9Z4yFSKC0n52K/hyzXn
4LIePF+XOsR2BcYGtcj6L7CrUEOQGiFAbzKvR5N/Y+CVGXQHUCsaBCDNZIK+llH1
sHduwTyACW+G4pZfMg7E1hY79UlXX5hq895V2co83lkC9bMRgFmHTzJt6gEhpAg8
GaIh350sj9t1Sf+4DuIj2ewBHQFYNY4vQGFGKiJxeJr1GSp33ncPpS7yOf8iu9t1
sNRYuSWWQ87fJcGFm7k2NeXrwFO3BnSmrpzrYVGQOibdHzQZv73GWPfEyuc/6to7
JyA1uBa3SJFxmulFXwypidgF7QxXuChkMn+CyOWgRAiOQjT6lwaIHxQhaNy8NOv7
ISPJMn2RhnMMuHo5ks/PX27l9ME+AxjibiTmYuDXq/gG3VY9KXbJwmHTW3HOowET
zm6S81TCpnqGFoPA1g3folcEu8huYCJ10zUXzopBdKOwfzeYBMmfj7NG9PaeGvLl
xGHueNhNYrdLrKBJZZ+XM9YRxi97xxCZghSy0WUwy9cezdrre/JWqTp4w1Qv5oiu
axncORs1YV7Ol27qeP7BtUTY4k0/25gMOBOp3UQLUov+1tncfeN3+UxyHek3AS6i
hncSYY1R6Ufn8WZ8/OB6SOzodGaowy0PuFo/pcOSCl4XO+iJwyRfFzQAvxklxRLA
FJ5aXkwjfRy0bfLkzXFBmg8wFP4nDQqlFJFn+gULdXWJp6ItIqDjDHWgUDd3u3n4
w6qbKbx47XhxH5XzPncTuZnFZhrMF95xH5JExiM4rzjEw1ybVAt/d3l0EpVfEihk
Alz3jRDjTexQVRu3P3xteM6vxwR50ZN/L4BdKdpsGXtSiFyWmzFqOE3lG38YkGyV
ZCpCPGUuJtIbteTiQjvRQWHvzZwhM70iPh2WOkldDiarWdfigdIDG1Ra7OOwHZou
fuqqmm4MBOk2oXbSWEAPWo93UhYPvGAvfeJIaUkekGp5CjMh5ijMCP7UwfuhzEfs
86Lmm66UbsDVdl3d+2y5V9O7n2Vb0vlzFteRKNoSreSafK1pV+heDNYYCJykqAw7
P/1TY0sUx1xCv0IWymaIRw4BavqEvYeY+6Y2qYp373WApX7Uan6NsqWJe+62Cjtq
pQGAAAGTJIruAS/eyT2QNFzM4WBcT/S0eZMdHx0xNVw8WbkRJ3dWHThdG/20q/Jv
A6Ca8BLEv7goa2TlKom3Gg9SY1CoBHhSYI/n9G8vmsI8d07LcLKRqcAlDnkcUczd
VHaTQuzCNptkgvJroj4Rp0Ych3u/BtlRoKPMH/rKSwnhGyTSbLNA+H+7QA3q6l2u
2kyWLs1F9y/Yrv2fSuXKaspfZ/v/HMMoq0pVSqNCbiIImky6ndBk1PWxhvXDPoTH
iycS6yni9AtobGAdRUsV/nlAUokp7XyRL9dvXvv1n7DA0G1YAu5UMUAobJZTkp74
kT65Z6fM0tuhRkXWet0+OIevTzO65wmNGica1SKGginwJJn/2J+xGR5Da9HLDRu+
mexcO1gKja/GQif8rdKebCZ6xkLDLH16V3uVIqFZbe3Qb+ttXAzdxN3/x2wb0Rpo
tCddONrj1Dv/HZcetq2kGtP6YyD6MWk/C04hxzkGxFi4oPYr/5LDtwZRpozNyHKC
D8qmfDZIdIP3SrwhH39Cw+5Dbn9KRiXHr2PHWoWOO4oGKBE17NZ9Ep48hvhC/r8n
gzPpV8cZZTGi1vP8lZjW+KatJp1Twr+Jhi0PW2prO+J2CsE/DNNl5n30ALcqvBab
/I9yVWGB0VL44oERMQmPIvp9JuQeo9sx8kJtlZp4v1swpvzGZIhZ5LuHjkT0QRRP
IhhJPcvXIjgclGdamJTrs/LZsXyPRX/eRbj7SrFWrrsV5ogiIeOAcwyv/4vRh5kM
YNx0mLwZlFPSaq+F98O+i+SmaL0phJWIZvxVrNuVqmTNiLFhOC/7IVUbAYcQ5t+6
btX3GUuh9glKUSZs5kdBhcArl6+Vc9xYHFFadwvl+0+JNGhQvVlj7vFWEYX9+er1
WdjEKHaZ5OCdCeGywPwdoT0grseXa0YvJQILYiWygplVj5TEu8g7Rf8NHkxWH8hm
jd+1MSFjbotm4wYHUYOQ17lkwT0VNbgJLK+MGUmFeLmEq9trNZH3VbIO9oYG1WVw
3ABX9nmmjx+eOnNSXuiZFA1QAIAwtTRZX+vBavLgFfFIJLcKYVHEnQ3DIog1SuTm
Eob1a+QerwMOnud4UlkmDjD/RaZTa6g/3e1eJ+5VBRIlBtiP/3WZvZhGShVXn+3C
Yy6yZljZGpuOtu9tA6sZpTvTtzLlnz9c33jZRMzMC3VjIgKkS2DI8+nD1wYYjN4y
1EjuwrGFBYendVk302J1/ljhxX23mPWYERtN2EbBydkm18zYh2PSRfi4Ze2d2usV
k/gH/aYgTAYq7947sSG3yJSkxBJcA7O3ztjVPYzVuc2poIlMUdVp+c56Hg6BtdSx
wDbz/Gi4hm3GtooKbz0WcpwwwfanmfK6oAUP+ryNJ6V6ECLbpxOtdasYzKyXC5kJ
sqYKxhkglRbtQzo4SRBu0xpUfKrwIj0hVZOpv1GtINorAHIThpW1kqcIQrXFJmpM
mRdy8K8lQZEmrByWBCq8kPm2Hn9Zoqm2EqJNfF/pSKqvkcSvcmmFCPq8xbSNrmm2
PlNsz34IsxoIzLtSRlEk0n6ybwuwCbFspnvYtrkq2d6AY79SQ+5Fgzje2gaLR287
oU+TKqoRj3vIEpF6g2QiP7+jwiTCxHEPgYUgsJnl/vZkowTTrTmk9MqLBOQZOzDl
1L9dEFBO1YzM+G9Dq6MmOIiJJo6/deCv/cVb3QGsIAUGBNEOYjv19PlnA/rfMm2n
opQW5WTS7U0VJ3P+tr9sX0EjW+ULzd0okei0coglVcKwqm4WHbm0cpIL8m+JWWca
5IOrgRqrpATG2KxFxjqOAUruuVKCN2OMhkxfLmDBr8GvCk10aXVV47hlIOi7qb9m
uNVqz58Sc1zKZWp4WIeX5KtwsP4Cuezda/Vfy01636aHc/Lh9TYa3WbJIiZq47Mf
acVTO780LQkRm+i0UddELiyEPwogqXf4LjHzvnS72DvLgfFgJy2aAmxzTOZd8GIs
c0LsK9qE6N/PTq9NMUD0pAkgpT0qX0Zoq2AqZ8c9RQmpDxRZzmppVjFyY/WIXf/q
pSCFXymuIkuSJ9KrlEXuFk1p1IoR+1gK7ijyUh5cpJ+T3DJ714gYUWHhHiOqbge+
aMX+gecATj78NhMEom7+Gn5DqioKLP1gq52tJheCP+KG8D/4WE9LFhtkTUIqdJgd
5PE0iPyjMeIwF/LuLmcyoYPsK6DU/gf3ar6MYIrdtSZPD8qW9p9MXDa0/T0K/ulA
/rOSZ786A2gmQ8k081CM9q9WRffCar06XGVm3/XER1u1YzRS35gUrcTawrxZbj76
artYFQJXjB3Mrqml8DQjZMvalPKGoD+q9Rem/uUMP5ILTDNuIV7dVvbhPDhH9gt1
iqaaLQcy8l3A7vz3FhNMJ1mklF92nq8SUJP4/zT0UvPNsDEDJVQGf7DFGnTWVrLT
ipWqHDyv4nWi2XUNbc4vcX0wNzEAD3qNM83vSK4pMzUdXsWEwYDuABUas3eO9kCN
OFq7cCHmk8QqvpUjqTN5qbnVoS12Bxd+NZMBcWXzJh5LluKeyFsVNK51Imz231mj
QGwJ4mRcm6F7v7mIq+X0F6gfc5X4u4bCgsyQma8zjjjEYwzEJgKUN5dYrBEpbvXc
lsN+9xroLNzTcC+1F8orx/2lD3j2RnFsd6NGgFnpCTQuUzZ3SDSUqytmRNtnHGy2
m18Awb4VypqtGuAwQvd8IEJf4Xng+NmAD/aB7DWcuUKJRyfWXXk14jnx10PTCPzd
xFjbtrpxl765UAnhi4d5AKXQ/P9A9rvlp0/fNhQabaypboMmEVYsab3ArLc9MFDK
v3AZW/tX6l1KX/wuVPxgObUbxpazvz1Tti06dJUrhyW3jPUe88y/JF0pS+gPRkZG
AjsMyutwa3Ia9QUB5UPc0jTT0qnnBbQuU1Kqgej88OwwOn6CKpWDNudaP/Xj5+Ro
ZJ7xWSv9+AywDnPjaBuVdtWT9OhTo0u34N8q7YJ8AK2xDlmgaLUBdIqTBQqeaQwW
C0J0vcyDGfjOXQJDhg1ucBYVxMQExTfcqkGRinmKan+iTpbKz+iDIDMfl8Zc+psr
bLGJALZwtCg2BmwhcwVQAvgaj5/oovC9hraAwYLTXuFQ3jA5PGEo4Xu4H8XxNSN0
kAHQgKanms+UXGQ7tg+dcfn3UkpmycShPI5kl9Wc2iF6RPGcBamDdO1D3+ONIhXW
G7k6noo3qUaIorKCCbnGX2iZQGFxVGoMM426tsyt2RJourIo9fVqLs10znDsLsvM
v4cFa4mwTXQi7ih9TXWsK86wXwHbmKQtm0npWZ/jYlGUolo7hHRf4tMw9SwCaKKL
V+3ig96bGrm7/06RDX4jszIn52SSqelphKaAec0Uzu5RHHBs5LyT3BS0ubaa5W5u
d7ZAZ7cBzLupottVZsCsjWQBsFQqtGHjboSiT+b5tXyFs39H9n2QnVKPax+PyPTN
8EFlj+wuKnvepJtBORZbmH58CBhFX6gc4MRy4GlvM08KOfFmb8BswwzJoZGB0VQG
N27d7iGr8TQIU2GPN8UBJUZGvMTXR9O75NDoIsiMR52igJuLEsb/wg060UvY4jrq
yRkPzWbPmvT7RC5LFkCrHSlTNEpDHwcpGbIS7n9sXVfn1x/vB3XphJdcKXnq8BIc
5hox+No+v3vJBkiBfqx6qJAto6e58KcVvxqKQzYuzSZmcAAndNAW3qv+H36kpd6t
HgAq3Of9pjsI0aULG7QEWdB+SKu6sb7PrZBsZPje5k2L1yel2WB+bPOi7gmOofJa
RmqHDVlKRrHE4vA+iQSHvoMJ8vt9+Beo7c9n3CEUUpuRWv7R9xV9WhdWfHlfeDx8
zJtZXq5rUH1aWvFjesbg2VicufpbuducXLumgDVyJNC28ylDQlcsPJe7z8ipn/Tw
aH4jACXllDfcrsTaJ6Xf3cD0I8KfMGCDDFowkXppyYINDspfyeI/k7qcthVl+Fqo
y9n5WMt6jGIQ2D2l3eV51SU0H+vom67UbrpKDHKfffwrXvXcFbQdDroQFXHbHrFK
7Z5AZ3KRvib9dzrkYYku3KjnXdS9IiOlTkhyPsStBF5CMeRg/SFvhm4Vk4j3327E
eP/5MqsldlAqJmloIi8x6gFWgZlNRkh3NVJ8KTMuXZ69x/LNziYW8LDb7Ico1t8M
2Yx8LC+lh5Vh+3Py4RCl78jWQsCeouPs0rMoYFmTlHhJaKXoXdv/nZhP6FhTKz8g
PA8Biu79MPingNM3SUk+ZajGYHOu/8y+BFc/LtMmtw0GTqLpsJxh5Z7W0ThO5kkt
L8Zp5cN1LtHmG03mErKHyrTWTwMAWBX9FZxeDAABM4bpcNCEpbtIFHK5IIgr5dhx
IY/yIypDK+LSUNz2wH95objvPEmwwxaUR1Lf8feKkufw/guFKfRzkabeUdeHjhJp
4rC6eJP5lZdnxgX3krQS9Rkan5RjRWTmN1BSa4Nd13hrvfLvh9/CBfI/IyTAxnfk
tsKFJaP06Chp5NvgXXJDl2HnWzNbqPdZcgqwlWrUBahkXATry/nfaU+wjwtaoYts
4XBsZvNPjJNGAfWd8Iv8rBT/WkWCUAdsGhvfwaHOnBb8lbSVJ/fSXSIbb9p05rMf
IgZXcKckLEwUyNZGxcaatBG576hfMp6tsKzZcOhIHbhxS90/BgLkuPM6VU4vDfGw
u+hVck9qc2xEqiqM/HPJrDo9ododXk51SwGQvBNd/QTwdmIJyqWw+kNpxuVGXfUb
1bAADVTjCTt8wLwS3pQLuviNgiAAR8AHR1xRq5t8MIp6Hd1udcHGPiLkddl9JWLp
F7W1klrjUtPv0EOKmvzryQCJvrnzg/NnU+2CC2afILYbP+iVsqFIcm9Y+uZ6bzzY
P5xYYthqfnaVyg6eFG2iXxNTiyy82uZT8e5ive0G45s8RTCo2PLjZ0Uptdy5CaK2
csHm0tGWffhcZ3YzGRM4X/3/H9gzNBvdhtqY8SzSogtrFocdxOBL2l9g9V0Xls0+
pKEsB1vyEHZ3bjogrc3ursp3rB/TVdutXOYzQTUvzTVJ74v/9ok66KapUuU5bgqf
1dK9WyL+LugH54ryRIEchcDqWGz652LRm3UkpduXHmR5pL7dyK4tVcWSsrEVh04g
PubJzOW/SMIUZL55cRucBcVRPQqHuS7+qQgSkPutE2G808WC1nqn9hGi1aFcZGLT
S3RJdb6Lh95SpeK5Q17tdhF36CbU/BebIAAfyrgh2s7QlIRePR/fiQbLUijqh1Bp
4ojZkgxunm+/tQCq1UKuPsn35cC2FpySnFiUmqqivrR7j+po6wL/8TL48bc1L0QO
SPsN+Ytai5efHfLVk6CX6p01X1UacG53SSXXClRZd+AJZNWPjAgXDTeT6AXJlehs
PwLPkPx3BW3Rzm8SNTr+TziF19ht+mV1B6BMXOuXdslCOMsm3jJDocM+CH/loSNs
/+LwWkbWuY7NzcoworzEtMB56nTAcbCMy1ziJCz2k9q0tR7pTKOZ0iv6yAmedfcw
lkG044EnKbBzbjCuGj24gJUz1sMZ2YLbttG56FUx8FS4jq+AwbUnOQSo0Bxru3Kg
rwCg+piiW2PZjdh2HyMhEDdiP+cnBTXL4QEFANw46HonGJ4GEOohoO/itqUJmQr+
tw4mk6L8QUqmYuGvz5g+V5YXtRq5NvdmMca/hW+ki//bBliCK2N7tqUd5KHGCGSK
t/PEVkU8nC8LoEKCsDNHozLawdqzjYmEKmJJDwvBcynBt2Ywi+GtENnRXy3PGxxM
s7EqmDwmurvKYEmZmFgDPVhgr/9LTHhSbnRXyrfBLlXwHTiUK9bvqTy8e2TsntM+
RWzb2SPeXK1c+y35KEi0Bt1ihuMhJyv8VdEpFoeiFHM3uhDx/goNLrKQpW2cHXLP
f2dA8axVsAKx4m6wFyyH+ORC1vICYsFi8SboAfbnRWd5wSM8sMphLHepm6TgXG08
QTZZ1taDkm9aCy1UvNn34yDOtO4TW7apm773Pru+Di1L7LkvwBEADDFNqjtyIcZ8
YS/+OUOL2/oMrBLnFPMyzj8suP4TxBPxwF+nOGHetrUC98Q0WxD2CMIcMWs5GxyS
AW66z9ofjsk4DQE7iBD6DlCCNfiu9Jbb6En9iwx5WgNl7oODBothCGN7SmhBHhcZ
CnBTZiZHXUhg9keqKZknDUvTqpgHIwL1M/cvSOXPJBs0dLm53EHfY3kM+EXoCLQh
mav6X8sl97QxF4AHyuy+8QPX/i9f3GoC8dAs63ZTOw0Op8Cb33fyb4bECjBRJ1wI
yCwlBp2oF9eU+CI1dLhIlohRNUIMUoeA0Bkfdtbxi77h82QmI17P+TPcaEq0Tik4
ZLDMbeOt/nl6UXiyH5QOlPNJBmqBqseIXOG1sK6o0bDXKnrlpai5qBoYhD5dDzeL
tywNJX4gjcCDw8riMfaYDDmbjt8iu1RSMRBYrxBz/FwlgORhP/Lo4ZTNMr/u8Gt5
udq5YRtPD8Wq9GGpiRfnAvFGrA/dH+OG3/8Upe9xaCLoV5Ro//rxDxjJDITDz3iT
bYlTN2oAtH+jcJ+BY0IEbeOn67JO2UZ6LgAMHj4phujKjwO8qr9amcxPOwGNQzzn
mOrZNjUaTmIftD8u2QkVoqSfcr7JE3l8GnRGm4N37qqwiUVTgozJ8RVe5lFc6vy+
UI53xEuE2Y5snQ2D1FlztsIilHqsWLnfo88wWntbuu/6LC3PV7xC7Ll5PNHbumSn
zEhAhqjvxRljBJ+vA9ffR/7kNXx7cY8HVsTvBsMke8VISxltJZcKgn6nvDb7gKjs
ZDwXWGJvJdT+SKlj27uQuLk7DoVSG+g8HW9Du6gbOF9aQOaF7JljV9yQQsgUmbbu
UsOlqgJ/JHTzq3LTr6xIiAd1YzgffuhdLUCTeQEEtWejaK5mopKwbmrSIwsX5ihC
p/2+3TEsPPRhCR2LXSr+Gw+AMYlmJyAhQrs3oHJMZmgTGhMhxRXt6vYz4v23sG9p
+0omo5/+tesJbFHp15S1XPnhXKFZrsFW0hTQ9zL5Qk7jJd3NYvnTW9bSLQGHf5aJ
EszW3NzoERqchhP+5xvC06dRCwvV6/hBlH7BcFtM4RwnkhoU/bvTMgGfFCRmzxLP
IhVjtnYKIIaJMCBeicvl08fM1fCqWsunixLnVi9VUceIbQXLCx66FRJVozXNBek4
SBXad6qRQTiFvdYgrECZpF6k9CGcuImlpZHcFzZNHGBqrBZaUdGdkYCVqV4Ac5VP
pxLGX8pIbt7m2cowr+y8vetLiw85eTfRUfHy0v1dbT3NtYGmMrCc6mEHRPxYK+T2
Nxduslxb2NUxOsTq/QhzjF2ke9y9+I9geCDjzEad8aeEhrSE8cR3X8KoZzL0YEk5
raFXhi+yfHUPFyR6QMjDKbpMutvuW5poJtiw0aJqkrn0/Zp1F3RwiXAaX2C0TgfM
l4SuUSPRU1g1wVFN/la3WmNfW55H6asx0t5gCbGmOKPl63EPaDZGFUDeKNCsH35B
IvXWWXdioGvrbUckSXE7npGAq9j6RC3ZnSneYZjBZmvd9UEfGaA8OawmFdY5SjKE
Y4eTIJyU9eFM/rm6v+vlTjWgcrh4VcFZH38OTo+vJvbOb54LHk6I4qFGyqVzA82F
cQJ67RTMQP5tfq4qmCL5guVas5CaUCEdyPWQLmkAEqih4Ts67YKrXy2srTIKj4pK
FELkKcks7xfkLMdlxIIbST+GkzXZyRk+NaHEFVJ/Hbpctm8/As2KQ+/x5MNrePJr
OARbQR3ebDs/cZXK9iutK2JViZidcgQv1Ny0Tmaa/XkMBH1MhvgeiJL8PzIyfn0J
FJtJ6jHbuNIZ9aF9Ue7TyLFL7TZFTQcIMXvvyxCY9a9hS0clGhGNQVxFKRKhBeEz
D/KVkrz3Z3AX0DwPTtrqHCxM92GkwZjgxVJF+YsE3pMszSHFY5YlnOBd9xwKYcj0
gejWxxxxhFnsFU5jDIW2QUAKOZaSsxflhMPRovfAVdaW5V/MpJ+ae8yf5DlnkK3i
vLB3Fw1XjcMhE436HjfKm3ql3uBi/pY/ijWp0MU5c78wfxgHJnoEzxiqlhogIGe6
7w2qVUIANhCigrEosHA0nrU0vVEEO37WGTXYDY6atimxBa8VzTAza1sU61Af6Hw4
y49uVgL4v/RBHNazPvBnJk4Fg4lholYdPingseBEeIZOGsARyyhaWKd7As84o7WG
0KJHIUx3jjT3aUU3N643+O3djNzeqBocLltpH8Ya5bfADX3xb5Uxo7D2+HzUQddx
g9UVhoyFl12O7hGoiKedCeRaFMpfz4kORua80xdiAO65Pn02jPHJczxZOSmFcbW+
+8RKcSbqLbLbfAWxfAVCbYPFLeu+3Ik091qz/2nqlPcv0Vnipf6H1hkYiYm0uprh
mARFCabVZyoxCDD01NzzHm+OOF7+HoEqn9N74qXuL9K7OcwH6t7eznUm9IiFJQqF
p3VPqQK7BajicWG9p0/lLhhHjUjFXmxaZ4iQE2YtYGOGxZBMnz4jPKc8MTtM7bHq
2/sPwEzKpkKaJVDhNr4kLL1iNM8Ub+L2lnmyNGyUwAHMGW+I8GX3Fs887G4aXchp
9wctpaIIb+cONGE4n7W+4AH8o6dStwhpgOzAxYRF2LvktD3MBi7Uc7xyGS6PDBpS
oFCCJXp7RnV7dzrk0uEIcW7nlsgsOuJu9ahc5a+9tbIVTNp1XuocjksJoG/Vc+hN
kGlgylE1SXsfJCt09M1U7EFKq420phFyZnOabP9D70dfxRaQ9bzalwHrcDuNSrEq
NLXW0yEwhKubUNnzBEzNMMHNzzhCSFoToRgloBz7Gr8bpcOdyFtbexcFuDlD4SFX
ZtUqOpTFUjnBEj71sdhjLCtwVnyTKtWcTy2CUxmWpM6/u4VazSyL7V14Ag+YxOmv
23uq4uOT4RhqQpWcatNnkjGCeOmk3MAkHnpjURMC3JRwWnwYzKz/PGO3FXdQv6/g
TaVatWAOuVt8n2wuT8rXBDQTLQa4PpPATmsidrsOMeYVGEW/LauyImYDxu6p6Dgd
U5pnR/qt04FZ7gcm66AlUrVYcuCVTY2tlKHldW/SRmcGcIXY2CpO8+yJKBTwNKfU
ohk0uv09/bTktzabcUD4KMyfDcNpmDhYVytkfjvIk2zl5OxM2HrVG5LBuVnh7lG+
PNvoLXVjhidu8HYjBuxW/f+EZh8Xt34n1yKVpc1wwFGBgfXo9Q6O/pvUbHkqyqZb
S1ou4Se5apuZk0oK/cY3K7EXEtnC+Eqdq+lp1qE3fRviKoiJ6faF/By2/PcBMarg
Y89KJyiqjPdMFxCIaOwEXqlyReCMCxqnX+tBThKJrb/KlMQWJUrgyRsXcwHK4ZaG
9E+N2/D1esUWs8tBF5PSRoglRYC8cotoSunljxbhIXwLvzRcpTMMArGu2ORWVcHX
zSgYA1olhfh2NYq+l2UuuLyfFPmRHKqaX4pB8Qh6GY+P/qUG9QvK035avBcn9e8Y
r1HPdNvgt5+l+Z+NGaIjJAYZPnI8v+eb6NMnAaWlgoYV5i1a4kECu+sWKPKgHfXV
ciRPL5bsWO/yEzlaEWDeXCQYmDZgOf8OI1YQz4Elmzcrrk24z4cwsR7bZIEomKKK
HSqlFLUztC94BtbKY/q2aIeRtqRZ8wTj9MlcgVGoIC18QJCUPgUKEGIrrEJ8omXJ
AFU0wlc6EyMzVpT/75WErIa2eYa2wGoq+v2RprTT46656k1dQuPUrUFC0efI6Hkh
rdzIhhWORgI6FqxXzkRL+jWTFAMmmkaYoRsfhSMzEWbeEe7/ccIlJUU8vwkBlfmQ
Bjqzovxat0iRhB2cjldBCREbdAoazAOucwysXX8+JrvMZZBykbvARXDxN4+F5CrN
Hgrdtm+19aruq8rbwOXsrVzhnk0IMY6rzPqOVRmAh/qUTKrP2UretCyWNus9KKZS
5cmCdasSd4MgFUjBVRiSKymSbV/AU8b7+AG7JIxU+P/IWiIFfayIuroIZIU+bBip
5o4uN/UEYuoxvhiZqUEBJzN7TMJbh8WN7dVHA2o/q3NxIfCmmxwLhqUQhC1o7Jrj
jFTx5BSotV2dHDzwN3AWlOOdnd6zFYIToBQlZBn5dgMDNgBjuneuVPtCTS7nhf12
FK1VgT8baupYFawKHa/sPj7Va581aOC0ryyZHCzQ28gah9NJF5++Jf/hFKcTU/8r
FX5WdTNZN+C34dt1vRosl0jFPIoSnATAAUVY2FIEz7mLZYXKI2smXuFz5L/iuk4v
YlZTMy4Mt+IkqtZE5dLci0GKc52WEEIkuqFl4xD+0IBnuQA67HO8x4v4Y9YelLAl
t+Sc0Uk5xUCYPwvKAi7nGtm40Hhse/RyKmXtHgtPPRe3xuD4SRaACreocDgJtR81
gBunXh2JXzZIsnNnEED3casYCYBzTNaA1PZ4ByvtRsREazHuWET+rSJJWjeSvzWi
MsQ7ITW22nAIY8Gp0mXs1uIhOcmJzJKJ1Vl5Sf7W5N9OybznbEvYhwemQYih2v4Z
NDhppLA05ttchua+sXDY9HAwkH4A8HJjQDhF8IOUa5KC0kFjy3KldjP/g6on+KrJ
z1lxiKN37nRzDKJYn9+RR22Da2IR7W4DZq4kIXU1Y0WZpnCKR/KA8+RHHCnHHWMX
4PTU7aLCMjmp8mfPFAMQEcOuYgk7IPunOAnnypUfgrOndr2QqKSLL4fMEEXNgaAA
zF3BDUEfkXXwTr9Q9RbJzd3MTPpfCwKEzehjyZO1hHaeChI1wFMNN4044nqm15BZ
reroXN3+wYoFcZ1fM5KCvcZGvx9wQ76j2PTnuJFL1yvrhW+lWAq0hQT9LCyFmUkD
0DaVIjMVmqZIiLeKsHapNMdmdrujR1ZwifjFr5tPONhfstIwGzDxA8mgMSLh4JZ9
c6GhIBJrdCVW/dwoa4HmCVwMLVa8YwaSuSrdwoQg2b10d8yV9iCqBAaKPwV9NzTP
ll9WhxgaxnErpXkO67e0/fxpPEdN07KcIa6kEWiGvGqd2VDLXBA48gXy/X1IKU4b
Qtxq6BfP7sBN97eSzL/D097SwdzS5eD0dVL8MhWZE+FnMIo3OaEWwTiL4ffwpPOT
gV+/SDBBV073ZJAaO1CrvzrL3GybMWm+N0QB5YBunWfgqUdhHY2C5iowRMCl0dCf
RuPtbEAobFwqYBPTVPipyBZqKTZem0GWs3osQngGCGUHQpDkV00qmr4NNydIZM59
Ji6gxeLkSllCYSuaD0Z1XhiCLp7Z0RopSyWSzZ4fJePYgV8JAA6Osp2zeWmjV4Sv
uklEu9Pmtr0FNOKzWwHWt+RnclcWt7mA5m48Yx6bsB5G9y6eUtIoBuZcr4RPHeR7
FHa0G4A9qZ6PzOVv+bDWOguaAzNJLy80JAw359k2m6KG5R0j+C2L+LYTJ6I/J3EG
AUMIHzt0lWkD5SnzTo5XOJUq4U0IfbG5OM186L8yoW4u23Cg3tWB+LnGRoDrkOjm
ZPrj5Mn58XacLi0EH/6+K30o9ZY8iXKQqsgni7qX+ttKb11wzBjGzT54yNw2x1fM
Zgb5g9+0uW9qa/7YwBGDUFDuqm8JXOpsk9sNk0Amp4vMzyDbbV3ixL5ps05hnIO/
ozuLvxf/mA41a0/G0WYxvDzZ7cWUBzzFAkAj8SB9DTaOrBP1jr85xwuEcghx8thb
5etIG7uYVRWxZ6bm2spCjGSMROeMpGseofmCoymVEcj0h9KSF0Gik3hZyWymsV4H
lExE0LFmIJogebWGWo3cIueeHNDbdeYYLV2SI5SJrt03+m7msS5FrwasEw+tgXDj
kHOiZNxClghyn00DCOnCORHn1/NkVkat24u9hnf+OVS/MT+RbU77qpOhNpqUpaWr
jzToqZm4qPO05v4gaO2QMDmKjt5p3adVeCaqJCC5b14+8emVmI5ygkeZK/1IeJoj
vUsea7x7DFLODs6dAjmTuIjnnFAtuDOTdPhFhbFnjNP1qMYBV7LcHjKU0MqtDD0G
WRMwAPWJ+srIGOij+9U58qw/cdCwJTZfsVYbQ6oRq5eMYWHk8LWyl2cYgKzp/eBZ
qT1p0pDOms8980Psrpixdq2anVQgWIt5UFiKYpGhd+9YE1Z5fzehaCRCPS9hHfvQ
xmz8JW1UEhll+JJkc0wXoCp8BbmgVs0Xnm5w3UVr0inBhbS4H7AO0z8J7kEF310a
N9iaSjzy3L2f/PpI3NrUGlvstGgjWJ2u9I7yMBTLINvYpppT8Kkfo2mAuUJ9gCSV
UpK4+0lLSHn59kH3cUDCaXkvd/cEKQLrXGHjmOrfcw23ObZygjKUNwsa73kiHBrd
45nbsDe5IJU1q7C+Awal3vu8iJKadE5G3F3v6/gwVD27lciF8wUWq6ZOsNihzChP
b96mjDe/jKtZ/o+RR1exmcxPuEYQNfGMMWoPNWDvKtHDf8NZpHz/uw6ycHCRn1oK
2XJS6NUu1o9Fs3GA1AmlRl0003uM++EUIRWuoayizidYsuurnNK7Sb3G5HCXrN9b
qJ9Gv0I2MuGuHfYIavgC6hv0eT9mkt+ikvrooNoy8LAx0N0bKo9lu4q48WWctgHa
jL4fQ1iqTeBuVpr0GgAfZH2iEATc7cyxvac5EqxnxA8Jap59NlZWcOpZaVHq0FgT
HhRhkD30raChTpKv/jg7YgOikB+C5roWy4Bl8mewzijejK61MEFmQ0+b9tPjdKhU
l+kNu2OMEcQLeOe3wHf0+H9+cygBH4+x9H35g40pj+aKiWyYoDaijW6+SzQgm4U9
uItUIOCbgonHhAnaQ20BMO9P+yOlRoqjIgGAFS5zxCKqmxEw2Tj3VVz8ouyMVKrr
m2pDna7exfq3KatNbMrelMqJqQ09P8cvsvsI6LC002YIW2YD1p+zrlecaKA7opFJ
9+yVeQdLBPtep79UFF/nrya9HIFHSn1kNu52t3Mb+u7YJDvwD1HVr/JLqLFSaUp8
zIWriF8HJs4xUwfdxHWHIFRRrIJd6Sa1yNgyTM6bPYCid++QVNJ+ytIhPpbU1v0O
C/DuAs6276H8tHpFqKxXGE1lCPew8HCU5gtfuajruk7bPn10uEcq8AFg9Wtnhu3/
rhhU6TXZ25aXmQtmztxyW+n41hS0WhkqAArRWFyp+cKRPOH1S5NdyhgsZKTOmgbU
lUMQy6fomp0GF7HlGQR0YJNEvrZJkic/njJF4DIPac2yflGQ0HweMp4pNF2ANag3
E2CfO2sPOjuOrnggjfvNi9Hlglt0S/1EQWoLu6GfCT0QzcsPdHcRGM39hjCY2Xre
73qTmzqTZkCVZ2pBiFyymGqVxIYVqIuVDjKLx0wqsAfsEk+JPLUP5sAsrIHq79ef
5w5saJ9ni0edG3mZiwu4ioedhtIeuVP6YHbrdup6rdfRgjbDAJSO53O4yvBqIpx0
fPtrd0xntREFJeUuOvpEHZT8tA70+Nl2N8kiX52CZ24fJG2IClAaBakX0ooTpHaB
HYnfws9tz4YMKENOOdVaHxFJMANCbmgLaQpjzTZYjvegak2TGMcrT11IvjJX0rDb
fuhe7A+0mDBoybQyjqtI9N5IpcKTPIohP/4Tboiy1k8nG39mGhnfkJu321+2A0m+
Xf9unyrqBhJTAUX4Nl9fXoaMeuxKsv8pVqY77zgf4xT6MY7k/ZbZ3sDtZ6ImRQPi
Bv5oq8pxKbwR7o1WKoXRLXYhbWMmOpeVAqnH0nbhJUlJNxOfxeF6Lbrz2tTB6AND
6iLzKSleKu3jKgXIzZv3PxH/dh1QDduSW0+M086PnHlxyEqIkfNcJvjrgUORy5zh
viglBUTHn5vCG7AbKLcRdZteuZlGVUsURTbeMoQE0yPfjI8Pld5WTAWsxEpPHGKJ
1VlTHaOKQuKRR92Gw4p5VwnaZhh+IDw+3bSey078pJXlXpxdGZtCQnD3AjGZRUkr
AQ1NTquqoDQBrkDXOWIfTkE7pN2NfSviAHn5Cdw7Wr5UKzPeLhl+DaQ6U2ZhFNcQ
oXrNmEoC5wLO26tIMVcdQDE17T3iDSHuIcq3qW0b8XkzObrsMyoR4oyzMfdvo7VZ
sPPVfJcc0/lVJv4tpwALUEkid9BKkcsSUXHCP/BVzXIE7sJC/ObaFHc2kZ2E0M2f
vBqYBgsGynItuGaYB3Rzh++vqaxRP/xmCXY1PGV3bhOR1BrLZc3WuwxZZAaIOUJF
l7m5R4UjDtm5vgpotqsJ3jIZem1IauWJPkBPJP4HUONUOVkQ49MVcsatCa2FvYy8
C73AYZMnaxRcV3glBdigdwxHmj2oMZMRwC9Xf6pRby5kAVep2MWsmBQkscleWNkr
NElm6u3XVYUxjCffWPbb+ljFOwqBw64bCgYAGca4M0MXQD4/JraZx/HpHeUEGV87
AQVE2jyqOO60ooljFV7cvtw8PoPM/Awen2OpQdaxV4xe9kwVLTBTHS6hzae8nrdC
AC1sJ+fLBgU6BgzGraRicnNdy3hlWD926GtpPxNGImPeSNMcrDW2WxyldgQpNrrM
N0U6mhOj4rybj5GrVFSzD/f88efeqcZ4q4pgfuyGQc12NITgXjNJjkLh4YEyjArl
52Y6hsWz0hvun8G7J3X1h12InWlLC2UD4fWycPZP9vRRk3+0d9GyRiMkAJ5QNkEJ
HN1ZWFl3hyy+FV/LJpnhpoGcGgo7GhSw0v2EmbG3GxVYH7l9qgWO30QSAi4FsdZ0
Pm5r4fpQEISbAsIQu7EhQPNqT++PwBVRXNQvZ4S8h2AYGjv7M91rDYh0/hdxJ+/J
LpjqC9j1oP+o5R+Esf7hR5gE4Z/AcQqDB4672QhQ32JdjAD3yaab3iSZcloo7qFe
QowiWUYhjB0H0NOO+WtmVL0fa84CvR41NaoD1QU0MRfD5ZDTXfuakhHYDHofCcx/
nJeo77BszpI2JnoVU1nZGYY+uvIcpbVfw1wVbR23yQoJOSNO4Zz1jJsRL7vmwtwm
EjHD4S3y6EmRqEoRWO4VvmkG3FfTBkorHq1yWtfYLNhsnHI5HlyKgQIzZ6LuXDN9
yf9230jJ1axcJ0YcyGbjRPoWrwDFmLtR+8AeJSPl5nJZdfgY8gMUm1gid6BAfCHl
QXOVEOUq0Y8SmIXpqy2U3Pt3e0HX8ju4bLRupkXd456W+wCMoJBDmPe+m2OE/Bl+
D9GgFxIFhiWo3NyNc8imSgqNRUvkMg3pNTwhFTekJcOuSVCU9j2PfYTEWkCrqjhR
OP6UI4nT9kxNbsw3sklFwrkJQWHhqRlg9m1nmQIN6OBBcK6Bex8hI7vXeHVBwtDF
zVMZL/GyHEeAEE2yiGARNvqr8Dzp6BMJhXVbVT/wQLm67hBT3PUdb2L9UBHmpgeG
J3N7rN9NtVZh8wbp6Roy/H1M3B6CJDD6ODTsk+kPaz9kD+nrV0lPzvz0dBw0vGEn
B+j6MO7f+PXS2SYrFwh2y00L8Q7xW8oE6ilJiPySSlgo4sJRBnPbvlJGeLYuaOXo
t1Z7lS+0cXBSi+UhAh/nh3K4itEYsb+Et0qK27zXkP6QUS9SZJBmXYOZ8umsoAbc
fs7axh5Pz7R1S/ipzWUsM4+kSrihWHzamx18x29WCJFcuni71pSLGuytjLy17QW4
E+FH4/mS1upHCzlQwGVTzxmTXaeqMrp+KWl+SnLcNPNjeYcuCXK8/fKbUixp5f1h
QAyJlEn6yZr1yYDHggJ1UoUfr5MBjdTohOSeh82Bv8a2l+4UGeBqCaQWvUlu+JJ0
81nQiNn2yM6Bn4lDUKFycbNc4bbCZEFrTB4mqc/kpnr01xLO/uXisb/8RuMioWoc
KrCXj7M4zEiqaTOoISwTlco1Kzj4I6bH8aHkM/ppiMOtK5pIVr3qAIgFvmP6X++6
PqhCDqbIfA/qbQjzICqMnMGB8zsRShBCz3af8emdIiVChYaubntThnO8pPc3DW8w
drMCRT354y+AfxggaXTZldmdARkgorpV75xDDzn8z8ffm+t55bdyRhbJ1jDKWYJX
aQRlDPgmsUkf8/8xsU+ZIrulm3Fc4C798OywJO20zN9ZtzkQnPftshGVeDXp71av
fEl71Jx7k8ErTHdtxalDFijy5fBoOVEsmxlJYYKM2FujH3BRIcbdy4QUO9tM3sRT
/b4930021YUCzQCN+gNLSU0QwDCFOtjX+UCPhjDBf3N9WV3R3UGjf52kyorDM+dN
lNp5brPo8LCtBfxK1isXID3WDGlXNOqMJBfkvAhL1ESZY3gkezlqDYpe4Pobk2eM
LHU7CtRn9eCxUTvAUq+xLewHrz8eloWP1CkQEPBvBHLo+5i5oLBRb6sonPw2DKPR
WhLksk5UOu7W2p1eyTyaQXqDzfOa2hJjtvajzbq3lsw2+/bj1F1GXNgW5fuOWjOU
hy4iZTZ+mMlfn1pltSYVUWGYr5xhe5rUEp3YC58jFABlpDWKb7IoUnhz60KAsjsw
gDaBAP+dMp115vVtg8fCIsxsP7QSXGB5x+lIG3iq/WyXcDLH/f0QAy2YNDZwfwi3
vMvdLnKeN6Psy9d8CD1g4gsiRTQAtww30Aq1hlmBh0AerKRH9+TMNag+/gvjN5CF
N0G7zHKb2tZZMsXeKUnyRWoK97Pw7SMa4pKjsrlQK8qaoFOAAhaa7F2CzHwD7DjV
Gsbl0LZvyPFiJkh9V/IrjrBjoX+V+MSfETN+ZcKQJx8NV4J70oPkNF+r7Mg8VxTs
JiwMPHEW2QDjIMxnF3ggyAvOPzT3JiPf9uSaIQd3M7SDr7UFDvbqWbKhNAVX0WSp
2Dmpbg2G6sg4ofi1AuOD4fSQna9bJTMYeeD60YQx2N9sNyMsQosoVWEgkKCQfa4r
Nkj6Y8RVe++ZpxJ8iEKOezKjIdUSr8nv/s++/+bHPD29EiX3X6iSdQnJoR68ljy5
tyxiS7CvRKATz7foCNkElAzATdNi6HxFPLdJH/a5S2CoYSEpEe9kfSTMDnkYC4PY
GOjHwlQd6yY3755aQ5rBVL3c0bZMfxJiRkKKdALa37QXLFHfSz5x30wShtb+j3x8
u4DP0cRIl3ctU4xyNJqB3udWCRPaUMfHAQPYoF45HscBpH1qcAU7K9t33VsvNO1C
rltCONcQAEwgqPt/8umCTjH4oRSQxA5aIeq2NXFxevTXmQPLF4Np0owQIVm7sRYu
Y8jdEQ8pJcRiXjk14aF09ze0ffDC5weEzwxAkROtpG53vkorWl5bq9oI5xA0Fv08
yb1YngE/4pl2EIeuK4yfsMSMh20WHr2yxSgvssSY9c6PDY8JnCfLOSWXqvAsJ+6x
rE1rOwDLP3RcF2xfBsZ1XuRAQFl+7p9bvz/in3TbJJAZUrDgjswYWW/5C28Le5KL
6RD/u0Rqev2uKLRaDelzvK7QSuhYDxhZjVmsPJ9N35Wg7q7pfDK23q+c2rG2scBt
8y4xuvX72e9tZTLXuuQIXA2HV5hFFJXSNyGyvhtKO/XJ7XZ/XK4vLeyb7xXFXMaJ
BIw1cHaP6ZAkQes/H/OV36dRVvXVbMRrBU3f6o1u20ncILVvgOhx5XWS2rl8s96v
Q9jYjq+JFIZ2Que0Fngyeth20T8kLAsQLlLQ/9lEoBqQTHmeXQ7HZdPGr26yICmU
lzFXnJF+8WxylV2JnX7T4f4/mBvlHm3LPrpeW/zmb6trX/9+wlJe4V692kdG13TN
KvZT/QEDiCXAWOvI7v/M1CvoCfe9lnzj5h7DHflrq5FJr6HRjNjdUrev/MP35sJ2
bpA2cgoNEZWMJAM+G5CmaP75lej+jE/SlyslqvcXMgzWXmgsNldoEQtsaTBycHcy
mpU8yRrtW7o2EFLpDbNW8RJ/zKN9eOfOugw5Plmc0HIA58/WMari5qR3FFxzIgxF
zl86nGm7i0KSoJt9/190dPX8wOOT1n/GuLs/Ptb1lhBSLsJmlq2mj1U8FIBpLD06
EX9OFwYSg1hd57LjNwJ/k9QITGYz7ACLG4OVPPZLsq+5oowjmbPzRtpHdG8LRym2
Q4kWKLg9YVOAI0PnnoSARLvaWUJQlcF2idnMkk3NFzH334cu9aIdMqK2TyaifbjY
/viF7yTVgWObjzAUyZ34Tnj/ZG1WkzOErnpOHQIWQIvaZY9YRwbQWwDHPQHDCbTm
u31MWskAJE5hufTTi0VVXCL9XOoI7BVIOCZwfVttsIZ/WeKbB4GwVgAEURPjkZdG
u2fwNUEUodJBvdTcF63PI/2MizJWV2hWvAyYEiHlygBiiBVn49gUb+8/p9jqqrkB
M60n7sC26seU0VBCXq8ShhRBxxQV0Sv9VBqgNt4mDWP8sqeDw2aoPY9qDyxx010c
ZgDd2J8tXQVSs9cyv8RMVEa6g256Wl79s1N1WLRTJfieV9sZ0oVxtNoxBoYWhhLp
rKgFechCIhOtVt5gaKscO6r0c3skxnwlUJpPeq7MVzeDEZ6+271Yxkj3xljOWEIA
TKvVWdLbUssYzLfk8dxHP/MEsv5V2YhXDZKg+MlM9vUCMQxe8oO2+CChBjQOE9pd
7rdUKN5Quzm5d7/eLJET2WhLAIHgjHfv4Wnr6dw9rKgTSAycTndUjEEXXIzbea4E
Gd1dx3FOy8jD2pDplZBzqKJmuhRBsefL0doTSKWDAL4jfOBcVAyTnCP62+YVwBc9
S2e4Dns7ZoLzgN6ueafvbV3JeqDwAIq/vOusr0FHt4IUK2d6Qs6ztUP4BBhDp2J1
iEPas3ciZC/k6LIux//RoMNI8meSj6v/i37KUB9qC118x2dPWiQGKxRqP6pDZ1jv
IxCAOWHXifKhQr+6n7CvL7Y6qR9coUvxA5sH0IefAC8O7TRU6PMnZdL+ewiFUQL1
W7vmbdA0oNAAKU96YavEb81evZLKCiPFdW561I3W3nx9OjIw95vV5gvgQgVyXP74
MdM4OEZs4yWYtexnQhuJmN6IXqNPGJUZKDNkD5r1UVY2emrNPbXP3iF0cH4vGtF2
Yn5HX6omeqMPvWr3Sd7JoJ99u+oKSIyRkIiOepP9VIJ9d6nZLehQ8VUX8ue/LuMq
+ebtNaOouP+eJS5apNHpIQ8ePQjiKytr/3Z8j0WjO0oW1OBJl0hPSYuNBOdap+iq
znWiU7DwbkqV5Bw/iDIrFy58PZ/XOBwYVoSFWsjunbeYwksnxMMcRwg8LBp54Z+p
f+aPdPfFqjBVfByF+Cvr8iPe/4DzfG2/dug6rq4B91uiAhQkiEk/XiLwFwDCThN0
bHapEbyjLi6u/6MtXmmMpjEo8PbptUZEAi5o7ab1Bjk2W3itHEfR4ARJw4f+p/gm
3+zMymJyLgHWKOBDQWHRUrJAYclkytNwqAIfNC8CoYXEHnQxX5UaxJ34x9uyA+fW
S8vk7Xrx+0TJzlW25+/+Etgp5Kc6elwOcX5FquiylxE6UKJ/WyYzsVFC0O0SAVBf
0NvUquAbDKfkdcobmLR9qq2IizPZpkhxMz9D68e8P7RetDwhPPerTbnxNTSSCIAz
9WVLNal5jU1oXLDJf7Xr7b+c8p5HdfrRuQLxOsi4lvWKJEgpE+mSAt+469CRXe78
UR8ErU0VWC7Hj3ryDcRfGdyPAZG0d0auLayeM5HPxNGXUHST1rYbDK7/T4wSZTIT
EhZ03Iox0Z4o6CnFjIMroVxGo9AQWWYYtWiz1tBbjEE7lzPV23tdWDbzR19i73Ee
PcE5BAazIhSp2VRc3gPBwj6Owqsaljf/jSznZ1rFHtXtRMARvcq/kakVGS3MPxre
JXU/pVVWLdlzrLEYnodkWciuuioWGN/c/kA5lFOVzexFYsnMGm8jUTZXlgtqK+uQ
cqERdo3W/bFDF5lEiyAmyQcCerzq/P2WIymYsS5icyci1M5P7CwmBXd+krWirjnp
i/v/TvtnlA1VoPLjJwkALKusoVfLFsUP1cUIjUbFt2ZIK58AoUuFhM4Em//ieyAJ
PwIYPGLZWWNuCnK7Y3kxNOoLOl/LLFaS3rpd3oSlWa02BEvEhofqrNgkIyWJqCVQ
/+bgpAuQHFrBGtSrCo2WAvOk+FesjSvAV2c5VvbzELx6QNu6KYI2AUFjZ0ED80e5
N4k9v1SEwgoy3dTqjEiNS+4Enmq1OlWuMlNHUfuIhTkHxYFe27blyFs2dKlEGABF
IeRwKfBb8I50LoyJWJsSrxP9jkJ5Hx/JZpT5yPMi8rMHVrOrGOr1AMIakDUor/MC
pgXc7Vk5jyGeqH5W1MzhK3H+gPiT48AzuTtTnrBsDcgWxvafJRj51XWMACnUAlBZ
k5O+x0V9VX7kBfR99T0L3yAR1CVDTtmyXW6xFhOMuhxHuMqiov+425yBAiaey3Lt
MjQ2sCltVIuaaYqtMpCr/yr4tZsKHd/pvpxiIEMVbpXK6bPqX6pVl601EokPCfxl
ohLutYpz9H5kZROTdABooq/e81YRYUBFwBl63NrfOYQD39dn7WPEUw5OaW50ALmI
B5egUfM9Pbjgm+ksArQqsWn85ntu4Fc36HGnaMZtejdf804+BMjNR5UvxatHJzyV
6wUnwEUFmwEK76CD2dLBCFKYEEYvF0yIkYeBxNHodvAmBrT31vjTkGoYlra9tF/p
uTWEASf/qNwjITmqcimEUsJMpzkDZXHMD4YrawS5PajV9p2YgKQHsaqhevZJWQUt
ZTN51UNjGr5TxoXi930gYJHkFYp+v5+l68QvssyjKFixBqG953JgRAJ0ozpM8rQQ
1cghTVhRfUNxQdY/DQKSfglcfnYH/18JgherWpaOWNUVT+xPV8/iWWUWI7s2gHAA
Q0r2H46WzHqtAA8U2fUU4YMWBEHbrLtzZ76Oq+9lVSZ4uTrx35vu4VUQixbkNekF
8gk7OZtNgFs/dlDsYFDHcvO5/v43oDJ8garqUMXfzejdtESfjGtQ3Zn8kPmlofsu
FzHwZo6FGnTO3xIl0N8LNMFV+pH70QdsEvshGqUzUuCoW1qoVIMq5tu/P4ipTRKp
VAvHzhlYAe6ivGNNv0rmr4rvrVw5mrt6e6jC/9cJ8NcvSiLtbMxnTstmm6AqwQJY
6+fYRw65NS4Mhe24eLDxm8eYRCc1yjKS330PMJwMIHbliBTTKcj2Lv47gS+zfeO1
7+5HPCgmv6nDNbFd4vhO3XonM5DnIEdNITKFNEhQKrFgwrpJs16kT9bCG23LQsVH
jACJ5jnazRGDH56MLpUlNq/jxL1M29eY20ZBl7HLRACh72TYvsYjfnPF8fxzjO0H
95zvNIrHKmsAjaD6NJLfFnyKXtD13FhJTcKfIl7EtRyvvnuaU0NotcYSoSXWDnOP
pNROyvjWoJxmvWwZI5q5YQ/IjuutveaWL9m53PgtTyq/s5X4kpdLvsY2jRuWu1OU
D9R6+UaXtMKkvvyI1PjsD9+ltLe2ebBrhH+NgICk680RcE9orTrAWRbaVrunmPJq
DJrWEpFwsmL9naEOmge/6AQ8FojdkB1WArkhjYzqKWyzAjtpQZ+0mwtmCKQxEdit
c9FDZlvbhaxCoslNBKewhnTv9f2CzXLLE2qRHvnFTB6L5Xlq0WUjcGjL+A0245B1
cQ9ffnWO43ANnnkYyOnnHd0qD9TncjF5cQ+WIHjxtBUdoOpWHGXnnxrZ3p45c8cJ
dm+jXyM4pLIJuLznxzD4jW91hXklwlx1rQ6SP6V0dvWgqJj5Hi47lTJGCuJVXjQe
zlP5p9i7wToY4LHTvO02vdexzHWzyTPbKxGWB9zhHdvQTt1Z+deR0ihoUgd4uHPq
u2S3QHZI1muYCZcwm9ZfEW8pHcLLaiqvgupT9fPFAIfdvzYq3L8ZXk2NCpCF5OZi
AAmZDkpKvoLWQ/CYp6fkx/E2DPPdTTgAxGj9mRa5Cf7C8Sm69d9mBRgK3ZrSIhWw
vvRyo5SfFf1OI6RP3ozRmyE0vKdsoETtcFwKojeXKTDYBssMeV4QQ300d5aRoNoT
CI3lebbzBc3eOUUyWlnQeSmQcwaDmncyD6neTxPpybpqF/oN1YeJlRbF77wJklYz
qclbBynEG7hCAPreZdbUKjlr5CqfhxTaN/oHgKq3kaT+TRzKcUxNQO+gRHlud4JL
NeD1tSKrG0BYgHC9L+n09+0p7W3zviDDS99ADQoeGnKRk+IzJ9iVEp/Wqa3HgJKj
h9K5g9pyj3uxzyBDKWKdO4YlSCTjBIpCI0KzCja/O2lIxh7agPx2varm4FIVuvja
ywbqs/vse5IP+8xJEPuSVW1AqhX4v4I6YhsbuaGLO8LZVUtWAuIXgEqsHZNi5Qlh
4kYzAE45OnLMpRjRTrr7+uUlfCp/yHnBQBXG1rxqpX0njnB2EvnaL2jPK9DTE1+9
2yQw9+HNHjBYmzQZglhrbV9GH0Js8cgyc/5xZwHLg73HUMTFw5j7Wo1FNrvdbL/W
NVENAtBiZPH2ny025tiMVaoDFdw7CX/ockg4bzxtbFAzCy3o0Jcv+RBx0Zsn2lUn
6WuDwXhpWknxPywqX8TQ3myEhyMMDtWU/0lukkfqzF8UPdetcUieSpeNbHgaZtE1
vaLZGLPlTYjsI324kiK7b8FzD1soD0BQaulgP3S+gjSXShr10lz/VbBOnGckyNvh
oAyO/JjUZYtjsFj1pJG+Bcj1OWFL88Jx/3H/vX71rHO1ASyl8rxD+7qKQQeX/l8x
pvCv5cnvKOc1to4+GUxDdaSKQuNMWHjLZknT+VtotoOQ316kMITmjF7a42dtKYOu
mQhZz6QDZxjRCXm9dDYMtqTNuh4rxk39U/cN4PotJw8dro+c0mHBTqUaBqLmcqEN
RCdBv8mD/MJ0Rf8eaMWa7SHPEXbyh5+2PCyu6Q7LLR5BJ2P/ACVxKojI1z5IilJQ
fgDWNOpszEmT9rWMWmLubKa+LTu7DjUwMVdwAWX9lCzEGPkajVp3NuDZaxKXFxCx
g2OKsnfS64IYgdqgL0fUEyEXrpj8tyjMNyI/DPchp4B/iK43Rx5meNjHgs1aUEME
k06hSJ5Y+1M70qg5TnaTd9invjrO/XsiZaysxwKAlVNel+GFYAO3KDlHiPelI2cL
iazrnKt6PRLqY8/CjchrFHCnHTJ5pKGfZgllku7Q6hJbkieeAIZAQlDOcSSqslCi
/T/LDagp7vF3pgY4Yz+duWnwpRn9rknqgb9sIA+4Y5TdyIzpvOiOom9em2ZNi4vD
N7UrsUjL14w0VNASbP3odRDkZGaiewlZ8QcnBa9R6eEPGk9j9f4pxCrvoLvSMkmP
0/xjZEa3ewPiC1KhQ5KHziAu8Hr1FeanjFgkgAlqiDhWD0TturvkuLhffHxfX9aN
9the8Jadm/pRYCVJ5wtw6qcTmDgX3bjeyNZMNHNZtUnDhklZR1V45HNyyS6yhGyK
VwKokS7Ewe2hHAhQzAf5xkK++qlB9uIuF9eawBkB2PcdziRU1i16+dJn+z/uPgBJ
ce72zWuBTxudE3nwOflCSbOM0EQiA0BVw7/svA17X7HNr76r6TUZUPU1UdMaNjPS
qcDU9YzRO5wdrP3wd7z4jjMn1xy0iIsgIUQPu0Tz9Y791asBIv4e1oFbV+Qz6mrA
rw4VTqEZjy5JfjUtGdyX2s/juBx0uWOd3KnohTu2Wfdve3MAmVnWozla/R2sz9Q/
Oq0g04hZO8zCmdPMdoNvUU/BtpSHJlbARH9s9tM4x/d/LnKdBihoDaAueWlfpHXW
lEFwGtzT4iN/bjrD5QSmJGPIucFCPV3C/O2E2U/ENAIXMof8rq/rXHNghTHMy8HB
xEdeK+EuiFoCNps2fnDbzyOTzBs0AcKnHa+inO+zvY+gLLMhuU/tqaSNvX1vjb4G
q7rRmgbRslONfGHwvGXDD5VLqZx+vJu81v/tT3ZLN4aZ0DU2me1lasp94LmOr+vz
vsy+DEZDA1CnmFgZEFVdHXqHYlw7/0CCVUnzY2TR9tn/TGcivJQKuhLDV9PR2DKC
2djqJCj4vwAgK5ya+EETkU6RhJZnGmaOpI8JtbbKAI6Y/rgUxd3R/fKlLmP204jm
cztshIgIpT76BUQPHaDwUvDw9Y2syXKKrjMOm3XK8XVT0BpikuFCQkKVuNJzmtZU
AVhPw1nXAy5C3CW41lPewKXsBuXgpJeG0jpnyHPZQxEXTKtwrbN4H84gtXZgwTwN
4vgr4KyEGSOIT/hX/U1Mn2sOT0MkJUtWUOmqRySu/DUjgwrb9T1RCq5Gd19/XbPJ
a4bsMnBSA969pEt0YJ8IJKmumM1M76rvIDIAq6Fhrd/EUzWlmk36qz9ip+xIEYgV
+PpElTt0raqBWw2VCAUGnt1B06y2vQdBDDZK1aCMsCaVUd1RAnNZUscSNaRH5vF+
A4KRf1VF9RWFAaD226SE8KaSYQ8lnf0upiAvJ04XoKy/1s0e9GIMXEI458Gi09Zf
ghANoY5DzSVAiwr83KyfahBZ8FCHOX2r50GZDzmhn16NwGBaLzMLJ2U77U+XcnbT
zO2ZnBLwOF/l2uhHCmW9rwDLZVISMee6RXhBzHgDYR4GH5g6PoZhK66ztE3iHoFo
vuG+F1zZvJTUic3ynr6RDfhV7B3r24STmb52sY2I2tRJvup47cJoxv71FP1VWqBq
2dXuZQxq0ZjswysNjDsbFRvfe1DttktfnxKiOn+f0bcCy2ADxL0jK6MAylEMeOYG
mC63cYr+qtNbh1kyQ9NVzx4BLvOfD2WrLRMJIvNgkDNXpMX939ypT23ffCX/KiyV
xe1kGfDeB8cDFHrVzoLYjU12FKTpVpG6RtVKY3haFvl4pdf7xfxB4+9EfMsfNCTm
FNypquKDe6zYqQruUnoeaNssuEzNdlu4RPscoSwX80o9ARQLdKxF65YHR3KnqOFt
PHLVI4qjnzGNgwXg9nx8aTvHcHnUbwKMoXQKvV9oQIjk8BBxNjNEDcZa46G/7zmE
T19DPdqKiorJprKWoZ5LQGqfyKfuf4MYK1nBNEvlqwhWTlUyfa0UOmtN3VlhD+TJ
tUsTacprHFzC0EQ5mgqkGg1w86C9yR2acWe5xWC35EhFyk6RmDDdPUsVXcIipogQ
/oiCy1mkncV49oj2+GBM84qYkznAQpeC5+eQ4lBfSAWbim0+Uc/nSw1kCB3E1efL
JBg30JqggjcptsWn65KPXaKRHCBwxCgTi8c0sP39trtwQ3mUi2RGAAQcl9luHCdg
Or0YALH6ggeiyPW+wpmf+tnHN8XV7kLo+KM5AWZ/+E0JcsT4yg8LEhLeZ4j5cXy9
FQ2uaUZ7eGMTJhSKMVXC7Z/xH9XQfvDiNA9J6Dso3Y1Ow0gZOrVgU5ugGYmjDaMH
u8Hcceqa1w3LuPFXQoR8tBva5rJHQYep8x8veGf6kF9XQxYOuw/9rKjVikJXXiOD
dwnDKvLpRipcrY8eMyMgyUuIiNYssxkDa5kdee5Z5gWPepOD2tYcTHGDT3UAN9Dk
mMoMDva0Jvc9UyWYwMmY8cOk9J9O4Zk+JHkFHM9q0JmqxLAzKVB0h67MPg/D1VsS
dfD0rQrAw99X5eu44Ju5h7Ff59PIhRyHHMilBrbe8uO0PiseMuImErqiSq1+KQq4
ZAw71DGiDV/M46rmXQx9Yg2lircRSQ+Eb3VWWKlO7b50PtytDLKqhxb7Y3cT04te
GInbVdqFd2OKwWLYkH0so0Ym3wHBvahEKvMRh9rZepL1Saoxk4TEgbCkeZyz3I38
FRWNV73/X6ul3DsQojORwzaO8hmMnSbi2dhwI/YcRaVGHCa2yfq6/38olb3bIn63
y7JlKhFGBAE8y5FuxGbSvL+kWtfJJvcqR5CXwJmqC9pAGyWJDKG0QAOlvYOVSomU
Ss06F8t3PKoVsKA3SwoG90cEMmmL781tm3v4x7/MVK8P5OEFeM+IYZoUmK/31nw2
zaOSPTaIbK/Top9M0voXC1RIbCJyub7Xi/PZO41NzFxr5uaJU+KDVJFHfeLGUMSA
6ojJB6qvVAVOlkDYkuWVgiR9hh7Rn+xnVRlPMWUwUyb6Omi/RD9Rd2oMT4vd5G/f
ouWwNEP4v6BU+SZ1e9udIVXcBWh1ZSEBxs+BP4kDZq7/S7JSRc8S8XHabHXdRA+Y
93EFBCo+g40z+7TpSEY+K074A9wwGCEGhKN3nT/OAv7oG5+53uIbRfCQIPPfIi+D
at/ZZHPomeoYam68BzLbOFHfLze+hYflTrOLR6GmRp750dR4AGha4GjCklr8gnc1
5Z4c6qGoK+KKF59OU0y/o+v0/njpnnHsvCueTQ4iT8t9hC7YFB+oY07Fd3yv5+fK
WzsKSWBNK21kJn6+Mu0Z1YDPlQGlwDBwzbLxNGYwD8puezdNXacmnq7XC2xwrgHy
dwbxTVLpDj/YLNh7Qe5MdMPY8+YdyCZGulDnUJUEmZ2FoWX2zENJ/pHa0AhcVtAD
P4SoLmdQmk3Cn1nd/CD+z8tUkfo5cL/JpzwHJ4fxm3u+7klOYTmHa+GXlrFF38QF
7pjbisKc0rRoYlKunuEWPet3FLzvuOZxm5ZdSfj1c3GiNjJmYBUXOIazeeE+k3xj
fxK6aP+WUxN53oxPHTauxjTDKbXGOqrce8dnbUENoxrSZfCcoMlTvmG26B0JcLEI
nml27yhIuF0g93eXxJmaLsywWtGVYdkNTiUD/yxjAKV0VKi2A+Azfg9FfqFo8zhw
HqeLhjWKz0DRHdQCdlhuFgGAFb+1IMRalcm6d2kQJAVJrVqbseypxFa/KK6kwkyx
9msZpXPMwT0SooY7RMPFNDxsDDI4C50PciGwslv3RPmEKg8s0dM+PTo/Un88YiYo
zUdJvIEWWy/kpfeiwRtsd1dfAxm35MxNEIytYG0LVlhAXdNfVBhaGAf5q4bedVhS
+eM2aMPdfQsqjz8cWr1D/7aK1uFLgKqF5/nwb2BoJTB+Pe1PlGFqQaUnKtluwwkn
MZUHmJ0ovE7nxfwJp5zI1mQYHOpHyta25w5rG6dtsGH48J76DiK1uHPsSXLo49GC
u0lqIfyfRDGqS6hicg423UCZa/qzZtTyYDA/jHGIpnO8PXPh8zNRtoh/gBGwE/3M
bJBVGY7gJ+6/G1gnH/tp+vPiwjr6qA1HEsKJlMF1OHpkhjoyGOqggiibNUwCRfGf
0nyeg7Np5f7LN8bfkhVLIZxB5t64H3mYusWfrQJfnBfmzN5csZThBNisopuNNyvx
oKTdHvJWz6x3ODMrXEhc5hedZimPg1l8/LkU+EIMSOWxNHoxx+Sva5iSAjNOhX6o
089Q7KcuDGPEZOz87y4sI0Fe+qWMc3U9wxFZ5ZEl8DBLuaa0iLuwZ5fd1WZFi+8B
FBLjJsKOMYzvzjjkFzoyPlrEJPJt9hvFmUoCuGOKDGh4Tz+r1Ht6DKauywerCMHF
j82ia1l0Vsjwgv52klSGf0cBkphYaMnNaRZ1jq51o/1YnkHHX4DFIzJugZVYl92A
deHOCOifDAlf7ZaUVgVSEtjVwaYl9xusJ2w+CiyFbASewGbcYvjRHUw/zRK8+gKg
Wf+gKuuiS93t0v0UacJI6CpyjpJkTVjzmtvAeqtBsPO4VbHdAm5SWX2reIU20Z4M
8hyNpXb/u1ZFWTUqknzbHOm35sGByVnUBmNndevHjAzCoEMb+h9AogOQZdqfoc9X
hbLt7IXjSgFyiruGdSFQVChgqkgwVRhaeE14BKowg9lTVHuuhlgX+nej4X+Y0orO
U2y+3r9PdIojXSFfPIFQzZnxIfRIS72/w4aUXDESop5H6DjamMHPLYTUMJGxAsLW
iJP7zW+9Ih++Olk3rNBmA5z5LGYJg+SBb/ii9tZDAKiIIanmNN7hUZBIkAvpno8F
9r8/P4qNSqzlJyhHWqblMVpcDH1uY8r9LIwAgii7q1XTKSMsfMYBnQjv1BUYQtYq
gyRt6ZRdcyiZjVWUO/Xenq+kU3YCDQR0vLqStr2q+oiaddj7kkBgo+rNK5bvjI5f
wvaf/j36dj2Z29G0rV6KOyDxG4WJ4XmFRSehie40yJddj4VSbyGXaqVPJNiqE5k1
5xWsK6LU5nqCJs195BKcTxEFg6K4zpbRFsL+huKdtxL/ZWPvdQP+IqgygGAuMTtf
QgNuS1Nm26Y2FL0U4o9uIvOqPN6KlFa+90Xy7x4NtZrMcFcoWpzoKCfvk5kNljWn
1wnzkjxYtEUkpPQd7sWjOOPEM8f4C/Q39np6N8GMByTO9d/Y4uLPgUAZArZsUQIS
/ZhBIv+0qVQpOBtsqKvU945HLgLm4vD+quMiVOsPp8MiaLWbR35LG4gL+01y8x/d
judLS3xd8hAJspGLm5MsdqcjHYDNWHGDQk81O00IhUnSL7SEqdKSMpVvKr0593MJ
mk6EVJ1lSL0j+QG0Vk1k3VPQjqal+fqXoEG7Oa13kEkMwq9s+gbK8kNmMAD6Uf2e
tQN8nhV6woBu9GoFz+WiSEEBC+ORBewr7u561n08/qBTb0TTYjtaMyx+sYFl3bcC
ccps0JWlwQFtGaHIUoyE+slhFP9QhbRZesKDvuR3KVDuNjDjytGvAqJAjGYsSSxY
8as120/uIkyOya6hW22apAWoP7+f7zP5scAkg9xhyNOai2Q960RVJjO2/43YQIRC
xSEFGlrkR3EKvEkOwYwJDLX/1HtleBoP+4oF8Em2efk988edHM/Hymv4ouAsvzwU
0nR8ASpxhyY//wZMfgKZbylZnpwgDhkDeiVTAhCmhTKv5fap+H2qJrznSCNxNCti
KAnXP1nn4xJXahS8BJy6B4+dDRziFCgOzV55LrjG0b9yQVHBsOzTVDzk6GsjzOm7
aMVTfa3pphuMmI5EnXcdHdnVuNY6YNBvzakSsu0db9sJ9RQGdww3nkEO5lsoN+VC
k7wf5ewXeX5Z1HcQ1T6hFHu7sjQZ2igVF5L2gQSpgVAsJm1/Tg94cPC3lFWJ5i3E
kXrMaXA4oVFcLiesiJUk9rBn0VVOhUS6BH3ugeDGUJOvuW6vW97Gob2+W0P75WSE
ukh1hg2h0GfVx7qMitFa0TgSjA+7257VwtamOuPCGdwPuxoglX2M0cgjLWlhFFGC
jmRWqIVTSasji9yiqeABdTH3p5fUahSKI6EWSVno/PlDe7i23LDDKx8rmb9M3g8h
WdtlLHBuBbp9KffevQRsnwMJ9U7bFscr1fLySRne2U1JzeGXvEkjH5BpgFyO5QUH
fflDlWFVOeMkWD2JnDK8+KW4M/E3XTX2Hy+hsuT3ZDvRcllhH7ZEUGcKaGB6D9MV
3DQmZdYdPEe6KTO/c6rCrK5W4+gIz2VJAr2GsRbmRVQMPqYvZlKbvL5DWWt2qHhR
YRXVD0d9gQe5vz8PzZMeBQ6VwSIkPMz9XJvHSqd+qoqp9fTtAW+PFCM6Zh27KIDI
mTYc1YNVm+oheFYMhqLdgil2GXpBZRbkwtDj6sABmEPCOyPuORiHTtg6OKEPZ8mR
hcGILq5mNWBJ4hTQa4SKHumwIkk3a1z51JE5pmidw8kAoIS2klBme7b0BVqKwvP1
ADg1H7hH+lpZZr8QUpYiQRnVLnT5Exh793Zh2uPkA47XnAPpCfIhL4mC5HE/+HTc
wkY0xky9dJx7MOLWeIFCJiOwoMptUohZZQLDmw2ZIaMgFI1FUsViypbXY9OV7znS
ICPHYLsjLUSKilYKS7U0cU7eoZsfykvV//I8uWB5lN50EjNPkfvNlnz/lHKQcQrZ
Dajhy5qrWxu6KW7eNOz2+5B8fD9soFgMMRG6QyHC0l0SseghJmRNDy0ufUD7VP2g
pKUcIop+8bxlcxjx8hp/51YVsSGjppcoq1OL+Er8lraZbXXOPVlZ9LkNzu3wKpRv
GP9LCtnwkkwy8AgMYe7jX/VMcmx3suvz5r9d359kJ9drtTnc+9uwWI/LI9j8PC5U
OqyWLDsHXYxSPTrSbuwOfg3bLXwqPEYhI1CGH85SjU+bZkRBBSahubna694DQn4d
tuNoSnkWQ6kkdqeC9MhxmrNJiL5lew8eb1a4QrXELHlNKyckOXn3DFDTLZbYf0fV
4Omvag9TQq201usbdPQpl94Euxo6Kp6gcOELrk0EEsVsvf+H8JB5shOJU80sfcSP
E+RFi1k3AWyDL1EBg5gMvC0JsjfR+OzIW6iVdWeuno88uJXR/ZYQg0zqa0F7N457
CF8rlWnwtf2IMK/fimpOjgU6owIipqkIX5nD4hYaNJJL65dfRru9RHvvYJL+z0Dj
cznKgL5uF7Yuj5ED22DeEEpdzi63VI5ATK0nRH4AlUzUk96BSBTUYhOYzMnGhulw
WqtvJmg/+ZohyCcKNRmkguK1BlRNKGn8icbkbzRO/wiM7B2GADts1jDhZnT2nd6q
pgJ2+tXwEA1LosJYIskUFSi5xwMdTtCSkAIc8wyviCo8zgW0gdTLOJgVwBuxxn52
K1bqKbL3glWT0b0UDBAfBEZtP4SIZ8JghSs1Md9yXmbLlyGrr+NmDv7thN6kepg4
dEmjYi+npQFN07WTe9yjgdX1rTwOgLr88gITMAMR56rz1orgzRhGYYELGoRKXqKl
c/6BK4STulK37+ag/bWHw85T03Ocn+h7NAcpd5dVKcPijQvnRlS22W76WfRPusv0
OWuOCsHHN3xJWay2x5ui0nAmySl4AvotdqBg8VwmR7cHuOdwBvh41D46VSvF13/O
EH1WmMYejsdFnQVRA/UnN54IW2EBTDzYn3aWSITYwIBwhINJ+3hHK13qoATfZWjy
pO8zoEUFLwoif30+jdEzHlqBZK23Db8a3PpDUOInvP4sCXjlxTU3+D+WH+kNOi4g
Hw1RCkW0wFGQs2/QjgZJSyyKcjCF7jQ1uHYQju6cJHPeB/mgL368rBEyaOdodzes
rSr8l1ZHM7Q+OpWCT+kOIjbUglEVrlxfWfhnVFgE3+pMdw90oQ6Sh5/9oGCi9h81
fmbUU5DDQX/DRFDAoACB9teFZ7YXyowsNERwv2MPj1Vp2CfdbwQ+Tkqy+XNTw735
qesWWmmjBsQrvN67ySFyaCCWLPUciWbDLGjyLQDKp8VfBKG7HRgL7UonEJcfJkko
R0CTK/tAA4xJVG6YZ/n2+VhaGQfmES+wIwHhfDAtPMCT5Jt3DuOu9EdrPGGJbFmY
S6rd6+y7cLves17O8HxBBCQzHdLCTh0bfC3V0RTMKCMNjLlsdwYCMm/KTpIjp97T
ME9H6dhJXDNYUOASOTvBy4bqzsH+uyVFvXzpYx3WBFCIlWITTYCqRtt2J5dvwcLv
ZB8WiKGPCpCG7TdPlFv9vNcwIphFMKORAzCg6OGD24ZvWQJQZ2t0qhcp9wW0XzBe
n3n+ujqSeVg4zfldPRAdw7pJE2Ders8iAdcQkc3yFPsWXpQVDPWeNkNGBxzOlTR5
dPUO+FbMndkp2yd9/WapfWZ72naTjIzbBpgSOlwRjx7XaLgem9IIuPLQmXCFP/Iv
BnGIXGvOM86eoxZWYTBCUzrlSi1friT8wXZ3in52tvrqv7SOLozom8hmEsGCu5R1
o/ELQybjMHgQlqAHKvnDqYQtjMkK0Aw6xctM6nsvhxXmkp5DqPRDqtLyVy2XqIpD
U4hu5pHN5rh3EtbdisvCi3Lu6kovJoK4SQbW42IlvD44RIVN+srfuqCDvNxt2jzw
pzM3G5m2ODhQ/fkZSd2W1MHGq9nBUMNP7lsHFMNSSOZjnt6GQJhY67nwne2bdYPc
m7EwFg2EdaRi89FM1OmbJVvI5KSdp8AHwYkLilEU8ytpfCe6i3P+1ETxkGqi8kqQ
XKBzGq5YVBZLAKVOjf4p22cgL+574pjRogNBM81SV98vk8ZbiQp/FDOW6MQoRbRh
U+KheOaShkeGKiavTpAVROoRSTP9GqBYKTy6Rf3o7sE1fOqXM2Mo/S/dJnR1s6CO
H4nhtatbbkEkXIGOuVI6zy/WpAwbb0JIdU/vgCSNkuAsdIYr401Aj2kYqoBMtbC0
v8/djBlgN6Zxk+12b9sgP9aJD7vzv2wRTrMBHghP0XayW7XRl3XLqVUWNxQLvej/
ez0Oa02hbh9YaazJ5ejQ5sbVLpBsTkgNcO96/bnT82FDVNsIVbrGzApBNmGss6ZA
JjUdHdzNJZFLN0r9uS8JkR6BhwCwilBFfZ4zsEmJ+4Fmy4SpnfC569IFOzZHrAY3
f2zTtBxdUH5T4gGEAy8Q3Zvpw7/Tpr4ZjQolkTZ2LADWjr/It0Dk5+wQrdiiU6/T
WaVZd9Cpbv964+lY9T8l/3CF4rnkMPkBburrOcLiiq5951wjPngw6r5UI2Vo0BaV
mwKLfJ7NmztTnOFVqoAp5g9nReBnFdtPHveHPJ5Wh6VpfgMyyuV7FwjKWbqYQc6h
+8GIzrxrD2Ew319/z08Da6Bt16Lk+tUC0ev6Ok6HAGR4c6Q+QGSGZgpGSGmI8sC8
1KUwV+1Co+IkBOC0mYbfVxPWSGZFOL+jvXE5YVK5HTGU4uufagCKbSWzuCqc1W4P
m6m4PUiqC4hHL7ZBx8mbJybPJK/s6H/zE8Oxrr9B1DUtFUhbnSQRrYqwy9mki8Qs
LOtf8nG0NCSBPzgscRMPivhj4KIqhXGhhrZlMxKQ7fH/+R6ClbHgwAA2eleva7zJ
F4kn2gYg6g5qhtQhBoOInS1LdfCkX2ARZl4tXLktjBHYYYX1jAOu/mOh6TV3fvug
kjiATBojUKU+M2vg251FYiCRteiF480+YZ20kOBt4A5S7q50FqYOgWnPMlrsHx+p
88R1+E8XrW9stJKUHoHlubSyGcFj71FPmCuwcey2BWatAVMejSNPJmuBXEMYSuLK
4P5wBah1CbudfEcyH8YYko8uEXeotzyQlxDs4VfPVklaY0qmnZdH4e3Yymai70kk
S18UTbSUFMdA2QnMDFY9mzIKF+h65cs0wZeSRTwFdxPPG7L8pyYa4mT5DUQp5bNL
ytHnAaJBXXPQLmw2x7JC8rcgvQW7r7BSpUHNl8GAPv5Z+GpgTNX4yA57pX5rNulQ
KferiMKd6yFCIG9Gm1Ty76Y/0gjhdSP6kuh6Go0RjEPXsBY3JAxBGH1v43zpwA2i
qfOSLn1Xp1aEQ+CzIE9RLgObPCTscVpYJcbZv0G4OmKGAkAoassNu05mD5wnET/2
zZ2ne4eYZAhhSeCCBtJ7v/4NUNmR5qrK2DFI3NpJnJs+HvemKvAKkCzKLtYElGii
pbHI42Facw/pvtMA8oSf9njlM23Y4PiR23zqLhLLeicSv9FSJiTb3a3oRku3xtcv
NGrsjkQ79l26i2TUyEciJ9aJqQg+YJk4Kxm1PwsoIvSfmWn/5OKDiU+2VIB8MAM/
34QFnYyUVToVqC2ovKxKvYg6/siWCXKussrhdPH+bp7+Ae0NjNIQYlleSrFE31e3
l5iAvll8X1rYR3qbx13QW+XTR+qanKunPY6iZV/OOqPjAjT/Q/+lvfXBeRnIg3j9
geB74FY4Dy7Qz3tzpNLaes5LHENVvlx+VxsoYkFv7hdES+Bcd3Mzh4R0kS/5Xw41
Kos9yYOvWqY95BzZXOPqxPnnp9hC4hggry4tyCZMbVuQ5VL4m/e17OXgwzWQpQAt
km9ISKXAuUvSL624O/zFHTtlTHndRNw/5ZucEfAhuW6MvcyhKrBhq3ZWVnL+FR9N
3PYVIM7rK6M0eHWp4vB0/si6argQvI41QERayZSnDqFbLiPCq2y1llpPp+rP9pXo
luMnP8syYbquvdQ/cRKMLhDtzO+BzU7XOg6G5h935sPz1B3Q0uSHteX+pxHdhIOq
Fxbg23Bq7m/YbD8VbVr/b8uPbNwvBw5u3JvZ9OLkJ3qFvVUogiGvjXsplbKStQRi
KelW/AckGYltVKJ/ADJywLV40SEWZ94v5228rAJj/ucPanboVZUzAAsxCBqof/DN
RNqasUYxGSs+pq0KYmVG23hZV815iGAlDZcTYGRr/ubJUFXG7Y54TAAVzetf97C3
LhomFDai92/5fEQNyBFO37ZA+bqEgoPicEHj1a5oFv3LGNuru4r53nD6+EUtXaFC
8Q8MP4EnO4jLk4XKHz9hUariLSoSqKKo3dWNl22jBsNzP37vzTc3IbFpqMyMleND
TBc75vljwg56LtvwDKvaMc7Za3riVGTRHMeTSV88oMEAxo+wGSaNGOTFl7/BqzCV
MeMasHrDJ/HBI/3Kd+eTt5Y2WPGScQcBKzhaXvGeNam53bCgW9nESjw5uqYR3LG7
ammcCHQX8bZP3unTY+1fK63GsEmb8EgGwf5loZV92hKHYSfOqEsSHH/bJhqoIgYn
aXfKkTzJzer2qPdPIBT2vgXRxCmvIv2jRJ8lHEF18eW9mQxaUHaoiJk+aoWH6mwm
Q9wj2MszXuujS8VNAjKQHW39W3UZggPJHJ71jjh3LNYs7jC/q49USWvPK3ZF+//M
jKdHFozSWQEaWCAvAH2VcqoVLMfCXGrBCS81Ef7BYcmRwS0ElBAMHo9/KbIbuYZA
Nq69Mg4GxqS0z6kjCt7MdHiAWZvFabX6R6Pn2//k2isemvyB/vkZuYyvBAqppaQE
keHIYtVY4WDWkhostzZ4m6ODPrYNYVX4gVaebkMyo03jmERh0lh2iZ6uMYunzzB2
Rbp/xOchpkHzcXqSOt8GheLh0ZpmpxgdHqKlYQhVTHfOj5nA6+qBFEzO8aEkOcYB
l6M7Xpt17DtGqry77UwZwiLb0fatVhWogjWKWCGAuzpqx/19VpW1VgClAaRhhE6r
0x1rZjYLK4pKq1j/D1vz6E3QxeZDHfk8iwtNmWYUekFuPVTiPKwBrMSW0Ex6pSvp
7/lm5BsMSDOKlopwPbzkAigvJOhwIDRgKHx8NIIDiv1ISzXYuj4l2cOfK9Qij9np
Rs51RP/fp/ccAn8Z8Sfmp35tCqSbBee1tY68J2zaQdBQL0fXI32znx/Fe2Nr6q3C
TxDSIG2Iv1en6uT+9bRUcV0ShKysRZ45kCQo1/Vs1XCVIINOGtLi2Dv9eCeHTxHn
DkmTHHDEaLjCkfhL4tNdHa59AiqUbEVIL9biGqNk88f+I32aAQpRbkc53PO6WIrY
GdsGEYf+ucATUtGxQmtf2wpliTUaV6B1hcIkUl6twgsF/FwcabtgmbntRnhvQB7c
yHgqz8pZWpXAGMz0/DD+yIjMx26jS2qladyNLX2vKden3qAfiedtEs8aEn7Oj9CA
0yfvEiX1qfeOao2UGHhGQLKhZ3kdfb57LBdo5arpVAa2QlHpvyXnu1HcHLzvuJjB
lDz5fS4LU/tG6puXpRxS2USOroWbWlEPGgpHc/cGniLt60Ll05ViyehPIaCFTTAc
4cVBctrYF2X1ksKbU7es2CICZUsri6GRlpGNZR6vlC1QqqcrmeXBPXXYahGsGnV4
ioq6NQRc/8ryYvIC+pqZse38AtOZ0G2OcbV99NrolQd314a9dplPC+b0TdeWPuVy
b2Nd2AJyfwlNQfmO/qyy7fMmgJ8CsyTGxK77BkLQcQiaRDd2rysmuG0H+EfWITM6
KzUV5v3szq+3gSrUeDDXIjBCQfLO2ZTX/tfw36y5XquuHTO1FviotxvFFTHCY7jF
9xyC6mL+J17CJKs6VFZV+N6+yNlB1DVGm4b1XX3fEOiZUXSU8wSLat9k3mvvXEC+
Tlei7aPAepELCS2vqOd28Bd1+19ATxfhYAtOki2ldLxzNmD037F09uFHo1edaozs
+1iuOD3x56HgC+WA5eqLJOEmvgtdaq/nURfwEU6OeakLQ8WD3mxaxSq+r21Alj7N
17A/5yFcOiK1PU4mbFPkEtzPOdy5mMM/jMI3Vrl7j5D0nQjsD4OcXCpi6MPsERja
s7nTkSLuGkYGNV+94rfQj4htcUxGJpZ4P3l7q4XXstsSm73ThavubRAKsgwvu9bf
9KltO+ntSinaYBvOYEZrEDnshv8Tqici4ksSkw3iQSZy/ai3kWOQLblEnagTv/pG
YA8lwSbHXUcE6/9OWdwzHjVPtkiCSizUtU5Muszw7avrjc6470WExvzqjW7ioZi5
BGW+6yQgV8gVBroprCH++uuwftE0F+UDggfEn2FMmNuB2jIvF1AABy1mvJTNG0Gt
eCqVgSggTdBMUc7XWkcbbTW3TKzvRXWhAxSi3pKOjfGUFw8+PuTbQ1lN/eLQK0pB
B1oUP09VSNGfwM9VmtJ836RG8UiIN0FO2DbgfKjk0k73WgimxWyn1ifmKfBM1TC2
VMKgpy7ZnVGe8lZEB+cq2yL19sZyeaYlIkvv6PjOCYB8At2RAljNVx6N/2pKJb9v
vPWF33L6jbwc/GkYjLvZiFiL0bz80or3z9GBpWDmg5RLBFHCVi5Lv8nJMEfZeN6W
c87bx9Ys2GoBsu+oroRINsqHtRROpbd2+4vZE+65TtdLWhv871vYy+0XbFZqVYLu
XCeGlqsMTjf2mT4VAPat9nPx97QLarPbWOfT9BjxHlvpfejgvjqjnt0ofI6S47hV
liIb9B63WGUHdu4xxl+99kMHFbvwsfEJcgzr3lxQ7hObmEZ4p27cdO0orxbwP0fL
nX7srSB7xt1F/D0F0Rj5FZdZscY4sS/8dTaEc9Y3Nkp+EBVLwpbGvVplaimnxTiq
/2k60p0zGczkGgcAT9JyPUZVC5bfs+FF60pgZp78T3Eb0F1Q0eFfUiPnN8HaJYlz
t4xp0WAj57pXQXCvuJVxhGe+MHSL3b46OkMI1csW47aF+HkWpWc3xJMfLMcKZV6B
vdg1+x5pbJ3Yq5ifIWT1ni8/MwjykQZ9GTcTZfZ0+t2kH+FSuUQgSkLQmvQr3rpc
IrIN9i+TH2MNRgvDyHN7Ly3y6BPzBW1KFKPaEv+v0e4SB6LoYt0jlJ00SO055ymO
gx23eJkXIoBrcRO58dWy7bZvgh3Q0bklKWUeMLXZn+lmgwPnfjagCu2nDqkxiDd3
oMCgkc5B0mdbFDTgHuF+GIrW3VFjaOPijmBW7GZ3+GHlTbieJOtdpQQDlQxEjPKE
JC17Klv3/4SRRzJZSTJMIZd7jMMWtcbJrl1MQASSid6x9ma/p1b1h17A0/fjZYTm
LRuG9JWQjsOAfNM6PH+RDtBaJfBiSWB31IQTYgRoCxqYL9DLdUOv71CKgDsoM43z
gGR5v6khzRLee6pcpiV9JPAMKk+pLD3mgdJMHZDv1psmD3Y5PTE0Hv8snraMUMuh
QHxoaHpdUhpEOEiZ2MsczB2/mmxYo/xW/tgIjgeakPDTfPq8s9+632H7q1h0z/m3
2rxxVkGZAAhmWwRQ6HeDUyLpvcmMdM3e8uELLcELqlJxhltoFvBACkehKyCacN8W
PMkoZ/X9qzVYRnIHePhkmyHgvxUzir3aAU/+C/3aJ/9X7CcPzkeA5dmd3QyV65vr
F6YESyDgfKrnI2mRaT2x1UPJDMKkrCG1ui5tt/f2Yx8a17XzrlsShLM83tN+NXUV
zJd+utzCncHWSL+Bc7+JAV48c0/CxO1mocRrA0EbWgMS+2Ia7OpUf/SUfqlOcYeX
26ehsU0KTxYdlLz1lhbed/r2C07dDwf3hEz4OKpCIqEXrFYOS5a84eFKJ3rqlbdR
GWRAMShtB0BatcT+ilFxy6c1G/ku3eQKqSZFMfNTBf4TSdhUKmW+H0sEL1AlfZb3
XAf4z6sV++V1u8EzOUgvqmvQzKR1PoVlpW7tRBb2qiUXsvwRx4vKqaDTfaMYtOLV
bNfLQClioOP9I9apsCVrIyZKIA8bEX26xf0p6FgdFrncJkSnRCti8AxYecowHYhd
blcvra7VO296Wqcsxx6ILYQuPPXSh9VG21glhyvKpNgxqtBfCv16kRxMWMgEoXPe
tcn8cKVu+VI2VdyyUXkWVukGTtCRV6BeYpslj3e9FQKvUQQtPaM3N665pqZDy18D
/+k8mqAvHhjF1nHq8iz7YQ8PFTybsY+Luau99ElL880BQlPmve18u6sFUWvqPD6k
Pi/Lwsgd9dWPQcU3c/29en69FjPBA7D9PKMEns+b5tmPycJU//HBQLStIFUtNYV0
cBCRQa/Tao/1fYsJgl5fXYGJkJHN5+T3pSv7c7fA9Bn2CrGO4CtHj97IflpUmt3T
OldM1kwiysc8iSI8I+brMDKeij5hRUo1sCZpNvgaRF2nNeT+ru/9hK1yQfDPng9p
3kqdlohtTVaCPThP9axR4qs1p8A7ZoZzwJhG9j/Vou3cW1QdEC+j68S43G8SFe6b
XSMQOHOfRTM5NC8YV+E2OT+xyYSR6+Xc0146IAV41JoDkvOs3oaxjrqGxfplYAf6
VMqaq1oIchBgQaxt28G4oMNXmbflsd2hkE5mLTD230xJ6rQupteogDGkOEsXK9JI
NHPj5gBUnwRFn6RFfjfxi5dwe/oXvWnogyiYuwNTTHaxAOFIfxeDbd83+/URUSym
phUyN03ifobhYM0PNYeqXDyZf/0Jm6zx4QquBUQead1AmHrUYu6iT23+B/v8N2Kk
FI4qBPWApv87kS0KjdwL9QP8WBIgy1mD/npTsL4Q5sd8QeGyCxtj97GCSOnBkJov
TLcai1DJmVAz+Lm6/DtmpKq0uT3BCV2XkOqgPg8OWSAAeAWVQcLih7oAOpdMIFra
M9enMLaSKTdMOgMF+CkgTAmsV77rFuvnIAJLTDOPhjGcdyIDJS20BEeIXjuNhRF4
jOtAyK0YytveaWTfiZ2tW7AuZefr5m3GrcMs2KhBkYbPoxnhu1kTvpwIiSt7tzCT
v6F1sL29pijzj8BRICFCefXla5EEtYg5JeFXXEI4d0H/kiFddny6sLNdrGG4wOu3
JheTKWANxQxz+DlISnJVnvhUMhFqfD1+yfwkK2OG5tVO4xMeetuugLIpoznUKvTd
sACDPnD1B/5XEVQkul5Ox1mb1qgXkgrF4USrluo8V5FA0++lOgtQWSglhG5Ubp8x
VWZj6d/Csub91yH/IY2r5V/Oj1POsU9bRnlMcqO6QFG2g94vzWJjBmFKL7JGzHCJ
LH7QkmdsSuWg3MRI0bvlPwLN7eIcGsztQQDf8wlgaHWABA24tR1L35U3iNrHP1Z0
Qoa3KM++odFVRJW956a3ez/MFE2+s4vcsQlnuLG1D4x6dQtqXH/H7uU4+eMKk5km
VZJMzM382nspOiX9Gm/5F/zi81/9GGz1+MFpi8vgwHEeR9L34oRJbgEQO950LFS/
545FBXAz3qZOSvicEfEwVuVTIxv3c2bO3aefY7KbO8i5opUp+8gmOrAx0Ovx3JOM
kc8WiEnaMXDgQ2clsSO61JL7Xuaf42qiFps1Q5W4e7vlOqXOOUK1U835SZIhBtrg
+MqLTmnxt2mxNWfscx1Qroy3EaT1/34PPqlR/F0IR+e5ioPMs+JPEYDMKYv9UOtR
We4Arc3U3ZW8AXYxoOtnMSnoQZ67g+RY8CDWRY3ee4uYwpcYS8Ex5ADEL1AyS0aQ
pnDFGAzCAdox+fQwP4rfP1J+fOlqebQRLPo56SALABqy9xdoQpE2J046uTBEdRg3
sfBQcH0BdYRVBv+9VrhzU51pk4G1/l/1XsL6aWc+07YvRWQhIDmIKK4zEvr+6WqK
6y6FJnFE42sJRvWiTbu/JJrqZJ2jlWscjwwojKHQgvHEBj4XmVgwBtGKjrJXkqL5
ioqKIhSkfKs/SW4NyGT3y86QGJC70WJBmoEuD7CPVpsDwQ87KMoLaCyGO37LtoRv
flw2k4VLs+svRUhBE2+aOlHD7lAHZzURTSs33EAbAR3VijASmssYLB3+NowK/TNN
CKqABtbXhxPiL4scJIc4UCAuXtUxEaQHg1zViAG2IaOV2jIuclwdCnEdmaKPcZdT
czSyM1o1DMgg0mTAYd9DqB2hWAaiCQiz/MoP93BKkEZoQffDcERvp6YKuGufFzXg
P2nWtqb1JSGBMV2wcJH5gJ4jKUF9i+zG9CRCSoEdQau/Frk/ARen65fHxDwLAYtf
27GD2i5ORpDNISKX5XsRtBLneo5S9a0WU4ak/HWqJ41DH6IyNMY9edAATs315bJn
xsYuofbB0IEwNoi/jzboOp0hx5yT6MuIPyMKB6r8FHXetBpn0ou2RdpA2BIKAm4m
uYO3BjMYhk3F2pYjPMmwylptTmdYrvDTp6HFcujb46IJAz4eUDrLsVAnjr3b5Tgd
r7Rc7GolJPU8GGJstOl1pDPrzBW5vPCRlF1LPUwLOfSoxvQlKfUJthkV9LVHet0s
QpCnRLwOXTFyGqvci4eTdxEh5QpRSYzMRfmUaFfLJWhoUQaUwd5tFC30qFVOYdUW
+H64i5dLb+O1UEPr0ZxSCELZ5LKF9d6rPRs635dlKRgVkwnV5KU0szfidUGNw0zp
EV/+6K80hDdoXEEv0tDM888z0BkvpHl2R2RgrucoTHCTHpd5ZPOHdfSJDrbXYFW4
3kHFd9/cpQ7/I1ai7/gL8qGG5w30zlRAiBoB1cRbF8sV5K5pzieEM+C/d32jp6oj
WbVHtsCKVgj8ONOD5/Mq9sTTgGW6oJkx6n5RnTusNezCHMtDss2H6kf1uVyBQwUS
YkroBRs/W+fNOUzn/rcOkJndGgLsC6eppDt23uAe8ZeAoPuIam4R+dZuj9FSPEMu
r6QxQwdoEHpulCbGSb6IZ3i9KkPbtWk9RIkeTi2EEB9pwiYemUQMRzRldAE+E+8N
8kxssCtJPYtcX0+jYGeuUjixHEoLdyLRFchJK1xMGI3m68OdlekR6EkzyQmz52/a
Mw6HLVP/mkwCDnTWzddrPRJn9F6sQnHJ57jYEJ9ZXW7CksC+YNag4WNAHWa8kzlE
8GqTTKxHUjQi1cfnZ63X5HDpuRCrH5gq2vcKgPCUcvEK2/i70XQndczfkywd0U++
YYTsOPRpSnKdWz6FoATCgBdin5zyg/aiDZQsWd7qifsqW0Gs48tu5fvjJIJUb9yA
rbZ4b3MUTSZGKjRAQO5ziGDD4N8bH3XxyLfLrSCf1VOFs5Acr2T+EwPbrAaXPw82
kj5To14aGOzi/6ia1jVpDzDMbotLxLRr7W0m1ahHenQ0iFNJ9TGxOmfCBn9X3PVF
HD1Vf9diWPzYA0+g4kC45jL0th1ir5f4OWfEe/+o9tZUasFPY/38KzFK7MkCpmYz
CWQMUL20jfwyb4lhnKcbhv5N+cId97AN/9VPHN4+1ISjASgOZGSZPa1bqhPOXxOL
Itp/KcN6buDJhMUEfhL1EZ86D/XbF0pvVb/eKrZ/kaQq6UuzKt27V2vYXfUyK/5q
2I1jqrP9FEPC31mQp4Nvh7ngu7gLGJv2wureQKTDgIn5KWihO5aEOZG944RB2kKN
dd2WJUFaZqJQHphJ9JQuNwDQwmpRGjYKYXVmFOWRllmCAqTQD4u50BnG6yZB3Ehi
mkOILcI/+Q1wzpE+5B3GmrFjTR8/K/ADEvMC7pVoIkfHkUW4QDcKv5k8ALCkrsYR
gMv9Rl3lyOb/8DrHjcA6aTiVYe8Mz0gyhgonWztb64Y8OZ15i/NT6fdysS9ZBDjD
Ttnuya4goihksn3ML2DAZjOzUhTU2Xd1xzl8935i8V6S2D5YEvA8utxJh96Y3aJC
HLjS/cxx3nsE9EPjnsPvjL74GotQyxo9YAujR+kfygeNhlQyCVxSwoC6teMOJzbT
UqPFwVDr+8Y3TFKeJJbVlTtOQGa+LjINDb148J7Crl4d2qBPpGHNeugn9Nrn9Jq+
vHCVNEE5w3gBBVcCp1imcwUb7WQ5k5t3RyWghIRFPxfE0TbuI86VpAMUjwuriS0X
PzVxKTIr8YLin9NWblj1C1E7aRNpMfKwyO0ky+4n2FHhTSmkfhLoqPmDUdPtlb+O
pDrr37xxXZxqm7fTknhiHXWEb7WkT8/+Q0KoqOFppNgGF51iHZLIBA2Hu7K5r/gV
oQ8q5LyfHVT3EZAHK0ZbY7rD+ld+Diw3uslc/v5XDEBP3n55tWl1y0crhlZ/5FBK
4AfiwDbYvf0GgozwBuC9e83e1Xz9qPtw/1BHAZ0WsLq4j7J8qZPBxQIfLv8qWgvk
zOfD68b8UA+Mbwa5tur62jL+dtl3EyvcGiqMsaoZWd0jWjX8aFJrVC3TdlvmjXxK
kJ8TNR82X8jvbpbme4G6ip0XkGOIvO7vdQwrkT7QJXR0frwlQAn6dKHlTHsKcFw8
8SNHmCvBSpQY/5t3sxf2Sz5CU3Ffz1gL9CO2OgG11d3B4XRYoZCTjpAYunAATeKp
+hF4TS/110m32GoZU3xCkHlpXGWTAul0guu0IPaHRMtnVX4SxG9lRcD4QVnLNG17
Mxvt/KZPVN9ytEt2U/+yDdYYysbWbPQ4Y+LEfMHk7ZjYqFdNmgobse5pN1TmY5m9
mMzK227p7H7RZzv3crFqAt9XMQrTc9qXFsA35l0x/ZEnmhQc9HRaZ29/rMkw0NIf
c5ggFQFffF6ey0AZmuyO7ou3ZtqaG2dJZxeynkdD8sZEC5TWKwlFxfL30L4GItpk
0YiRkdySHKFwc2p9Zr++eW3VADWNP8tj9zVtIo5yq0Fm1l6P6PL3lnGW7K52nqrv
vKwHqgydWW3Mi77PCqAAZNm37Sy3c13fjlNndQ7L3e4gCB6TDjR66nkD2w1M+RTI
WWEJjkkHxXeZ03KqKXZu/Nnlw2vA4X8EJtdGjdHlzI6Zg0WN7zRYiXZG2fy3hw+d
Val73C9GKDeFvfscD2xgUXBm13Wa11f3OfN8VDAdNJolgdrNQnkFt2mFHptQI/90
/yfl0Jh7lrxKV1r+v/Fq4Kjr3kKDDYT5YDvzmRJXkkNN0Cba1zko14rP16uWo8RJ
+QV73byyA0JTx6RnzN3Tc2mAoBaxpLbfTww4WGX74WCzv65CI48sk/28sUJZ88A1
LiNg66pQTyOM3/z5ZYLHjbqvDhEYKqMeMMF6KeMn6f+f4fwKCRpeSWkzbS2ED383
Xuh7JyUcVNXCxB1PmrMu2SkKNyToTX1dntJHP5b1JDIubVpxKWlIAHu+p1krdqVB
uBDsKEpZU8z4g45hG7UdQGiaX92p8x75wo08WKulm60W2cl2vpNu1wH+n5ZeLNA1
AOe2DnplyBT1pjsTNZ2UaFX0N7d2YXNaTTyvbg/KlqAd3da770oF3QGTY6Up/yv0
DMZYTYuVtxhv8RuFAP3fj4ZJgVtdV725SuT+ejrADBF3r2GcuI5fRuZxowmCWxB4
kOgNhKv3WE1tjrFG44eolvCZtU+Il87linhIPI/BATc5WaMQ7TZQCNS13Jxff/B4
6OBU3X/nphNVLms/43ISOPk3IN8aObeIdIJQSd3IxDlRrLQd5Vy/0ftSIKC5tN//
oeCW49Hk41mdydSiUkSBQn9kilRu+sY2LBWQEhIK8SO7NvH1xDeXTWHPug05RWP3
nDpTxUrxeciItA5LTbNhuAwHwt3SJI4Bin7NsX+Tw17OInp5ncsUIHgK+nifBCSl
jOW4UuqymlrBbCpuEPd+CaVYd0yaY8vghmoJ/LQH5PUwBgQ+bDrR1xHZhdCJviPp
YvyDVeOej+vTPkoW8qgTFC3iZcI6S4+d939/yDqdx0U+VocuQomE8V6uv5qJolwp
afGRhZTreVeOdsGYbH3QeEqq4qau80RZ/9n3Zq5Ra06mlwDMF1JoOJzj1fhPhM/8
/MkPrwTkWOKCWcNOPA9NCBy+Do3FUpMpuWmB7U9sSZI2k/ms26zswhPYTLldOh4J
wiorinZG+NIntl9bc6Udlk4jVjjcU/ff5Kr6ncOyWiKD53PEnZiqRBglJFzAR7jZ
CsU6azCjZzGlvOFjTLCuZkYXBDngW4lXb2l8tMwal6bYVRI3ifWkYSyDWVI2DZZq
hPXd/gJ/uDkFESK/nzgq8cAhfNjkXVPQkAfzDoakLzf+fyJm+6Tb3PKMUQ6tznIf
oxX2EImLihc8DryDzUR/RNbtX8koxwukLOfwvHqOgFDioWsFteOiIrstxuegPiT9
YUrhOXTxRWVWLCpoDQuFU6IwkEDte24GIyRN8lXx4AV1Zznieh3+6eBFaNmt5pYF
RM/OQRutCqyvqfiM6dCQhTbkMfosFSKYmyWoC+L707yWl27RxysrIk2jof0ir+4K
mUr1ejlJXKoUDv2Ug/tkqKyrRjb4Tatcj+JwlL0L8Ox2yyhTHWDtILjDp4l5Y/vZ
1eRCWPU67dA5oT7T7TfpLkxdz9odgDPsVtLE56CV2VtIx6dik4JoRINm2mkmdami
gmqFX7IC9X26oXRMe2T57OLQzHbZ3KVZn2OhvtC7gDMHnFfdRuzBV7XW8Fi4HAEn
9bILq0l7CGTrjjaKSCAusmEa00a3OOxvcUPTCowp3sIgMnYqc3pePPy6Kl8a5z6d
3s4mVbq1qjsFtL4pYbiBt8kmSopRHsPxDdqH3hPpVID5+KxBEnrSfyQ4GkBawJkr
PI7lIdR0YyyZwfFpD6NtUKBcOOUsUMmACBkzTiDN7V80d2mUBe52y4Bs55Y3RodZ
viV7/mG+YUEz2K8MV73dumv6iU4rFi9IlW8nxdsnTX7uLP10POHjmyntTNCiIvBi
/VKzdNJichN26rG0+/zAI6TiBHC2Ni+saJ9S/Osi2DD9D1c6XNZe/hXf5mkPgWFa
0Y5JmLCi3EVGmuMivQ3x1IBJVhE3nKD7FB9YgnnOGTu08TjktxDRWePYmyhVXXvi
rWBu+ORuBn5r+u39f+Okjk5YFVZXAYzgYfHPsBdTJqK/zRL8cu2nDNs3j/o3ELaD
8AjcqcItGVT3ALd4lhJ6kCCjuDZPGf7JL6vSlhpgH9bv58SBrC32mXzi+hd+Owpf
ilIyTDmTviVF8AjR+IRjbXxmn7awOWHnYH9EBq8uWDXzeRjjBjQusUq+oqzWavmF
uQCcxhPQMW79ZSlCuED4Tsjw2dh+VpWchiacdg91c25QTLs7wNTkCwgGJ85eS5lI
c10LMA7M6en4rSUThfSsVAzVbnDfc8kdIOGXOKEVGmCA/Z6gaC70xn9klEoY1jcK
xRZahSjcRi+M0UAWWMlv4hI6TeRexEp2wr33qOlKxGlGs05ghydp4JAHwBN7H8G+
d1BeYYQPPDwsXKZHNESb9bTds+rddLKbHQnXRjfhnhDESReiJA6tvv0Qq1FvNQsw
XUOoNSOHWQa9j2lE7wFK54jODaRVuAcrHMXzlUKdGrl9bkrIXiCESKSuge7EVYb5
JDQyIpT3UntBBxoXyE9QXrMTzhr5IrnQzDWRjOPFgel/1vtSRCNn++y4lBZUvAu0
ZPkO971yOlmVsMoiMYsJTYUjQ9jeTuHoleD1D/GOaUThlDodE6FSIKtUIV/GVI1I
t4Jq+yEB2/kw7e9FY0cAZjC56aSRMZ49avtCIChvtdAyswNgW6pD4YhoHr0TIDoV
A0NdoG92rLFbCKBCgQnTCXCQ7yK60JFt1rmEL8SeDY32S5MiCFbDn2iXjlmq03uI
n666Eu/IQH8vV7GyGGmtBPInYamS23TkZUTH1aF97xFz/OrNiyCKeg7Fqd12tE9f
fgujjo3mMn4uGWYtd4UZq4efop0LSdO/RhinzLodrdKJzcHV4qbpd2IDgFGc2Rz+
P08vzYjrTm1zZkfaeMmFGNXgXM/ELosU3eBy1cXM0JLpLj6iRS3e6YmUppsMc2Su
waRtFKIi4Ry9fAgO2sxaAce9qWhrp1Zri89RAVvq18JE3yteGURGhlRjbbUKJ6Xe
6ZGqlf4pWu4MyVwks95V/DIUBlC8D1AfusGuQm4KlDkoXF9MdYtTt1Hc5w9bojCd
uzWdYJzG5+1Re6LNn4VHiPIyhUVJIo35/IlXQx2hpfUFzqzaEq0Cai+pUHcJAdvA
fxblsgOpE9ISw6StRMiX3VhBLmks+jIHIb5z2O+g0t0cWBvoyf1m+9Vr45VmoUQ3
N28LTRZQyIbODCaDFSTt2k+2i6LMISzq1DoovbEFkspbaSIjZAqLExeD0cGjA1HV
uJUHrOWOSNdcbINqHKxd8BbZcnX+6naYuZURsF6WPBzFF6+AMDz8KTxWSRTqPY+T
nUBhOaFqrDdklpjw/tOWlC/GxH9bHqeHL3w1wsEyA09I27aW9f7UBQNCJBj6Lq68
PoWXLUxYH9B0zZEm9msn/BP0/RR93oB3y/Kf5JoELbrJySrw5NcJ9YOLHv1gFkju
DUh675wvd98PJEUif6UJcE7cSp46h8UosvDn3wsnuA9Ifi42+OEdlectM3BpZP5b
o5dk+E+YCHJeJr9YbPfJ2anr7bUqEY6QGYzzrw23vUKnDyzh9vy9yrVO16HLqyRm
30CQ2O5+wLnxQNz1bQQB0KPHmZklbcQ8WGSiGN3X/DQVdQo58XRqMsLiefmobr4v
iGONt9WRB34oxdKnApaM40kxSjf5VzWCrahSqLO34bG42yw2Ej+ZS1gKncr3G9Co
P/v8fWUOxJGQPoy01pMWC5ZcMKys9LVWM47SAeagZ48v0zi0Xr0t2Ahi9ALmKAcV
xIpwQpzDsvKfoculqYo8rbUcVWwJXd8S3DdTijxf7OX25kHTXwq+nW6IbzSdWxDM
rQPucnHinug5rlqEp7MqEBLrPuWCJOaDDqG/yI/+ID01TLNelF1mlf8MJncWQOjU
4cu6VHeSaaVj9om0qstFlBdPpQfp6voc3flRbT6tW1dZ2h9tShhTVPnLTwBeH5ob
Mr6sPB2diOiuWlpl1PGkVsMSNELAxKvA3vn910V+dtYKPSVsQ1rR1pNe9d9F7nH6
QD5hvrJbg5R6Hrvt8ysU/BPgExMz/AYsCEtc5/gp1f+51iApjztbBAXFyZq3S9Z1
VK99JOPEQB9kq6wdzNxzLNyF3tVS2U7lvkDJqYY8d6IphnG8+8T5q1K/QojYWyq5
b6YB5r9uPyOXGRF+ix9uBe02MMC7ayx90hvlsX3LIZZbIJErU/hltOwpsuD8cLA4
k/XFEHg9KJMbdJNnSccXyak29FGj8IVeZf2/fFL7QH65x3T/IhU7NxDJJEFlCBYb
NYRNydBPPfVw3mrVSTxDFfLzFyIoTF7QB+kT76hSmv+mHZuuSG9iE3vb8R99OS4Z
cwJ6qlrgBGV0S20VCZZg0ZjD0QGbQD7XA35R2RXsuVoAl9ZTEsmI2WfaCdv3Lbdc
DffF1ePrN2wrGvIBHBa4+OtnNAFU74rJnFhHUx2wjVmEaPuHYpeC1A6XksX6FmRx
MxQHV9IUAJvKqv5AhkMmQyV5MieOb6jef0NnkDeZGJoq3A4jwtxeQjkjOf7tKX5y
Wb/qUTb8odPdThm5lLmLrIfs3bvDkbWbxDqsRt/JpqGM5fTqX0w5ydte2ajhPs/Z
rBH0ZPMpithGCwSMdCK97/1lkd3B+JbEM3DBKKsbW7Xy7+dVnWpFweyqRebDC3e5
Hx2C7E3EuJz/oiHGm+PhDwXPpzgghxbsnomXhinwxTXcGDWb0dfBVeWLb4L6XK6n
jR+UlXNNSHeAnIeP9vQlB328iJ+O5go0G0QcpdOsZAzV3ejU2ng8yieRJA6YjLXJ
MTrwstR7VxoKBz8DydaNbJTw9OnreHH+OMFlROpOUfQMPgSKnldBV0688RaGM5yE
nESlH6Hy8tApxSLch7UyuCQtajBCwiBda7OJS7pljtn9R5qqV1kEyh1209ktVy7u
8SuDCNlKVh0UNzlbOIn9JnXd7LFqkUhh4bfgjzoesYJcfRYjh0ZI68EDgXw+B0RO
2J4HptPEaNf+rPr90lq3j4Z1SqWY4zqawWld3MGrKpAMoDm2TR2fvDdaG+kQvI7t
hNxphgiuPWxp0tyVW65JEv6wH111ZvbuWuYKz5RbkW+cFgwGwruowKeKWTdq43MV
Z0I1MCa14OX4QWQkrE1u/h/x7OCCFMWmTNfgze5Jaogphcc3dfpqhaUY/u/mStE5
i+DYZ6iBi6JOuSiq7IX1lMqDAWMURL+a/W3fB0chsuNmijv3xAl03y/zW8rNI7Dk
jfWlaGKfnSKmh2g3UUctr4z5VvWfpfbsNw9Heb8GtOUuk53i/f9wkVu3bBQgiL3e
ztJb07CGvk/SeBEn80iyLystagiIgWxPQQ1M0+bb+lM7LJ8YMFFG0X6mvqWRjc7N
Bli43vq64MKyXTjx1Eo4RmaIQ+W69qoFC3ACYx6kRyDNSVYqv1c1HgS2NGi8dR5z
RMbd/kcP6cbLl3XmEPrrCUqZCIgLhwgzua+1WEgC9TzjhGKH7Y0h41qov1Vn9Oti
oHDoFNVSYdj8gH5LxiLX5OU+a3kKEUmpVyiP/a6+aZ1oPCcwSGAHW3gV1SKjdB7F
zGCQ9scaa2LrJkklxqr6DjXEfCfy9v3KIdqhYPMQ4NJ3euchgcXx6nORMFKfiP68
I0/O7F55nLalEkHhJzOkW/DhPRTYCZJPd5ApK4SF4TTq/Z2Nbpj8KSwSTxcOnt3i
pVEgtOAh030dDxB/i15E/f6m61LkPbCO/ooOCAFdOB44NT1JjVy4sO7MT16eg0Lw
JYmMGDtd1Ld4g5Vu14snhAbdVxa5xO4PjzxpVNRE1LbNGeruGxUh9LwQz/Hh3RAs
RJy75zwsREN04eCvoVH2qhFqHJMzSq/H5wJBWtssFa4Nx9ndRVzfVTKwZ8GvTVVs
wAZWQ1/FE4+zIxupPQSMYoNBukKVUni2CV06zRq+ZzlYvqSeD7cOM0I8L7g9bHVC
C9TTIXL7h642NaMZKYL04ACJKBN7baCcbnd4+SqXfwOXgoIPwFTHBFfFiO8J2iK8
T79qJMPWB/ADnAB9G7WCsB8iswZdFKbTdcUFGsBTxTkZyBh41hPk7IIIKL1u9GPA
MZ5Tdr1KPD3tpYYW2ZpxohcJxH7fj326CrZ5v/fksxTqtWceIGAojXU56Dn/p4L7
IZqAcVgNDX3hvHNTg9gDg7ESNYzBepjNzTi6/FPvDOdOUJcKlA5yYNgRbSr8YFpk
ea6099+HBNu2NY6xFCwhJrM1oKfsGzeUDfNtJUruuwLhCrmMgGaBXbdql+o05gMa
M+tSNzsGmCpH5qG9Gl0TouqCum8i0cXwXm0vMCg7lSzt7vHcFnaOhKNLvvL2n5wk
gNIaQ2TRyKgWP63mGeDwYJHJUWBNh0IR8SRGMSSf2rs5Wv2SvgU1cPUm9liuB0IE
SaD5w6Y4+J3GwyDBX29JJcisyBoHR0X4ZAOxFxkaCPw4UDX5r73+aU/1hvxwN+Rd
P0J3qb0KS414uP9CJ0NOTkS7TcpFOXZqMJ0DFr9MkH8uUpmN9bunbK/PxK+ePPwV
DnZC/rvt0TKyOCCfw6D//I3HkHaUSf4Bri/0FNJk1r/r1PlWlG0o/XSAes1rxoMh
e39Ny9w4fG1bXk6AJAvlUbnk4cI8FL99dL/z2Z+LPYHh8uyboH7vz7y0FhP1vLmX
lTlPuQHhc+PGarACDInjixdP7Umwjvddz7FBAAY4WE4OLYB4zyz1wM8kCzr5VXUO
VRWqcg76/iC/uAIejsZUwxWZMjbimRRJMCAL4uQvDzMUeLdo7plaenvkheAd9i3L
FEXFjG3OizvqUu8Ac89DmamK+Kz9z4JDyRHN6pQ9PK/j7zhYg+Zz1MM0pdWpl1Hk
sMCxfyEfrkJx0XnZp63D9xec22gq9VpP1TMCdzEx60CN0r2LTiok+GZK6SBnGofq
cT96ytJvEhybz1PNaMhARSB2goEYq9jFbc6pDQlxjZqkrtJQ0/zk9anSAzDS52gV
8ZtayUVOihl3HyOLXY1etu9NNrxbmq7wG+sRyDQ5IAYLOrKlDi2SjSnVef+wRiiD
oblmF+tQWC6fgmTQqV4HuRYx7RvdlpNEn68Agg+BtOuh9xZZ77mW6daFNYX1MQkc
v3yX59J+hKDozMjK1+3Sa+ZfmAPbTyk9vgZd+8P1+syUlijLidGwbFvGGuYzN/M7
Z47kIFHVH3UbOJYm+u1jR8E6mQIp6tL0VXcHI636ee1cGAkkmkK/QTX1aKDcjALB
Uo4daHXWa/zLCnKlmmjbyskGQBwNF7pTKIYCE5xlHTn1VNybshEtFC0jyaaXyp7M
03PVARPVY6qjEkhTcJ+4bN59HW9hwjXUbeI/5o2Q03jTuZfLzDGHAXE+Ky+/GN/8
cTX8vWwngP2gxosRf6POjK4azwcDeJM3dYmIc8YLPhaZYC+KgGTG9N6BIOqulnh0
ka2OqCzKUtLhvxHxUsKFVBTkda8Uo1mq9kySJSoIBK8CHBfvlyVHaGe77o45ZZFn
9sCChAgjl6V0NLb+9ZwB/nnCVPHU3tzQLRQ7GkWsyRvhLHLdhe5sD2gTCCIKEcvQ
Ww28NbOSaODPk97NATDVs2bdvb9dgqfhABmV/0EHaXICkByfjhuW8wij1K7JgYbI
qlHWmdZQdKrMe2FloQ83T4aLEJ7O3d4Vj41WELYKpV83Ho8erQnuQRRpdqStcK7h
18Bv2HjFM6TGKQE4K+iaJtrYy1CGT9LGjwzO3QrvRJ3yrnOzKYxNRrUzcNxwotu9
z4+Jwgf6tAtr0RroOiVxKhYcT3+mto/Dus7aBJHqHTuDQmU7oNAB2Kcmg4FlH+6I
wEYWEQxULsU703x4ewNYBsZ+XykWePRdXgNFbmPVr4fs3VPALHGBsVCOJw09tw87
2L3tiULZ5hUhakXtmhG+LhxbicO6p7jy8Ws8od0LqkQM+f96MywTs72iY/ys4Kzv
MH8tAAMBVc5AEGNBP2jDRkMb+KEBOBHauBKloLcMIVuEU3DpjRu8FrCsff550fEa
CTBIYnxNjMWtKkYYh9p251fhPkTLAsiUhitOtffmr1TGyxwbmtxlUr/Y79OVJLRU
ImlvdZST6AEhJUs9Vl2tPWx0agA5lbAcTdNPgq7nTKx+qrHNADJWl48ifCIw6fw9
dawsX0hQSwzARuOVPv935IsKUPa3hjQyp2YOAVUN+87aDZrZnVUWADGQO69xtEbK
2ihHRcHoKB25FWYRyImq7QgSFCsHZMW3erlurGOrp/cGCkqYQbnrMq5E7xvw1QeY
kq20aWQQIulM2iHsvdyhjrzufJvbqr3CrFzAiq1PhZVmG8+jUdentiaPEH1DmLij
mVktL9eMpMW+aP3m2MBIO7Xka6+aa8ioUZP8vpz/171ykz6sXVtioq4y1kxXTdj9
NqLZjx2tNy1gPW3abflltakKNPuu/kJxcAk5HN54uFJnwwtNE0sdP5v6bCh1Jm3A
OI5/9JM+67GH/d3PpmK61l8ljPuqDsRSa5RLPQmiDiWFRcKN4O16MnWBLo6Hyo2z
TYL0Q6zHmg00p3NM6pSZC/HfnU9TmlnEnISuQgPILlcdzpw51xo+/3dbq+APpTku
9KvqtA5si7i6MNYjN4euopu7sGJ/V7ZJMDEK2qp5XTcg+liXVraNaLsBOKzCZTUe
Ou0eA+ozTc4L0c7ZYU7ZYRJ4R6qIqKt8BCmKnyzdSdxeBK/hcdY15PoZVmhp2e4T
cvEmodt9i/SIoCOjRYCgVxgjG/Z/WlLNNjN33dJToghfO8wFxVtHIflYCBrfyPMh
MuWFIhoZdd4ayNGWncPeoqq+G415FkY70pX2ORsc5smdKB07IMRi1UcCqH9iQgGV
gAsa5dIbP1z3WlN1aMxcQXczBqcUcUxS5ODU3fpWOxWhIgIjrRu/t66fU2dVh/Ir
MigXzb6L6Ev6YxzCXDV/GmHO+pEDLSZuPRg7GNaEEhSzS9SrICu6+2jUs0JZukEQ
iwkF6fI6jHpShLM/GbGddkzBwG/ixESd4dNisj6UUefC3kyIjX+G2NgXWGwEmP8J
BeqUIrh2YoYh+Jd8YhsoXG5XtuQzi+dagaC4tJG+Ca6H9QwnWRaAjvrK1iLyuhMG
3F31hEu+xpI+2noD5Hrwfa+e1siAQ8Ymd5ltxe/MnB1JZlanwOnNu3H72NYqWylO
f7YvR0GK/NCgP1OFXCmBc1AwQwVlLzkK3rS2jgTU2xIVRYPrB+Mi4p4c6jX3CsAA
pIiF4rEfwJohSGZybXfV0y4jyd0oVnxMx/9YWjctuPl/L5m7IIZdHZqAWVGnj0Wd
lvjjdOmVg0ukFzsybt8vIP6Q63cjmCPvSimMJGvFX9Qy0IvhhM1aNfsWcaGeYkqx
Gp/ImpBvSCUssXpKNNtYRRzyLyoE46tLeQZWuCsZxnGCaRwfRBUQp8kzyRAYR6J0
oQFhtg5SYl0kPr10l7GlHcwpz46Q2dMTlx10ghnGxZC+seSCVGGhsl1knBnWAGcq
VpOoGfW3MjiNayZXyzqtUaXzav47o5zYILrtHIQai12exwgKHcaa6F+noUQYUYol
NGM90XdmVmu2lDjuwQVMGr/L1/y0GEE5ZLlj26prH2VaP4kryVfntm+TBfNgIK/z
za8vpZx6fzCM/TyZ+7k3uqtuSmqaccdq1cjmxzX+vyX4eMSrZ5qBTGXs45d4viUi
L1WpWDJKqyQQm06mTlUzmY41P32T1hhRirrO8KD25C1pdjeljeR05OMIe2AEV5lu
m5yL90NyHr/71CxQcyCFuY2nIx13zLu7J3LRAhU44oSK2OlhppJ5ik+blWmV3Sdz
FLYtQ1yd4SEpUHo7gpG0ETFaiYn/8PdQ4iLefI6BoIkGWzaz5yj9fQwBZNp9vIdh
8ImjUv7Ql4xFjN7bIOs7PjmRRvExv34AqHSEz/h9jxlsWiW6dqTR0pZL8wtUF9Hb
7JMHwowRq+Fh3PH6eBPUPONWtBW3U/gDnKAzexbf/b1HfOYTDeMX7JfGJCrN3w8R
qEbLLmSXjscfliYxww4s2C137LkyGvfXd/IXgR5dUy/Rk/QrQ2IVYAzK30r8fjpH
3PJLDZTMnNxuWu+CEUlxnOHwSRwIHxoTsHjppQSjqZX0ZlHd2cE/da+oIKclV0U/
NIOg9xXvEdDuJV2wzQN86Hvw0nQ3+K5bQ0nOaZziO/aKXnbqy/t4VGvso5OIFm9N
1+B1Qot84o3jMIkyc9pm0JgOvEteuRXpcFyU3JPrCGT2ySAvZ69FiE6eivHML9/w
zBchq99l3bSVwXiYEx31uU/OFvSDExcDuEACg73NBsnL/da8vMyoEpysbHVraHSr
pVOPp+4ZA2WL87IeWBrhBRmO5XC7JL/5A5q1xN2ee51Z52oYZQixrRSjtw/a7ja6
qjlapzMhGCQckWbqJwGIf9b5ytfzupxHx3erNTGKEWiQiQ5QfV8PctDxoIsCADA2
6UpYcnvjUgkYCrgfk6YmMHrT1ER49OCdnsv09QpB4+cHnv76X60e67FIb9yniTgB
egmHw4OribHjCLLIIwg7Eer4X7LX1gNI/WE++TdVsel1zPPYA+NlrMFQKwr71ygL
mFZYC2AY9BQ3vXyAlZ8VCIBWq20r4xzYrZilosu/doFAEkwXwK0+QrQWKWydZ0BQ
WbQuB4tLp8X1tP8SnA/qiRvu1YlQ0U+mLIAILdPpynzyA1WkthLaOG7SCMvDj77A
jbM/WpKwoCWybqEjzV0ASUb7PgWXfpZc8bk8NQFXw86OkthUhGY3f5iZkgus5O+X
5r5zJxbkAayYk5UJQtwys6oUSOd9m8DF0lVu4dTKDjJ1Ho7QbqQBSi2MMgsugkra
oc9OrhLQ6M/xV5Vm+yFgJpWMutW0QdeWbDyMQwvOUMols+nHrcHNefSaRDHBPFeE
6PkDnNbw2Vbvt/bfRzVNJkZXSSZvXXPyac7yjjj86lEL7nf2jGsww9u0EGj9rbdC
CRbH1NHIOgOmCZuqKtD8XfAvO4RUp6YF1QiKg+IT6a/wITcstWsFCgP/OzGf2fQK
RvU6oat7INu2hbL2P8AgT1sB9MnJCxEaoR249Pt05ZYTaODiqyrnmdnbtVgILnV2
S7xHC7qaHjwJ9SDQtEV7ACN63hAiMJ1zQBhz26Po2NXpcvgYkviB6DHfMGo1cQGW
sHPT6o6z0GVYOjeaud4k6ZjCq+HyXcxaB4w1FdfoT+Z9xlbZ+Kxyk4xC8SVgslib
NCwNCS1Stzgr6Z8raN/GKoIRC8eXA0CN8kkoSAuheDpZUXoU/9ndgggIzciNr5Qk
SoPdrTrUC6ygrmLF7V+M22K7U6xlcxrJ6E2jlLoPeuAjCRxm6f5ZQMUf7sOInZ+/
98y9exW1l5xpfAQGETt6tiDH9TYr9Mq93A+VXeoNbh6pmQXni4WiXk1PRko1XXWK
g6EpBwdUA/AViW4LpSciZMtLXtSQ9XssDL92h/amympOyY1a5FKW3UtA39IoB2Nu
e0RSeTyIpQ/16V4Z1m2ewxe9EKQHlCDjwcyqt5uU7cF0suVFUCtrdrULD+lysQ/j
q2rnrDaGQzx3/z1VgdsasB9+t2JD2gw9R0rM/+Py0R4Jq4IjNyv8nr8sKdOAcPn4
au55WuoaSp88Blyqqw5YhqX2dmzR754fX1jlTdnBUkdp/AvM7JXbWQ/2AjQYXWqw
USGWi6339OZy3zVf3JMcQnfcS31rtNJp614aNJoYaVy3hrsxoxOhRw9/sTnMR8i9
8XcNMB21JAOYy3gLrLCTMW5RuMli8MUhpNHfdR0t2nnwB6ZdqEqncNr2oT4RUrIu
k5nLXY57ipeNN2NQX4+sVTy5hPF+gRr06uRK/IQRyLpFstfY5n/AeBJy2AvWnJe+
m4AZa6iTJ8XFz6qrkyn4V6uFm6Eq/gtNcZQmtB3GWWWfFiZkyjPvkD01w7jtJJ8C
Vdkef8SEVmQclS78YHkizMFg9AVEcRwLGFrhi4MxPIPW7jUhQjOIofzgcnKFPg7r
Xd7je3Y7QAhcyEoLFKXOLCtdCK1lJFsgS+dQ8z7aeVImOdpLfiFzjXcpmdr/S69C
TaeH3AzUXgvnznmJ94/wt4dA9BvYMfeacUyDzRoo8L5/Cy7LDD8p5RvsckfWC24+
KdqZ9D3h/pT83ydYw/0/fP+8rEesdrT3EgLHOJqxQEOTw+9pSUq7Yho+WLa2ZMiT
i+vDrQ4SCMMq3IlIhtdFB/FrC/uFzGexBEbvqaEAAKR8etonZv/E1MKoDiMMIO4x
PyFIrhAxAB6zAGtos64Sh/OvhsQmj7LX8JmBtWKAdlK2Z/VBxCfzOeIPKfdwtM0b
lU1jU9zLZiHav86CjJtwXzbO6aDoeo2iEqAVrcxc/3ODfbukShKYrNTP5oHl/Xf7
Hx+wou8/P8fErV7RFjOBO0bcqCSiBB7HuEHtMZ+fHufUD87GRxHiblxw3B0BI9rK
brpuOgvm0WHfyUZUo9EauPsWi0bBLcXWa4lY0TH4XmXXw4v0L2o8tFnIaVsBAiiQ
oLttXbjFzJVDYWpa7SCZ4cuS9JTsyXMLj2TEYOHKZwK2cGunjhvzJIjwkT1nffiM
36ut4Ggt1sUUxpm0AWDAx2DJA3o0wKJB5FIgVoSYCWcnctu3x6XzgE+fl+TPUsUb
98g76tk6TTbrb9Olpk00u59MSCFzPYOnVwP6S0RvxXuN5mYwfWYt1/Dd5BBNsx0b
bh/RrFqU30kPVQlmmNd72mbfS4SriaRraCMqWe4hNHjPmjskUON/U1RQYElL9XK4
kdlImGynMXuDBTEIhRo5jBbBmy2MygAMFnwHfF2pmNeH1lX3lt9hWHnUvxt/oO0Q
h13bP6W6+sKd3c2UzSgazb0UIEcINGIOf2Z3v2mkzPvtlxhR6e8CwAzx2yCW/+cy
ECqfQ2fLHuf1ZhU5mpnmG1EQeNNddSp8hce5pRs4RmTQiemnTkxzU8utD6iKCFtM
BmfjGz64rtzjdgeeDi4n6UjFHx20mu7ptnZuJZerrKQ4zRyMj98YbVdkuxqGRmjI
XVBRtAJCRFi+6LGrA2oOvoGtLgP0VlC1H3FW+ubjsRAwNTFkE0tzTfKrOfj3WKsY
CGgYBqFoXB7Mzk3/IytKNHiIAHEb/BwVNHkDMRdm4io+pgOmP1CnxkCFsWdNt5+d
rtIpa5JlxcXJpZ2Rhfm6XlkcKwC8IT/tyAAaYz1jtw0uTHd6aGTJNriqB9/cdK5Y
RBtAQsYdMUUlDQDGRmtifVKT+hba6G2Wg/9fDxPNpcwuIpTpohroOJ71deGXSws6
KdM8vSnwmte4KRztwakntRyYgVYkb/DYc3hwO3CwXXPFURQfiFOX4CFYLfGGNU2B
c89eJe9F6AdKPcDIDnrBKHgdNr0rd2SeAoUxaxbFPxGWUR2/KXrtR/vmGcx0UN1E
OF3opy8fVKKbmhyocNj6HefNcjqNK2lq7dVAmAq+3mMkQKpObunpDVD60rn9RvRZ
FFCeQe7JpvUJcQov7wO6Rl1/U7zfB9TA+t501DRHZSE+bt4lNuM3TtSJjMHXeASq
gn0LwZb57SGO1cEMNChEgSV+cAdIidl3hjQ/4JCTANdg/OcyXJgYGCTba5hXssbC
plxe/YOyFak2VPWGsFIVpherkFW6n22TBoYPEL9KZ19QBvYoGacIlslwVY5gqn4A
S+PQWgWLjBvfWnl/M4Jhz3HHEfltibV3dFnJz2Xhq+h4DgfK9L3XfpvTxYHjef7Y
TgMSZ+gPJMf2RiG/zPXB2EB66lNiOZc2WrULH0Ju7TxUrxVTZAzQGU+eRUTGpALA
MZYBHdHNUMr6BklT9ToHKNZOW+TkOrib4l8V9B5r6LUPG5Qkvv2msMDObwaO7cfz
6jyFoVsUycEu9KIVxgmIYk3HWZ6oNj1i3Z6IqItT++83q1pX4MgySdLKqGzi587Q
EK74T5PVCv3lZP4082Fqv9eOYzOuzkqrLwYTiMd63mroxclkDc4TN94DgtMuYNBj
jJzK6su4FB/okJikqoiaokQyAnGGfZe9PGHGsT3vp3+kNNaSNJN4fb4+zzBkKX+E
p65flF6UUnLaD7m7xVvQqsZfkQfB+JzhIRCDrEeGPvVCuyd9xLC39Ddp/v0cwplz
toiOwziNmVGhiLnCnKS6JPO7/2cUTFHikjfasCFaY4oaQufITSQMhXfTo5ZTuil1
hPuggLW8IXuWfmJMg/h9ef0EkXKI8Zy8AZJl2oZsd9EyPzQtuLZSzK+Ves8b3Ip+
77ONQF2qOuYbl2Y1MB8+gI9PmBQ4tLnKVTdcDYtWMeXCwV1nuw47/eIS9gwn40Pr
NdmD5xTdVGWoD/3BSQbiK2juJponmPqaCcHNoA/jHm/dASHgxQzwxEDMihwWPhKi
EYlYOwSYwM+WGWFVKN2uDrQ0jt9N89HgBIEBe/7kyZTZFCHKEu9ZtkUJN+8tIRII
WLEL3xETP7+HSWBKYJ3Qml9SzAOy16U6CVxHaxf3oBaEgHl45ARun8MO6m6/LT1f
Mwo26fBYxQN9uX7PtxsPLjLmqR2TpSiWA5I0gFODjJbclpdIjB/Anh9GK0vVdJ/s
MA22VyusEK3OnLPUTsqA+2sbL2Wu+oUsEqNNeKHpvxuxvbgOILqvylTAGYZXIaQJ
tckvLnklzDdg11bJM8p5MHtCwyKvFlJ8hwEpHbpwj7GJxd13pG4Pp+MDOKe7xkyb
icFxBYhNnZwPRLFFJL7YmT5fjscnBoKukPvyNhX9+6wbn38XXz+2V/GUeHU4N8sQ
PLA+7hPpAwhdHGP/OjMVQfoeOyQe93ywmnkNnA8PX1F/x91YJwksDWGcziMcsBtB
hUY2YYz+RJ7fb8jHXR+n/CIMFVnKhKtMJD9CFfmpHifeKuS17ThESLoBliGDGnmC
K3US7n2iLqE0hFA+3ZwCqjyUh0DPB1m5Lttv9A1OdKJQZDvaEYMDLD+TTuAFaFEK
d/Xn5ULnjNqvr0pqR1wMd+R7n4XnE9QDg336aZDtDGghp4J8O0i2bCSDlozV1fFj
s7WFtSm+13dJDQTMLp7cRXKK+miUr313VSOAEnQEb0YvyNYiWEZNjzhhgdmsSYGF
DSkesNtAob534yUyFnGEVYzUpeiNnmqBWTzRQIJcagrEeW0YhMDOi6m5FN8XCalR
+Hemjhi//t9DIsTdiyBEuEwfGN84Dhzccsn/qbdYpLfOdcidIPkx271kCqlA6CYL
ujsKLFe3g4LqwUIrczF2FD0G7ePKy+YBeoj3a5ZyeThG7TAQfzpqyFBXDcRFKbAu
01HZ7jfiErQnelj/RQxzjz19pAV1E0jDqX3DjYuis88i09Dhk4mXRYUOZM2StFbB
xXAcSblsmN1o9MOyHXdBy+gVKWSXxiKBxfaavppZ44H9tAgnFz0BjC/oNW90vRh/
h+h9z09x2c/Cj9tKCMASRpLSFYVoSmWD5VDDk/FSdUHYnpnl9L3bj3pxWsDfKGVU
xw5M3F9AHqYlOEpsjvdBkt8cJK8SKMPAOwNdpLfkxpowDNG/AFKwW3kt5k3OVFKB
XHh96WY7IxuaLvVxVNuGKLdED6DoC9MUzgPIcFS49UccbyiVtZEiS3GnfqgSONV9
lmGZyiU2umotvBkjdrO8w7zO2k4nr+iS/xFJs9VvUaNXKr2fDdal9/E8Fir135tk
b5H43Q9c4nijg67AdX0zmoYiwB7M9LcR9FbVeGRanB9l6b1lR6algYPzTUagbtO4
jWofzTwFeJqaigQUHBEDjMQV7uSded8yy2ssK2PEAY2ClaRtYgvW7TQdOeWindg9
0aZtv92Dq/P7ovBTntTQXuH/wXvq7/3Lt+NloC1rmXHuHNUmktiWwX+ClXiteP4L
7Gg/TET1wk3iEAcX43sNexbzQV1iXolSegp3tU33gJ7ivciM32bhR5IuOR0v4eOs
hTWslkqyaplLcqbtxB19af1z3KtVuqIMHN7otxU0aaUceO2rvxTuLq3fBKUKanQ+
SbPxCHd8nlg28+y7bWdR6X4nmgo8Ng2Xd+SARaiatLXRIuybhx2ilYfBWAYCYT9B
ns8X+/hlUPgnLhjZeRq7tgt2Ujg0/yNe6rORtO4lQuAiclxAo+531jPZsXcMHekN
PvfyTBKP1Fx6ChjAiSh/cRsEL9h+zkPXS/aHh6CJM+ITSXAC+1F7MHRba8da9m2/
NMIcWRPm+u47/JLmU0p7YqJhYYE4AG/N8UW4i9ejv74FwF4L9vjK6czUgIsGSA7F
rzFve16/VjTyCowqXq1gtLBeAjakVfgSpYSbiteiKDjU17gWAzp/kVmgj4ilyQAV
GQhBG39B4NxrIj9jGnESAK0TssLBMFhPZrdyyzGhZbqw3bA3jUAcyeqv3jeUUbIr
YBny+UqMCS4MLQJLtGyxvUPG1DFFJN/Gpt/UH9leDzkfC33wMTvx7cEDeKZXr72W
TWQSNrMsKmh3o7wl4sWDB4UHGCODOpordg1UU4s7lrQx4sbEH69Aqq2C0Enbmskv
LpHSvCw80n1Z89ehD+MrDgd5/YOl0qbbua7H7UwAyT/OWK94Nt2jpuZ1eqnCzVdL
SDUbshHgJEJZVg5DzI8DgYBU7apyXzALJfVxqstAIWxHQK8lexnKWAH+hb10/cap
+UWg0hm3iimSb3UWZ41I7HZ0o/ThfCtkheVBiH9lORKlJXnh+1xx7Xfj1L8C9niN
xz7bf6TDNlLod1/bK7BVccidndfx3SgiSSRcrULyzBJwe9J7+qPLoCKgOwYOnfSx
+scnZA/m7lLeehCDTD6WW8R82PZYPLhpAKVuBlLuuvsku239i13hjwZrvZx4OWk0
m/Ex+71jzVQJosA0O9CHHQoXo5TQNAGAd6/2G9ERkRpk7IBub8Fv0rGDrc8NycbP
U+DdxagmT6wEOUjiWq/yAkxyXL5PDtPxkRDjuxmlU2ciuPyPaDVVaYMfqvROOm0c
jGSebKF1a9TfJGbwW/OSgnxXsjWPdkHpkVit/uXfI6cW/wcmzcpEJRUJfDeI7GJt
ebQf67/k+/Zf8HvLHXzdcK66o3fShjdgFqb4XSCNkKsm5/yYOdaMIISrY/jHkvgg
9kfeGE60Zox2Kc+afgLkwHsjFyeVT/hjI9OBhjG9PSo+b6dCAu1xb5aeTjG4laW6
CG6Zs/HWCLiQU12zX8Fpx70oDpavNgLOK6Dh5N+u82m6gePRj6fnXKEp03Up7Ve+
T8tvi1jZLHW1L5B355/RYLx6Y8vTXMA5OM/w5tu2p7AR+LzxgJ+J5elBLvssP1tD
+XreDIokQybGLPNQwYLfh8RhVGEjpCcHDa+EcGWGFbEON3yB1v/kkC9Nmnlam+Gi
ZlJnN8yi4j93Yvqlt0WfwRwOmC63Q/dPQ60CVf3iF+Am5knUClGC5IE25jkUE2a4
27KVACi5JXoMeemi1uqvVG9/cphS+GdXijfUrhGFmrCDAn6fnb0/3NxCEvAVCksg
sO+abbh6G4ltf+wdGHDV1kuyPeT4b27H4HR0rSU4SxP7Aah3edT9KegRg1ltb04C
WtsWLyvK+J0rFBh16vMnSgN0BiTnLm4QA3f2n5OCru9JYo87Wvw1hOtBifGY4hxX
Rb4auTx8ZDKvUYlYGOGPrv6nqVuubuUdgASXsZqwd9F924VcRTIxuX2bZpcKmemi
XyjeoQ0VMB4hkP6QkOjPLXy9T+9dzueOdkz9C7Y6SVnJ+ppBrmOLvftuN05iA5Nl
XmmRb+aKPV1XEESCmHK6Aarej6LfDtZY++zCwnMYlqP3dZnCoqx5Zpwvy7FIvKly
s8uYoh7Vrn3zNunRXn96GS8sE6bcxSrrCDODqXEI7pagrNBj2q9BIiQcqnFisFHt
Ii4PItozqVjeO7JNTGm9AqnANqswTX4l3Q6h46XCBJDrU8rREWABDqSbNQghhufb
hNSEQTDiHAuHyzSTO+cdC72Vo6cN7yOqRjXmHhiDKuef/p1aQqEZGLBlvzrcfCZS
VROX4AYVSg0hOkNARm8yX9cpPejrT9hgNb+Tiz19prpDRelpLMzUX69OIylcGg7y
NqFMdMVNOjFsnnCWuyGN1Kk1OqFsWoKt+aJD1IN77J2wtBOz6FGHr7NOt9XSx2tY
gm6wl7h6JSCgZX5I/aqrZ4Rkhp4G/r9d1ZJ2nWTfNkn04lERtKQEYL41OhrAn4aY
ySQqBe/d7mSRrfOicnPoqdAdPsxwFfZeT38RLVZeGW1o3epCcoZJ7IBy18Ych437
o/ktSPwANwrBNXaXQZ01BChoS8z4du8jfh++n3WBpTSfgANdSTrHuIDEkUhTUcn1
JRCwPbqTmGnVPsQaJogFsP7SnHV41eh2jRn1pCFZhKoCAE9Xh4eAcWVtZKbo6EVP
uw+RxxtCmJEbWU4shd5fu/B7N/t78ORVkQ81NRSFbDMvjHyejMjuHVY0+bElpwJ1
ozIerdGwX0ZGuueJi4QwxZFg7OAefzYnN702usMz8tl+2f9AYRo5Zl/UaHVW0Trv
TP71+8OeKnzJ1OwjIMxDWr1swIqj8GyY30Pvkjb9jaQSt66FzNivQvPgsDrMtGBa
1S1AwoSCzWDArhU0Z8hH++ZA3HgSEFhRh+uCmTpwc6YPL8ItslLmWIuZcutCPSqc
GM7QKM39A2Y7ym5XkTAJ+jBgk35OAESBly+y/mVE43Xpsb7P2oujE5V+KMF+OY00
Ra9KG+nV3ro77qErKRg6iTnnH8Fzfom4G0+BPvufuZYv09lgIyX5CpPuVfYZDdP5
gR9u0sqlpyw0sjKJwQya490+rWgJ1zk2vqQWN7cJGlyG8PsrJo5QPmsMKPwp6Ayn
YjeXTvaFvN5R4scEEfGi61YPssDYut6t6hNv0P9ptXbKyJGoTH+aKda+Je63zTtB
45tOKLDsj3REJtSDJ0DgSUZwrKfQyjPi+mjyrLblEHkSMTEIu8620dCyLZc1KcxV
fnPiMwoJvqjfXKfNN1J7XvKCuNWUrmWadBllI+BvKg7nGyPICrwhB8kgAjORcD8U
+QMXS+T7uRu3E0G4mgxD5LY8BCLiQAbTssOD5+a3da7CULsJmMu27XHQ4uNOnQ89
7UpfL0X3stOA/yZ99Z8kHypnBWat2e4RGOv7ImP5O+0VMDDqR7VGcugw7nQpfmYk
Ki3DX+B8gRtBNltoY6O5tn8/tIdhdPuIgH2QcAMbwyTYatEFsh8jK3pNwrMMKehz
W4O2SawLQDhj1IWKHNLqZOKDmBXnq4hnWu3dSjGkFYK32EOTNAiyBmKYScV8z+/R
xHu9VGh7Hn8R+W7BT0RCscn2LDoIxOgfl3BGU4nWKdOJ8riF17XPxnyG7ZvRCKZ8
1wsdCssthCynMxcULCcw0PnZN+84jYIYC4rSaDa1DbmW+p4pnL+JVeyD9CgmL/wH
GYEGfdo+2nZ1HT8EKasVoGPAnNTBb+azkvUBz6RZBkB7CAVVgkDEAKXsZDiCtiU5
lNQkgOa4iBufvP5g2yNjs8x92B9Q+88xnqIrXjW1f8/15G71aEOlWmGYDedfa+U4
WlbKxTv3v2s7irRXGQUPSFM3K8Sp+X/m7GBQcgyPjd02Rzc7JCnbUrsRiaFqamKH
E+6de3dtOTxMjsPJjKeWPu2Q+X9TpwuXZ9ig/2XMM4p+Z65qhFuMiUqU9+NZ6F7s
lb5cfKXIZep0oLmi7TIovtJEg8Xn4WcIm1iO5CHt5usUIGic1Nq9vOa1HxnarHZO
f7UObrdLyCy6zHklZ4jWUIS2UdbudALVx0sD97FTX1mUfekjhIeV6LyHaYl1mnVn
CCs7v3HDqJtFuSBIgtUD5VLcMC07l1V+ygB71f3mCE2UkCAMeLUvNiq8tQKAgiqe
qd4WDRfN55I4mx0+P+P8myZ/WYCoUbsWu8ZFQmVvr/XAqx0Slcu/K4IERYWBKveY
8pnLP2/6YFMGWeQqfNOHCMUGlnU8AwnWpVWlu+sp3nY5VmtVDdhrXCnC//4YuuQP
+ox8qsseSvB4YP8T03XW2AgYaxjRAFQ9e0CpqQFbRWxjD5dJ8wBHt9LnxJK/RfTr
myjUG+7lPQBGGWubvuHvMlMmWtRNJR34Hx8WlZKrsATQf7HgWf2L7w7Ow6KTGKxz
Px6t/4yWo+aMZjxqD/WdnJATGecA3A1Y74DEEJNOjaJqpSpHDs4BFFEZPF3xObj/
HvfXGBHaT0H2bNNV5yZocrY7cOfpqX+vK8tfptzIprbrEFPGWAqb6lt5uqgM/4Rs
OksvhaWC8q185LRmKB6rRtytY4GIF8jwNTJ0sBvbU1x27BVZquPMeynFNQxByJxb
tEaCaF7HNXjd4S3Hl9/PdvWlvjbJqTBDYCAiTMDT67EBIVqVY0P5HYf6zFjCXu9c
b7MiZImjTxn+75UmrAmE1OxMoE58W2PaGArCJzaYagtHJkUyBK9otBGj0zHimczQ
ksruVYGbphnngxTUJHio4rZixLWBM9Ee3YC6u7g99qfCXoZDo8Oq6gL0e7x9Tn3q
PkmmmwTzIOX54AzXoHTioclM8R4S5K5Y+QLYicdjKwYsR5azf0miMbaSW85iJALT
Zi2JRxnDvt7YLlP5VdGw4OrR06vY/TMtGJ/Mznnf5MTu0/BYQrM5kZHUTkBOC9r7
bkEoSASTaevN/e0Lw4CgGW8GPRPUqujJt5vpnsFkTEuo/mrjaHlIiRX/s9tSE7+c
TVQagI2uvY1q+Dirc7lkvX3B6mR6Ret9pHb/ceIARPlY7f3GPndRz9Aan0O1A/ox
KDU/He490vpq5d/wKOAmi5nRvDH1cYTmNkQJ9iwH7e1r+mDFHMD7Dd9pdwBRdSkQ
dCwMS0cd+y3pj8pGoXxg2/tX5muKjcw3g9DxbpKAOUtvYNe2sbcSYfpKYY3x0oE0
1KFuoh671S2kxc1/GrnnxatkzkTGaMx5re/KWkjQpWXE0VSz/wGJ9BnRsE0DFI2p
jcsoq8XMl85/5Zsx4ghsLQe391Ro+syUXIjSrMLcuW8cZqHGgxflsPIQklMXrb7O
SV+x9+C6j4l+TfTuLjEOwEQ3Q5Yql7RmT1DZiNiWVd4YzSkc39dMiMDX4/RJwQoe
GXuvZsehuQj/QtWdXs5j+aWF3uiIf1WwkcE0ppTYQk5cPN55yqyYEB8DQgDzwDHl
Qcvqdq5s3qUel27iu03H3w7/HX/cgS7LPL9+uzgSFDXfa6a4p9SriSCEyVGExKTu
9jne0kAUSWYmT5b4FCkJvBb4gb32zKWIkhjmSvuVh62wI1f/9xNPpe02rHQh24J2
brRAitzyNGBhfZ7BvP/vXExD4PklLKi9y68h/5y6T9vIT1XKvFrwT11d45wqVdw/
71rSfW84bOW7fT+N+WRuL0z9TvYg/ueTZZt35k20lWT9eYn0zguBGHNy6WN3nABc
vkQF2SGJQdkXKS6g9Sd5SEWTohuJOE3Xhi99oxKeZGlqpUTHO0IGmMDbL5g44p4d
WeOqrmS/rZ1A4ldCZPPwbdJ5FlYV16jq6116nmPurxAYmnl2oImqaCFz6ldzYUzC
3s6VpR/RtK0tTdxpF4R1Gwf0/T9FEjhz5V9p2zq7vfHiTFTTTauctsaLLZE1V5+S
R9UTHgh2uYBJu+kcgfqimsp5omu/AHJ1mDslXYIyc0qALTvfGofSs3KO2w3iTFBY
aoMu4pXXdGSgTH0vvxNgWEK6WKGnWd7jtP35Gwq90dkMWk9OBAxbRdb6ETbpKPQU
Gb7KwIyFAagrsm6gchUoQDU8gZ+8z0FkDi0C0xBtCgKusVL+1hTZ4iS5mx3JsBqf
cQE9Z/4VnnzPgobuX03cejaSBQv31uEosr+5QQueVx0OovwsIn61paNZ1hqgV/0p
uO7VloBj4urUhlIzz2bDZCB0iOLntvSuAHd7xrLE0WbptYrpUPhMOy34AHWdcBcF
e8eMJXiIbHVKYTcBxCA/BZhqRUlENKCJoDF3HpFpFf3Nmg9+UTFUtqijz+1S6/3n
0Jn/kuE/Q5ETXi68ZofawiZBzO6fHOQNbpIZKBXBc/SftL6A+JCgVRkwrAGxOhCI
tv7VSQ/j72n4AK9gdvzPZclKseN7pZlfFQ/dsmmg+tbH0byL1Mu1nmKoaq35akKY
KuoeHT1idvI/RLYl24FZ3a56YSbATsSkHJ+hdI0pkQZTJyA1wr8gg+uLCxKEledi
frBybuEE9RCiDOK++wwdQYr4E9HJhrR7ckLdCk6syCLy79O4wWMAIsOdt4hCGlIA
qqiYduwF/MSnL/3Bp8WpAqnyrRRZbUC0i3ct9n7yDhekHLKZn2pcjcmy34tsfCjv
p0Yv3EAiD6lIQaYtoPnu9k+XIjeF+P4Fpvxj3o2m2xloFfs24yM0UFiBG3FDtDYP
kgSNbYwoJwt1EeAzDg9LkvbmM8FEPS9I2dr00cHOJiaqCymq9KbUmnUns4Xpw/hh
2vrQbVSLRZs9uN0L8NBA0DHan06fPD8T0JIakYwEY/FAPP2W86n0I3E/BeuSef0X
VsSRut2z+MEZi64AtYvyYq1OzhR6Fs2GzQH+x83l4BCFjJHqpaz5Rda/OqlOosTr
3DnmxQYjIKLUjlDVFZEmnNZP+bXsBOZbXYKoOMBI4b/MSzBm/ldaW+YlAGoiU/Kx
Qor979GFuWfIcyE6v9v9/8Im2Oq3VKO8dMZF4c85Wjo+2tcI3i2F0uHkodmwwd/B
sKF3alz7SLRplTD3GJbeg4Wmbpq0i2gOWDVMkC+0hVJKry3Rfm5A5ZQ4X1V2Rvwh
AlYI7TMn4LFmGAKHpSJhluAyIj7ko9oUMRRHrMkLQZMO++Rxg7++2Ru4UtCHcl7m
v+x8abs//TR+DuUT3Z/itkOOVPs+I90/oFo4+4Z+uvwuenOkwO41lCZtzIMVBIck
B+wKhlrdWPsQt7s+aL9EMWHfYlqUSEozRBivMKtVnec4XqoSiANi+BZwigilS/xZ
3Sodyt6HRmrWqeJadDR4VrpdYeFK6hVgQdNmy/UDAI1TkCUUktM2lsRSD5b6asfO
OhGA1hDdF4r0pUN3vrbhKxXmhuEtgS+xEppNGvCujog99fgVQeN8fdTjpojOLZ/1
ayrNIeFaHGoUatCehXCJTo1WpsaGfKHeM/6/kp4cJREw3f1seEJiP7bkeDGHL7Pv
6zUyncZlIceIVdgzpg/lDp7vRUHEfqsYa24F5AUzGNd2FU56XnkujRGp8hE3vV4c
nkAgZlAyuA10BDXw4IRksiD3dNghDqll/4+WQwpwplXX3jhdre2D7g243xLDrbWK
/N82SmEYigczkE5aaqzim8vXaTrQ6eIdId2wvgRRxWZCRPtOP7ULx0ldqqaNxXRt
b/jyoUn5r8tIm/L+tUjwcdKKnN2K5quV551NcnnlW7/88TX9UkxenK9uzLzX5BJp
uGEHSJKgRe7O7EJVTtMMzmSufVV7Qj/X0DWqKPiVzvgYbR+q03aRuPa0FM72Hu9c
wS+sZx6y4XcEzSCKsKT2A8tFCHErC6mogIemaaG08sJiCv1RSWomW5ns4PN/6tER
y8fiDnHaP9zbtdzmPpX4aykvJdm2ej9a0lJvFjMU0X46WH4hsUZLIg1Mz50Yg7m+
TawGvtE7zrCaAuUqCkcrSuRRrs8NcH/lhwsbBkFno9mJ/lUZt+lN2q5CzVasjz+e
cXuIbFQl3XUHZD2XRTYMiv6XRw1J+nVF0BX2XEJa+9wFMZybMuRDIxMGxWEr0U9A
KHylAjGXKrtv7nPktNaFxpJIE08kYY7PuOGA4NY5eMxZDoafScAe/7X4ULaAXTru
vvSYfncYNyXwQtiBE8rP4DuISjdSN/xWvD/w99UHRGYQx92k+3iIdGS4ZsoCRJ59
yTMjw0L5dtKgn7CzR4bYUSYOtQsmybq4WVE3SEiM/kgid1rTJlHdv9YfZ4cuNZ4M
Ub1Iv/WwWFNAs6AdiMWLX4VCmV3ybc32R9kcMonwLHOlXr7oWTfxRXgYtVuNU2AX
gHikEx2jdNqRIBY+oyKz8NRfs68aOO5Pax3s4GA7BTor3ghjwYTdPsD76K1wYtFT
SivS5xGbxS8MMrtk7LsgeWD8INGnMBXq7amEorouQnKTqZnPY+gEUI58bReNlC46
Wft6VeFa1Y8pkcl8775o77Rkx6RgXJu+OJ7ZXgl0sHbt+Z20fjSpO1IrAFESb4ya
gXTqNDDOKTfU0unEu2S6isrlr0QH9LhgdblW0OtcAZ9cu9lCxWd+T+vgHLBsj8p3
xd2WAiic92S/pGGfdQJ5uMMYQhGt8eCw+VXMjRDCVQJZZCUhCGrzzF+LussGnHhD
HWgKxOiP7+XCiLP4TIU7Uw==
`pragma protect end_protected
