// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MuIgT374nwxjA6tUbxz2S62iWcJOfkkSqW1D5ic8bdywyfIfKVRM68p1fw2J/rwP
miV6EdpIPWc3myatHqZoSzrQby1IFh+/eCOZiEkEKwoTbHAYQjVSQAjPKi7YwSn5
uwN4sJ6s/ApVQhZvu43D+tJyoBvklr0E1uxlQhWWTZE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 38576)
QQbxM5OO0V3OxBS4ZW1YCIVtocKMLtZm0vThEuaiZoXVVeIcfK4aDtVGv7AFCyXU
6EjGEdfIwY5l/Mj7h8X/EmJ2wVWvYY04R57VLibV3oYQlwkgzvFzwFLoG1/4lZhJ
59g7DPGc1gR7aWLjwhWybxSwwNr6RtHYFD6zhYRfnJ13/vY/uSL8UiPJgwxd1kRG
5DyDGdAA/p+J7HUtOyZjevf54uV1vhNysOEi6sVJbiEM1hAQc93QNJqDzRxUV0vz
8KfSogGzmgUTOXS3r8oHzxSVGj9hi4HOh04NUcKhlSpPwslonBrrP6DGz9L0YvMy
oSS0iFDN04bUFuZ5L800kFXGKEw2dU7/M6CV5AzIy0RelNEOYsJmmN0UcM98jSs3
wiD/tEy/AjWD4wesxSCxsmD/HyU1QjE04GGls9dX998nz4a1DLGSrPyJ7MxDhEFy
EU/7RmB//w/FoHlgqiZnTvSJDBrCkfxHtgSSi1ZEPlUVknx1V2QCg/MDH3jZPpAr
P+7dczw1PREaH5HuSfSW+zk7dw1Rc2q0oFq03Sn5LjMIFTrVwCcMgTr4yAnVhA68
O1C/DxLgQEQWNXnF2n+DfreadscxKkd3Ntog8YmsWwvU9/G9mHO/ubhUf94GXYuA
36ASLi7elW6AEW/is4J5sUgN/EeIhwnwq9BQJnXNsQ58xur8PApsmOK2yejtTd9L
z6L+z9DAc/jSlFTCyp9UckDU3+WSuqOPAVZC6UB14y4uSVzKeQXxS31d/6f3zmCq
JYXw/aNIlxh0oFNPkGD5zNTtbM47JAfZg5HSsS7WEmdTKFYY9umR+WYg5orn5q2E
CXLaUa8Eb4jTnZtqGQZxAA3OM6tzbCfHqGHxZ6zIM28umOhYhOyEM/XDBFC7FF/K
xl61INvX5NJKBF5Mn8uCMuLCFytvgovQAJ5NEir5m3ootq4pJo1GQsiNBRuqSnmr
PnDINu/WfXqotliPyeYUSkZQvcoWSLtOAFXWlKrQ+/uSWPCj2V19e0KskF1nnB+Y
7QbE/PlGRuyCG6DSOvXL3Sc3ErRhvcTsR4jiAwx4jD8vIqt2E2QotF1dzQlPlFzs
7yrTBVQxVuq+0kF7wmdzeNTqU711yZKkiYAn+TK2VH+6wmQBsahEs4bSA5gPQJ3g
1oyegWn6+lBE7YoBNFjMQJ+Mg6wIc2UgD5wIyQMpw+pWT/Nd9xjD7STX6rottQsL
3FU953/b7ISofTsrkTnI+57646ToWHR8pw7gFaSCaZjpPqydwKOOfJargMfrdGMt
P70oSLsfAHpK4SxtLr3/jhi6gsbenSCDtAw/hvPIWRE1uPp5mfNgM8JaKOkArDYw
2HvdBWjEisoWF0U0e9QIDKLXmIgEfFQsEbgEn+oXqDwgc8bg9fJ1e5uqTNyFJQik
Zu+gPoM+ecvwRhQYu1eovFxU7Zih1uVfBYLw47GdLTKx/Xk73avsW14NA3/of5qA
K3sD2HuXM+QFx/NFwJzev3DDMos3KWPkZEc1IO/nntk2iJi7V1xU35Wxw4D/J0So
aNvn5ObjRHqdRixpPWw3odJjOQv/vDpBmKXF5HVQzDebX4mjU0ceOfixh5y9hbY8
3rskRgeSG19wC45Y5M0NIvoKxZfixuviBRmqe0QW9mwBAMRP9npOy9YPH4eUMk55
5XmSHgoJa68XAy3SEvOEDpwfJI0DTdZamPWCWCakL3ZfSAahbkRxG3AMvghOlKWA
E73ZfB3KhEhM3t51tx2Pc/hwOmh3IIrPB/b5C2tNXgtk3t44Y3xZZomgPm2SnNhT
sapsk08tgRWZiLCYMwo/qDU+m8N/jMRjPi0AWqYiTFBAwCMHwUF79svAs2or6C5M
M//fAMHB6xVr5cXYN4ezMwyT+f1nmbGxWLDsRBsDu4sgS961LfopIPJXvxEDI+MU
i5dO8XwmU4rzcPydXaHCOboAVur5Xy+ucDk94/o+lYC++/4+qnAEAzaJV7DZeiWP
6otOcOyDgOgCmw49xwpzf1/PN0ot4OB2SA8PuTWYXKVkPK93h77KJEU37UpGc3Ad
0QYSNPNgJzWHoqYq3PN+UlY/xqD5lFnwJ4rLUmKtUDJCQdvEH87cR/gSo+e4DWY/
JMopKG9GSNpShmEbCTXcG/ibOvZ9vNOsr5nvmvdiMCyoB/pgC0WC/xNPZ51f0tLq
ahKovXGZ34L4PW/sgKKLnRGimbV8qzVW6+UEm3p76Hc9/onWAvl3nnnvNYyaK0pk
BnEz/ShZ46Gk64LjvYvgGwXtYKKMwWNKNrtvU404fiisI0aLzC/DnemHFloadRyB
FLyy2yjOrcphY/ZGyjP/y+TVkLRkgpvPxuAlMqZaQsDy+QW0gHoSgChVYbjlrlTd
Is6/KdVUmG+4dk3cICEecXhcLXsKgKxcNF9F6kDCQ5/TdIT3sFFjXcglNVRyN11C
ipos/FeSI1+3lt6YMF6vam0MGfyU2628cfLKAV94+P38QQn7mQZZ+dX/gVkvXJBT
k5MNpH2QagcAyByEOGmUhBEYjNA7M5nkfGxOXWr7bgM/zCvm0vC6IiIT3EHwQFoO
T/ynUw5gsR4xFvHWltqjYdyQaEenUt80F0A/lcoN/2AITRnvSey0w8vGFQdsSAP0
1jzLRz0yiVSTPrEDUP2WyhLtPbn0NoclEqNChDdY3WxDuD3t7xouAqUUj940Yjrm
DCJdu5T8CPvVgUJVMsbj8tAxFPuSnVyNqEPerplVnQM0/VDAg+9V3MN3wUA3yGWu
rfAPiVdAqBKViIKGHJh3aolTP1ykOh69d6AVhMEBT+8b3K6XLNySnHDFr16W044R
S3Kx2LBknZlJB4vf18Db/thZ2EYKHYJ/XioGyMqEWHTPg/1wO7lcrEPPcRR66p4i
IDEYx5SZ8xviHzekFHrSp0luPz4V2MY/pPYEK+BoqKzJQogRwwGs5bfD6EddgZ/L
CDxCDt9yeu5QJjV7DySaPK5XnBtByk6C+eG9hEfT+9DzPz0CBRRolhsnUh3HX1/o
TuUs6CONxNr2iZ1Uog5AGdvp3htfee9ldf0w1NLHpul4A1d9M8kEA5wpg5lNlZ/1
0v5NikhwZ8ZfWiz2Wn9HCl1PAefNE3D4LvA0zNPCh4Ucv43qwtHVVs/ISxayX3zR
xUEvfFCpSg8yJUnhm0dDn3aYObr/DGi/SmsAg1y2w+OwQfpyQZxCpvGmkFQHoNoQ
LpUfFv/JuxMZIAgJ62V9e9xg0k1bJN0ds5eWlmxHFnsBFXrUpWLVohToMq4mFWSP
w3eTXkfsd8W9HIkCEerLFsJ913JAyhbyB46nvqjtoXEd7zx5jmeabcS4x3kRBqug
fPWLnPcbzzNSnrI7V8zYLPoU9jwaeh87ALtc4Eb5NkL/wO4uqUK4z1VDsmsO91w8
GFd0TPKpzojITk+5bVcEW8Uxnwpk1N9ORbZ33wJ6njn6IT1QJz7RaeEmNb9gg7Vb
AS0X0XmKeij+kAVpiyhRc4h0btv1et+CIzLZrgDnQVcH0ZmChrCBycUSWWLIshFa
B4n31FrWmwfhxdeKxuejj575UIlkFRYRvXI4aYeozlGeEP6HxjSpq9y7oadPsyZR
r8lhMPCRvvyE5rItjXfJnZwRFKuHMGK3z1A5Ok6TrqPDAeWe8f5tKrFQvxrIvkW5
49q3LIe3xkhF2px/San2INeiv8Xz+ODFHpz3Cu1TTdW8SpTwR6GIyfsbB5zY4Wrj
sMH2/WNDXVQqFiRJUVXbkdaV4KiG1c8kz3lyeYWEG3yWQegkWRaKDkEAfN89vNmp
ZOC1MCaBfAV6n4Ye9yxH/G6N9n4szveFrC1n+5jJAZJ40z6bpIxbEJrtrtqjD/wm
e191AmV9bF+CxflM4Dqxr9lxK4FDGGraPyzvALtEQY6ADrdeU4M9j3X+xxmoSut/
e2lN9Eox2KoG8YC5aD32oDpHHTsu6jxz86+ruqOo3sZ1ccVXliuz4Mn49ukTcTr/
u9kX5FNRvja9xSfLRf9AbpfxcfKxKws8g6PGS8t/TCbARVnlWDokKAtP3kXabAHe
Hn8l70bDQPnQBGMW93hotUklOsD3ZShHBcEMZ5JyF4/gmqzFBJvJy8exm5lyv0UM
y4uleeMiVkSL6DuFHUqMC/CNdtBjJSwi95OUkALr+fWb2JmZCWM3WIGN7AuScl0/
odPTSIbqCx2yIrstymkeOcwNETNM3vWk9aQuqtYXmHKvoGcC9NCDfL6Rx2GywLx2
KhpPBV+HxhRZ48IfB1aI9MIWFva1y1oi9LsmMbrBe49qWKt4VvomZzp6850ZCUzS
wJzvrhVmhLv2nMLSr9cjOGVQOUEwqUiwkVAeHetOFAl4OYH8V7FPCwNKMb0/d1cs
UJrmdux5J5nGRO6CXVwSJ9B2W+uqnwCfSVBC8tLKNh9NApkwSmLl7RGuOhUtf+/c
ixoPzpG+G3wVesrAOafAdT9hu2rJs3dghwjDG0k2b2H2cgE7lCFfkEUYj2oHtzHX
HEiLD05f29nPIXCHZ6iRhU3YElk1IQvo7VUDEAZQz3pu9X/K9ywublhHa9M/XCXG
936xkHTIVFfdsfWu8fXyGHUNLpO64oHJP7/NKJ67xDEiJJBTg44/At1oQTCOgItv
eohpALRNeuiUFbwdYLh36EO6HSSV1nOMojxPxT/U5kBmCs+PENbjgiN3oQqRCHqK
tdSbQyyZ2fxgThJsXBzYs94r89/1j3GAsj8Juk6Ww9aowgGmYp2+se7vEODfCZ2/
sP5/BdpjgyUHfWHHQM3Lc7E494X046vVee2QlI4QE7ooqRnyo1pRL+Gn7DYu9/Yn
mDWoZRHEx+P3L2ZxsMCjEe2KOybKwmxBlRToWOFSMwSlDRO6QHDfc77nHcE7oLU6
7LL5lDh/GuPSSe0O2oySVV2Z1UEVhWaSUOVbMQ/QA6fD4d/OnfkArnxnIY7TCi7U
lIhxGATb5vZN+Nc502wU5KZYz7kJvpi2q0hwebb14fMZn9scgDtsUTZK6ZFgHiPw
HdSrkyHFkzQfUiGlY5/7ccObIjzLdZLL/qUMA+tVtcfmlROkG1fj+5ZLRflIhxda
xAyHMvv/B3SeZNggx8IXnQdV6P89+oSMpiMjYfnhnYuREafZsmJhmRVARX9ksqXP
4ihJSouDSaYsOmSVtFbg5lXkvtJKxjN79sciWL+fTl997aRI9E93KsUlhwmqcGIM
32Kt1q5WXOGe0WkCvsAaNfeIzCzby4wC2hWgEM1AGyLZYmNZWC9fIHjr/ssrmgIX
wXSIZX2qgaarG+JriNQV8qDetZxCUIz0PnFf5QX3J4WrJP99GGZBj7N6e4UgxlyB
tIIL7y4zVnUU1PhxKpP2HSvzaYOJpwdn0KsL7y1mcDMJW3OiGN8SgMMokdYJSySF
XgJbwReXGcDsKE/6FbgBBr7Y6Ih+rznDFGfdyxTy3B2/9y0aA+/omweeavmMIp/8
Fz6PCapnpTSUPkRr1PKIn5Wz13M+TAsPjgjeiCjC725tiBkxSbCwdUGv6YWxQO/x
lyd9irno1/8h8oSqksZ+PujjJhjy16QizF+W3u3t7QnxrWpCRPoLEFj00fwbZecB
lJSVzCc/JiGtdsUJXT55Oy92rnvDPJEAL9reNE++5n2ivcWv1Ft+cLGxqiZgrKdl
FuctNpDyuC/VfNxKhGMoi4tE3YxLXZxM4mrkhW2p/ZcX3SuvlC+GtwC8sgvv1z0O
hFH5FCzkAo2xjaEldY8jb/AZ9GH3A5ejdtP+4I7EHi/E5ZfoI9cftdTBCNkSwcgl
FuAeYbntvWHdE2bVOvFHDKOavL8DDrp6LI3kTY1NsFR5HK1ouUWYrGa1y+s73d/O
IcMmLimzHo53mE1QLON1OOB/kJ2kelGAygr0bYe0CG3e6QOl+OrIGlvkuW9/YmVe
DLST7Fl21hXQO6G6VLylxVffodSs1s+09GRO/TuJ7KW9C0CbMFkNLZO/OcxTXL5M
B+XTKxJuzbEjqpTujHkOUgehuCdYk/wcsHw16M3BFAZ4foVr2hFBA0n4Hx+v6Mpm
Luxo2Bk5C4fEGHheilPq+J4x9cC+PFSrj0Ubpx8KytGmPnRM2XNJ5tn5VnkxeulC
CEEmSDnr1kUFlVZFkY/YaeWKeeVhfXgQt0aBA3Ogk1JdUZhnkABsiYR61n956COa
OklCsPBOn+HlLbDdDeAHvegx2/eNfv/JNRcB1Jn1bd58Q6NhuQ+hjr+6w2SfgxwT
XFH3624vfDgmrTU6JafbOLTycukvRVnaddKgTG0xjJIS7VVr3tblyTC1tnh592Vx
awmJV724hxI+Rz7eea92W/XPpx5byNrLCOvWma8lFimZjATRq4lKz4njdl+E2pbT
g8f/v7Oxb0Dn+h2VDEAe+bKySiVcKy11hYmc/him7Tj0Cmk/DuRVakONNbQCo1Wa
kPy/sOYvjdtuHrJ0FGSs6q5+MWKWfM8sVERyFf5nt3326BfUV/tVqMpRDwmqiYJD
43RH4UxEfVQlzWIxjDRKFMK8qq95gAzftV0/KSzBY/v5w4KrnvuGNAGWVMXVEalx
w5cF6Y40b/ewjKQMKgBwuCNe44t0rR4JXQqidvAh0X08XcdK7FlCgfB55P8EcmGL
ZiKo6Jk7lzLIoyHdp9c6xj/jeX1D8uLYFYZO8vXVdP9mJ0pVfboVvxUmQaWHZ/WE
oJlyD3f9Z0fLGlyfiDqTNoxnYEr1r/KriqNWkgyKRH3+uL9c8Y0lreHYvudMceiS
EPsho+Sm2RKRGnNg2u3zI4DQ9JdEr33yKr3msIwdaXVAalz9d5uAAIAXF7npg9+d
9JV2R6eNeHiGf71VeJ0YcCZyiB68GK2Fy/anhHLRaw9/JQTpBmlaxqEGpU/rBqZq
OM5HBPrGSHjQa+8VwRZRQ/Ro3eHKlADnQsSiwiVn+7hFrsRGwR8Dzp2smRTHuyZM
6jLGt54yZh+FceZDO1ng+sPt/p25f3uLGqPknphgInRhIVfyaE6CO9V3AofWCt0M
ZCUcQlfpZgYRP2umaCauiqVrLn+7HB7vS5gdHKElAXDws6jtcdYLCr7aX2/mOCf/
X7baycENjQIO4iSlCvjF1U/xKhUHGQMfl1zdqOMuyiAxx9ni0/HNlSpyeVzNGEvk
qRKm0+vtZDzmPsKzaSuEGy7AMEdb6GaMu+hz4LI2HdrAdZe5RTNdQVkA90HF2hwa
C/wH3yJmVUiqNO/mVvQrYGhlbWPP2AVRZmfgtc27qmnFEvnm/oU9o0/uuSnGdhtP
GleqPltni22nMf74PGYlFeiaquv/a8lmYlhnnpqr5ekKLHM1HD1op5WYCNE3Y7/d
RIohGnma7pO4DYACzno1PkRW1O5ZMhk44OqaGIcksp/uL2e83PiGAzMEDQG95sow
7zB+o9h39lrYiWJlxOhGuc0dX2Je0Vmo1P1KM/BqBnan5+D258vFOAnvNo2F29gH
zcGe91qKy2sRjZPO+g+ZfeBo+Wwin+bVJaFeMbCTj6pwuyAuMsIYE1KXtKxaM0XB
TY9FbZQmkXJaw18xtwwWPdNdpYdefTHgsNPbgu96/D/thehzp6TRngLaL5sS9X8R
+EzfuvS7SUEO4m7i+pGmzkdVBkN9GpK/slDgfEHr+EtTfoufAVeXzhV+Sw72G27f
FCH+fI/enFnehGbDEhGfRgHdnmvt4DOwUog3D2tDToyLS0PP+kGmUh5VLpw3nUe3
XgTKbOnJNo3ZaP/2u4Pu/qQiY7Cx4hWUHoCRNSjKXG9RWtV/9WuXrRLCvH9aO8j8
gMIeblLS4GdBTLDivisfUltzvQokEVbG3p9emWu3iZjC5PYvGYeqB2M3loZNTIxS
Ze8gZNi60dFZO5WXDOr/wE6qdHEUfha64gx8sSmCzsmWJTycSMyTLgI0O8C7EX5d
cRfKjDXZPxA5VG4iHFl2KoJ33MFI1GlEaJQdRg/iL2ExKLhf+XgXKE/dZd+kh5lb
B06Rvu43a6C3+ILC+uLsCBb5ulRRIBRDe4QDfI8mgUqsPbFc3A3sa+NYm9vn6/wP
7ukfr1Vj6NVUSZ9nPoKIbIOI+Aq4XALFOAFDD4sN/GnwII9JQbfhbBcJ/sLkg/Pl
YVEu9OreM4dcvttFMJXfaI9bGjV0KRUoCWWKegyzjHlN1nv1xRbNiD8FhK6UPAUD
YCiz8qh9RSChwqEfqAgIZjD1678V95RZzyyJcqdBluCyXfALHl+ko7QVQ75Iw1+T
4DGNRm7rA8jol1Ctxd3D5XFSQczT7WxwaGg4RpiNqYzTAY/y5LHsQlhNm6YaqI5l
rY/0IDnrBRmAGwuuV4cMAklfTzZxKw+3hvqskWaWqzp/AEphmYL7k2gv8ae8i4E2
bjZgtwWYa71A7NmapGDPhulIJrK6eDUxYHBsOYqe1movrlKH0elyB5WujAfPTs1C
PYrFEjXGfROxbRvIwNSJKWX0aD3aGXG1f4ajWDsUrQiFSP1KjM46nrHFSG5XaeQM
k9MpwvfsT5VOa62KDeodgxWzPL71a3/J/DL4fScq0bU5eXcMUQmNTisQzcWYlOte
ictkl8WJpgqE84f1nT9x4Qy9sPJOJpVEa6k413PrIJQXqy3gWz1Vxmt6GYaiXNWR
whFyAElID0OflYyB+f+F0KKWomSvx2ZSHlRb9+PPMQj0iXX67oPctLZT45KtCVkA
6XxUeNcV+lMUPPN7DtjFlfptYVYwyYXY8jzXKLOmzFouE6olCtoSAJofOhOaORls
arEaiRz554uVh4IV99c9o4ruKv4WjUD50MhgiHqUYsLvi1oyyFqbeQIk3SHVl6W4
u+bisybIf8qeFYsqbcrZuVoBCv0+0Lb6cAKMvDoesXxJlJA48uk9Nxw/U0dln8QN
iMoaSj8zFTdZMVjCsjA2+I6tMn0KGhXPeWx6azNMn/dSCtFeGLbWB41uG1ntkZSe
2Ly8OBYOzaPKl4H3xIVdl+zF8VOdIT0vW5x9HI63pHP1huCbG+VpZNgVu+PR1HEK
LlEaUrVKUXGD6DQvQcIHoY1vEdRWXyengoFuObXlzXUttpu07ZXj/UorSfbfFQSb
G8oJfePRTDsXbFFrPqV4ortkkcawQd9NXVZZ8dIUMg08DOIQ28TRUGLfVzjpRlQ8
EIN9YjJCcqFbBPnQORJ7gELHPWLGEHy5a2HlgwfLkflRcZWtpXfvqUPSeDIOv7BR
Wmov3PDeuPrJAGUQm6HRgwVuY+JYsMGkKheM1J0t/VljVhro0oWKpKtpUwnuSsY9
h+QHvtULbSG/c/qTDlYkFS6Hs8GK5Wysx6YvhPJjxaFeybEDjonM8fvuJ3dWge0U
2b4sBCUOHpwDL9gM/nWi0iDaNFuTt3YUt7lhb5crlTOTO8znfWeDru3exSkyHIBU
tlt99E+J5FfO5XDAtWjdNqwUlhj6e0DKP0Zl4zfirW0PMkvtwmwbPTvbrPjtD947
auGxvxZGXbDGQ/ql0JoUM9NSwhKnCnXYYYheEj1qe9U3i1ELO+Epw/BqqgylYRG3
77kEhDhhkN3o6MYIzeAk+KuB33/8FBFRrw8lWmD7WaXcoYb1kMQBRm1TPX6sK/xA
s+fYgF/U9NPKKU+cSgFkS2Rk95NxqB6+tiKIzEVJxEhU3GSDeejRuKWbbVNcIJQO
VAzK9PTbwsjB8W9JfLX6kJ/UfDLXLzdIHBkNj05JL64TB1YFSdI9dyDEDVYyqST6
rrGFdxbCSmbxCOcOm7aHTQn/0Pl0fJty/aAHRCoQBT3KTCyEqXtWEOtjsm/grolX
0wVUxhzNEeQxX40jQJrFnoLk0Br1n7gF9mzDNnxOfNs08CcCJ/4XdoMEIcrKNBn4
pnvkP1tn4Lgez+vAS0SXXXsNL3kmers2FJjdKZJ4wp9vx/DtEPE3kXBzLFkKhkax
WMZWM3vjXA+RRbwDaRUsOhIsfBVIGnVwrNfajwQ8noMf/ReNlw2p4+dCblv6W/9T
tS88dHhq13amivNot6S05Oy8NKkdVWQQ9RfSjM0dqiE1qHfDgjz1QOvvZ6av6tiw
EmDaUsS1LeZ5yk2qnknmApDR3atDVT/RJy7ZssgwH647RH1b+CDvWZ46AlHGTgMH
PRwylA6UajOGjMWX/LVAaEiVPcEQFVjYCu2IVpv+PyHJqpAVGH3GfywdVCgLoyy1
jsb2IrFo56Z4BxsbbyP5PNal/wK90R1SCozbNNchjAzLzh3G94utlFzcl31rj0bQ
FxzUQGiaTXXZdmigsB2mIiVjDPFgUmAWp2lp2dNdaUTtQ4UCRGOuZqzVfHhslScJ
mqWqNNSGolmZGTVscjWy6k1ljDzY0pQHH4QJPYvlycblaWUzl75PCuuerKdFHsGC
+6AkM05I4ifzJDASzS+cExXWPZKDs4Cj0BFY4BXNosD7rro7/IDnScivxkozyP5u
TwWiCILlkAfxFDjofOqgNDX3BUKN28fYOXOFzmH7ipDhG9tDB5dWzqWTeLrQtaLh
7u0sILs3RgDYagLySyyoRdCwnF1FFl8sf98OvvPxBU1SaUi4OMg2aJ7QY5tAW01J
jKpEAljaHjJz/24Vrf7yix6+3uO3FchNKMdhbM3RVfV9gy2qIs6hZemi5dLU4wOE
JGY736VdVTqFmhDHrg8MnTtLEzwXaIWieijlJqWuOM//wfrQ1mJ45svBQ9SPHMG5
7maZ6weaLxGZB3bUSGBy93YSJ2hZw9xEXUA9F3SONkPgybqa2/Jx11Ehaik9uBqe
F4qOZEUlqxmr9rkwYNGERUdF+bu5wGblLh9Ua1jaolZ7etuR/R0HFUhY6JtczB4b
viMID2aaNAa9lE1XkpWYXDFTOJEfRIK/mTDQJOmuDOOsUYZgR2ZB6xbGdYYY8uDS
5/DJIfciDygshlgjfV+Gg81QuECKGploYYYea98noAXVDpzqwM375Q/OdvJRg6iD
lsGnP/PkiNM5H3tWsgfu0dDJQSuSp7AY4IZiKIUkYwSKRKNC7XK8JcpgSZ7OL363
AQbZ/R4zOg9D372M69G2TBrghfw8CZyZhKrN8tT3CBa4d+9HXB1cX1gpkLwGmnof
mIfaY8idjCTYNTmxbfIKl7uLniRIG0WiQr3grA+jFGdHTadckFniI8x062uT1EoZ
FuLVlSQHggWEJU+i6DkfyMqzQgpRn/2LGeM5//GR0sPZTIYhEFjaYlbN2cMdGJoh
CchWdzvlkl7zZD/UqokRsgpk/hcVLtMkefJlo2NxjnbTdRSAojhxBSWXGCZFIAaN
36dRfEnqhhIzNiYWiSRuoSdH965htIYi3iGAEX0S8B4Eab38EugVWEoeiVHRQ+FE
29tKRbSk7e4PuYdg/8oe91lr2tBjV1k+QaVC2HHW1IBUVPG8xoGUExUhykdfysRo
BOvCnTyrx1Kimfp3+7KvlJRJsCn1uzuEJ4IYg0AODFnibtcM+S2CNTDdp5Ud0BYD
oAO+KVG9sB4MQpJ8pBYa1ete1khIfYKyEV7Rn9J6WvFUQ70QQlJtmi+TEwGMJOlY
KFdIEx1aYOu6jioaAhhWQJ1KLbqXXkBIcm43KfiDbPmSymy4j6BCOpJwCW9j5Y0b
BmVaAKlq21y54f37EHOl1GKunf22a3pVtqsglcReX0WsRx96WZFDKdo4oSk0f/IC
/Ht1xJiZbVTCmTAT6xfehD04h4w++zIIBrI2JTacKECPzfM25Hjs/dwcV/NgTelj
PkutMQQbVYzwLQrzQD782FTO7uUQC22BQdH427ZYRYvADSZj/X9eQsK/8kW9CJf3
W1c2oy9/z6XY3QexGLFJve6v7MSOmKdMGGa0nZBtrqLG+SX9VfNQrkBnJcmc0Eyc
ddJHkBDs3Xbzjg9D9z8kxN2q5ZljyjyS5rukmqPJlIbQA9y2WtKtpiWAN/kUQVsf
FNRpG56qo8lfoxsxl4rw1xVWXQ0Vs7mUuNh/bzTh5fnodk/Ig1RhY2/ExFR5IxwS
1uUxf6CX8aHT79oEtt5ZdBdPa1QL+vRBjdAkbvPkk7PWBZpqOgDwciOoa+YvLqH8
/GaecZCO0tVIqyi+NsUkt7a3VlIy+szM+nAx8+gO4A2cRASRBzQoJcLbW+58NxWk
mQrCPCQ0gzdDK2NTXb+5wabg4WCw9kdDejrgjpcS8hXj8oIecbRqmT/6LlP/O0Nb
sg7CpcYF/2heoDQ8cQaLz3+4LGgM8MXefsL02X1/K24BboW8d2hoD2+0Fk9q/LGr
wSJFgXOic5c7pRv8Bdi6IT1CB9uPt4u7TSaKIxk82RY4VnuLO26jj8JmFVYVsNRm
d9aLoTjNpwLEj3GvpLjzH1h3gzkCNCBfJkt3p5L2w1NixOX0Q+/TAQhPunPkU8H6
cyN/oohv75FLqjdBgl+A7h47Pjk4o6EdmR6NctJqGKOloZ7/Y2EmpKDJk9ycVCO5
j7fFnvUdl5kPl6sHGsbcqC/8q1YB9fqoBS8ixxdJC+XicggkBGZHDepy/rD5ix82
svZE8Yj21ad9wgdt8yzIkDMwX7EcnNHFdszR4XQ43Y5X1j0U5mHQZIRgb28IF9HP
/D871xh711MKPaZITBRutBN8ioP3BCLW1SDM6FrLLEl1Lr40BtsvpA/4qbP8W9QL
t/bT4pbtMsHTrGfAZXx0d2LpnjyiS/oe7Ic20ru+1DWOaWIqNja2ZuyDNweeKSyq
ikpA+50CQ/xB2NKi+4KPSLfE/JyQA+y9tvnxeE+Jh0m4ZvEr2gSCRYVNEY5FTbkl
yYEbFqxxofO9Trs4v5D9mAfbW7WTyJCgCZQIDlrm6Os9KiT1+THl+SNfqZfrvoEn
EN9Lq2Op3m7NeXTUHOY14dwhidhGwbWA4s7DGQTNXq4mcv1tx2ISYfKlGFtMRfIT
cl4gHLUa1uE5z9TFBsn26d+Q5gkhKpayOoWg9Th4UTg7bWNDdbr4kSe+RX02tQT3
oCsm9tgyQKNPFXP7boCQAiGa19fqpj5HBZpvyCBiB2ZDQuhkDXTgAArjP2yGKJ2E
4gIyzsyWbWHVjahkSAhOdzIjKRtjSDKrPzUtie3bsC6yjOGgL/K5aD7XWRp3Iyhh
0ok7fmW93yuxQovD+bvu8L9O8lRuHwVJbrhBBj3Cnwu9dkOjm0mql8lYkcjSKrtm
JJY8t3loVDXf2jXLYLvwT4EAUwY3FsZrwJ2NoSpBp+un80dVT0yccKjAnTJnLauq
cxJfHvmo33tYicEcIX30SPVlH1Z8V1R4fB03/YiXJardCPDUQBmhdwq4b+NE2Ug8
HXtcdm2rX9XCqcyo9J8x2k+rKQdok5kL0GNWxCiBnEC2IpditJXJaPx31kJNHrVo
ZyVe08rtn5JPnFn5gsirxMfbnNv0XZ5qcLt9XxBYRQPKAnyVHipqgmU6Jxu8ZzLI
yFR8KnT5EqC6loRZuT+aets7o1ZRG/tt2nAkwixHs/nyRj8gx9cfD55JU2QmXiqR
TVf3aCpz5vkzk7EU4AQb0VL6CP7x0D22wajuoTGl8pq87y7tGHK7CbLvM6chJzSa
orJr09suYXJQnWdYG7uoCqc+XYuj43N/O39jCLqNdgu6PYgCaXHql+BwwrTtCHGo
/DaKkJ5ipK/YYCHElUPpudCK2F+mPbwsKfnPwl18LJnrk2JAX4SQROACocdxrZZG
mFqsLiPOZcW/MhvcRX/JCClttgEnTSH7Ov1BQC0SG4e4POYU4eTXtDI5XNiwyUtI
X14spesFbDJdnvvCZOyuAw3oBOjmmeWa3ip6WbKGGpTiaWUigf0OyA5Mma8z0bLm
Vgyyj8yNEgUJVoTHf3Wfw74kUkN0SRTx3uulDYSeujAMcgtduDEP85jT/XmhleJ+
R88aHA2CgHn5fsCIIm6t3kVqXHovfg+HcywfEXDyhcPup+R41or7Nftjc+gJIO/1
Tb8PozNCVlRX3uqpzoZ65hVbJwGjzBSFAJAtU356zSlFXSQ8aaQdIiQ8nWpqL7md
79kKmlvmqfXur6ufpgIJQe/6V9BO6iM4V4mTxPzvKkC0osypBZBDiFbmb4VTpFwe
YgPHov/6seSVamgtG4QpEG00JYCA792Yy4mJ8AWWDomKnFCzgoiDLYgc824jFYHm
/7Cql+UibVQ7ekjtdioaaZQGMejWqUEVCkYhZYTlJTThlmkB9ElkKTG0z/ZAydll
BjAKXmRN9StrnA/UGuYJX5+qYKkXUhcW3vbJ1RPGdgn5LPxPZyyCj89Cn9FC/WWK
/orVjaM8nUKKx4R0vqeZpzYaj6Qf4QGkCUDqdt5SYjp5+mIHfpF36C5R6QygKjEp
tCabU0oGgkjCWmPAIXkmjy/8/QC7vkFuvjzKxmNU14l0lJsxO3jSVpL+kitCAF7j
/dMD3GSCyI1Y/TGcF6SuJg3H4LPv+AwqxYwM6nqW7EGOhlBkaAK1Y3uGXle74W3K
6iXjeOFeAWHU2crHBElZUXmX0dz8VsuTpKJ1QzO/z9ATaJK+Z/cmRB1XTBeb7SUm
7lFOtOWzHzz5nPHMBOKgEI94xhBDrFAmMNhJH6uCbCWxc1Z0McHWUep082CVIxI/
qNtazMMgdQB6x/HZzhOFducyN39/2xwxGJyo3zjPnu9Xms7LJxJezATqhv42krlZ
Yt0CLUKVPCbpmSal0oAi+WOEen+q70EwgnyA+57VKgHFw4baqOPRmoqfBR9KFs5W
59Kev3/5UnCayVRTquFGVNZGe8F/xz37R0GGx39Kn3yLl2S2IXX5waR3OnGjc18C
ruixSAv9kNgVnXVfF4/v/0WYN5w/aNVhTSM0GKUrbP6NLp8l0Y8wVkD/sWZ/VtV/
fLLOCVe7nA6npw3hoXjs63rS/K5zk+A3qmC0VYrL72+gka5lvuky1vMIf7eZqciR
3wL3YApanLvkimU6KufT5VokhzmW40Z7hi/tFI+umD7BVwUr6zmoSlVPl77wbWG5
o9ewSwT9ygsrzUfzKpk7780OfdO9shAVGIMK868zPxrD6RX07+4k8LwUHN2J87JT
uCp1Ex7EmPsJzVdu6i0/fIrc8Q5Z3ijrUPuWtlPxhRMAizb3E7/6DJo7LE+HbCEH
ZPYYzGu70U1Vm7Qm7yN8/HqEiNzlrC05Ej7RnlbHpNUXvCCw+T5NOZ/v4hqZfNWC
YNPJgJ5RCvI4AQlYtLV/mQZDCBY7XS861leNtZkN5LVSNnEceabCkR/BylzvzIHf
Snk6Jh3vpke8vQT2QJNvBsY/g7f+0uY9MCKFW31CtX2VhzgWzLPfESZAsNueZRNP
HHV2D+uubjumjww/2nc0Bt/5+N1tN/qzOCcDU474f+lVa/pZ0QcXc94eJa+4Hu0r
MemOBbZPOzKCIRb69sNsvwetYVI8MDVKFYkm2HtZhHRFEGUphK7Ao4Sp1foQNNf3
3dr0oUhNw7D88ssEiL3NS9RSNiE4iPmxPhHtIv+mFqQzR5y9JsJ5+B7CQ7jsOv8W
JWPZFGuZfDmFEwkqlV5uvpQBEkIHouUWnTQb4b7+K7WUOgmw6BxDioPPH98ZPJOr
QQIDEnIlXlX4oC6M5nEgYnYEH1efVKT+mRkKJl7862Bpj+Cs7y3at7LRcO2gnQ4H
Rnz9e7dGTqJtEBR8PL7W9umA/fzkBYReZEckC7W4Zct9454F1Jv7SLWlTc9jIPz4
ZSHX/+WZ1EhQE6thnSMZde4EMXnCcZeB5cN3n3nLR6MUuciV3EYk7KmJgK+CSvV+
ufxQSmjIlaFXFRhtnC2X0+jOJQbS8kUiHo9Z9ISSZoeb5QkOE9CV6wI0y7RRNlxM
8nlgUUayISFKJ9uuk+4ZBIgcmZE00VV1wCgM2y/ZHUgnFuw3sPyrjxUnQs8d6l1N
xkH23z0iqUGahzl9lpAbGalupIvDFrthOnDpx1EDKBaFvh9mUPiWdTAFx7zzxkvq
Cv4dLnFyUnBiOlk1sAebTzkisFdLuXFpxzkWOwYGLNtZzN4snI93JNctQY+GPnV0
fv2Pl+pZMAw3SpjHZxei0BMu3Q1bbVCyGYcQfhQCoD5c2/2Bxfw2WO5WNrD8dY46
I+8RJCbN4IlYxkhbUoBqRtJeLOPTg0ZpUSYStDoi6ebeqWb8ovNiUBFFQEWtiwd0
w3WUR+DFHJPEUJLbq4EWbfNBIjfLtcLy01D81IdGoWhb+w2KjHLfnK6+Epdoqq12
/6CXXI9A96aGikeCHGnbv3YvdTshkAAlVl8R4uMhp/ZKmxp8WcJTllfNEANNXB/G
USSG614j308WfMzew9I7HUEC8lflwELya23iIRIs5jgzibi7tkClxp/SahoU1T5D
vSrakBgRv07BrAjy1zT6ZZk5AniaQOY4u+I6IB2xEVD7yhQ6Xol9a/CMyp7fpjV1
DMPUDNxmpecD0Wr9WDAeGCS03kZuMHcIqT00kZmV13LIe9bd56dZBHvLFnKyfUTG
pMdc8WvuX1H1dtsBk/Z5Hl3ZG/cW58cGpcI2B3vjrpFS92R/4a9HPtQrG5+1l0fQ
OPzdm6L2oHyJ7CU3r7WlLPdJsInqyVEjArW0osiEUhVflp+IBSahZlm33eda0nau
8dIxwkQOZOSiInDwl8r+ow9Er0k9d7mHG5TEe0xSGzV9wOLk637LFaGXEgmAnlQH
Ntqs74cMK1ZzswRaZiFNSW6+FDacEV4jieUdlkd8/3DJA65WX5mjXuXV+64kmOwm
caD8NVjEzB03Mq3y80eL+GU53fgau7TDhJA0CKYApTTzvLti8WEZ8XB4vduXfmmk
6JvByQ/bX2QmVHSM086BvXXjm9AYDHFG3S6rWD3IzJbhKD6ubSB90Ce8FdwY6aT1
wne5dwRBfsPLBi1S+2gLyZ7jDx8uZTDc7YdFKC3aQe33I1xOe5BOD61PAns3j4YQ
Qi6Odxr1vnNgZzzdMEcEWMhvJfttt/mnCldWwQqkwzbl8f6PXVBnERCkxUbpuvnq
AzfBl0EIpwBMLLEu78QwRhyLsJ/+R60U+IDLm4i3WxVwhKS+gLfyM+e1R0eAZh6s
hHA+MutwI5omUpnib/QbsSbOkTD8A2az5Bpiuka+HQnxMiCv+/YjLyFENF2yLAnA
zfHSKhtrZmt1JHtQpwjlHUGfrseUdqB+8D99CymR7omdxoVoMXrlgzzitQN8FrrV
s24cclwvmxwygKBG1jSOm+5Gm8aB/yJlTXp97/1azLLmh4QWOizPdSXa6hm2ddKz
CwdY4zDmwEU3omtmLBpa6LudtLFf4j1yhVk5/WaVG6yOCkq0co/Jk2+8FMMgMROt
90cPZbxFLMtU5YJUvhcsmC1Iqe9KYwYZNCk+2ewdZXYRtgM3VIa5z1WaTUg5Py4J
iPpDvinID/HYmfP57KPLXJotvZcxbxxQYMQBH5fQfWgTK+5IzdxhsE6bFrwkT9IE
080VmH45c8sH5e9FFtV8v4v3QDHgqtUq4bo/YY2Fj2zSmowpgYPRFZ6YFEb0RmCa
4R9tbo0lGNfwh1aXgHTAJK0lixwYApmUWcvGsvD5MDShzGvybVBdd08PNdQaV1Jt
6JlHvsqi52PP9esFwX97l5AoXcPCvDSxbdXV1RCrtPG5bJr8LhU1gK5yMa9BB6tN
ZwSjP7C0dv2rsV++MkkNjwM1YKegGtQFM3W1S0s6R5Gjoxph+4q5M3Qrq7CIbRx2
3F+tusIrzYRLR5tHqqmpt9Das4v8eR3pWI6+r8CgjRL+Q/bc4lVdANzjMIqmrpuN
3XLz8WoX/Hn25c9xidBiYJDBKaYIMCSd2PDV9TCK5T/3oiNvaP0+eoz+/BAhnYAD
hKJTdL0Zf+BjvSdQZPtrct04k7aSmAfy0M3TNRaI4FQC5Tyc+2L7XOygMUijTU5F
8WQZNz95JkNLDZ1rdlfcs3te+IiUiZaxyH99/6U6efxLUw8ApChWAU41pCYhV5s4
thQbsbF2KRnbGcyI8nuX7v2PFdr56qSOM/m8BLbEDIqO1c+Pb9tqVmw+ivYfSg0V
YiJQGkSUBLETQkfA5Yp2+u5HpS9LGzQLeBUKiDLA6shVlMPlbRnGXnNUsGBbSeU/
Fnnr7nrupEmKycFyBiQIO75ZqT7vW67a00a53eo/Hwr++8pR4Oz2hCw5yQX24wZ5
paatRzUHLFfWMZUojqFSh00Bg2BqsKSztiiMt0Q4JfMsVZupAzuv/8CadIkML9SR
Jk3a0PytZHFn6edgvxOYacYrN/8XS+y8hNDO8+G5IaOJ3cXXiKRiA8GPrfg2wJgb
xAe/GwywkX8rQVowQWhRJxTEawezs6c5pAyqg+rcpr9og6beBXIQP+bJrda+bONv
HGD9cxVwn2F6ZFFIq6t0L+3Q3Xhy8dY5mTfmtN2j10c7IgJbg0Px7CruhkcYziId
pPu+vQck+k0FhLEp2Qi0HtSC3Xf7Eu/UU+xGoN3PFZ0smahAeBq+3cRbkWkCpp3W
cLaqZq6Oyo4qyGrxzFpXxWxGUVqd6kNR2ilkDFN8B7xb8qQGPxfgsnWEOIg2NII0
9mtoTFxRlltJ81BjUkneW6AFt645L/dyN9mkYqSWuO3m8SF/yUOpJfPnOx4qpk2Y
6Fpjy7oDT6w33QjqOtlDZrQRUmWsW7Le1Kb0TlN0OMovAZYnO5joolLda1sOlfDi
JKlzMo+MFJjlh+pamvZChgevFaeF7nRoQtI0yycFiqvAevdPdFNvRbjGhSuEZQrr
XQ/p6bUYio2YtvVZe9rGejaBEIsAOQF0rtBg/y3OuVfuenp2Z5uemckpbNSRwuls
EQ3WfGdlaFXa5poCVRdr1XXjk7uN0L2Iahd6ltHmnUjgub3IUL8Wi3mQhMgAYCmx
jC3gCIfdjm3IB+P36SPQT1v+MNMFA+6AjdbQcF9St6Ud/QV9x+pET18d6WXpcMAP
WkHwb1IOl8vQFLZd9uneIUVqYw3dhyvVBNJgKutGTNB44h49uwnOSD6gr5NVyI+J
b5SMVjUiz3zQOJXrJuYR6nl65652wYHgjyrPk0llw/vBDBfzFYoarulNFcCstxJB
sxgfS2qMPV+qAJH17yLWJwtlSiVM9dehfy8MgdSXcJ6tc4mXAKXK7I43yq0cNHKg
xqUTXka6nYFhuAxI94lSB7cPm3yLO4GxLPar3NGSn5D9irk7pFuDIAYO1Ip41Tuc
0/437qQN/US9O9RYbXakTv5WG5N1p9X7NzWbitFB7PGnxOQcuvnKTYkS4MXwPcd3
/qggPy+7vqj6n6GLD7OH0kHlPHD2TsJ+LL/qEwe67xOOqBL9SKGSaEpbgZByfuAm
Vp4znu1FmT8bCzL0BBsISKkISBpzsl5CdCFzYG6+CGiuX6NZrV+fA0FWuIN/SYCS
4J8fqreDgVKuuAGyk+UEXyPWV6VFu0l5xYWQo91jcYcOwagPqQ8zUvtR1xdhflhf
/+JR7aEv7BM7vocTawX0ahV9VZsbvPoIDO3OtvV+ZFTJT8KdV/MwgPDShPFapPMs
bmDAAPe4XkABsrPWJ+qZjxsXE+RnPoU7ruTi39jG61Om8NppVXhnUH9DXLpRfng8
+IaLRzR79QbcPJ3y+exVP2ZDtqF4OC1cyytzPDxAPewzjb6I+KxFuxLbAnZoJoiK
9BfrmZCNbR6abJ7WLlxf4nUQPZ4aASpRVORZtLqlDAC08TiSj3yBQLsd8zy9og5f
8ZBuYLBx/O371xao3uZHEm/YGCLZSptFT3b7Kgjrh/2p1frZFVHPxjgQGycCJtoZ
FDSi4WR0Fyle0YZDrIwSkjxB8O5J/f4hKmelENieLx1Y9r4SN5pZkmMnsrZSgMFE
81odc1hm8AbW0zvnEzvkUO5aTyTNvG/oNsFR2H1bZ7npbLg+vR3aPFEMdPGeKEDa
jodI4FtplOV4+TQ1KG4hJSIT3lnM/dD/eQaprXnDgu5HRVzbjTIs3TlnYHPcLW3Q
R0EVT+LFfvjJWnnv6s9bR55rsto+Ok1wcOaPgteITUDi3itPRqgJw3/NP87HfuND
k64ktNoxES0W4Yf4FLgcVfC2XiLKSGl7D6BmZC1K+T5XDMSKQoKFNNosnyMW/mmv
OM3Nr6k+4PCKWeduQwjsQHdD5RruHExeWKL2B/rTGLCWrZoPfPOBEWK8Z2R1QsDj
9gZFsaHceeq3Vxa7Mv3hS808BMZA14OkMzujCW+0UaNz0FzUg61cbOJdqcYAJmD+
Mpy8cNEaAVcW9utk/knk1hzpypPxupuiy31jWHUFeZjQ8zfs4dg2YIp1Ve1/YP7f
i9WXddP5AwJ56X3owj1fQcQdNT4fvEB5h3tRWUNb5/T1yvITbBSXu7zxswS0jf4I
q/q3H+BIyNgV1VM5BwIU+e89mMFxREzeG1C5jfmpgZstEG0TWgvqCWSCpqanRKB7
aSUNm0bUTNaZDxtKN1r5yBz2/L6mBn1NM2wnvJC4t33iAs0m/0wNS7lCJbOaXeJf
Ua/x6lN+KUIePP8yWD+fcmK4Fa1EIrDnJqhWVewGsCWLPtZtgDq1ttGjjuJTY/06
P7xH0yzJAB2LVDlh6StJ6GFD/8s+DHfQRkZaeoaNr2N8MfY29wzpSa16uRmLzgk5
gB0uNXMa6AFkEjDj304NOay50pV8iqYxOGnSaaPD1kZecfXP/aLMXDjSOeK3QfAf
+X8EzPw32QNTK4mIQVCsEmzRjfmMn/hlR/5KSCvCZCaM+86YSmntT2eB9jbRvHIQ
FEbdc58F/RAqb18x8l2GnRkWxaht/uUK6vCOhDZMJR5sHNw8lTl0uQ/yQHnI3AGS
bjvpbQcR3OcckcFXHxoZ8pkc/CexW/AMjEj84sFyqRMZzf0moOJQorHcli6R4bG0
KK6FXg/1VmZ1wAZF10y8Y0UyTYEB0ciBCI6S4ULvNvqE6KYURX3q9JABUU6VpL6y
8dWjDCo+Bn+FoAMaZCfFefiN+TJiRDYZKR9eSu69rmhuOzTheRiLAWlCvLA8uzu3
1rk4XAKtCNCYbpt1b/3wL2a7hNGgYC5kqgOtBCkMJ8cQjrv/FwX2hK2Oe3arcV+9
m03VIdRKcTH/PdJbUKw2WgSRqf+q9am4U/pZrqGDUHf9W2t9A1IzirxSBoCOfksT
Kc9rWT6LOMg0XkbcJWeVEz9w5/KI2OqlLVKi9FCBMtml8IKdioZBfRQXaIRoHKuR
Xs+erJr0tuzdUKHjYD0n+3AmUGpMEvl+bArqc/+Xg7K9B4ad3rhrub7n6rn+OpCx
zmZlnbnfJAqoQZduuMwPAtt4X4aVdRf5KZkMg/r7zmbi4Fbqp1KgMQROz9iiY9hx
VGjZZLUUg6yEE3kcAV8gl+gfQM5l372S5csi1CVDcInD7U5Vi90YZYz/5PAlELyd
gWR/g4Achyam48vv2WA/tnHHy/EXKmL3PEaXsx3ThSGCQV25qVxOEN9SkpsHphO3
q9jnwL0vD8gbuzN9SU327WDOHKE6cBVrnLaqTN+Cfd9/LOc9DHy6s/yDUQ7HaMcO
tdIIfecMWhKzOKUTn7kAqJy0+5M+ytqsYF2zo1K1ooU4Jf5G9ttnsH5q4yCpa7TW
Wl1ng0WjQtAQp4Sg/zkd16cBBEwbnvsCQU+WmJfgCEnZUrcN3sCLjgesjliYlvkq
7t7BGz/2f60av2zYdYW4bU3mNhZSrRTK8X+/twXEVqRkr4TscenaJvkFfaGDqZpz
PK/JKIL2HLwxSS1QRoQGoDw328CGXa09+d65+bTF7fb4cLBCKKSXWQHilAqhRfqE
zx/MF5/8Fxn+0GCmoHU20d3q0mU56ZydDyF7hO65SksCxybkHPnT/UTw7WYQ8ocZ
VNGx7mV3PyoXcUCW1dQuYOaSXbjXkIG4QY7QpSKuyLDtH7WEHG1Pldxf8lWM46B6
8x9czyUafGNvDW1bYwfMR9NV62qRrdR9M1G9K8s0kD6MzXsf96xgLhFoiEK2YFG7
ouWpf5NKOMkesavi4Bzl2jmyWU+jTBa4lazrpnZThN7BimKfpkCd09bgXy5wNZMb
uwfm5vw9kVL1aDZRtsPxXF455HYIkW8IcdDu5LN1Mq/SbW1QOKfKybyRfTlZCkNC
cuABNayOI8myOYYxEVOGBBwIrZUKqDlQIABQ5XmSNVtoxyHLZUazBmseokKI+H5v
CaOhoPIuOfbQdPRtxwANmV56xf41TZBnu0zyop/fIPCshh+mGmrF7yt8sMrO8382
cDCMbyzeFjkTfBwT/gJr4LLWtVoE1nTLWdS//PBI6w4RH4XNg5lDNMXVenfflXOa
fr7fb2AJAEAm02NF4p/mqAK9p7OQ7PyqDdKeeMJDSxmRaUhc+tHKYIIKnHqHexsC
HK1GgbYJPAr8htzeWacOFaPX5u6d9CSHHQAMy+tYjlnmPfuVfUYDy3IKuGerQbkV
HxghOfquLXtgF69Km0Iw55An5taGXkN1SLVTSr4QwFANRNZ0RdGcKsJ6ILZ28x1T
QRV6aDHWXGnbOUZQ5TWwhejlLS2Tl7NB6XOYlfC3VhNNXSXGkWW+JaGwTogJHzad
LWT9oonC0N65D/UF+x63HYWPnbL7V1JLK+Ao71UI1l4Zymw69cy44+PwEE+1zWke
UIyehzl69ugsbK/TksFRf5DDrdyEF8vRs8msLQmBot41eIfsLwJ4667c3CuQRD1y
WlXa2LV9uLeunv2MDhoHHeLfXXcBoK5ci5zaj4ZUAVFqWWH6TWZ81Vv9kFP66UOh
3A1pd8lBLy4YCaqvOV3Br1ahMJZZfaB2neql0pU7fJmt3eqtNETzz8+gSLfD5pQM
bLQYe8bO6Ozhvq/ivQPQsFM0wjIi51io0FBqmrixkUNwcUCWFjPOX84BgdWU3YCN
TYhhaIw2Ym/k8wkDXVPAZU67h1IInOCHbJV9+OIVIrQf29hVdw0Q4wz1Ef0eQWgX
49+f/xiQ+olmCSsS3e1xHxeJIrex58k0M50jKX2nUfm/ve0PaitDDLj/pQo3zOpZ
cmNqTuGLyuKVW7EpJMIqM0LptaFC/jyElOJFzZehRpayFTK1N93iYC9LsXiocS3V
ysleEP2W+P0XYlY5dJxdNubrQ5hI1Y5vbFVhSMpWROolHbdFyv6Yea8mWaJQqqcI
9NUL6UNtzmHb9/ZAIgOuuTzZDMqICtoFXi1mUAbIHJS7hO8sgeTnMBiP8h0Bxsid
ePA5OVoqt7nvqmpLMl6X77JlZLEFvysBEoAZfRrmGSyoGJQh7uWjcDgtVmuxmLjU
mnbw6he6/pOdl7bhjqqKfrTYo6rWQf5fKQfUavIPEsdFIXA8Cyzdrj6fdvVb+BLf
LqK+RM841aFsb6dmuLTILPob40zziUzL7eltFXu9wLZahZNQAH3gOrdAm39anAI4
aIUaDruzBuNyswiVBu8yCiW0FHzNnsqbgtNufzv8YI2+nEK6wY2dCrW+pbvJVW9W
Zyg8BhI1YkNZgxXGhq4XPnY+34iFlTj2kNsczLpmW4WkynPWBzoJO8moRhqh48IN
l2OXSkD9uwFMVjxmebosdx4I6Li+eESjIyWq4DTigPfW3ZRaBA8JptXDAAGWFPCQ
3RKXEyjJb21HZOuydEqk8mZQVjZ8H7DIapKCEPYaMpc/KrM/b/HyiGKpjWRpYD21
BOfy4RLTYKivcWsFg8ur598lq/Naug9icAIa3lr4F8URQkynz/nmc7AWBm3jsvDX
Lkckqpe/709kQKvt3l81KZJYqaj07KJOMbQhUANzUhHi31116gsAu3f/Srjswvia
rNZDPNUmE0PWqc7UDFuLTvnqGOxal0CGqEKAvktGrrCVDdhuzlyTu7nkVa/ohifz
rHoOFvitlJvjHJZVydnA8Ef/VphK2GMzYYmlDig/OhrFSqGN342CT4R6eOBQbKKa
Ot+xbriK2SMbxne9/YnAK/oL82KXdvHnQyXrb2hL6tVkieHiyVLXfBF3iDn/qG3j
EqrBbIJWN66PESjBJAyC7uVdMZFPIpfTWSQXY/bkdAq4h2uN9+HEh6PzS4rnhgZR
Af6vNxeTK4GG/uMRXT1OQKTDwFDrbRm3lrfzKGztHyb+AF8lH3qbEmSSpw0Ea8hE
SSgfDNDH7gNUDqj8Xdj2sD12iibSZleBS0ZvNGWoVg2SORFwSEXYA6olr9tQWQ5X
qp+6IkwKlcG2UTTG5bNhbauHoZZCwVtloKP8naiZZM68FS1hRtcBjc23qlOiRorx
uYcRYBEAOXqiaL/I9J+IhbpT12vayiwI8LJQORRJfbdQ3Mmc7vnpb119NOEqx/b5
lXqBG4acvDovtBCu4Ne/p+D3Z5sHDoMWBT/dsiqJlbrdPacNvmWmGlnDkzJVdW4q
TeNMqzCOIOBaaO440oJgmdJHIKPBpkS+ZAFPnvjmO+f5EvxF5q9IdgX8DXFPMfn1
Rb9UqhoKBIGh9vnLeXjvcukPPWTWczAhNO8dIMJ98yV5gOAZuegFKWkLV1SkVQcL
P+eSdZIsp4lrcLt73rFAzrSvVs5rJRDoVPo+/0eLEFSsrzYX9U+2T1l+ilFpqJ1H
+D2EuASXmavwybmFTTFZftDEQiFNBE5MPyZ2/QgNH/xPyDmO6eLnGnQC7Mc5NTmh
wVSGtbCG7EL86Ag0BiIv9vlhQjgF7V6/YAL04MLiiiah9dD5vyIC0liKNt/ArXEw
K4bJyrEaFBEYcBdTdJPycHObw9RHGH+IUm2diMqPnQeDaBSdO+B7rEF0UWpgDEHT
8Z79JKRjX6lkhHgAsKZaBbROANccY0knCvUAktYfLPPBkwe2r94hofvtKDJiD/np
6qFN2RkwICYGiCJk4vGi6hV9Qv4Hv6UZvCKr+Lq+iwLK697VIKwweZiJEIuP34ay
2DufM2M9iF+qOkKkVBsCTfROsapQkG1+KCnPSMXF9/WE3t/O3PY8M3D/jVJ94MqQ
8OOeJ/aopNUiLDYJYPx+LtvDNjWjbrLPde2LYJRuwlgI9LMzBirsScHisbZuUPjX
4BgspNbpOVp/AVMAF2c0uB20eaarhmHGeXeDPaIWEw+LTSUrZuZhNhmYmXZGFcjc
zSbuNND3w1ag7OEsF6y6O9mMWYahtPPUuSrsBQCOPHKLuWEB3I19Rl9/WESQdUg1
+8sj4NFRIqSXBXj69U1CMnNpbsKDK6b3mmIse3sgqUBcD8KDR1Ppaq2Z51RvwLN0
sT+/atpljzSvPB0iVjIywxU4HU0JJALXw1ch5Sl4eF3758ri1qW/jiTrEpylZkHm
rLLHXms8L238WePrV2raYMPPtCK99RdECSOhBPB07g3H4sqhmzd5D+RdoOFIA89A
oQGzVia5JJthigkRCZVKDEQpz4ZIEZBhEzsazaXqSB50/FTJnbWoFHFL9h5yIqGR
BsKzYP3ti+s/Qyh17gUIAdQdwvCoACzh4qln4cfwK2yC/Mm9G/IpFlNxlKhoCnBU
dE5DM1ufWN86EYE98jh8u6yRtH0Ks5e+6l24t6tvqa/9/d5DJQ+lf5TynOf7rauV
VXpzDD2FMvFrJABfCtuMr67bsPO9e9vmEuZZWXKeZHAYjwidj5+4IXQ3wQJvGVZ9
n0oJFBvHNmI2fsVk9E7JH0pWXxITD55QKQmJaOrfFwPaIHS1K435xRxp1lWGB7qm
u+YW2atrQB5/eePj69t2CGxL/AnvTrXAtnAxAS7uBB1ivpny8YqHHLan3oBjlTyV
fvL9lZ4zH+UurIZpQwqW+Zp+Ck9mDKoJJmkWD5xPZAGBVDfB3b+RgmAy5VVNCg2Q
DkMcmXeaww7te4NUpy/Q8i0L9eDzoHM8PtnmXbfCuQ7qUWYF+E5HOgCAZSZMz6Yw
DJVjtoRcAFnPIuFqJEIFPrFAxWzHWYj+4biTuEh5W1Zw1QFWUl2KTM8a9gJaIm/f
m1txMIIjKFgYmp5IEH3effYaQ17+/yI49MnnIBOO/UIaeqxDXE9psEfSqKUjq5XP
3QVzYiSYG0uCmOS7bl8XsaYQORy16v6GkA4/pwEM1ja6Eg9lzS8M+DEQ3LBh4Uhj
6vntNizYA8Qupf5tQ+ZmJGZ1YYFxOqxW7KSOrOpyc1pExoOg94BJwTlvwilXCtuy
ewqpcFNgpV+Fj+czmg1n6ZezvinyueOS5R22L4Mwh4C7albNToN7STnzbSXP6MOm
dAYYoqQ/9IxgGxEM9n+V7j9Z6niKfR4YZZnssU3f5rg08hdxM+S2H1Oez9KKrLbD
cpysYLMmQH6C4qNIhddsavrly+MJPH1B7HKxZEJosRk2fKK187oYk6Tar/gk8cce
As0pbRhC7Lx+fIc/mVgLHN72DRxVoe9vzRt6pBNPqs6pf2rrTanGrmIXr7zgEtL/
ulO+S5fvY/cG8TUZSAlrmCWa+ktNJgZSJNueV31jgFCfgyLNvYvbdm/1zSiyHB+v
c1CJJ/cfBYPAvr9Zdrjza4Xk/t1ZFwocUYWMpbmauVJ6HJsg5kNaHKb10VAxjCqQ
y8f7EgJIUYix96cJaZi96IN3RBOynlWDgd3iFJOHprZMo6+dSmoGMhg0nG7OUEHt
F1WsZU9QzYbg6DV4spK3EQwmLoYIHJJGLPJ6MzlQCW47JYbFzS9qwKGukMhvO5lY
e9nCJA/PSgRcbT+SSwVcc4VbX/kCok7bcoN9JLGEbT1ONWB0fIfwSLvn11nsaPXV
aBUAFIK55pStwLOBARm3toY3Z+cUVBPY5eGW9U6tmWsekaXBbugeohsCxkqeVZA9
je1nZi0G3PgrG8PwvixmFpNrEE+0T1HgER/BJWAdHtgBXe6UgFzZCCbdRZRUe3PY
mA5TAWW+bYqy2BODeQqJ1qub+DBtGeBfGZy6Y0MWr9JHZCiU0POVW6QnfWMbeekq
rD0sIj1N1PDOg6V/zZm7tTVL78miXp7SxGB5ELl9Sutgc2EWquY7sO0ruusnf5RO
LXx3Kxgkes7TeGvvhuCSQHwZjW7kHwIQ6ycD42tiNUpABzll7rK3Midlk6Ofl7ys
VdyVZOhTr6Agr4E2u7uVl1c0EeIztkZ9Fph8unaRltQ3RX81ChbhoYIlG7uaE14u
PUAzHC7nZjRDxXNuiXjyWWup65EFGVJAAJOPsRy7P6IDD/z2pX/mJ5Z5ZMx9igc7
A6j+GGaaCLNhVm+CysElRHQWxMVe1TmvgnlLBVB/7FEq5tri5eJMVpiTxSsh2lER
eF+08PbWmNh9OAYBo2JnWZRSn2P2oIQQSAEYxfKLtuI5K0OkgaFGgdwJ3UQeM1Hk
SPPB3sqyKyX6ski1xPMIDnms6rwOxXZYktlxjpOuUEQfJxfGP6Nzq5SkRRK9Ozql
DixC/QpRkxxcZ7eWH5oLtwX+uKk7halzD/F5eYEpi+1EjyRF6cgGnLSOkeBM1qla
9B/f8U3d1K5aVyFYjNYO5AYw8//uXc+46Ub4GPEQIODy6bHm9VhcuZ7XOfik115I
SZNMA76cbbqrpe1AzwAzQXO9lV7ZiHd0lCA2la6FqaECXYSoIuWBVoDchuLOMkNX
rktMB76gLwbAN8qyJbyiQ5JrgzqCDRWcLnrpUwUjCq43GjYF84AD2AdGVsa8YU8R
SSN/87tX3exRsN5UtCHW2O53P9cUGXQBqB0f+wW56Vf4UWPji37LBOPCn1Gi8aSL
s2V43TWIcUXgLMy/vrrcWPSjOtzWR4cCu0YTxhwVhOWzKFz64Xt6OofzwQUrPkQb
xgS0iqQlalNbRfdQkAhCaFVJWbyNN58h5vXY6ryquj5zrQZ+vWLnOHFZ82XrDN67
cYYYF5gr17e5yF0GUUmOi/25wvqzuKZ517OxH/aKHICV9TC5FmNsHS3NxsX5XeEP
LcTZY1uSNbKt/rlsJN2JCcye3HKgGpvUyJX23zB54WbWl/3413ZZJfRwpUp5lzqZ
3WRcNNorMPRKBtSOe+E3RPK7IqgdZTjEYXXaWnkieS4VCGpMG6EwE3vJ9XNwoCpI
PgEqIAJdck/9znhK0UkI3E1/V3IwUB3E6Dd0uHRgNKcjjSTDqwIYeGsrItE+BkDc
/40/187n8oc9x1Vqp2CFTBSr5Wzk6BHysd0R0YmM+7vDCsyVtCQ0IIIlOUbb9kfA
cnD9vxF2ND54r+AT7SXnfPRbGJzWA6MwpN5q41AcUR1q5p51eEXSnkhZd5+rvoe0
vdpvg9SigdmcmNcwz+lOST2qy3PSqWdozFKljeOSE/9BO7F9/3X1vtWQdCoCDdlD
e0NPUBlaZy8WPuHWB+hrTAC1s1GaS4PIE5CzGzugfUVaP5rS/XxGg4KERjsA2frZ
8hfPgc2Yk3ymTNxYOKd7dn6hed7D+gd9CXAgwWkT9iFvrKUHLPK3xWMywCPcP+kH
j2LsAql4ftJI7Qe3MjyxjRM02NU/nNsSYfzEFlY24YHMIeR8r5RDt3W/Ywq6J2Qe
iYeg31CVCa89K0xpRxHlkaVWpSn1a/yLbdfgn9mu6HFPqbruSbpCJPKpi54ZVLqJ
C6WZSx/rUZTb11xUbIANu/IHSWKVECqJL8JPBq6LYuVNJpFI1zqkkZlr6UZKzhcQ
A2kPZ+Qv+fJiAWo/X4RHjqxyVg6QoW1Qb4qrXOIOSNvo3YU/YvgAtrTvTEo36a+E
5XS2pyD0ywsv5cLXSskTmN0nsw6hRf2CWK3sz+D3C8VTLEcReTeuJk+INgRcSfF4
Kj6VojLcn/iI4pPmFLck1eXn25182N/WqO9U0wnDBUrGg27XtJjiKHXFiLX8Xljy
+Blf4Iaxzx+rKYS+tuWuytaLZ4QpQqnQm+q2zHIsrH515XWX3UgjvQr+VxzrpkYK
glRxKyqjB5jpSWPDViFfdAjsnlDooFKAdsbYvQK24VHmLEjfBFw/nR3XdSxbSNCk
8NTugLZLXv4t8zjOlnVuQMgH12xItGFN8neGHmhBvU+nhHhT/gZhWjPP3Q44Q3MG
e+ZPuuwRVzg2Alp7cmH7GZl+/EnRB5Aiy1JLI1DmYiWEZpbrjfba1xhujhxaTkNI
CyQGFUWTBMcx2ou/zeNtx/RHh6EhQgEk9++nG3+31f/lZ1IzfUczcVWRpQBP0oHE
WkPKI2TjkmytSgptdwgoAnvYrvRpU92G3jEkqHcboUaw1NdR49oVxqzN8uwmZEhJ
AZtI3d0MDWF6scmSWzpfcXxG5CcKlUwrQ7fKHQfJr09W2fH+B7ezBwZPJ1MmrVEU
WJ/teuux8FmUXR3SpgY1G3Tsv+VI4+vtq/2NCe12dj165z+EZ6Fr7SQiNQmL546W
CSOv9au1iWBVHmJ08ojtSjzYPJZEPj3qg8ho8sz33vokZGqHi2vjqwFXhWuAf0Df
g0yJGAX7exMBXuHz1mLraVunZeh6iliyAHeL70TbZSkOVQOt/Vzj0kcIaeEvJqa4
H6EcB8hHEVNHIgk1UR6Q2ZQ1T+gKUnlBtREfJhfTU/kfgyWvWj3JKAVgKYasYocA
ZmIsbNd+L1edOuodNu2cLWkGF26jxoOxA5/f8l/8bmM9NhJ3nwDYHd+aRjVM2PIw
Rc3FkEnmOZF/TXwf/eki2BMRVYSv+djtZ010q4cAci1VOxlPmkRw+O2zB8kvStgs
yBdatmDZwqHlfah7jC08sgd2mSZpvqUirPIFeme0XrnmEcmjqJrH8eh3/Rd2tD6u
MptRhWK5WSRqKA0xBqPiahMNswEVc0W7Nezy36PsrKXt4CAu4vuac3C6xgekjbYp
N2JKwXLudP9kP2K8hBdgKl1RO/LnPo7krK6AhAmaXTzWizvwFqSa/iyPvY4dTahs
Z2N1NefLknhCek3V5FKhhID12HeVKhXt6S3ISC7Alx6aUxW5TqrzOieaqVXG7I/w
39JdpnQm+GP+6vu1aZytSa8cwSLGyviBC68u9dWc4IFkuTNRPW/knhmJo2oyBPUr
vBMviwRHz0HMP7bR62yY6q1lD/spf0eD710nKQ1OA6uJzDSvmZOSs7ABxpFb+dEA
5s3JUxt1hMeT+6FVKQHhjmhIVPEGMCH73ZViPZytOFUh9SpSnbouc+EHzm1r4KCs
PfeT01TkOOZ8c3t4J9fCcoqYaUdA+Fp7HeLuTxB5XHa5K4l5tmYGboRP7GCa/Xil
6OgqdtIDLUMj0K4BNGKWurHhVVyA1anEGgU/mc9/zZm9aw6XrgLpBp7CtGynCQdW
mALfpB3GMWUafQ+2vnMOZ7dYFj4sqHLgYBOP8ShY8J8J0j4AV2QF+dJAnoX6WT+F
P58IJ4O8RCRRZewKM5ozcpYDrREXYC52TtoKrcR7iW1cjXtuFF8WPawFYNVzZB8G
m6461LWnpJH7Oy+UBUNxIpaBGcXHTTIJzDZLgTjTn9HKGgBsXIau3XM1oJfSjzty
1KEc6rzhmZP86o871MAmTCVKtxT8OyeuCnRoWXB0gIM2fdGvxudVUIw4UEl3q7/C
55vX9LGTwDHWPmVMmVrbtcSzlzgRPmXMGgFRdEMaATHOTftdF+6dFnqANbfg7C9g
/8XLhciokjNIFqS1p2cg0Kjaoio+lApWhMrI3v2x3u8UxWrIlakQeJ49BqgErt11
VlcNUuJAXi09UzUePZEHLwIRmJ2PGiVJbPl5i1LFvBLU+g7rD7RnOC7bdiF/rQzR
Opr+aHXXdTOPQWCtewAk4TONTdNpQwHiEFAvE98bbSaohcpKYvDH6sAZTJhCijzK
QBXl97mBSFqNmgKhdNXc08bvb8wQo6YIL2bdSWVIE722JHajPdac0ZglolzdxB57
amuv4Z2FnrIF3VSoAUIzQUp5P8BrYl+4OqFtTkaslxyUdwasngCWvoibdILn7Edc
q9H4+iPCrWvB1xfYqoIyS6xqIq5IQYO1ePGNdRzKF/KSyjvbocnPFt0VLDljQSBo
gelEsDN/MXgEhTFN7lbisnfKTktVDbujd3YKTVoIKDNNNxf8y670qzbLvbHxd3NS
pZNjJ1SHxGJUvJB0aR7mPZ14KwDUoWl8WeS50YhpBTTbMg9B7GQ67d3TPp4YyMmZ
TvL5K21SP52w8jvjrnueB5zXvbopBgflQVr7R//Tx84IW2+CPAPvh1FePDjmaTts
Ec+o92GxbX2vicoKVbBm7RQxRfoz08nMrYbjs2Gx/TyrHMn7BHOBhDuYNtCOAcbb
CQAPPYDPgnCoDt9NhUXUUks/miwAaXz3YPS7DWt/8dfEZhhKfaWhg29RMG1mvGOS
tBSs8HM0i7SOzAeIia1Utudwnw9nUyeRmlAN9ZTML4rVINn+kalJwOjArSopeg1L
9kcIlwQ1g3MJky6/vyea/wWsFDKalWxNd2P80vTxailjx4U3LR+qmJC3Ovj/j1f7
WRxk6wJPHKj221ALEIUnx8V7i1D/zidlPokWddDHwgAFk1Ua5234EwBB8GBYd5vr
DIhfyZZsF9WQrroSu/Hxk9Z8IbQXJEIzfU3/mp0PElJKa3CDRcSg6m43X75qTbCd
CTvXmHrVkyjpfYoAXA6Izh62qdnOVBt5ZJAfhiXepafLQTxYmII3ezWbXjfC7pu6
lj2RQtfHpy7nuEnoXeODCR5RwTD5e4yIhLB4zWF6RZGYykAuAjv2UjFv/q2XU7tx
JCYWiRvDdtGeiBkAPwbxXoQNqNR1CBZD5aGohsVU3Xa3Z0b4TsBe7X042rxLLaF/
naLnMWuTeOetcwdxLRGYd2IbQu1w++KCs3KPN5+ubNJYNSW6VG84MolX8aBRylQY
MSBr7obuJ4GgJuYluTcr4aW4AeYdzmgydEoSTx+qJbnAQsY4v9Fr8IOwaCEcwlUr
rtZN1ZkJJzShC1xv/R7c9/lFEDOuckkMovF+Y+yqFgWtSk5sq5VQKw7hL10JFvox
9GtLvYP8dG7oIgUSVey7NQ7jfic+Pe0paRC2l8WVBmJlY5ND1gooTHP6+LcmirvM
Ofm80FGtJV/n/Bil8TDn9w5G3aSrVWLmZBqb3iIlLLNE9JJIWRUJ09+vKNxVuFYL
wlR8G+RA3jNsa6ywLvKldHsomgDOmZxzjp+lcs0cayIgVi1SJpdJScdCvPoNZ7vR
3JmQTCL0fTVYrNHFxaBZDkLvVIYYnH1ms34HyS+PMn/hpxCl2PLK+xGcAimhsBao
umj72m2Fb0h8CvCUhkGe2Xm1pOhhhnI1a11wPmB1lmvYPN9wgzGA6kcShQ+XsPCp
TXer7XiyJBKkzO5Z8sD3TVjUdoeVPG3xHDYrqfg3dYL42CXzG447FgJKuuxC4BSI
lJXD9PuSfPnHrNcfPWpaGajSxnQkTIr3nrSNqo9opu9BdEo8msdWOhVGEdG0eIRB
aQJK8f8lFZpS12GYn2ndNA8T57VW+Lu5rupeXUSUyaNEZmE5//bzCn2thevoJfij
2PGqEYFXx00hD/qjlgS0I7ELWX4R62/CsupvSGj1Uev+4uXwTm6xcpzLXi9i9O1j
93te/vzQNvzux5CKTZmp/+tkb+rwB+LFs3CWO+hLxrOsxWTSBBe2iSduMxv6CDOs
y4Ot+sIy0trHKJwsofyEV0l8xjKgytVos6rrK3AlfEGL9hlPLgdxE82cGr2KTMjw
3xo4ZshaFZz4nVlo4JMcfRZRT3bwh5ZK8iruBsxhCNnChAfmQqTBgjHGGHV7V2A8
P0Bx1R/XgNVhBEZGeFj4FHgGZE5Yw4Rb0XXwJsTafOSZ2mAgWUn5yHYAFkaVS8wD
VVhDkVyXyRZ/ct13jEafnf2dZzlq5Fgyao3qgBovwLD07d5Q/Hj89qU+dTeRayy2
hcAW9Riw6uYGcp8n1qQGXsO00/HgkJWdoPpojXsgSRZO6yZ0dTbvwxveeI2M9MXQ
ROJ5UU2LqA+NKRwHtLgGxbAN+wJG+HWWe+UawLA4rHaxF/GlhSAP4E5fE9z1VTnk
v++sD4ORJ/3GSCFoeVvhZXg5ibGglmOhrTw6whaeK3bpp99NJ8GTaK8Urt22b8Gs
PQdJUhYoxIG4Yybx57H12gJQ+jOOFsxjFo20RMTL+u9PH9egwfC2eIqwyvstt2qE
j42X3phgfg9zfI1Wkx7kDcDk/1Eh/mTD1bbBKuFKv78+8cUqQ1Ydq664mvT1srwv
TsxPLO/n8GW8XnBtGut6gbD5q2plQLJ5rvG9G1XckywWd8mcfhaGxbFvLg/fyw54
SYGYCOXJ1xHB9dPsEzQ6awVCBHatlq48E9BV30DAkpCV61u9c/nlkVGwOgdOhPxW
rBroas3M+PVpixq0zTOcGiimDj0oGM9lf8PPOgH3EmMUzUgrfcJ+bo/isNgn6Ctp
eD2aEYpwtQmrcXd1G842AdHZp4qal0ycva8dRFlGuATZe9XIkVThlITVKQWc2mRj
5+hiu3jNvpcArTSYw9qERZAetnaHECYt2hEIHu+K2dbmicljipOO5rbrZhAcEVP7
a6aTNBtHUA7yFwHpND83y/BI3i5wL+O6/+vs2V+qvz5vrnhhwfBxVIyzyamlgK5B
6Fqgf7WxjQlBvKycPiaY4avFgM9yCyWZBLO1dGY5xkBSakojdBGrPzm7U8ytZYCX
itjyrQRab9bF3VdlLjI//z/ZRr4jtKfreC0rTmeiGFGLjSyKEd7ZHRUgEe7HFnfe
gR5Hmy+h/mkrzZHgiMbbGbLvgfoRDauRYPShnYOOLZCjzHonaaA0Nby9RzT3mYIx
8n20H8shAXOt+u+zLKfy/HIHHD1r4iDbjdaa1OdssEuKjkvp2nOXXIbYCp8udgJ+
tVHOtV1QbEJwamFpd1CifwWlWPjoB6bhViOEaZCKXP7e2HX4yzUSXEWD9v6egXiS
ck/4YpI05WB1vQwNzgq7lPMNpIF97bnn/hU6IbNNnM6/o1rhOj5y6fshykoWPgc6
7gN/JeFmF9ObyHgGOoVArALBzTV4Szo71r7grM6/074OsQSzgDxGLHwFch+zqkk8
yKcbm7YObAlQkWymHQlkeDMCsVXd83p5O0f6qdygS+MVReFCwbPnjMhZ3gsxZ4O+
2/iafv1YmSxGlWVHoI37b7gIeeH/CboZec+k0H2/fe94BPc+bALv6EpfSE3EjjvT
rPjl8kTv1NtVj84BDKDnsKlmwk1ndqHWZw41re1D04S77ai4HcPn/FLCCD7tkQ3m
S5uuZpUmvjTq5wKIcxLIof2vZ+MQ78vr6Ze4utXNrkXgOBZnAX2q3G07rc5fewid
rqTH5XMszF1bXHEM82jOXU+hUfOXl5Z9YWrvF9S5h/Y51ibzg+g31id4lHRovnnq
i5oIP6Es0Lqlzd4sd7pVmwIRdPH6CHZj9cPbVwUYEm1w40isbRM6Ky2Rwi/fIkj2
6oE1JXlm6T1SGDBHvCIPOU1/w7uTwKf7ySrzj16cwmD7JnrNN39QKxPx+xkJIien
8S2EfG1U2A7+ktdsBAyn9EdfdkYShmrz/kRkRxoYmeoh/PwurDvqhmRTmlvf++ZA
3nMRra7cu7oR+9nOFqMcSc4NV2XnKBM8xbPaeLpNcNbBgezEFJjrtHwMaWzcQsge
pmC8np+Ru0UoTewtLiNcaFaS9FP2T3cWlmYr+ZSSFxliDeDbjAMN8tvfykV6L4Yc
hIuv0ReHDuLdNVsUSGcUsT4wPenNsM7n36AW4BQbTRI/IsyRF2e0stwzOXco1N9J
Ig1IuxqLABOeUOigiCimxlK2TKptW0tNXYmq3hJ3BMGyTM3qslhOueP2oGiDIBsP
sFlcIcjdJrQawsh9pmoSh9Ge6GDg8RtDeL5022zKFo3GE9Gcyket+QTTpkUF1wFX
xR7+ckp6un6KruR3nV3nU6L6rsHofMkPgV7nJMCyvNrOEp6Mu9PvFVH9c2++rHZ8
d9fxfqlmmL68goxwGEAk4QoznAZcbn+3r14f9qL5XSetpeSVV5stQoaGJ71p9sdG
90N9GJ/IuhtD+S10YA4TYyNf9avGTks7016cUsK1iFkocWpC6fDzupgh4cV4hHAY
NPoof/oRLqlvN4hOem5RoK+QodlarGUoMPmNJ31Y3AqE7+Iin8AVIKD0hYP+XWWv
lnhMwU78sCA3A1oTMzS/VyjlNFKb9SoeaQ09wHnZSIZDIFzM/upHVHSepxnUMQvq
mClhlYrQM7C4kms37ROQzGm01mYgK9jUq20DUcQSj+4l00otZ/uTmj3scKr3Q+yg
iCQ7mTf73sCeDHx81srUVbzTXLA0xx5mNdtBdX6AfH8DUj4FkHxPkENjkTCu7/RL
0W0WnM1Cl1Dq37dbPQF/w2oJfepoJFyhCQcbbQuCXjkIFUkKVXlHXSVE8cnovGfO
LGSDv9ixX5IsL5bvH13knPX5SOGpir/8YbcGZIAIbruwsAFL/jNbaGvIGKk1Q25f
4hFJAGOVt66LPkT20LbqQn4ZNinDn23wFgC3+6doB/C/8qaC3nG+QsNjvQjC2YEi
3jMwWXNXL5aAhOggPzXa61JlKgTMncUJxFrDXU438CG+qB5obcBSddUFqRzrBtVa
Wf0DzE0yvN5kkppFYI6anlLX/g8HW2lrZubPl0MacD6Jat1D4z0HNM28RG3jDJ6F
RVTUEu0VnDTJelBqYFwXt3oryOHlb8PQkijIMhWl+ciWmkB7GheqJOaw+6t9RoyB
FtJNdOCWl0ErMUb2vZr22ro/d2e0EMEU1aXLF9wdwhgluGSQKX5Ti+Qk+a4illLc
Qbc171SQiFp7K3gkpndvFYZmA3qJKsCifqLmzWLS112g4AsJEALWbHYt/BXis1hh
ifQqBTS/fRTf2jrZJpi4ABLSH5NT7FSq1BZAsYikxhKMVp6L6nVrmXq1TjoBDfox
fKTMJBR7SkeL5bnXxvTiY/Kl2C5d9/80lGdUMRGhCfrW+WxYCenk6GNPblTTeFdR
DpdsVzD5ohB81bqaI1JfRsorqvnGak1EnUfZEH2G98icYJNUZQid1PMWEcgYMDj5
RxyDuULT3SYOFSqndPqgnOV2EBgDvSQkomOLne5jxzqbyGc/tnCAfsVnj5v0tE6L
WGkVXEbqhmfrVPKydD7VEYptMTIcbPQ7q4ZXtIV4klOltPHq5NvoZY0jbm30adC7
SOOTNHBizozO9pNa63tHdf63775qsfC8KKM9jO9IhGmwoF8+fgSLCOGJfR3nciUa
E2M0eQaQCYVnNvSCAbAGwPhXnpETsoY8mTDVeSCUoqWiD2qKss0OxczLdGt6BONC
euXwt2bVKrS7XYy7H49Dlxhs/jRKS2YU2TjwPlRbChw3K6XhuadkLBWlbtNmPotF
JR5ROs5aBEoDz2x/2pdTn3zuzdCbd2C0nzCuv4yUDDr6eTttTPapzoFi8Vjiy21P
BG0GGaJBO59TqfCu+byeBECyXm37OJn08e2EeplFuILYD5Oxks2NPSmf+18XrH7e
bibZG9kO6OneHak1zQrN64gq24DJR1fu7hFw6pZL7205XIV/WuVU2kkKKGAFS+wG
zhpCrhHRsFPWyOXrMa4OVoVdkZ38DraWTINyInRLiijAuIOXUOTZjRu171ynne8g
z34zNiBhPk6QdHmXjfQPiKASQHOM8iHH3ssM0LsIw8Ox2hDO8gOZFGvQ+Yaje8Yq
YUWX+D7oBxtZpmjzkteUyi/vjn6ze1/TeLpAFARTgYBKii3HOV4tGO7Opj5TqfGB
0AjOcYJMzMZvOLMP78CksAeRS2ZKByZRxsIgJsst8WXLd3xh25H49Wxt88JKgeEn
na37qkRkM21yWdoD3JolUONWrhBjiCC7KmkpVGCXgjZBmWtqpcntLLSu+S3MRHhc
bm7pznmnSX6OgNdAnOt20fRrU/DJZJFPN1iFdNwfoHf+9RY/B+yNPK6KgPkPm8nc
OQ3de4rszo59RL1xwDsj7w+I45lBmDwXa4y5vOE6Ij9mqFjco1MWNAjmxbgKLc46
gv23hlNBjtrwM6nSrBEs/ViWoNUacChEIaFM3bppd9uB/mLhCIsmm7uHHeI82vbr
9eRXN5UCxaeui0+2+gvNX4Tql9Oq9CtlIYflPkMd1DEXJyFXgrseOwI1jHLYTHfH
S0KKdAZhD1JgEJFz4xRt4NExES/mXA7u8CzWPoWy/xOIm2/qMwJDM5vDS9k50hBh
2SsPBHRQ0DjiTJcUZLVT6t79YK2ypZSbniMZZ7s9BDGyeqk8kBvjjWc195WNyzCk
GAy6cjZsKKqwvugnsvD8ByG/R2O7WYgm3VTN5YTkpvaskPWVEyu3JoghGWUq2jV4
Oco6C+FZQkp6FWE6U0gECr7r2ZH2Sai+IruI/tBiU0RbjNj441wqHMX32EJ+tvwl
TA2IzNZR++TiYzo/X6NVFbixLulk+fBzl/qKNoWWnUdPcgf+HeTtU+toqydf2Dir
7i07wBC8Q73FS+3NtDRmqSvopdiV1qmkAVWH0QhkYib21WBxCGTKNwyWQLx5wQ9X
Pd5ej1cfA4/hJPu3Kj3zAbrhOp5bbhynzlQy9OrCv9CrWf/UmVZJg+U2WoJI0BD7
rFklzKH80ALcfJk3LuMFQa0HjJZdU2Vn9C/+EX18NLLdlgB3Ki/Xx8oIK6GGzV6/
ZrNSdIn3YXUM0JH6e4lEEqa9T4GQFwToNXKTnciVMG0Yp/rTYXq1nz9M7lYKoeD5
h8RiDTMM1W4Xuv9QJKt1YygKRwXAgGfSJ+7vR8BfW4Y2N8I3F+PkbNc7YfQmk+pc
JYnOhTsT1eGJJdO8iAgNo9H3o2VF7D19zhJdDG7JIuMp3Fz0lPhgW2ahwcReZ8rc
szypTw4Hhm7jw9QdT0ZXysU0IplzPy+bnsFOSF9gkzkrlmeTAhjAMVbgdr8UOMMe
pXDlYKUuYJBYW6Z/Jbdvw5dOMc95edt93Rt12IL866H34IsklvS0XGSS7fYHGkGg
gglGHrz+jGsMUotGSSe1Qd56q722uqrGPamuy4rlqn7K6SKHsqF9U0WOlmAtKZ2S
SvsckHj4/juIcbxu/k+CXPPmR0djZgB2FpLTN7xIQfZxz0B714m1aaRDcr1q+UPC
EOd3gNZQD1tBgzL/RHfUNI3GuWPoQ4UGyxqtuKJ80RJ8isRgwORMoPooMHxwZxsd
CT0v3l7zwD2pFghBTEWcDDR1edlXnwU9LxEYthLjGwVE52fgTXRViT7hZKsJ48B5
N/bH4fAih4hTMlCf0LQkiQW8MJxENY6d2zZpDm9tt4+VVtVlbmO2ct0VQIrDHJhh
O39q0E33tDkQGAG0qvI2EnHMSedPyAnd1ygVmrnj4ZIBjdJMIl+Ga519K/GbMDHR
2VVeEdXkVFYLZ3EQFs3r2ogNd9V4dOnit0VHfyye8HF+J2dj+kIGZtfwWxf21dfi
bK0oVrTqg2MJUU+pFpwXPm70LWMxaoroF2P7twKYtNxTXHsz4973Z7IwYcKX3xaX
lQCIkKAlvCK6rRINBjIBxzcMXa7GObD2NuF2QVNCilWdymi1tpQECeJf5Jj0hk8H
RzrgdWdfGENJLpvK8rrMiYqGvb0bxaP+oYejMbvqnZJAOmGDRfkrD2OpFh7P2mJ4
8AxASOgHyC9zRRwRcNavsBQ+3v3RW7pLi/F3NLk9y2Dm3CXA+RnsXpwXQX76X7XZ
VdM6VrcPyT3DlNC5fMIrqQYV1mO28XJuPDvOn/tuYwqr/vbFFNEIr0RdO+rijurx
PHSj1DecUo85KfWYvQA7iaqCzs/3KcPDX9LYTp42vyij5xmkNovyBvTtPBAjglpb
2D99X7X50nBukeGyb21mnb4slHcU4GxRNZH0hYvdsaLZYiUrzDdRu3GLAAmg6czz
wrGT3/x5fxXN5AxBlc6EqasemAvng2sCmo4pDOwxDOpreRzWQ3r9cFYjdZ9YAvmT
gHtU7Q2dWmDQ1jOldWoAR8p1D3S+MCplQTTCooDrIeCm5gWawuAixtbvojA5x/Z4
1pSKRKPppTV5we+mK0hkF81lT8Qs7NoZrU/ROM1jmgl4YC6JzgY/VTOrOmNoajSV
g2Qa35qOX3zVFasDJicPCrHnvj/W7OFpPgifccgPsAd9GkxTWSCHf/vtVuM8ALZs
tZPO2LB6w1ZjU5zS8HpMTj3KWorkMmsu9vTyQvE2ywMQaUb3GLQsaf6Fk+6fYAoT
jOdLnRiRpgODHzJxSG9VpVAiXs5YeMZqOBkrFx3XTvookSLod6UiBMzgfWoELVu3
3pPpQhPYxM14hXpji+8g/t9+gNdk0pRH22e4rdqiUWThNEr40bBJ9da2+8oaxlVi
7aBZZh+U0jnB7OSpDbxiYxhN6QfeFMqTPiyvqfcoaG+JxghFhW3AjGKCRp0KfNlp
/gsFgIq74hDGz8Ldskbbcu01HHSRZLYg8Zg2YHdRpZpUgW6ekOsGUkfHLj5Qvuzo
dbhHBuZZPlvSlJCz1VygOW/oJPYM4pwTjJut4dKLbaa5XZ3A9d6cbH1ojRhvwVwS
cKKazYW+5IpMxqACaMXOJ47JLqWrIAlvAJeiEHFxHCN+x9Sy8FVLFq92GjWUzLUi
7X1NsMcCwAHUcWAuVUEqUnZOXhKZjdO20AXcxl/ojP69HfuUSzwANtFkaaJG+Raq
82BcwAWhlQlhG4R+UnA+/lJWsZXLQFMR6ftthy+27brpgwUVSk6ejSqrFFV9DcoB
N8NoDRg9xQBn/6qGI/suUW0OB/Aclvk5EYC4DVVYW0YylwWwfroOslxZpwRCOWsm
5o1Px8A8O32AXoAYHYB/4+lp26sEFD4OST+OXunnA76GHbVR5WvuY0UyMG8XGv5b
q9eILkKjxF58z37DuSMGwMACuDODqukC318fakdepfN6JmDzDx07pGtLBSncjd8s
YDWLYACR78cwx2F/Ar7+PdyPa1j4wqf/x5C3fHXn/UrvkMfLxCsBqYdlxaI+qLcI
ZegT7z+4HHdyQH9UOXHoGqTF293zpVEfaoqjjcRasPlKp4gZCumUs1vTS5+VhfFk
ER4B967QrsiBPoyvqc8yMnzgOruIUDp+nCXkRCpgrefHeE7rsQaJHDz81aB+EBfA
huK3VOgoyKuyu7zwwwzXUvQv3XFHR2REe83yFzmyfUg8MnrI8XUqthfFnNMfcoap
9/zjdrQ7XqoXlpEnvRhJr/zMj3Kw3Tyv/UhSRDG7E03THseyO/NJrJ2xPOMlOtdv
HBmNT5qE1sT8EEyGAFau9y0f3ZDtjqc60ArPyonvC2FjZwwcloCqzHi84g3oB1yY
XUdNBD6uY3J4sJkngCmEvmeRwytro/3u62Ln9h1u9kcwBvyyiJjxp0Th70q7Zeiw
sNSsOrappECK8Kdw7mC/bDCVX5eS2ihEXDcsbbNc7H81uPTtvMdno12EKfp6E/0p
dm2cXROfTioviqFuGWIwFRL+qTcwRUNCPgem8Xbw1rcD0JcAUlNVeedMwzHfzeni
EbqdMiNf85gesDy4y1CjwC5qzC/Czo48k5ri6a5k3IlIwNeul+X2CWsjaADFJaPw
/bsQ1QlLir+922UD/XODV/xvutcFoSaWCt516Hxe3rQuQ1QXreM77Oh5hIj9UUeS
pi8Z07nuA8ASjQG2gK6lyf6GUGMQRp+RK3zqfgSEE232U5j8rFqwHdl1MXfrLvLO
tqkaFstXZjcmS9F/kD7k4tgFEbmxElKDwpl25nCL/MtsRLr2W/9k85iVVMft/a4d
YsiLTLxIpi3N3A9TId/W12QF/gWFyjPG/s9TOgciN50syQ4P9pE+IoXqLZpiWEhp
/M9YQKS9ANsYzABQZidalNmvQ77TnfV3jlcSZtHOHh0ocIxN2uSl2k/lHXsw4LaX
3fLF2MfUpN+reF6txZXBq1pdsT54solBWzkY+0WqllvIYSglRS92CGCdlUMT4TNy
wAC2Y7rdovUF783kjJhSGlwfjwOYS2G+uDE6aT5+o4yRIBqxeDFjA7ZGRB66DKqT
N1zi2sPak7o8mBdOXry2qEaj2iqeOmXKsWpfv1IUrZwsmEq6DwymCCLXB6jw3F9Y
pyLwK4/gmVLB0N3wyoJBdLA/MUSTRy+tnVN7G35NgY7G+P07m+K+bGosE23R4RC+
+MkUeJb3/RCV0OsBwbjhoqALbmwQxpyPpggObbOu5Bwe8Yr+Zbl5/XzOtWU01SGB
MuzVzgweqQJdi6W/cFF80KhpcsE27yQU+uFNGAbmPwbBgDxk/k73hSTWjVcHk9vI
slf/Twj9cl7/lw4oCeFjgCvD8MBpZKR40LwV3jOJWVP2qcIwpRQwGbKrOiZ8GjgZ
byldfkoQbE2YWjxkNQjmQV6Dwm/5PL8dEziwnIzld7N5b9zGQ4bgjxmE5kglpb6w
YzVtMLrRbAyNIphIs0fMJSIQp9QwtEf7aPHmxmQ0HSE2Hdk7lgtFkEnQT8NeOZI5
a9c9NVJANwR/+n8Nm1wmF4AFnli0der6vmfplQai0xteZ2RU8sSkqGsPBOTjeFBq
aoCW3FQVK6M4FngejeEvsZxUmaQrb4jljgjN+4N21tPQBvlM9vLvr/SVzZqlyQ26
PoOaLmB1AyJb5JiOqcEcb5OrvShfaVHhySzcTuIptIO+vsGiufTeCBuc3D6DXzNf
i4xcAcIoqUVXOL103w5R7oWD2spBYF1Hbmfe7vuTU6VbJP43PCUbShUmwafwWGOB
EthZq5j8drU/Od6IrrKiNmK/qXjVkOvecP9MMX8QEYNJMLKB/2MWWtKjWqEIHjtO
TwLP5zTBq0MjlOoagK0mQlScEwH2o3D6mZ+vt8otYppFfIzFXnvqAqAfBmA+5iCc
L79qsZ7NlaKH1ONlwYruAXv4NSEMkl/UQlwYDPBADon9lR7Onz5T5Cy8Y68qcAu6
MduualW4DOz0BFdQJomcH/84IETfMTplQgrJPCzrlHgyHOcN4x6iHwtaymdUi09s
9snz4oyya3sdmZDE/1Qa0wNmB4WQJk+spwRElM7rHmuzMyiuHUPFJQPj5w9scf+J
JSXakL67l8vrzkkqeTb8BFY41/pUcpiJO1NhwIXkettRPt83pz4S26IxRU1p232M
lhpva0mXNNcHdvNPVb3X3dlPoT0AMct8m5t0b+QgDCv0JLbyij/U+zN/L0PHTMm+
4auw2+OJwJsMC3uh6akRfszYqnLYsEy2PO3xuUO5QgF9UAagIbBkfg0AGCoyGdEq
BomqR1wo4BBmWtKEYoH7wIFKEoV5HjanOG8ZV8U6D2PwaQXlo38V7e5vOF2x+9ww
gdWrczQiBzP0oyUS+tan8ugCGhDTxI/n3RFxt84wlwkrB9N3A1MSLIYvLDuX2p0I
VSvhtMbmiAdCcHL6TkAOLjPafOMiKEoVqO3GEnKkTfnPnAOLF2g+k+dFEsO37NaX
kW9vuZ4SY8wA1hirPSOwqqa4lH1i5EkZuTBKdPaQ99sqsgUor2VSTfHuHx7WYZhC
QyMp5mWwfr+oGh+OZglE9rV1C9rvwLF34WkXNzScE898m8WKM+LUMPdH6KRqwASF
scRZCu9RH2gagpjmU3OhBDPSwLmh3PkBU87wkeqwNXf3OQl0fWtSYNFP8S4/h8az
T0m6ZJe60fwefEHp0VAkrl04Bh3trGl2ECMWm5dByBwv0gJ6SjDN2lHg15saIynY
bfsNkAosxN40nBES3MGHs87Dab8imQ5b3q6tfLA9XT+9oLpciAyK9UMJilfkR1wt
ZZUK8K1K4d57XoRKohZZwp5sWsHEWeW2TNc6LH50ai36SmhRkVXqkWLz+7+9rkrX
wUsq37dTWs8nB13BkTbSJIC7vN7q3sF8FeasXkbNaEfCoPmuBmrg9b6BO2b6/+rz
+PghCLPRFuAfoFb2w+4Xink67sXcMldkRPwU/Fq25Is3xTXZTb+qQvlYvLv0COer
exwtDrTDGWQ+5l6BQv/8UQAFyUoH3k7NIKAkuuVpOs04Fwx5T8/WNOEZFmjgrbdT
Q4tcs0vI+xyIL4q5yevbM2+lkmnYnp/dXZ8ma7P9BYYOdPEyqmYWc057jJJGj5JY
6CNp9uA/d3b9ZVhHqq7EPSZ1Zv6qojEE9wVBnPPSwG7NaGSZstw8i9XR5RENeZzB
JuieSab83GilMk7aUh4XGszvFHyOvC26WAPNsVU+vzFAcqUUS+ury//9mq5fcatE
IMxn24ekQ2PViGnjwI8HBqM2OkoWHkg7blBBl0FysyL0BOXLuHYLZOhj30eosJuM
VPGBM9beqbuTrDYqHL/7bX1se4ZQSekgXWt2qQpCmI7t3w/+nmX7NlkxhjXkn3mW
BoDMEwB12qvctLfM76Umx/ugHF1xtGqjS1R5y0dgUP/YCbwc4373ZEG5vdd3othG
dxhsm1P83/KTfL6Wpcuufmn6e/W6ZlWTnggdW6ISsJQQNTs0fx/ALDM5fZ/Rzz4B
UmQB9htWOOZLe7pejydToip17q9/dUjSR+iaa64XXGpqxrByNHYeCX3NAcseeAai
xEI1ksfseaYy33Xr6MH7LJ79dZZl0ZwZesJWoCIkFiwoZdlEKXkEpsPcU5gmXIQJ
i1w3l8ccCscqYVuuRHZvGuZII1/btxu2fvK3nJkm/RMbbTCjWqdiT141o1D4gNve
AUY4RfsQ/Ekrm1cv1KK1riJQ+e/BtxRxaU4ZmNnznZrc6a534xV6WXZGvrkunggk
5QxUpA2bxPCe5J08NR6c78r0yWYZP0dAmb/jTxwcP7jEg8cW5Dnv3gwxJZFk3Bvp
JWJtFoPhGS/jv6jnPANXlTCauo6W46hvfWL46QOJfG5vtRWPg/MhvM+5aK3XhaiV
0awiQ2Iw7jf1alO6+rfS5ZMkTLxeQhvYh5j/CAKdRUcKYoZIL/TINYhfprxpU420
ZN88+1LUR3OTG//APAwthxBo9ktqsW4ruiOVBDruGWRWEmc+FMoHYFLbU6H2z4gb
+H/Ww0sThAAH2x9Zv+lVeRBdnaKnGr5X0b/pBW8iqFFGRWcqmCaKOZD6Uul/jFwa
Ak1wx+uzJNKc07gB/MrkfMQ2GUwbnX4RWCd5NrxfJKIxCsM8WO7wUtp2fFjbX8TF
AxK+HHK9NQJTpjrC2W7XkeVy5CDqAu7tMDK17E0ePfvMnuHAJyG5DRJ7AP1fiuuD
XqEI6Db7Byt8ZGiGn1w3ibX1KolDgGjRO8nFr5fE8HlvjHSgC8TV2dMeTWX3R6wC
8Umg9TvL556Zt2jz4psMk0Ba+ArrCp/W16wAfA3pL3aLnDa8yHwwRC9TPQ6Tn6Bo
PfuFajFF8MUc3KJGAnwm1f77QEYmHUIm//vtsrqnWqDSOcf1dRV9tWTIIQU/r/8Z
L1JcBrHCFy+W2JlKL+ciBnNeqr50umGLEaEY7uvlJlA1H/azXVLhigWJkXaCBupW
Px8N73xNChbqUfCCW3TNpBTUC0YeCTLdFmayG5gEEnKPE4t3DhUYHz95OWUi17JC
gg2DwXM0JIHy+M3w9nHl0qI3FPDVFsSQK/APxEA+6n8HmqOwZkNEOX1Uyf5N49q6
Yfht5RHAdKDpNkhKEhnVRRcdCxeX14t2Hk1zS7v8uX6TaxmqaSQrZDYsv6mcwbUH
wZQiu/UUjJ3D2SIdL4sBM+/mIuIeiQsMBoSq6GPrD3u1vMT3msM5kjGYTU/u1KIp
pJjMj0L6j3BQf5vxRj99GIMW9lhrYgOBV+aMm+L07gmwiubVxfmjjHCyokbt5Qu+
Q6rHnLd+gg97yjvXxCDdlUPEUnzdG4/2VEAfiQQWfT3AKWoFh9BeD1ceYIKqXHP4
bXpcZaY4JNBPBHhBa/sn0DS96lFxW7jtelHeIbUv7z/1TpbzI8giTiB/UmbGsjqp
er+DlxhKAM+ckOarHsEY30pjkes3K2eITuxgs3qDEwxnjFab0+BiJ0RaxTEuoa3n
V2Y8vV+YjNnV44HNl/r5bboq2CHqdaHCtZT9czenCYijrnXaQIMOkuc+D8aH4weP
wd1wKwA27z8s59AhaLo78EaSv8V+o9wWqlQpNGfkeUzJVfnrpqsD0wOSnbE43tS7
oIm+LglYa5/MRK6osS0V8mS9IFYYZvejo4fqQcUk69ZWgZRVhlGUc86QncfclkQz
wxxhz7SqNt+lEPpiRBc0yRv0xwdpmrTqT1WeOkJalRuR3Q9Ajbhv4InY8vYKYIVa
fxPyTi793BlkGs6oFgRPds7Exrgo+9SA4rjK9ygRa4C6zhDeo5xmTCfzsOFrsp0w
SDXZijJcmYz+GnZuniSY5z5hAISfNoF6X6kuHklhB8/cLVpoAumI2Tvk5OZXaLfU
CbbrZKVuALVQOUovIQoYPvwsRQEUpYxXYUjIlJvHbrulozT3mtEWaPpVjVGH9Rux
NLqZOOp2KczyWntf20bD/8ny21rMXm1AutyY5VGvQRLYV3b6L1Ecsbb2HF3vsRJK
+6gYc5ancZS40uhMG/Y9FzaGZHbr9vRqkGmFPT32HEkVvwjfjsVL1oPoRDPE9XgI
Sg4MT+CDwzCsQbgZbqCtnqj9d/Ur6SAeG2a1Q0ckLyNeprUj5xQ3KGYj6uF7/5j+
gbNSQCWArcvp11AYnBsOuGI16/kzkZ0UavLsICXAA6u35VDc1bACJYGpwdTmib+e
LObpAbdbJCjkF1FcnfsUOg1BbiUmpAjP9WnYYzmPK+9Lvnd4mOSIsjxnZUxBokXH
Zjae89DUjzerpC6PiQLvFGKeRVs7OdbyohSvwJK1frp7AbBs6GnrocjOUL26N31r
LaFnI/ak+lN1OdnpPIaGgQS6py1mIKZQxgFNIBm4bWGxQOPfX07LtqMMDAGbSqCM
0dQCjymQxkWDpl96QjVpt3iBdOsVpsI+H9JaltEU0czFBSCvexM7PQvPKWdlrmR+
51ddjLE6mREhu8rRfmlCRQKkH32Gvruetq3Xgqrs6gGlZKyjM3KF3jx+jGFGDsCk
49sYOmw4tejbrm/+E2q7ww81NSidcXgRDVAaFRKVCvKa28SA2VENMIVC9ssmSON3
XWg1pY+K51Dbo5/z+lUQtL+QGF/84QBqGjs1SYcuca5ZuTHwo88qERGVa5hcud2e
RLoy2GIsON5mU7aCYsmlbo3Oz3A4ukPo3LMra56qCzEkoeQCR5YoYiLmZ5mLcUJH
OQhNWm3G3CKLouHMTHdBHJshyaRv+qlrCM10GIHBPeecw3uWJEBW2p03kJYkrYZE
+N2gkObE4WK+ng9H2ELlY1Uq7Qigr3RPxxJXgZ0BKNI6+jlkv2v9o1HfRSuMCdoR
rUt0GPkkmVrHlsTNalAgDlYuNvnpraq6fv6HbFSxFelFYsYp+0CU2VleK/wTAYNW
ZqpJRs9PfWOlamHodCLnpwN35g65X0wfa6zIjacXqYgcVENbFcw58voMfG4BEMa+
ptp41MSu1komrTPMMs9gDRkE2lDxm+rttZ+d5CD40oLlKkMkhLCK49RjoBpe13HI
9PUdk3g+9i3zw2m3Pecdngz5wb7xMu/qWISVAtdeZ6POIUIcJobiPSd9UimyAaEB
YR5yVDqcf4BRPUt78IespLBIwdCBb3hQ1dMIP6RiMr5s6t44PL0G3DGp4zXPLjrT
yfOP9YsQ4Eluaeg5D1C56N5R6izKqb7ovZSleVi00wPfRmxBm6qTjnpNRTkM5zyS
e4eLNOtyVEzCW0czljdCyPL0zGI7Ud6EJwytEoGajRIDKLioufnTgis2pDG0RSc0
VVwaF9M2uC4MuEljSojtxazJeC4UBKjhUC8cXNdUyhZV0zd88T31dbrUiCzaLY2a
TJXpA+677VZsLGVELxoTQcu5ky5Mc+RAZIrpwbNjq9r16auwBnBRB3AkurT/d3lj
zL9BxMvvVGbvDb++qbXIq5J5LyK9CWng0A/VoSu71rqOP75ZQLhBVFpWUYAQvk/P
56N/u4rJ/vGX7FJEYqBPBnmQS3/GaDRit91vrppMB6QdScnJWiHXtSuXB3d4MIU4
QNaXJUa9aDJq08v5kDjqPuF9up3tRHIBK+5/zhNBFM1PkjTlLvPx+gRldgXh3rIf
W2Cm6jyk6eTYjCNOInY1D311VTR6IY+2rNlwLUg0sB+7BJMQR6i4CZJwU1bMV9AN
SdsPvfeUNtw6Iohx8sM+i4N2HP1HXJXpJsdQE1GJc3/9hVhyi8Qn1ZfVtDjm7mhG
nEQ/NIPEufCWfJ8/sZuDdJr3/5bDQOJvMzE5Yxr8KFZDR1G4vJ0JL7sPJ5Hy+Hbl
vHQr79pc+KQhc0R4eVAszcx/fzvZtYT5LgMNaHfuisfxW/tubOKpCgz2GGIo0jNl
RvIbqFqtoIA0mIKiKA0ryAn9JbV/wiVTZZW3ErN371+qSsW64cMkutAXTG+PUrQF
cNds+fKpOnSeLnnPDPrIfHPMdHsWPddBrl/xLF/zCib3ScRE/j9/h8vSzUHgU2Zc
ogX4fj/yDdKR0NSRHuGB4IWyEFQI6/1qj4CpyVfM/dWc9yW7bRG1l7W0EQrM+Wzb
VSHjIZF4vxynqPqkkHg8LMXlN8NnAr9ja/m7H7Gky0IAemTdnJVhYJzaNyxmqytX
XskLKHkHECEbCo8CvgLptbjsBjQGujXqOtFq6EQ0WwkJpbSn8IzyEEy916ZMdqWd
5D+EVXbVDTqJ91JINmgSaDGPljtuWzT3Ug6DQdqOIr9mDPULNCQI8OTx9YoMIopY
P5TLnZmOkEqitoBiY5jFx3X8nmHV60MzzcB8A+ZY27BI/MLqJHBJwEJfFmpOvDtp
Jeao16U5rZWx46MCGBPqxw7J47PkSgxKKnNA4+iTeugCl/XJCzmjGlZgK+mbFb1z
//dp31ELJuAamEodH4ougVLwhDTzCq/oPnfaj9IwXKfrW4Th2Le+Ud1jwogd6cWF
5pmNDEAag/ZMfAiIP6ET3dtRimtRWSDyfIMMYRqWCFnCbzDYQ2GY7WmM/4B+h1CQ
a6WrwxeVunT4xqcSoh59Egbj/vLoxMPerw2QM5F3Mc0OVUhvtdRfDW4rapHcCdfF
vHLt99ETzWteQQZWBc7EfovPMfmYbjXmTuwypQgdpQHPldYEdu1lmRamdXx23ci2
4p8yrf9Wis/2lkrhmVo+TcRyTQetbR5CMQUZP7nlrHsq2K9wPKB+DnFfYIZ2JmQK
nm6C1inD47qOCPBGCgc8XW1LhgUbDPX4n7A/BNOx1z1NBWHLXXKY9RgINqDa3k40
LLMXn/rwq4BNvQ6QOMsjXtq0ziaXZa45IueMccrJJeazE5YAxGk82QCGDldOYbJO
OjNhaJHdlSTRWk3n9p6hoINZcLF4ppxKXGaRIvLXNyMfAsqDef+KQtknZEZ7//pI
UF8kOs5iVAf95A4JaBble+g0+kAkNpLNQkENBz4x1oBLA9Iywu6hqyAFPhnCY1YY
F0OqkmT1AAC+0QuFH/y2ZQBeGvo9E6hnnKzOpa0SeQOA2Omh3yS8uJB0XXOhdj4p
V5zmMZsRIECp1ZRxyx4S71RWHE9uzzyrkiuar4vuOhgKEl6jDJJbAL1otcFkvino
cvChNAxJ2Sp40IFve7Lt1AIyB2xQcvJiKKUmDkx7f1ivNVA/9rgXj7U0hyyCqSVG
PusDlfkhSHrQmh0J4CcTKBjFm4WSmpGuybIcxr8G4rYxz+7f3TrFJkuQJ9tpesHH
N7aj5nlq9F3M/iN15raT279m6XE+OlKHrA9okiPRbwwaRK+g4SGuWAZFIlROnH/M
l6/8Nx3wzjsON+nq1yCdKz4/GhdACmiNG1Veadn26RR0uO1v+erzGWgo0zbyS6DH
7zmPjsl6lC6aZV9snKrVWre3UhLc1hPo47qqQKdjawuT2A6Quf3UP7FaP2NFlXf4
wzPqlQkOKabfeEaKuoMwsLWQWXXwb7zGpVJ64TOIDVI1wdohOvTqsRUCy2b2Z1T1
2qNLNahnHeksnmzzZ+576JhLmraT7oM3ib7OGUqtlvpUE9+d5zJrr1+Goq3BM9SD
zVXSQcOqTTIEuDOAZ3//UWnJTXkQHHpXv4vG+MoCY3phJ74IF+d8jnhDt5CyYqxb
TwW3/OSGc+dvR0HlLjAcXt7OVf4+Dz9D3yNVUJEZ8GoKJCAHtI8WpjOZp6gmQ8Xz
29HxuBnWp4SHRaqWKCuGQQNk0ennnqND9RX65YsoOVinfC489Q48RM2jRkqn8VB2
iHoSyxZOUi8JKARd+tv/pKn/guyyEi6FYC+RFCNUK3obJ0QYtDEAkF33EKUhHrYr
wAZk54GepTnhkVZRWh7Y3Wc8Cho9Dls2wTu9BU9rVYRcXN68YIaCbNIVFj0qFygK
1yLzFs7LDPWpdDiOMjYDApD6Jsb6h7sugVddg2vD7/OnP8cj8NK4Dpz9XvxgSsBS
iYBcsrudzcckAJX0dT8lnT76WFf2l/AjGaBjqeWg82RLIlO2caUdTU2+hZx5zD+/
19T49FykXigBAWD+x+EEYOG2BLY9NI7jMx+fIgxQ3nYUySpSQjeHADUE+CU7i6YH
FtYyd0zDm7A24QDDddJ5sTP18IoPUl19ioOU9noxy0aZL3eQEmOuXtjHNqjMaaCa
YM871dBQ132mKrKthMvhTXwm8PhE3YcZ2Hrme46RAsa/GknA2nNeRHHJJ74/7n3X
NFPmfZq77QrR8FUXJxv616T9eemVNCOzbfOk6XWM5CTrRf7Nz/bxyOiZ/ooxTl7D
UDXjX7+i9xKKK5Jv4BvPNcq1qhjlV/2px0o3HJ58Ip++kDK6Ejai+YLE3Ao3TE5Z
UW18VBkYfPQxfitQGaMuHJejUgURZnwzsLGrsRSY4aUU5T64Ok3nF3HuXQPyGhE4
KeRg1mqjf9GkVbg/JuPD5gW5UcyHmRHsE9ksfRuqD7qjoZ/s7ECTVsmT5EYx3IGx
81jw+YGd/yOI8nfmcl3Efx6yZNspfvbCdjucykKnY9h0Im//iZ0X7Fdr1HMJ18fH
cZ8AX8KOLwqFj3pQgUXE1uPO6f/sY9qJ5qNdzV6H+JncElLqolsRUKmSfhQVW+WJ
qt/QOQ/Ej9GU4ceimJ4JglNIAEIAGhKz0HrhTG6Ki8dDBR91b2IenkIwEOAtMd+/
pNQPoH/sj4Zl+NmpDQuDcZMCNapGpj0VeDe6/yMcBtbWUOlsTKGF5lAxdyXf2Zf2
oY3TYuhMfxc19mSFji8JJMnZirkI3VFNbwLG+HBDnVUNCemhUeNC9nnfxuAE6T2M
j19HuQM/eLZtXgJGJIATHWij0BaJgYbd24rgI/p1cYUYrVUDhvFzudnq2QK3/hVy
uKcNIy+c+iReG7m6miqJJE2bRv40pgNPWAWy4CajM4zP+ZpbGcx+JSpQa6inJtOe
xje6VWLuDxyovlYIjSgpKM9f+qBo3pq4t9V2Wzzsq+0/4nnokQZVx250co+1TuGK
nnwCtwQnq7c5sQnQdD93cMw6ka73rjfegvwMkL67J54Ew2NdsCP8wF5FxHuB+WJL
/cMWvAo5SbFb7lBhd4a0cgeSwbYY82yzhDc+ppgwa4gzhgmXXBM3MaIRLPCXMIY8
FmZSAObCg1gXsJCU81U19rVNc3Gtwy+QClmlqpkZtHcqp+4QT40rym/W3t58KqoX
ibjnxhqqgEo6dB8lcN96/mEB7WXJra2p2AVZH0D/g1j8jKbWeb4stmQtkriRD8mU
XW3k9ReKJx55M44bpCCwafKoGXL3J/l0lQICFG2XMEacWwrcnuD+eA/I0S+BWzJY
B61CeN9GMIyIhoAwEX7NE4yhdynTirRyJ7XfNmtCjlEZfl+KHVSypwr9uGcq9sss
o63JFTGAx411s6GIOGypP4Z7E7OMjhINrXk2DKL5scvAaHAhlkimg7WVAwMIuArf
7yFlMRln+BgSeG6v5fSNF7hnxoorculwPlgsUOIa9Yf9gsZSACQqhc4s2KNTLRwo
T7o/BtpVI63RJw3aBBIPVVzBnD4ttt72XusOMFuvFfBzYVsJnDIJFhOcMYSXZ08x
jrU+B8vk8ik1DWpTzSrQtk6w6+C0PASNd6OHRxt5lWtqV46bmcqLSdZuEgpP0UsG
Hi+gpLHsYDcVephy4MU7SBfibZzbbnKXZQNXsEc/2PWSMrF/osNyB6klwa18Qc9S
Omm2QFHTa42TCUe8KWIC+1O3N56hx1T6SVzoF2PL/2c4RlfHpHzIprSItbqEoDZ0
/D/LQqsIGKb9kH6w6H8vHgOZ1Cs8zn/ORPB5UHSXbj7/ueKlH4uEe0xUXG/cAg5X
HGyEPyFQ+n4TD2WbtwWdisX3nViqpPXfxJO3NmhzVTMj589cTJke6VmRy9ws1DbN
I4dO1GiAnmR2Yl79linTnak9ZA8WrGdCDxLLKzuq4FvjOQ52hEN1rQJvpmYEtBSx
/LIBN0mcBgl0JLFgipXr24AcgFzasluvGo1tD0C+iUWdEqhcSzTiFvu8BaJDVArU
x5pQ98ynq7LHU5cbU5EPwoDjE8Kq+mBW+JOYF72+6Cf4obzFUQ+ODiMvmi7PY2/7
oyu90fXojQEZcnzybsfXC08RF02AvTSggtPHvbLGr++vX4RvtDdkTvB9RnCNhvew
V6OxlMJtAidnvCmUXKbcf4mb6xi9HYpaUSTXjkIv6ZFloqA5/dpprICi+lAzB2+C
ieInCQaKNC/kLuCTU12gghl7u1kC93UtH9ye4VTP2fQCL0B6lzpKcilCmsrTg3zO
xHr18vHadXIwF5GLbbpnWLQbmgw8oxQJdPGQ49Chac3pXyiu7kv9oWZaEtPn2vde
/jG4OFikothPijRnRHQv0SbW6tFoTCGasyQcjpOr7Rphurd3ZVFMoi/PFsCKGrq8
DAgYbPSZA0yun/ZpbdXTRCfeyMA37SEPqT69yu5Uyy1LDk3pgCp0uIvs4fsGaM+F
/7vPTwscOv38Dc11yo6xu5mMM7NQCgv2/Dyq2bW1pTjDBVAd8B+gQlXaOJmQX8s1
M61YX2c3z0fquQilli0tUpE86WrGzBf+ARuYxlyzTkM=
`pragma protect end_protected
