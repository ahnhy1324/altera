// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SHjgU9gwhllc2cYOLwK+zX1aGZqY9KO+rlSRQSqXaQmyl1po767/zjMlT5+FdWJa
i+uzeoxaauyP6+xaVcK+0XmS5IFJYvAehYwwQuJN67Ll0nWOCmBEgTKKxBy6wdlO
Qj5izwtaxBjCjDSvs9QxOdDhxcetit+oMHbOaBOMCJI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 62112)
SdkVsPA2R/cfBs9PMT50WAt6Xe+bAxgkLv0oRYR0FnulqWpiVFJLf4hfh742nJpO
3t9l5qVHirtoZigEuFxpZUP8osZputHFqYV8gGfFDX/1rgWZVccnt+7SIAjKD1zZ
qBEWZ5HuT+B1KB2d9O+WAXsURQtLSkkGzG72IKWNbK8Wama2fPpQbuAj/ZFpCgE4
oS8uqbhB1R3mFJ1r3GmV6+q9X+lgwgNcTCmy6euPEIo1J+tuYR/slMvxc6q89NZM
VForIIGSoGGs6igiFDEzDCu4Yy2hiLJlzrmV5HXJNSyxyyYKWEjK6NyuYtjFaeIl
OCD6uFTF1FTEZhjO4UHv7xi808YExpi7PKd7i6O48nxuOi5Ny6Y3LdEycd4EumPj
cheq2FJ5tMUY6zpsTZh+Nlt5KstH1d0CLQUIctkmYHqQQ3bDGM6TkYw/nCuUlPoP
7HpbANjppsUPPJruwm5hNggzpQ8upn4ryJFV7FiHv338Vv1e4GAqKaWH3fw3LOjM
erGfs+zG+TWj1odhpiRjjjTDbi/t30CGlKCnxbrs1Sv8cMvWLl9H0gQbyqcSUb5m
YwGgcWpBJJyCM9byxo9FSBJkJZaStndn9dAgxO/H6RZInGrWzKGfvzYGQlK0oEUu
JIGx/ecknhbzhVCGlbcBEuDT2BGcJhrHsGUUkRZExyYSY+C34rViF1fWUpB7KGJR
fdiENMZH05Pj+8LoP/tCDnK02/pbHAKyn73LXgVJLqYQwHPGl/aTGvf9wmr10kS+
YsdVgrw3eU2ZqekLN27AxJpKqUgPK3cGxX2EHSNCIUIMyMvYKWp9vKIQbTUycGOh
BfGIsqcRWmv8OVcpF45/jygmCCBtSLKcNUYb9z5CBK7s1MLIFv+bzLAXBSuJ4ja1
jof1Z5UEXDAdw65+5/vM67zbLSPovlALhbk/eS/l8KV6ATgO0tk1267UeSo0xN5S
aL/2pZDfUJn4qhL2dKSDTuxjaNygfrGxk64RMjC0Z90GC9nBxR4XrLSnvNLvr59F
saQ0EGbIc9VZuXGjnOogNTfNlr46lm2ESjnVllaps3fT+o5Wm7hopV9tCtrvi7PF
YYF7pwF2Tp0kLrTyJmoRWAPbuKka4WJS8LGmnPHGVtQsCOAb9Okqg8q9LL2lfQXu
dlKPi2WOXT0+L9rpZ3/qUn3NJbXSm7TLtmcuaVve7qLY8qSAEhrFR7y9tv9eVbhW
nSOu4+QLlIF4PNqAXAags2VLhHl93X41zP5SGtj4aYiXhJtg22JZ6t/WSWejPGOV
OxqoWvWmoBNftJq56v7rF45RWChE3hieul/ibzAkZr3izAOyXU6WRTzhXUohYoTl
SZ7IVIVlTYSfBgr8mZRRNgi4ij6CVISiq0o9W00KQgoNcb8NA+whgmK6qxNNLWDm
X8eHoDYe3n8NY2AdQGoDTbPCJr+N/DcPZODDdE7TbaF20Pn4GiuCaIEq5nCTWjx+
mMjdBTpcFl38CKOJmm+TbvZNF8kpFFJHzGJwQufj5gdkH22hcbk5ub+QIw1UhsWX
cXQciD7y5diqb8yOEMfFHPE1zMwle65F6dWdSwq/j0VAssfIausYi8SO30SAhGLT
01vDVY3R8sU+BV8WbGsEXv5S39+37v/ZfBVGX0JEcXQ49B4bUxblqrTHiP6UttwN
W+OQwByfy3hxaMHgm80GLt1ZQXrxNxHY2k9koT2reAvIFGyWCxLIJ69iQ7l0uZ//
xqEb/0BgKls7KbJI0/EMcqMFgZ0Pp5o0N3zkABU41PycotqY0nn1vlIikLZK4Ct8
bLDSkA3sIc83WEcxKeRsxTasPHMSPPLADSu5/uH/oA5Lr7i9roIp1qL8+Lbc6zcc
ptl9AUTfqi0ODnL3RQTnaGZuDgHzS+knFflgJcOKG55Tf/bs6fiGqFKjqKsJ/FdD
hGF5vo9ouB1W9p0hS/HZI1pscbKG5aTqg3sbtiguECyWVGyhCw0jXABoPFXFUQfC
PgLwuA1GuIGMD2Xo2KkYaVFwLFsNxYf8Fn7HRMltAbD0YdWYCfATgD2OoLT+huAX
KqWmSUc5fopZQUOFFjFktISsr/LSGkikEqZJ7E11AervXzK4X9VTJEXng6Shv9Bo
DWSHZb9TI8bgGJCngCEAiZizLMZTnVtl8w+e9xizpULAi1SjCZScm1QLe6Hf9zpj
AkW6FKg25ogLGSCWU0Sw5qvb+cM0aw93G+5om3RpqVxzP3qSfcktCdmnHhmTw+O6
WTnJ9A4sRHtI+Aw74dHbTGYK5aw9ii4JLgUpx/Q+oT7FzpSja9B7aOHw03OnTJQI
N7rTnvCJgwm7QtRuwEhVCYrhJtFNMTEwF70VIURww6IBal5lcG6jFZncno71Y8KJ
l6J0QLLkncH/pOT1I6pSc1pZLIzQYQD3HeixM1r0or2qrL9mHy5QuHFByPaQaT38
cYOVCNptlpddRCn4U+L+jWoGmZrLwPS8X46p218X94ODQWrB1F4KoArBqMJCoOzp
j2buscFaTBC1D/ibfay/A5WKr3a+mUtmNnCfensVYmFsxHs+jP8Nh09e0sMqxnaR
MHgdKOx0NKpZ0pp/GUVkKfO7sSQXJlxRGzZXxqdAOqQ1Vub8VNcxpbNr1tpTN2l6
WTQKvLuip2KDe8TXui3U+i/T52a2RP/6Fkfv84ykhHn6pXExkFFKOaFWuanNA3jA
xZZL2e4k6u/99hwehe4kz2W8yvfJzZRyHIYM+mkuU/WLxB1Ap7ubFzpxgDALEBf4
UJ/iDTaHFBdKoDaq5EohY68oGcpNchdaZ+iE1fyY/6ArOqMjKooRLe9romEMFpm5
F/CqzH63CKJ6FYylhl+OEtGGR9x7xdZBItk67VL1epknB0QORlXuZ+lySrV12se7
3Cb3a+PCk6uj2cEcFVesV6BlfDU+qcMKn/AYBKBvJ/MNZUGYx0CytqJDusq4xyiE
ZqRZFkHRBoLu1wpSuFotwSV6afi/TVgTzxg1Ng/JlMOG99k+zI5ZZVEjA/elsrm3
pa2rLq3F2GnSLqJXmY2D/xY9upkWWySMVHpgvIdwpmGUEbOIt+fy25anHX3Fcom2
Bx3OsZTcnxVGisst/8tUzMmNx5K2PmJXji20+FTaYmPlG+pX+qO+obAtODaM7lXH
9uAsRtk0n0NQM78Aw7UdpfMaWLHJPLtj1Tq7AmaPCjtj+PlwZaZCNOPducK72y56
zZHpPmw1va+UnfW5y+j+E4wdMlOt34eN9LCE8bVytcXDMwnvQM2O79RhGuFghLlx
F4fcN9FFagGlJRUy44dDR4FZWCdCSMw8plkqSRzErO5DhnD4o0E47BirmfRNZeiY
w8Yb4BwmNRoC+9dvQBKEyyRvgCLOUC8AFQfDkjxmrJDXtVRjobEWVOluUIu3wiv4
z0/FlmlYDypP6tLIOT0LuuUMk6ORRZZYsl1c+HJjuKls+Wxu5nBWZJr1zwXc8bWV
u5NMSAsjYW1AaKovMg3CnpGcquf1xnwAlYxVBg1/wNwYzvcfCUJW5mAjc6NH/bt5
vOK2pckImevIb8FHFW/RtTBq1hwe5vk13yQUIGowDPCAhrY/fy8tiF1Kiz05xON2
QQvsqoCZydM0V5i2l8QFRZBnXDY1NeeW89BVNhwqzZ7ji2DTRI6EiP9fkP8HqEGQ
sOCkwJvUEYIUFWJsPrp2YZDhzi5H6KwqWT8ieYmg5GVyYUZRksFHGl69E5iVQzF0
XfdO6LZr4CBPRr0EfI9O+zrzOz5QRlJsB1QEUgJ0n685NJ5IHGmNdYNXCmkYa0YY
SaGnbFnLJ+4T8U8YBmYE25Ev5L9ijpfBWTzIJOQihUqnk9oO1wzf5jF4YrIv8UXZ
UTK6Pb3jYHJ5SpmDnWVSiW0wqKY+po0iPNrwGaFgjHY0Qhz2p8ZokKLPIiZpzoG+
Z4KoZiAFkkufLTBBxOO0DsLpMTd6pzj2ERImv186qHZhqVVFWFNLrJ914KbNUW4O
sT33UfkuwK9bDz9NJC40yse6KTr1CNM0lp7ckULcJiDOJZv08ZCYq7Im1OlUicPg
YGoMTLblN8WhpHMWRzECcXq1q+AS6wuSi9dmUi3IFVYplH4sFRbSdMNrjCVcaPtN
fagcBN1lavFGs4c4vJrGNpp2V2Unmz+Mh+DjdVJUSIAq4xW4HbO9QuEAlnYRy/g+
oV1DBQpiFtP/S9aqWTLOcJKrVH2VISreZ09DHKEJ6f0u8DVlvj0wVRXPVd75jWQB
gkd/atHCaMBsRXYDtOTGDWaQw+NQcIZp841HYQQiP6qJwWSYmuAc43VPGQEjlAXc
+srGp7wHURc37pa2c0JiKhwZM5/zTcDs2uEYHl8Xio2QiSFQKFd6WRFiXh44q6qm
iG366V1nM/SXdrw7xd60XWV7gNY/hHqwz+7XCrWHOA5Nd0nqLt1pHalh5dqSq2+m
e9H2a81V+vx5JNBeU3ZQARWCcFrYuowNO3z98aXl1YHb8iSFuXHnIq2+q6afJ8Rf
anxqe1xAC+FMbvLBUWF/eop3e00xAZSMbCPj8FwXhbZjAdbcsOt0pm1L3B9akxX3
Y9rpGIzJiMtcq/hhOWwnLohZlTHpq2o/k1iqIyqrQ3LLZD3afevCWzM94u8SZKE6
65USRwF+pCy/9IsejbTv188hHQmQ6qQtttko0us0PzvVLaBwk2I8pJ8jJb9PYjaO
mtoJJWVPgL8GKl2lKYx+DdbUawlIJpWwOkIBgl2ZzzLxGjEkLzeZDlAeRbYxjXHy
nss5pc6uQJq7XK5foIMcqXydse7xdsvNr74V4zbx5vWlJcZIaOmpMZtrd0c2gkx+
rNd2VcqaTMbim4K8WHLP5NTGzBaWiBaoh7tcRPcMqAwrtKUGd8AkvNLIiQqO3Ye2
/D1bpSDnQLm7c8qHqFircqU/9vavYNEplXg/GIrqSfTVsMLXQ0EP3wvkTabhp33H
JBQ0TgwDmWQmjSg4SGp9htzsjxA9MEKiYZPMqZ8MGuT36uCqTOj2IdmbsMlIfcQ5
+v+qlpU6JK30liuorkp64BoahLq6chhsCQ0NGKPspWPx7vjlnQBGEB/sxVcHrsFy
DVDEno3BWWnqhmiurl4QGw4EF+5cPFLnC3G3v5vA9d7zMlPz+xgOSP74l5qnvLlN
v9UNsoTBHdaiQPacaSXN/mD51Kc0Bf2g5v7vuuw3FCdTWIpipz66ryQW1cLTYCSi
j/ybjhMSyAlX6GoD/Q2EUBwUpD4iAs/txZ083voUJWes9KLwU1fRJ8NABsKhr0GY
qpO/eW1RgzVEsaxS7w7Vd4ptgOxneIXxREenYOJgC7nghbemsSNJGVSM4T8p+aiR
Hoiq543PaLW6olYeBa/xR31f6LNtS75bCyj7LPDWpvMMS9A9Hcu+Bv31aqD/9bTm
i16bOlIFdnYCQ+omxqlCfh8ycCTbZmiamnXH89HSBz4UPGCcgIuTAl8TkR7AnPoD
qabzfK81BK7E4CajQm7WBWVPOSoQgi+LY6C4/pWzu/JnsBQ+T/oNehZW+3D9F8F6
8xd1yERFd1GcnQ1982jXt9bqh+ePv8XEQ9FhGsHZnA5P1EzVGKxFebgYgqeiz0ao
pE189BPGND3KX8vtv93tR9iBCPhPf8T8o+xEL8d5Jg9V4YM18qaU0EbUqkH9IMN9
XFvZseiBiFjYzmQt/ERhOZLKkA8soezraGF+IHm3QQH3xj9yGQC0V1ciR37mnM6j
+CpLUbroJwfBEVcwj5dHP5Zmvv8ruULxouknN5XXNYSq6SYM+mMR0MBoycNrUQyM
K7zDJdh9xgHP0IDjFY+N/GVaZvjk36hFmiRCGnsPrWdwr9DCJMmqq15aV6B8Tv3L
YV2HAnBph23GJlsvExwypaPgOQKtCJxI/jpPMTj7JSGsH34Qcl/lY46vI0/yCkDP
0mc18JWF7s5J/AvimVVNVEZdw11PAUN9k13TE6lHvKNIow3D9Dn0b1HK0+LBRY8T
VzW3mQVHmZLGM99s7aslB3BHmsLmquXlrJ1nliMFgn9B7L9HF/MQQ/harCa57C85
mB/MuaWoVy7KihdJNrsIbremYSXPX1zH221caTRL4h/HAzrrSjMJiqNFgVFMn+vk
idS7jE8xGwCwUF6GFSrfKD6MEJEIhqcrEYkc0hWy+rcuJ9sTe96kuaKn1THFw4EX
WpPc3LwGXylq+AyQgcUBCiOg31gEtbPuvHVxJZtMEpjhGyQhVn3qF8hWMsLj/TKo
fp2dom/Gv3i/um3uL4X9BAr/3TDz5xQ89PCfvkgLBUUVCugq6VMvnLKu1H2YAVz4
I1o1nbr3yYvnPU4C6y9K2fgZAEpB57c658P3XbrHSOLYOW7XoN/ZfL3wywF5UIF7
RZvQBbteMqOjqO3eeeWrpZEGqpgkJ875tp+AhG3vIbRCbnNC9txTOIAkNMGi/R+T
OAlxGEuqMyAoLe3f3KBEWGovGF+It7GtBIhSFpU7/b0xh1OgIZGZejRpPqr8Nn6Q
eG85PwwftyNXo6e43V9LtkJQnvZFXesfKgqHyQa+ZjG2yAN56z+C/uuNT2zjMJY6
W3ayoF/B7dqCMxhi3sFFCfHZw24GKw2Kf0klw88PB/jlP0GW/ClgLxBDFQq5DpWz
b0lNHkTXoFqycV8qYgJga9RrDdVOGpnbmWQ4zf1xk1k0HrNfyS5DSlPLXEF7ppac
x2WrwXk2gnQJqDouX+uEdu8mRFRKHlOnMqK3JWfJoHeR/UFoh5w5HPw7GSSYPaoC
HObl84zhsmLR/I17pQjlJm+p00FDHjpMYrNEhlOsxSNwnwfKGfTwkUUlLvdqmmo0
gO8YSADj1Tv0EEIN4ryuKhNtlwqWgDq55+HW7Zn/j/zSO98giMCSLRS7g2TYLwki
YNy4ipxnGlqdwS5BuO/qdMj7QNKkGqN56LK0V9FTa542TXbXvfIjNVyyW6HZrVSb
0L3/n6G5OUiy0FNww65Dhw49IjsJpCWkRrwakkh7jNZl5TV/I4XmOzDo7WFa3okT
U5tZFS/YcQ5nh+W1aL5wqGeBf+RIwKU959vLMtN01O8OSf57zWkCRrThyVFFf0ld
WexicIwyIVOJZ3/TJ5sogH1XILh/d3T0dmKTtqbsGQZrb1E+f9JSB0BxcseXgwnd
RlxR4PbCt+dy808H20iD7rYy8yFRpyjfRcGzgEMoUpYmgtuBvuwuFjKg4iHVSPRQ
I6/jfmRuLwXJlxjlodAcM6QLRC+DQGrarwyLjQt4bw7g1aYsBeg68lwdFRqr3rgC
FrXuFZdr7fRXRmYRL7p3iyXxW1WjUM3sdCROVabfVAkitq6IZpbJxfJbR8hTlGyb
puaJOpk7Gnlbw4O905b45VU2xnRZNPf/lWpErSbxvJcvO62l8c3d+xYk/rf/6wG8
wL1L7byAhlMt8u9KcOw82wjOadDVHIX3yQoQ6vAvdkg/vUuscSAs/dIv8MhQjSrX
gxTgMzgvuarkY2nhMJei2JMppRGfDwUgQvHGoFTKvT3yTyiGbX/5Wv2sfP0V4bFq
ZFR2Jm+5df0y9IOpmNyCruPH/yNv0TgwYd2U6npcpwbJI4GjR1wN1MLzl8W5W0Wz
yJDgPtHmip3jZO92gW3e2BBHganeLfxq/a/Al5eYOzlaWMAcbtdptiPFrQj9H2aZ
I9D7YJAQreJGA6QyMYer0ruwOLq7W+Nu7mzeQjtjYSN7YkC+5z7nyMgWyhufY4NJ
beKN4oRvqb+LpESNkFKLdyNwwwG8NGWIdY3PFRwiJq1GGOpYkYdZaz2rFAfy3LLH
k5AVuJO6WHh2DiVImVrbVqCFuIwjtBi0j6PkZVp59wuRcL2h1W67DzDqHJZkSuND
xbrd1oNTIjsEyAynRdrU9eUyYagXd5nhsL/9A0P+DwRs40rwIrX9s3lKNJarcrC6
FXlbWIWaoC8I4Y78vFdf/dmtZ9bAHYFe6vmcbymnMvqCnpby++5aUCWqBNPwav5C
PfIBj8V2Y+dSGmOcS5xmB6Kb6kq03oTdch/5+8BDSqkPhWv3F0Ho59HuJTKHETdG
97WRSlNHdb2t4lquGQPC90uLXGXqxtrLzM+7vqzlOZZt8bwEtKBwzlgzrRd9B/1+
rUgVsO1fBuYfy0DC7EW8Lth+0UEtwXG1AH8dazGG/xwF8A/Z2tsCbsrsmNF0+9Xb
08GxFUmECrDODE+48/cyTLNYGpkTdftQbzy+RyfJazKwCFFmDZ934SinyqdcVuDX
WOwg7MC2uYa++JB/sQymeI5+tWM9wiV7EAm5OsqAHn0AF0PYjlQ+dbY5jpmxZ7SE
JtNMPTfUla53PtDKkYPXh52RUx2e2Ruc1ck1aML199LDVcSFOW6zZV+hF0OAU5rC
4jvegwKEckBoehl0+KS85KSA8uU5GxijpiqFahHRqFlL14ww+OnmDJqpEnjV961Y
Nz2Oqz4D0X4WjARVI1/YC3n+UXKlf5nzK2KA2YLn+NLq6w9bfCLiYNtTpkEeBfj9
9TAzBEatu3q0qur+/av/NXZN8W6FyRZWHjhdREbp2Z15GldCmzN3dcNFXXY73xiL
43ipNFxdRDdfWwFx7DYcxOojiiYD4lt6dvIHlCrLE6p+lleyqEcetzRbHdZdVYLM
Os7240cU1sXNzFcvJqIV/lEsQUOForwXX6w6NiCUkPrB1DPWQ8zfxglumdrDqD7S
V/3epkq0HL1A6XDs3EZ9IlpbfN3zBu6sA+N8TTrNPykuAc7Hnin/qXqD2iDXmJ6G
SPLo6pse6nX7rYAfXoN/Iqjg1aCIRuBW2srR/9e2dBy1e4E23sfAGpvpCYh4Lk1h
bHBClKAGIDuT+8ws2OA1jEfCJUqy7RG+flDQt/iHYYeYkFn4TO46mH8a8/ver8uY
b9waGh7QOQyYxXQdAg4cL0XaZ2mcNWTJg4RMEJK9YUiCTF58ng11CMv50B3FONNv
+HYWs1hA0qym46ZwXwrAKI5CGXAyF2h4SBFwhp3zD/qYt33PBaicgKQ6x1yLULH5
xqixjXfRgf4edYo3HNoB668eyGnNRqQl+a9K1J0gg87sNRE5E7UNoyZBHFGVkg3s
gtE0TN4iufzakYflv+HlhPCVXlqujKWtGRYv77TszJl5faQL76LWtZGEnt9IpsP6
FjWUZZoNaDO3tN9YrKwEzFoQUha9ZPOkO2/0HPWxSZkoeUtpckVjFJaYomPfZpKl
GuOgB32nfqjPvZS1DObcYwhimmJFJr8Ls5iyWdk/ukTS2KTDeyIbu0Gsa2/yr5hD
2R9SyIGKU3hPRR7koqODuN9CCzfmX8SKwd8vJKsUvcmz/khyyeJGsSvnhSEV8agg
+djtIo6ZugsbFj7mg5YKYhWql7wlsDMP4huGjTSjapU7L0GMYxeGFTLrfLiaWb6k
bJ3T/F89hPmsT2Brysgy5Zl4xddxYFqQ1oGb6iCM7nWNIhaKDi7In7GGseE4a4d/
Y993UMAZ4WJDvo8I2cwUdjTgx+yHFoTuxOKh9kSVoHcmixip9OR3UGomWBFtvl5c
7T6WdskY1wQ45IyVbpvr+aIQA6BQWvU9dhkCWkR6akaYigvf37cMh1pv0UdNcec3
q/oHqclTD4h0LGT3Msvkgg88AR1tOTxsdMFdGlpjvcbHy4JuPWsi1EccV/SaRlh5
L/j14zxGP06HSiNmnD8Z7S4f1OHVz4LzGO2MXT4c73NrZxpVIt+76lpoAaoWHtJ1
8NXXBM5GY/a2O426ljRaJTrfHMx8drYNq5YpNExskRtBdhHWCBmzBo53B6eMZJEx
iP1XZL5Bh/qK1Lenq/ruwpY7bcTypxyzfx0ta6uVu1XAKuOow2yqqLj6Nysrg5id
kzsDgM/44uMtPdX57lX+U6dh4Nr7nbXl0fmlxknOPipLbHQEmcZno3AqKR56+vn1
MDaCJTieKqANyj2CaJqbhkKLcdeFZWlyPkkpfnX/kLsLo9SNg/01lotWoIM7MHBS
enfcvR+0e9yDJgSnqPFUYPWQAB1UjWLlkZs0toOqlDbIA3DPboaaKEbWokPhkfJa
y6dDEHHgswqlnQWHk83HwRn1QzV2yAxvte/vNUN978+GV3hgq8+nEJLa36Daz74b
mQov7UQ1L+7hquyU2gcwfr045J8TlOdCmhzGlApzz32kT976zRENNz1C/nIGc74r
Qig3Kbpf1IC0MBs4AmbZsP1JQulOVZoD+MLt+v7R/8D/FtrhEHmDBUmrUT0b5vXD
04TGBaT9EAFjqWLhz6tyki9NYOBjicashxqRpkr3gk3ftu8SsomZhTJUq0LPpVHh
TiM97fDCyMtB72jp8eLCxp/a8djftnAmzBznYxj9TL+ph2uLYDMN4V3DNiPfzEGx
pxwHBYi3OagTl2bj0+H88qT5g5HyYrjY7WvO9xfa3DUabQTKlGmdUcA2WwVPch1l
OiiEXHPe0//qYtw8AFU47ox2SSmb7G/VP1oMns7issq51NXAWfmaooAIZ4TGurkK
VmfA+HRvhFlyiR+iLoPtvD8/4RS0HvTdLPgxdzJNsL64EtI0YPdgREnyHJ49/0K5
oi8XfHH0sIqK/7gfn3vaSFxOKRocGIsB09w2W73A1n0u8OFr8jmal/aqsL9Hj1Xg
fUW7CcPFGHJYLXn2D8hhMMbxchbh4gLMu9DrXihH2m9wJb8L7vr3X2NgLU45PZ0p
fY1PTjFtv8wWVVdpaLBBFbECmIQRsVjUU7tYqwKPDR6z/bjDxTWi1lNUOz5lyH+9
wF+dyK/nPkIqcokbAWQi0B6sPScC3oedQJAlIomPLFnfGYifmq6d+ZlW3YMl0+NU
f/E3ojYeSgQY/liNEVPWvPhTlAW6HVp1MqAFSQRflB8p5wPlerRsfiAKOcwJceMb
iybH/nQ62tgtvEb+mnZZQ2DT0QnaP0EAKkDLWu1JHXtW8CqRql0APFW9wGYQuH7U
4M8JaoqgTQgWq7GTW38FoBNCNaKypGpbu4aDF0KWEtIzb1i4pJ29OZPPLJlLJ+E6
15Ceu3w1L6mhKmv/A0dQ0IdlxmJs6ayZTcbj0yqeGRQ0IjMSGEdqskj/HH3vDs3w
e15uLqO1+HMAfHKfuX0l5EKd7y/sU5om61GvHoyDITaXxQhjDa4O5XGerNvCalbN
V1xUszmzHFX5b2CI0b7evd86WL58GDsWlwo25Inagnwrxyll7OUVuzkSvl5LL9YG
voWGnV1zRZ7NWD/UaO66G6aSthVDfJCE4lQInqJDf5Yg5PLH2V+XqFCEfo033eDj
S+2uoD0IvbvKRSSm8eMZ5ws5YpXwAFBJC8JnJ/bN6Mu2QBo6wTTPB7S9WtvJmpSR
bkJU1PludnAfCHn4mY9jDiIoIlylsMiuyFWN3soR9PWLXRR0MzDho9KJSkH4IqR5
n+XmizYbrsLT/C0kR2B3KNzpvWZZarA8o9H6597I5elbkpjdYwimSz1jfAMHoug6
MhmpWCMOTLnt8Pyb5ieWXfxqAnUrf1PcZC+SQpBER5q44FDXUAygAC5P/vmktCsk
AvQ51NhdUN5rWfnByk9OP+B7zsq93srvBvPLMs7U958l++KZhfDSFyYEA+We46PY
yItG/sMD16zycaeMXX+bSBZRHAJg0CmvO6MMlN4yJNndOGYk6s7e8aKmLBPaa00H
wRUafVNuQb2nafC92OSFGOkzevnam8cxdzLUA8TOi/GSEC0GS/CC+VJ8HMvGQWSr
ZrkiZilcf70zVeObCsD8RA5tTSz+dWdSK+UqjM4+27MxyfF0/cWG6JSJ9qRF9cYG
pHWWnoB3erjbEezMI3LpBD/XBNq8zjXikYVdzxprbCetLP2GdjePcDoTL/FE8a+k
vUSqVYkZaKHa+k1OCrTDvyR4dazF7lnzUVkVRuZOMhEhvYq4Q26IiUvbAGQFUxaf
QXIXTqbwpZDzphD+tWkjP0uDa+Lu5LCzuiImGluoli3zrhXfIpRG3iuPlaqFRSIu
cM8QNfWVIPaFrn76vQ5vu5Rt50tFqCqsu9eF6FvRRkDaCODUvZOIGc9fi7i2KAgg
I+6ftr+3KLqoJ6xhNSpRjXn5BVoS+w3WQBk61zQONGbbkgF88MwkJIiWRDB2t4uG
GRiek6nxwJL5ZctXl1/fJFaUmBDDOVGrq76AjHRNFXp3EKbpwKR25HwG+FSto/nO
vqeIgkuy/oO+piXpQYn3rMzgchGpp+J+Ss96Kcr4dnUCujtZRwypwGfCB7xTYeAr
LEArlDy2StAq5FV6OplyjnflDCaCNA+EP0199NdZXqgCd4XG80ee8tf4mcv1wuve
zzoCAUAf++1UAwUjbIB27zmPAvn4mzZcIKvARWv+f6NOyUGpvMnulNctmTrKTC93
px6k+v3HbMMSkPD2BD/aVe0rMPodrfIezFZ1nGBELi9tmjKOybeBpudvUvRerHQN
FoFmp91lWkdsqKsQIwFqHpNQzqBzKDT84ZtL1xbzGgmNqStRaWkkTKbZOQxCoMJ0
uOPmYqV2NjyoJn7FlpvokqnBqugaOJVlifh4Yf8lXaQiJe9tBOlrR437P/F+i43Z
FfveONHUjhFTI5jfNDJ1v+HCVFl1YHe5dJmT7o17wK9rNfCYbYsGTkSzYV+gzGkb
0nWyuULi9YSPWe2aHMcol6UWC9H21mJrQcpNZZ7oYMw24dMRSGdMGX1O8En2DD3g
hd2tItCeH8vnptKpw25kSfa0s9D/P8evWjHslcz5Y58eIYi0HL6exsVeVQ+QfHDw
UWJ/bfErqV1z4e3iP99u++/94D+eH4vs77lKAvJuhq0PwLYME66br7MagkECNNDy
k9nO9SYHLulb4ex+iwGj+zqnkhXR0chhZuCcuXAYSZRg8MmRCy94Fi3APQVyCrQW
OKIUOwviMkOKZC96ib5NTGGB9YMrcnrR+AWQIIqJqa8aC/FXGkLqjDaJqhAQmqQO
YuP2c5kuNDBD9I+ayx6UEIgooKlJeKdMAEuQsCcl65Gc1q/9yJJpoKPbxPu/+soB
/oVZynWAHKICiBm8wdmPQtr5DsFn2ORBH4kB1Lgot8Q3qQoHOjDGR4v8TwvaD84A
iWpAOEQ9Ox19nszTCGUwokexHF9sfxlECZO+YVsxwZNGtC/4EHAAwdk54BYpx3Oc
Ma/cbqVKQq2qJSCEkgFDwi/CzWmvr7cglAhakswhPC+M2uJ33i0QQh0Ng1Qv1Bn+
G+3tSyd7EWlPWm4bnAE2oL4cRlrobHCIrrmG1Z7XHpWv7Cpfo332FObzt4H7bdoe
B3symC3GRFiLGeleuJptEKbiUJ24eq+h/iK9jcfL5pJByIAea31irmmZBfnkDvtj
sMDHN5kagB+oiFUMk+etulv8UJplwily9X731dYacsWt6VmDMy7JXqsgKAnFQEdf
ZUedRYtbzJuPmahoWzSYOFJpMiKBVqDP8L03PLtVFQgVTsKuZ7PRqX2sEzxtqP4R
IsK8ruIwrdQ4TisZaJKjrwe6PFm4uUFhQNiMPZNG9h+U+tERCWGC3qoOVd94QB++
vFOqgDoDkF2qcFU/D4U2cNe5dPJD922ISHa6x6WLD1VNKBxZJ4N61L8eJiyr7Zxe
Zdu/xBOcWVEL7BidTlsBujR7PAvEIRYkBk0ZUx9Goo1qksa0lEknDUlfDRw9lFAL
nMRAUZdh5x3e4REepN0SWKms3DcryOQSRT/bbJNtObiqrfUOdFs4EdLl9glP1BVJ
l1Fh39EoOWN23zEPUEQK2Sz7DY2Kn/al2WAlQHK/bOCTSsOHvXDEzyIWKXXQ8vmL
hePtScLgsfCzfmxS6mQseuuBP8vzQMVzwVkAcS3Iuk/+s8JnA2k1AzCQJcnU/B+a
VBh+gnox7JVwTDVYMYIjoz819BW4Dtb/kihIsmxbztfBVcTBdJRP0V3Y4Ci/kxh0
Xg2aQJkZtDU2GBQJOK6mYIToaf0gyw3pLlTzwDma2396BksBE1yaHbkB6CQ65Kxl
jg9To2iZJ0bHHuLWrdzKfkjr1XymnQzxr7WLkVd9bHJnWGeHYddqB0x9TpQs8UsH
CLvad8oHNM1JuML5LK7oKxLCDHNqMeSYEEnY61G9fjBBaptfx0877DahJWoURvb9
GFnPrltosuaeIcFfL6VgWuKcBxmM3G8a7sa3uNZCFP1VV3QPX/Te6LURSJKt5/qI
q8obCkPkTIHPSesYuUPu6Rojq450MYlI6k0OpaEDupdraDXXbcL9s5QVJUXFy4Vi
YdwUvplh6JO3PBAzjdSoWd1iByfMAkJ1Ou6W7K/0imeCcmDbQrV2emcqFhxBGdl0
Oib2VlWpeAl9LTzkPJUmB0oz3JNkE6BiiU/ilj5c3SFbequrZwbK7x3to0py9Ksm
dwcP3tvEOWi+Ksv8cWSBEticFOk/s4vh3QCbgY1vjKl+zWhbKujscbgHpqb6gH9S
9APtQDrIk9kFjrUmdxcFO8gIoAQYPyf7JdJHofkrFFgkbhI4pLnNMfmEHJhPPi/r
A403q6hFwoYl+Oe9BGBVfrMqFMIUIiJzYhfIyitshnai35SATt80nuVC2KoQLzRl
s1S5WkRnDHnWWg87sS0Ltbb6cevdWUV44y+zuxeshXQfJ7c+pZ09d6WwRRJOnwKu
b+b86t+Q/dixZrIpWjs+tdDp+E6QHZVGktyT1svD8iJ4VDIZafDq/cxTJOr0ij4f
RCbzWnEeEBNmwyg9XtuTfYedyjabKhf4XZS2Lt/ry5fGr9hbhXNPw/vYbO8+Omzr
KyL8/3+bz4nBc/wOMu6gZ/9ujaXV0XrZSj2xTU0BGGLfwj2wDdUPI46wrv32oPhe
WX87SFOLkAVuLiRxwJEmUUB9RmFxBzwfsUWnRx/gtrqvX6qF0HS71Km+7XGHRDjA
EMph0K9Hnvun+l2e2B6UAfoud+O2wJSrWgE94o6GK0lUwAlLDAhdFuvw2rS5iG0+
JLcrIL2Mz8JMuAws+i4H3ASDCRHRoYeC/dO90kG2wIPZJQx7EvifW/wahyv1fotC
dmURm1b/9BWbXmb42xQZcXieKGW1pF1K/nsL+rBHf+bLcJPPxdsCLAT9+/bcIk/f
HsTrIRr11b2KRkR9jLJYLcGhVhEEg+7zpZULPgFOoisp26B6ioqOTZwOo9Z4wu0f
HWg8HbQWmXZ9xOYZcMxd0t74sWlRdNARAiQYR7pYQ02JS79afEwTsrvgnMIRe14J
Iw+LzJPFZr2uyDws/BHvUbMNRHe4/zSCjqJMbsuaBFYsl23w7bh3qRQ3LbRibFyy
ZjsyS0T+L1/+/SzV6Y8ACzTiAtxdsiBe5fDl37nxLTbfn48NoLKdvlapb0pn52gz
m1kYK/EicnXN5AfEOHvS7U7C4Fe41INhHxINwjpHYmAdWsTXNXdHKn9vB4PCLez/
72r7H+3YPCdIoSQnrlLxQPlufmGulh2L+aDcyL5W+LqI3TMVrfkTySw93o+wcJt2
rH7asRgOCu2AtWor+1n5wDTvsfY45Afng/aZ8wx04UjxNoz/LfoIO6UQ64SIJKFb
rnmtqPpK7DY7gV74IArJ2Y0YaBW9Zw5zRWgjGLbhQjqzCdBibNQrKKD8VrpHQfo9
aq6Xg4WO4GQFJ6/PT+AHn8bbh/XZ0Oo/DlfMhTpwc8bufihAsqQHRiik4OD+6MPY
nqoGPZB0ltJYDxpDFFrmYtUgyh7CR4VBdm9pTNkVeeuuqUUUNfXy1SHu6nR4SRBU
5zMFU4/58hKs5PsecaCoNeFNbNKlIhwhBRQ4t3WT4ChxNY1AaYZHrG27f/JKWF5B
FaVrZ/82emZV5SW3g2+q4UIuXQ/T5D1rWFnMc2jkkL5L2/WxWScg2jt4QBMoUZK4
i+VRI6EVEf2Bf3demE/FzwL+2IDg9lQa5OACQ/BHaz0Yfoz2MxInVwlMkgi1CU/l
ZdkkbMcxoHKO48x5Xozzd7Fl4h0noQdtB5rYZ3DInj/0ogyLrAZa26voYsCHFKgE
rV+igWobkVKndhK1Wax8KIJ9Z+3Sy7HrYoo8Vdm9sexkHEPifulSeSosyDj19Ob1
Fu0tgWGgcFr5QRYJLXs+4I6b2Nn4B/aY1UtEhq+dadfIydxO5LgW0CPgquwp03Zu
EQm+BNhpVTtMwCBynwKPnosU7myL4nKrR15snLvwJfNhjTcyfAS2poxXt6vsnjLM
IAz2pBnD8p+1BS9P+XTCcmjR8LVBfTkWYmeCyfr801S2hYjhGRqlrqyPmUGf3FBe
d1Hbn1KBBV+jHWImNnss9/vZ9JwAAs1CwhyPghPSivWmG6l2k7OPgniO+RRFsYE0
iojrWziJr1oD7U0/tx82UuXdzfR8eQeV0K0jCT2SsGH1IXTugI0Z5ctRnQDoU9tG
PoyVc/tanFD3U9gJhrO8NNXWtqvJP9tEfTtgP61Lj5FAxHa2norIonLTMJ0HTmTz
uOdlAvFMd1yZNFj8a/ubjRiIbD7zXrlD4D05QjGzrdr7LER2s6cG3ZxkN8iQC4I0
ZFkF1gL7etQftv9wgyyKYJLOqRCsO6sPH+HmnpCqp4ULERcg5K4qOX0u/tJn+4OQ
C0Gc+xzwHKhdyNv3cywzHhr0LwPeyPbjmzYXy8i5YziMrrdhCRoruT5m2X9Etm/a
g2GquLEam033tFOe+lkroyELqBRhw+LICKuUq+lRjHXsUwYPb9E6oyOJHaFzPmUr
+UHaaQ9QE47iXL0IKjmXuU13awULtZFzBggxWXLSr3+X7h22RtuB8H9pInTkpc9h
2OyPneTWwMcemHQuWwRfeIriVTKh8nHpqvWaiV8XcsYUFcLW9RC1kAvzHJmwB1mr
1wkzuMV/jFJl2z1Up14CA9PWLrG9MEttqymPMC86L9+s7KrZG+XtDtd7gDyyXfVW
D8mnSRnb60zSRYuQ14WvH+v5qM0DSnoBsS/Rcm4cbIiebO5wUcfbsZDWVbbFcs5z
K7SBl0VF5N4SoI3EMOA+c5V/+OEJn9ji5j80Y1nfJ6lPRuwDDJf9bg5stg4ocMfq
Rm29HHVvCDokDtyF7a5LnWLRj0l0N5Veojm6RyJN2vdwUp+dVbNZV+4HaIyUyRrs
ROR8H5mXjOBrQQXxjK9Es8teC7YOdGQBaRvxeXXRCd83JPccUA22hQBE4t8Mv28F
KAx81I+N+S1xwXXTENgxnN2lVCF3pPmWyX2ee9qMiqSYMhkWot7WS696oeNorSdE
x/TPN20TeQXtw0CG5NlOjCpWPOnledTH0BH518Nt5oJmAeYDBsCtCAApkz8/6Yry
g4609El5jUIGCUeTthBv4GCXDUeSQpvNM2G8sA9cbFblGiN7RmGNXZy5Ak4C6+zL
InlvkEfLsRCnZEZx2u3ERoF3F0TfcwbLAqL+/eCqx0xZIE+pGYXYXTPJwEFfBPML
yNOO0+yWpCek7XeAq+jeMOKZTw9P4Xp9B/ebpNi3iw7OqEudQF4fIoy/wrH8/t2O
Fc6/JXmTBmzo+fHlwJmRLsPStdiXIYH6vkjB5+xATqjEkNxJlhu43Q/Qv8PB+Fn0
UVfTcHsLdx6ytfLuOoLtOaCJglWoHntECWR2SWdum05ReMPXzfJOWH56x8IjOnYv
kAiyioGHqmtakltlHDLblFXZv6xgB+OeAcGHocPA5nuYKXaCu3kAk4nuJVECeEgP
TiItFxDcd42RC5eaxW2EEXn7vgwNSeGHe10//D5n6swz6dVt/XGLGa8lapXJxTpx
BJfdel4+WyGEm/mePh3Z9g/EO1uSXpAQF5QjqvV7phemfKaP9risDc7sft7X6qgS
i3aYdpGUICZnb6JBaza2qd+nHNs2chvAsgMl3kqAfIPCwuOA15eQLDHFaiKq7BSG
t7/bFkKou9LNOD6tjbr2Dn65Q0jX2lULJvbMaVjsxmzpqdeR5qkKIxoA//lkLbmu
OVgwG6515LdEWlIySGABHW6aLUICzC05EQDCQJmqCiCCAWYpaE8uklKYL+RQZMll
3VAK+Z+9dZ+9Eb0mwYVT66Zqzj5YMFFTor4TUF90+tQwqo+HMO/1GYKNvs2RG8E9
5uuM14cKNvU7w9bU2xOKxwNAVRnKeXp3IfdmtvcxBojW6yzB7RIvp0PlKKyo5HCC
DfBXZiyuKAfAv3XmnGg7/6grM8+QLcDWtFuLVzZhlXgkaXSL5w6gJXscqq7pLOF9
q7Tg2tngXLC7M8BhFTU3cQthJ0KBbrVVnh0/+PD4HgMfPy6svcAkF+2ghIuiKZAi
kJN09ncWLnEICxfoZvGCHkSZXpsZ3v5qRgybjY3w1c8D2t5InHSEB4YZXCaDKFbE
aB6dhwpk2Z6rsG2eipZFVuIVQURfPERKuyVJo5MXN6WPc67poxnp/eUia2Vx0Mzc
hazcFakw0MHQhVw+Cle58HfijXpCztb4Vl1sBjOkIAnwRIZfutWV/8duMN+7o+5D
RpzlCLgiOuUp+rV450k8wv0SCnR+2ABV5KjF7eegnQnCCthuSpJE4XsV9GlZ8EbT
Y4O3ZtipLgkp/E6ByF1BsRbac6YLOgld6Ftdg9DeYkw9fN4zNnYBYCrkEvfHxg7i
3HVcSA1//OGCxzg6PMxTLLM8C18o9CqD2W3Zllyivdp3WGtmBQePdI4NzCUrD5qa
Q38/A9/hd6mGhkQ+WthQgSS0OP1AKrRu3ZbIcjs+i5P5QfAqvUpWjBBgqwc57sMc
0kdMS5Gtr8xMzQNN+Lt9Om52v5qiAttI4NP2v5NBd9WgSdBW1pPy4I9uFUpARXZV
uVn7HU42d/QkHazXk//JLCipVMxxNEQaZtvSDj8D2ge8krzmcLC9Q+zn/rilTQlk
8ZBvNiHQkOvC6O9i5yfe15bt9Ip8Ik2fCi+CHESKXij/JoOJ8bPJyjAQIscfl5DL
qwgor4B232i2AXYrzPIXgBEPMisXTXw4XS7AeYnFwNZnTSe2NkSX/qn8Rm05QB/W
tYLQm3Nm1P7rbfG+ad0GcH0wy7NSmXk/1kXL3fvjVqDTW0i4ANYR1sks09dI8BYH
YThZMTeCk7fCbG13pqi/Oci8/xhBhi038+SYB6virbje7Jy5RrFoUZVQ3qHjaFba
HgUen95ueEkhmcnH39x3CkbGzsCLFMO5ibleccSJh0yEG45TEoDYWTTK8Cn1Hdf0
ORxLpPM0yQdZqpB9KcGWY0sUGkbxtDCDYV+u4oOUaPAh1/Lmo35uGcMVHecOaybX
EqqAkrpbloXEWbpTsDFyXKGxDDK1jNsnr8sReP8u0WKrE3QC6izPTVrOBqrUJGzS
rJkn4ZwHEwnaUgbUxknvYZgX0qowsaLDWZA7NmLG+kAMsJi00kqDlaJ+pIpY4ce5
7O2PJdMPLdLomQZFXJ2iD2nsxUsgdWsde1Tg+nO/50knDF1UsqrPBzSw/cOZ+7P4
nR2zMiqymXa7qaeIUXu/a0HH/vN+XcITwxQnCbx162ouXHKvdcs+b2L0OoyXjfF0
YdL4eEC25nNPilX3kIvZFE6xIQqLjb63sq3nQxpvmQThnqrYjiHwL4nzM3aVbSag
yNbJnDXTa4hBMc/n9EqBKWt1Q/H7TD9RU+aJsnMRZMLQtnhvlqU4Ep17/c42dlXc
aN9hzAyZ8sdpsbYpe8oh/D67u3QQrU1cZUcPp6GCGlZtyoWWvtRTi47ga5zlCFUX
ScoQ5mx2WU4p2E8aysnPQQHWQJ+Q08blXgOLrIJ4NQYsuUfvwKjzWYAMjuTvJUM1
uaiYM9/w47Y3h1isxY4bbeuSLcAER56Vl5BtoLO3VbMmGNjQX94Cd2sJe4ZAfxgC
FAZIbRKJoPYyMkfCRZE4XBt7NGorLbjZbkxAkD+K89EW8/29AD7PVXy3RHGCbxmB
YO+KKzlEEB8sPJvshR4Uf3jViNRsCUap57+3GQPIn1/fA7G7uP3000tu6b7v725e
S7w3NihNsW4Ap2VIU+zHRePIlIb42gpSFpWujspncBPCscDnbH8u+HGDMnt+Jhy9
EZPIiMU4UG0JBzGMMCw+Cbk+T+Hu1pMqVl+G21hgqT/wEHqer0192fKjyHgwvRPB
v9Y17byd9PvRFbIqKeLTCQ6GDqyT3blb12qLzFTTo+ve1hLhV0JrDmqDlgChWSQz
XiJAC5Z6Tdf8utGnDZmI2TC6+tOqd7vlbmmhc7HIKeZtcOWdtDX/AQR16ao9woCH
xIoCi7/zErvF39i1CV+rnHfaSeqW18Slx52JZ1Agibr1daZTMO5OeY6WSoibr5eS
+03sAgxUNkyRoMa1ZzMJjznYD6iyG1EERrYMmfPNOib1n5VdfsfeXxEVMEAsowig
lSOcwjyi7YBSg19LRCPpg1es5aYLeMJghjvFTX9uVnAekk8OYiDQUDdxNu/rwkpi
KG9ETQ5zeELRDPVHTqa6IqZ0gzBs+gwnyhQLt/PLunvw+ci0AwNI58t4xWMCVz7k
P4NQ9GLIQfHd8pq2Pfv3Rt6fwZtg8WVLxb3xpGSchpo4jvGyjhjry8ggdUtQmD/t
JLjPeMo3bURMatPVcxTYG83sXaiS2z4QSRPmiQhvtSy1XIyi2dmaLiOcr8Wj6stE
EW5/bbVZPUvg2pWYQuc/YUz7/ek6Ej7UVvuTlkdlpcJb2bvDsNb8ouG4GDYNTvwQ
QrWO/g2HSG96DablwreczN/st3YBieh7NH6iD3T3mv1QcGwYlofI5iu7WOBPgTf4
RFa9URTKrKfHDiN27+N3x2PchYw1FZFNQv3lCB4/+ctRwVKvg0U+fNAKZ6fl++Hu
uopb8Lh6eOqpq2Wc3q6NDDIeBT2HUg4Y3HssVchxz960cj0UXn1ucedK+5/l0dpB
PA0LDlhHEFVEZ3t2epChIE0wLadLPNQOYgzIj8nLQ3tDxKwjMBc88ZIscFc4Hdh1
zuUWWy+ZtocZ5XFf7aMTz02xxAl0uqpmPADN3fFHhvZv+ggCWGc8K3Qdk/UM0ZbZ
rdWz3XOn0os+I535k0YWOGNilmp9R92f0pb2sYtxPyuajpWzuFhrVqhBCfhWK9QT
Et1NwaKWub7JrCMmJplmpAh2u77ENeCq41iVqRClaQZUBRX6Nz5XCOjanTriXOwL
Q/0xgnUqJmrmagWrSpa1WGBvikvRNC3vrym8616rTb+DDSL9MSkBsojkcQmuoR5v
WCKm0fHb+EEleMe1iKhRgUqO0bJmhhBIJv3RtphJYhgV1ENBKJXRJOUJ0OnP/GzE
n0HUTu1NYZX6XDUiTeD/HRYwzdmj02TOmy19Jd/OV8q0QFmzZ+sGPK1Tc4VcPW6c
qSAz2mElcy5+/14B9t7+WcJZzrmsR7SqY74E4tL9CtdAbVlZ5eWzjz84ZGL05U5y
lH1cskkmgAlQ0K4CB9L5HnBv9FE0uV3oVwetFN1bdw1D1cd5XfURC1W6FQc0YAKX
nUWcxOs/GLZ6iE8kTXKw02h2yLy3uL4psCEaFADOSIgmj51tre1Q4JbzRHBRh6md
JQM27BJVrgt8Us+njl+9Z4yNegw13q9t8+ZVrws0Cse2FWSUXmqDZDmaCXzMukEZ
Z7OEEfDuzdjWjzByZI9mB7SkjpR1gxCGbty+PFaPoZcO0bvARjn0RlMEllot+ryU
5wb/prdzecCe+ZtuHKKfJESMeMUU462NM1Seoqul8TC5mVtfT7xlSDZq/JrRloiX
nZIeTm9inltFQ+ZYJ7EGG8d4byNRBtunPgL356YeBvPJH1tWQd7FOvpoB3emyGbT
UcleootXLbZ2+lwTGygICsVgQFnbkgDVJSSYHpsSf/KwI5rW9k2oWgECD7PZXuol
AToVwMe6WFcquyUo2Sxyv/gER1whyH5ydB0OH7X+jw86hLVv1Nbsf8eG0T7XNEDO
gxM3nCYGnUybq0RdiXDeqFT88CammSqUG46FT4rUgp/z7/skxXnhjUIelLNfmpXu
EMKLWbxTChM5RASbBmSfDo1gjTy5HGVJJUm49KnoAkZCfIdq23XFIiyMMnKK1Yd5
+T4d04lBDvWNh77pcOBuloziUoiV/tFYFZCtXyxFoPxucdvwFfUvr+CWacaqTr/A
jHsHTjyGTx691SoYP4olmZxmVff2AQrTJOgTuoPZknWsqn35HhEgd/iiv/ByzEMT
lZ7ufnpCCoKZcH1F3uS3EOmRHWbMhaJRmxr2Aeqou6agmBE3Yxwk2hAYdr0lb+mh
uMukgtp+YVltxp8dHdVZpAdn8CR6GyGW02CXfInM+359fntVftHLs2J9zkSr2pGF
mUUP9te9NisWHJbscvy+FhsMZ+AVNRLBG3iDnvvJW54T1ELBTlEIh2SC5kttj1b7
l0Aey3dLHCtSE4tKiryssGRcNZmDwHmMnp7rGVAO1Qg1G7dBiBtdoKIJXQRjSP87
y1Ob76lWj7S4ljP6ZkLgAScvzakVVYIKRc5oLDsIklNWZD3QzoBfX7dkzxWDvyTr
ru7mi/u084pTPp0HTR5X8euBGWnL19ZLRAXx8RJNeEciGNSemIAHyJXPm8/aooQM
bIbmxjbSyhRfwvj67yhJXChBSa7EnagxBXR5y/qJ89pyejDlkPoi44JPm4ahU932
OBR6TKstT9ZNeHYqg1M5OunhMKY97mkwAvrVQK1iVbNWJEEy86j5JGowA3QZwZ7S
g5QVHd8+Wj0JapQu5yG1IZ2rLeHGCyqgBq2+05yVLf22M4xQmJctg0avrjger8Z/
6FbIxUG/Q8F3y0F0GHmwVLulQ7w2zo/E3Rii4f2uvbqwopcojk99I6m+GpfsHZ2H
XZvrzRDMvWt9/DqoEw+bFI8B6SuRYKltLJ6XYRqd+KuNCMZmDmKCAedgqamSS+HN
oor9B+SMdVy5g/CqFyLQDxxZa5fMs3qS2sFznVHjjroW7ghQrP/LwhzLXgGSFBIy
GXztwZcadwdn4GgOjzCN+iYj0UcMylJ+TFuh1ox45PAHDF5kkwhEV6UGUjnABYZi
0yRzTTJ18p7bL+hStXFUY73FnbzKCG5+ZJ2qFBGfIeY4U8e+Zcx5UPMStq1q6pyN
hV2kn0gjc6ySxFhjKW6NfQoD2i1/urecUYBzwOe49ic64t+kQvER1M4LPvoWRQqh
m6tD12eTxgIOm4c2bqC0LMEhCUiHMlO0K57fiqsGn/EGt/b8Vn05Ofb2br5OAkWa
ygEEzXR5quPTKV8fQEQy7NqJ0t6oPGEBRMRUmjHcW20wq8Yv3K6pkRsgnZwLJByG
vz5Wp64A2MFeC4NGwvNyhckBH0R7L2hz5vliP4/P3VAWQatZV6KtpC8KlL0+ixct
hXpQkHFkZjnUiBOwbnRVn3Y3jgvpJda7JnVsQ0UeUtCMHWaOvSVpA0/RXlx5Wbkc
+Z3097tqpO/711rw9kAA5iNl3df2LP93XLrqxW4Q+SHjmbnsDMUHHSIBZfaUDYNQ
K1Jr/NZmMEfFVvNT1owa7R482yTqGMhnhwY/NmU1L1wE94g1SIct+UCkUk+u8C4b
Rp/JX+O7jKYcwJlO1Q3WPFWW9qkooC1A0Zx/HiR1jJainjKtJZnMgcZC7AU1GrRy
m7rK9Qgk0oDLrgzeqtASTYMi4JdN05HYnFKNcD8HDGE54QA22QPIqKNcY+2kgXbJ
om5KdLjNav3so70heaNelb2uGC/XsTo8BN8oj1b7VfdP7B8hbly1vR3RlnbQ7KCs
LX1s4v7hTd3YkDllO7FKoSd2VKgWPHHEG06mMtj/nDaQN4F1W7LviSFvTJhkxG/c
qI91lMsXqy+YljX3XOUh8Z+hVK8ED4NFeFTldRZ2mpa3wmPW+xIsyBh8IQHIGAUn
qtoO53FMHkuMUym57Qwrx3Wdh8a6F1OD5gyGtmkQ00UrZ+eJlrMa6qolKoRkpmRf
VK7yjfwygWJCt+KzAwnCyuAkaFgShY+EzM8pJ5qPs/XsYtMMsYxCL4Hj98fwHXT6
7pQ8MmFasCbdf/XMYIo5ATN4aI9YX9GVu+nUuht1Wr3eQ1xLKCW62ZylmzSoR8xk
CGB8pn3FxVA0Hxsus8I344H0rorRTfr+jtpFrDUDZs5+Wxgm9AgSW91z7rh/cMy+
tgVl5wKxnJltm43yGP5T1oGeOj+3p9rxqTkW+9TIlkVyMAc2y9SmICmGrr/2xoRt
5axDg2rZqVMcdxZbGug3AdT/GGiJmgs+fSRScWg/eqhM21EJwiOwb1oW+x9zeSiQ
PO92T/Fg4KLZPctR658jRzgJJTsw3HqQ+3scsX6qg1YXUhtzfdnLMMZtlJzAq3Kj
eSBLgukD0WpYgQ6BXoeS4RdTNVQKNT2Z5uF6DYeOezAYunTKS+dPJBKlkezm3Suv
5X5+85wDwpgYo+VV2xUdgJa5M8As3gAOh3Gi0e77X8hzIxLc7rsHL1/nEZbj6f4Q
0f334aZN3cQHYmRFhMt3EYwJqB9yjApy2wqKTreeB7VnPCaksjrvQwa6SCy11yFS
JzK+NWPiM9LQaWegJsGPrDneTvIE3xT3Y0T2oNoueZsQ8VbAbhvc9ltCkGhsrxnh
Nqp18LzzhssZRDpTYuRDknfhu9/QFCLn7jw3vgwcNUhNikuTWgKJlENq99NXYbSB
sLPDKIxAP6OQe+ui8/fQEYxtlKrEkLJYq0yVX19fsw4NrWatOphmcW6LgePmvSoi
PvkQCQR8ZCETfFz3QqjJ8zC01aFsZIh5TzTfyXd0B4yxiuGRx5QcBpQS7KYy9h8j
Xc4sgfhV28xLhIAkBsv3km2lkQqW8KpdpsJKg6+f8mafxrj0jOLBaflgCb6vr25q
3UFy0dEA7/rCEr9K0HhBahXUdJXZDXlgsQfQfLtVuCPUwH3Arx9gdoE2PKdSRC4z
tKkr8qnsRAlQicwaS+nbdkS4AYQp3yQKBeBgpgNKgYDWp2GFj1kxgyuMxPu/HWq1
HMoEtCqcyZnCGnJuFrVh4OIOTmnQUa0N5dRfEBbs2T3EqMrLBZ1X/P9kGT9L7jxH
JEwaEMFn2eTQwgQ2HXP+lEtLUhOOy7NMnAjtcrGUy/8ln/RHqXli88uryLIKIjTs
/+OMXEJNx3II0ebRNuUzrPxP98Rtu55T1GWxBqOYqr5faaWuPGL0U3jPmrkxoc2O
2culZk5SjqzW55lYWW7hl/8bQRihvkEqSaiFN1l5YWX9GXUkSxxUwBg5YOPZQ4WM
+nrBP+PBD2+DSoaD9wxmSAQjslFKTtuoVvK8ziXPWVJguDZSBHjdC3LKTMeDluMx
GLWFpxzdrc16I2MYB3qiFcCxuMrtWHNu31S74KVaDswjcqxcrrmC3hxXbCYPmPgV
xSc8oGzOSL+zT8msyfem1xPvmaDWwjm19Sb+nSGamF4OzB1+VZ3yXKH2YDdKv1cA
nYu9kBMbHOnULxVwZLOEu3Nov/tQoDLz9bU2IQKppYs8HXf61DY5enKuSS/+Ow4o
KjoNdJoZkOI31JdI7f7mTqxWDzqVmLt/9ApASSC8uRSJmfxxDZRViX1jY2h5Uu/m
5vp4N2WukC6XAC65qimNa2wexVitaiSam/Pmh1PifA4iLIDGFWavPw1KQ+DF5/TU
8sEldpquF1/4JkJipVoYktlRTlLG5dzMtINAbAOWD1AwmYL2LHiC9WgtCS2ATd9B
kWy76+GkEiswLbP+0m40Ws93MW3vOQUtjZ15sfBaqI6SyPcsQCm8VhycTRUtwFXa
9R3FIShcjxr5gvBB3sXoCWdFlcUQJXp9ayN6DdpZywyfDI2aquj6FVcjfHyFM2yA
une9prKyoJTqgnZd15laDyhxt9H8S8m7rYcObIeIphz30NKJcmRiCROVyycQZYFt
7kk8Q5hwLAgPZzP+mmq1hEZMoI8C54ej9pazE2lFZ2Nz+Q3MC42S65qK6/kStFmz
BXOa5p/kGZQymPA8znB83ftzHT1NMftI7hqs0ojiyqAdYsUnri9EnC7j8hh+CVV7
+v00brZbOirjdDDZB5kJ+AZ/GHdHdc4H5fJ/8SJASoCaef90oPfu1wQjEGyoLuvb
E09mmQBcXxD+R94daMb8C0XGvT9hBxA2pg967JuQXXi7JH1VKEiywuaiJEJqYeP7
r3JVhHZ2W9rqmr+zr9JSWEIhh1QfXqTyDAcbYfvfTp78wm5STXkVWOeaCZY4Tk+R
W5i1WtG0ZR3PwMwoM1TJki6Nmf90aGXtVTZDKohxErmWyXJyI3+JrEIU4AOJowuJ
h9DUbR/QTVYOtoflQn3PxUYyu3EbZoEl4sDY9pLBe1oPsInNuSisF213XJ7SHKX8
e0729l9/U2tyDFN7gPhdMJPi6ufz0LYMvSJ2ohQ2AdHmO2eZuVnfyTgsnhW+to3i
M8qd1qcxdNFIsvAnbveIJPm6uvnKZwQfrTAjre2BGRqa4WVfd58iG1SOSVzkGH7U
PwkMKHLvFrdllN4P+tGFEeMO+yZ4si6b5qCZAbWJ7SqayWviQZhNyYQRgTZ7v1eA
ZzV+FWBQjqSlnHxe/zKSt/cuXRcVZ9epCE5lEpj7/8K1/mNK18kIZ+2WoVch/KFu
4MUy6OTJ6zmLqFvpmXHMJQAMc1y+i2QShp3h5xtCb2yHLNj50a7wUZSUg2Oj8B84
EuCGDryZGouI2pTsDVodacMRLrz6Z0OoQKDyea9mNI92FiNymTT83rlaXbR5bZBz
EcuCtvhvl2q8X1Q3nG/Fk5/oxUgtGvj67Mu8NvVwf9eYCqQLcytC7Rk3KjZq7BA5
nDu8kOZ4qjewSq8qQ9ZLqKXJf7SNYCGQFblJpq6L9yX1+HDuzbomtNugnIVTqrj4
kmWhXT4M8GY+5+ObX1emgQ6jcKAVGD120fHp6lyXM386keaicl2QI8LFRSAfeKjA
t0NtNsQ6xRQc6xpRVH0u+8iliohFuIyig0We7h4VtPxQozYrbh6t3ofRt6cQ7F+E
IHYb/uBAKf04RO/WikQg/kNWs0Qy3gvpTPPcERgfQdaDGi5o4udL3Kk5Ld4Eqkdz
8ci7oF6NW7eQEqcSuHifn/Ndg6BbAKwWW7yjEBD8zfu2erS3wupyMrGCQnXZIDEF
x1AotHfCkSyuSxqIFUaF4nuCZppHZuIAMGF1EZ2lItPDlpXU/69QHa4ipSFkXAwk
BXfCNuCJdshKdGFOs7zEy9dRMDPA/dvpX+emvpOqQHJyfJMBOKK5xduvMfrKJnzq
N01t1nQCVXRi0SGpz+oRoa94D7SeUvsqIRBLOT3b6hd8lf+mPB/eGrQODaOteA80
6rBnof4kKfbKcv1lEEgqm1Lj9HMbOpAb2WfUvssdc61gvy/83UWf3sFKqGsg7UYt
InEwp0qCfGD+iUMLlzoZ2BFJn6Eui0NiLW+ifjWlIcmrRfMDRTHMvA+WlcMjUcMo
l7Bi4D1lWL4wF3sgp6lfiGKYTx6ktqKLwWvE1F98m+I7VDMNZ4vdogR2uURTtzhd
Y+aD+nf5kY5jELbxfY+/PLmeAH9M9FFgVEQ+qmTophvBvHs6d/6vOVTWMRBjyjhQ
R7fl91dUfKrys5Dz7IovL/3dIZqq/h2706cZUA4buI66b70t2IV9Lv3VwPcUMMbs
k3cgZM6Hm1mnN0//a2UISYHVWJz8ZWkSWJLO1dD5I0Vo21xywo9SWsC7Ac1wjk+9
N/lvEWBznhw/r/1EOdmcgPinVjUVh1ItAQ5WiPXsMyGHFYSbNpnM+XmVgZECFUc7
cx5ZzI5s0bZuQPA5RYK9U64GH2mhpFI4d9cslRN/SeEejHD1iJId6oZydPE9Rynk
kVoX+YBVNLM4xOUcD8GA1Jfv3Y1VArGyj9KKy9I4W4WQl73JYJ82iAP8VtLntZGO
HzsFQaFgSEpDRKQhQ9O90RGhZOsiHcrgGUuSmRFuLTfBQNpXFtlN1BbkX4eBoWpp
VPUIkAjICC5IzP2TE71GYx0Hn3fz4UbortrUMiJeQcCHlPk6HpFZ5/zzXQLnzA5U
2eWTY5yBWQkDuhSdprDy4LOOHHGfSRvyYrf1lfpJ/9Hrg3DBm75Fm/QK7Gra3blR
lgx523iVrSWzLvEpVtv428OhKrM0D+vsQQh8PE+zjJH0/sBBEKrYS8kYx3vY3kPs
8UnJvC0H5oSsI/tOZVMU0a36gVtjQIlNBLNQmefqwe7O1u12SedG+XKCap5hPtEI
WOIYO2E7mbql5fia8Sx7mWegWJO6DDqM9pGw3MnPH+wcy9zxvFBSuhjj2spXd1ld
PEVtPhAtM9vhHFwSGswkrMNSyNIp/zxlQE7GPl9HqnEAHwikY13IWiUvxCEjPtv5
ETiHt2k8mbgJcZClCGSODYPQJlyoJ2ZRo0TjzNiGd2U9eE2FBD3D8oqZEiGeh5uo
LBmhxPHqDkS0Ld4SIPlBRDL9Lt361Fv5j/NniV8alRPP2h33+VFzz0kjaNm+asi3
8q4ab3qxbDtCMpg5B4NtpApjPidreX6it5HEvy7UZWH68jOMyBoU0auhYlGirtew
UbL/jNLrm33KFJWmSckHVP3yX643BTt6hA1ZdysW4001RC2c6TH0EBhSw/zUEHyG
vFH4mM6D3R3N40MMV2bOGhta8v682ZaU9k4G67e2whzRnBm+8WekeV/2Gmz1c88S
h7Ny7DItZgS/RRK4eatekWRZgif77OPylH/6/qBr+uobpaGfX1xG9nNDGxyPzE28
m+F0fq5F09l7v7qeldTYulMok76P0CVNLD55IHDYyu38hhS2DZj9WptHtkdncyxb
d3Rhs5iE/yYd83kA/hzuoA3v/3XgspYu8ANlpumq0rS1+R939H7TBSzByf8eVXMk
bth2o9F4CwRfxyyKx/neBHkUDe3cBgOAz5JYwzeu28tyLtaS9ZxVEae+CcriniHd
SdkIbF9BL6JHIMktHdSlzjxcWQvvGa7v547nzaVzqF/DrOBvHCGW55RuEILDw3g9
DTH4rKIwlDcDw30YgB8DIMYQJnYD/qXvP26EGTHaVWlPtCfvJAkGIiJy+FIJXoMP
9Wmip6xpAltEi63HQJIGpd/SchFiMoqWeMLJVcOjJL88entD8FZM2PGSxWXT8NIe
/lILl3O4t0F0vDw0/jXAl7bZZrOlfdkMfZZD0sY9Mc+RQdZy3vJQOZa3A7+MJZtd
EMiDmQTDJLy3XPGHOuIg5amwk/MGz+78L6Tm9Pb++XBd/sraP7IiwE7GYjDdv1Dd
hy5fYKSbnkA8QjMMciD47EtZRc1Eahv7xrAKLZXPySOKH9tHS+IfRIdAhgwREPPt
fPqwhdr50g/yuqaj60G1DwT3X2BhG6Xjv+8aq6CaVFns3JoDDCW6eY3/vwO8/8A/
HIyqe1DiyaGLfqI0QS+z+TnyTnpgzqLfj4oCUsZuUKXdCTNk6Or3M7GDlipavgFv
NaDDwPUgQGPf8EHP7cYsTggQtD7GgJIBEDUdRl8gSW1/9y5gRAMsu/MHTNF38FBR
5ttB3MU8fuIvYQnLfkDyrUuF9ZIHS6Xgtb6Pt2HKZEpcgm2sl3UtWnR71lhrFtnL
iJbKmwS3IpfW2XnxRgn61k5Mf27edeVgkokIV3ncIf5VwFQlo+/mr8zhsJygpng+
Eo1cP18aB59XS+llIjvA1ktkGbxHVk1jO6a7vmMwKi0QHXeD0SJj088lNZJ4wXiV
9smbQ6Xf8vcpktPEFyuCvBWvU181i1U2jApt7qqQUqlgkyrTIrSW1tLdVPe7yaPN
F+GT5YYA5Zs1fn9NXU67nNMWo2IR7IWbIdpJ52ozzSQnxzv5HZ3Hs5cGRHMdv/Nh
iTlEE6S79bGbh1TsDIjIrEP068qpr4svX71Ac7no3PToYseQSXFO9K82YMaMbAbT
uVWWuGmsTHXyJKMTwhqkMbrnAdU03I4lUxwa2g3mTBbvA2LKoo3c7hT98zTSGUBI
rJfDj5oWeNATnXijOGA+Geby2eTOaHOpzoXz+BC3/mAzb+0cArdMf7WtpyTpaaQo
kgzc1eKJ8UbPJIcPp29fqpeQBFLzElQkjebX4/eW/vqjndkX5os1B0Kp5JXjhDn9
pYb7k7WhUCiFrDJZHrxvRE5cDpRbkSTBxKMFM4cHyjxIX5csO/7MoLAR7z1LH1yH
7JkkQwQF9K13y2PgJHjMCJQSNskPctATP7S8z/bqQSBX1CoADuLbRxck5AIKSxAP
TwY/IHZk+clONCYockiETrrHhiSvZrzLBK90EEQaskFZuhtaAcjtQcGZmA53zMT1
X0p+sylQf+ydfR+IygMMrzq2CHUAgKjr/jGbdWbmpoRO4UuZHxMYsQdwb5UFOcv6
x7fyCPvACOAyv+dw/ijJeYXcjjC5i5yFvG3sLIYDZvKpoM2lCW7kwpmF/WBh2GXA
ImwF0hlzUwVIQVyfqoW44ZFuiKJVB2u0kECbcHmf7In653IhQCmNodaB1BuCAAEZ
TbBt3+NMNHxKoUdNMNI16uptdQhdYOkQk/dF4aBajuAXCqsClPpsEPAKIoyQn3/9
rr9GBa+nHGinHGjD9tPAPcKpVzGQlarqPqPDnd2uDKOhle6zllzUfKSlhNnWAmd6
LX9rMjMXYkWmX079qDCtSMyxMjD3643QPEKS9EzcPLi7vz4I22LBahhmawyEdnMH
c51kOZqBHiVRSAxnhwmVsN/eKkxYxpR9HYBy1k62gChAXs6lQcfgUSmR2DyGqxxW
ySfdRrO0i1GMwy+lPW1RDlurWIAMkdwWAEmK2MT/HlLaJb46LYs4KcJ96IYmt/D/
RCxA2mqyHxxCmNgY7Gs/F3EUa0TsBy+gJXchJDLR9K0tMYYZQgA9nOiUIERnXe4q
SzutyUwCR41J7c5B9glIslUUd6e/Zb6cp+XOrgnx8rOCHbA1qpjds8OmyLWTvStT
Nwqn1OSo40YBEQmgltYbVK+pd/KYyZdPz5DK22NOqh8LpSiGXSoG14JpU7y21Nxl
OkgRnJbt2mohn/W7/f7Tv7CUdGBTpmUe3Ge8nLQFHZpxSXPqXxKTWv/wZc/Br5lK
5PNLKC38pP7T1M9svshwJnLyV8q/q9nT6Ru3QYFN7eIw+g0/Jt0t4IMw8ivnXzZV
ZvC6hBJN1ZV7OXF7GRGae8mOo7SnNb2LAuwtVCUgPQa/3o08kYM+6S1J8lUtgTj2
DqN1srqiz2iRCjGomx7tsPY+B3C/nHXKZtB6B6AEyXvWmuLKoxPRpY7C4Y9SfmJB
wxIWtlZ8sQgu4UblOMNbePrLtU3NtTH7vUKLDanM475EKqgkNY+/cLi8pg7hrO4n
DRe74GncgGBaJEMq6b5q7d+1cVT3/NQg/7k1AH6rivRs5zstTW3aa/NdAiVHy30f
0/X+Rc2vcUsj6VmsMbDtSow2HElSVFUl9Mo5IkruSldrjbJNU8k43g/FJokdS8B9
KYb91tWbL60M5qA0WccLm2/Rw+FRgSueRJqLLB7WrNTdClrTDi79Cr3WPHrilh4/
lbEcbLE1a8wbVvJpoorXR/lkqhG7ltRMeRrNid0n6bH04V0iUMwYeXHTifIYF9lJ
fsW7h3sgAKVpAlWv+glisl9mjDdEpV6WxrOyMdR1b9GgKpe4cdp9JR1ZzW7NnAtM
JVeDUM8rb+Hsj/hBwpvlPHaY9IzIoBHZ6Ngn1rr4FiwFCq/KNyH1wfgeBHgMtKij
CxM1umrtwKqwDhje3H2PKqHOTHkOVP5gmR03IO/5h0uAREvHpfR8vagycjogVbeS
lGX4F+Iz2Wrb8o/5adYe5Q1IAvp2S8okcnhghjjTdYHtCx9qPYlv0Nj9gdFb7C1d
Abq6TdCPtFzyivDrAK9BMrnbvvuJi/hjhVCnPVOJkIkwbh+FbMiNdmlvV2cMk8Nr
DZzPaCMaNvwTdS8b/6L46Cr8od1CbhaQ5BHhxVQAjR9Svks42my9nVBsLbk4I7Ph
egdwhOFqv3F86jE0IU+7eH8skECdZs+cPyj00lseUBXDNhi6CBewks8ej5t5Dz1K
jLA1YwL4AY608L1nAN5Mi3ZGFrw3jsTnsOqerrIK9Hxm/trg6x5OeEgfdw+7N0Gu
ib6YEF7R1J3shAl3YlDR5/2ctzfUn9IVS+7t3iUWs8wLRONK9bbi3sAks63MtO2k
uAJd/sY0G6z0eV82+JB+Hsl3m2KfMzwNECgLugNRDNa+LPII268AsoaiZ0XPyWCq
xEnYuKGbR09gecN2aTt8YHFys/YAj3/EHDqmSU22ZpLj2Zowz/sNsgOsnE3ueyJE
4YTj6o4gVngF3WoJIK6GNncrxhIveJRlDnFCyRDZKqQwHGvFDyUQa4F2LMnhRY3u
QanQ+UTR5m4qKoTjXrqsDsHePlZ57gVu142SKmgFILMlVmH0EJEPDRS7npk9dcoG
PygDD4vxz7UNctNfFlq90y0kFHFkSDsmgnJq8wePHcw4jbjGWu3lTLza3YMHprrB
rRILM38oUQU+0F7/fvuqXNPPcUV10B1EB9ooCd/L9AkMzoyVgGBZl+Vfx4fBKsM1
KuKM+vXtvuzNOQY6ONIjj+XnL57GCQWyHNWkjv3cn5yXIThTGn8o8QjQN16yZeJc
eozueXoumU460S27G5yauIL3/pmlV7VIOwT3AssuskY5hqg6Nklh6Vi9N/JHyDoG
Vftm8HDXLNZacXiV19xTeFPkA8dF7tD+xLiJja6TkanXGE81bBmJhu3Pjipwv2EQ
+Sx60aDmIpHsywPX6BlKxB/Cqxh0w3Oyl6hRN46LgNcFP/Cb2MVImKdBN6dCZZDU
csvikGvyAFRwnukL3adCIZhYltJf64mTwwGg294I/ipfE4IMMy+tgBaXRM0gr2/u
OuRFU251gFywPfG3eCGVUoiheG+NDphZuv9eHpfXJajVXKB5oWFxPKw9Q+ooRXsS
mK77dvm/ISvD2jYKwm5Kl9pPTs24rcbVkVGOUmdHUPwATxlon050RkWcu+CsC1jY
dI+sTyMNV6JTviqFXFbjsSrHCMIXSKqh4TU+dGKCuim47vQHtKW3ryWWWyijC9XA
WnChnLv4B9xy897sl4Wq5OgDAAWYkzCkF/VtWjzdXnM4QE1YQJ77Vs7KY3FyH2gP
0T9KkbkXhJZ1kzxooHVKN0s8e80a4u1TE5fPXvngEWGWqn+zKQHqjkl8or8RVQB4
SKczo5+Mc3eWCbV0QmYgXntRi4KPn9O2M+OCHZfRJJk+DwkKqQLMRctvEU+BMYM8
f1CmOig25rbYdhNek7BpC9jayTFDXOCdElyDXKkcN4vnKnyhA93mE08ovBh/6yRi
DZARJASd1W69ZgO3PzJ3cF7f3kQeBLjYgccGs1qjoLrdiZpxXkdvImi5RFMhl4Am
dtd4TgMVHRF7C0iF8FzbzgYKEMRSsxIuc1V9JkSUYYkl2pv/3UhzFaAvLjVXz3To
2KMI7IxUSYQynIEKX9OIiQFMMwGSLIzHty7TDPwGQ9LHEnpvqJO5RWM67QGa/bLw
C73zs+q2Y0mudj4/Ulz2deTh1U7jmsrsm8s2EI6FnpRr6szcR+hqSar8SpOrs+IM
elrrOr5xDsmNJ/i8jeqUgaVGaZuGSVAGAsEuuNYXhP2CDFLRrjFxSh05kqT5CYLW
5RjDH7QLGua/gZ2tVrWIbviJJhPsi4FCanzHSNMjSWrDclYEPdvFt+s0aCUr+eFV
8745GcLjnYlYTzTt/1S+4m5KPWv5xQ3DKt0daQvjZwfOU+vGJtmPH+4/a/O1vCvk
iDpStXKvjFREwwkbm5qJiejStuonZVhrPFaVbD8j2vPexhBx7VZ21anJGeYHJwjS
gshP8U2ljXZsQ2tizi4ucbvZqstp2XqV7y1HULpy8IQCXCiezmITvoGhUzbiOWQ3
gHYTjPN1mcAj70krTIo3PoS90sZuydqO+hVbK8WY2HMLJdPbsIYe0FJ5rCxto/sx
cNzJvD38kd0nGwa/9Y093PZL1xTw7u3edIbmLgpQOfna1lybxKX787DuHnEWYGci
QUSosGJoyjUuyPxLt/6/1j4nEse7OzWTAngTpjgStBpCotmLnW+qKoua+dwL+zRK
DK2OgVIrNV6zurDvk1eo5RfcEkHj1vyhXFihzM+He7Rw2Iha2ax/yFOkSgN1EpMK
J3lp68VKjABb9CGTFyLRIAS2rGiG+qF1zPx4MyFjs+Uyc/n0AzL24EZpPHqahydl
Dfmtauf8tM03sWq+RshAa5NH4VSccMx3ES4JmdtVcEyly1xL7hKgkmYGNDQs5qGZ
NIV2IJHV83Rcetqw0S/vPGB/jzX+75hMKqt4fAbdNX2C+mCQe6t8EbyFRM08tXbJ
N+bRT1YKOwJ0tKv3KXm21BGA7zNvhMgx5toAt3lkEA6pBE3kDdbvluPmY5zqSe4m
QN9bpaTqZamAKdYRSIA7OLOftenqR5onEUlB4weqnz1XOMJLSN1oAx+27R3G/vYJ
xkc6GEFGpIivAVHqilm8CIrKzKkNLYrDwE5GC2qrRyxv9P/xEWjZ2Csj4vbiGzO6
a7rk7QF33B0YlnaznuFoM2Kg4P71h0CwXXbpC6+ejFrimvwc8XbwAYGCNzXV18HS
9oitujvtrkPX4qOtmxRU0Sv8Zf9CKWxPlVJ4zxoADuUfmDOg7O4fbHtPSccl1L2t
4+i4YXP85tcLxvAGLQnD7TzOkrNInCXImB+pXr2wE/f98tRtNmSwEDRYZ1ZoGoee
GsdWbVSs4C8J7xoOnCAQ047q5j1JEFQXRYgBP4Mx1OH9S27qi5/qJYz57feVFfs2
W7LKJTgfB3wTnZDxPDnkeaUqzz5b55C9rDO3pHvh6gTYZ9Mew46gQFvxGua7ubeA
dfkvUVeL05m1/GLMW3HkIgNyJI14pJ6+zVjbCZFoonU4EynT7hwaYG6YRiEHHnmb
JMezvFj7sgL4aXRwMqYrbnPkFj4aDQR8RBdsU1wqn4qFqZIUkGErOWjHZmdXVRqg
bLjoxFznoWGYSmD5U53y186FsIpSlSM4UCbMCpbgFxF8UD+NelB3m3ImSri/tS8s
1b/ZzHlU0nCWpwNhfbbtbwBAi+ww2DRWOUf2265Gs1KhQw+fX2MH1nA00ETioyQp
WcoHdcW3BbACy1wLrSaNeI6QVTZUvLDeUkysMzO7ovGOrQd6L4d/Y1wuXDzJMik/
hPC2MoK7eynJY4gBCcH/QaMG29HTJi/ONI21V8lOPGz4VhihL+3Y8Xhhy6hGpcDn
XgPW61QTiUvxhMX9355mfiCs6wWBsAyLTzITKM5xn2sbTVnH7GL3jjeB5c4ThlWl
wYr7A9Ep10L2ZCaoL3eTN5FhR4hG4kxsEEJ5TXiPyD2jwibzLYG1teLrNAa82s6+
+DYjrLbB1y9uIOTFz0eQ43KwdOffsh9Ly3LiMEFE8/H1EU0O5O1cXNE2LadBVVHk
kaZc5o67qZC8XJu/+0pLXvH3OvqpTFMfnI3oLC3bKpuLSe3LiUsVC22Vii7PWySP
WWdjzaVZoByFX9m4UDpOZiltAJTpKT+4PSuWDk05LNLXSVao07pe+yrI/SBdeJtk
SwaMqvWPdASMFcf+Nbyu/x2BzXHVtkkxYTvhFWsW2Jr5hnXlFE/lOkLUzL6cwrG+
DRkl2EH7f2QWod4r/pMgFO2cdrwsGTbR1Qp1TsY/W1r4SegkHQLa7OyU/MohtBwd
pQ0pGlySY6OlmxdFhM0/peurn6hYGOQNxcdQYBDyERosrHHdxgL75R6kta14A3Ph
7LnoKrSDfx9+MVkwrH4p2dWPwO8dlzwWrzYLbLSG6xREv6elq/bpnEKIPErSS0nE
fZ3rh/DyL4o9gThYfp1rfjuzayEiTjsj17dftIj+ZLyQigEFUt3s11mRHrRdpZ1W
RMXmVPo90d+GKi8lop8//CvCisIQ0N/f/g22RBbEh8UyWsQOGb42CtxK/mcmc+/E
SVnok3n9XNmALfY5KOdyfBNJh/97WdIDpIMexwlw4nyEJXQBroDy3Wi3wMOFgjfL
+nHKNpvdF9kC6mWlMyyZgZnhwIHmnLSaAlqn+5p1ZjrdXznHLwbL2EZZ2alp5LB9
crzZQ06Pyma5YsI/WRPBvhPou7fZBYJHFLZMvybGt5MDqLj16fTIYHJU1twGcfJ4
tdjMpStrfH5bIm3M2YnkdYQXZ2M7yE+cxwQ3EcOCrT0nHoFIK06Q25fXmfeY9GVZ
/LQhGXXYu0F6eyG01QHiJbjsOrchj8cOR/YfGBUeBfCjQTolI1iEzHn0fzl0BedK
ZH5pvv9+6Z6FKBtWo1srHtA8lFUp4LxzM5+Gp+Oet03e7B+jY5GjXA40Rjz3apZx
yEHQjkDzajmgAoIyOWMCjCWozU88iliPrrCnNrLC369zZas2zh75umuG1yyLABuo
Pb944SBld9AirnGT8I7MJUDncOWry1OyytMQxCnIsdarFF6IExi+frCb5VE67+Z/
F7gTFxktaOdpGy9MTSRk/s2DsiMN9LR7gdAe1njJ9YCgY+F/4HpsP8C+kuXdMpJp
kieldWghHm3CztzbmMCdeaY5VP/zZroGD7IHb1Dw8I7wBn/qHqvWrm9HYdiX0HTR
/MXLwmjZiJAPRW6oQPc3Gw/kUqYOBoT6ZyH5RuemXU1qOERiNtXiUAKQc5aYoOUD
GcUVRVXqAyBaGsIZs3VCL2BlqPQ5bt12KJrm0eoOQ80qD/1+qUWmUB7fbk2BfjRJ
8HMGSUEKHq1ZoB8p6fZ6NUZ0QktDdyLS4T7xVxAdyUMwioRAJdpRWZ9hBPphOVBX
g5IrZb8qqSe9YKWmLRh2uxB5VEZZtJUG5sShMZXOm6jnTaAwDn51LWdplJzTncvI
hVuWhBmkEH7d1WZwXQtgDMqwIvftuzMnPRhnr9oGlDdIIgUIL232tmJZv7XNz9HN
KdNq68p45kzYzorzDcESnim6EskDSr7Nmk4kKnS44cS0xss45lhF91UW2uANVuH8
R/N//6dvbLRlgy3umxfw58al4OAprF7O7LfIIec02ichEkNbx87VZSq0dT9rwS5M
vR/VyatijqMYw7kSlV6+TRiBEdtcjaJa4jDp3bckwPSvvru+PB+A270LOvTqve4g
A7N3jfN//XmynW/5SD7bzT58pE/aQsh1Rx6KSvSwizUg3aXEfG48xA6OVpSNrM3Q
Odki7kaIEIZk7KoERqEQcvMdRutYrP5KItboB392QgA05VeiRqFmQ4Ru/dNzgzsV
u6V4DBjBlBLd9ZsV3ukhzfg8T9ZqHWyV3UclKnq2K/S25agvCmRcftxCofHu7kDN
kNN8xP3r48aeqNXuEzdg9YRywWrqNBKWjG/dJQ60nOyQrwi+cNKQ04ClfwxZMSca
R9chMedTtBA+nqKS01rhw3C7oy6FTrHLfQqEW0rIyVP3TLH10k8P1Qy4vK2lk9FL
E+U78jGzU+bz/dfkvdFbiq/bYHdXorolFXVyf61ElKy8zkJ1WWZTHh9kItWglaBG
ofM49m8VoSCiK0HUNocWUpNynjvo81hre9y3SmXfGzo98B2kamEKrFSUiFac2cMP
2uYo/XCU8qyHTzwYdFHq0caRIx3RMqFNFX1ckGHjnfPXAY7o7V0ZpD+LXb+vtYPC
QsBQ/1YzkCSpKoPxhSBsOpf0Q05bw99Xzl2giALKd54XgFiAxKcsKXQVJjt3xhN+
rHGKCULw376txMKUGyxFdxkAUjktXavrp/SKljtQtUs9q8dkIttQUTTbZrpm4Y5U
5hdJj2NktzYh4fW29cRRVcd48oe9K1MEEPiW0MdxtArb8++ZUYF+TwMX6j+1hf8O
6bnfpI6Bp4dClegwBJHNX72w9TOAm6/vXYcktMSPBISeSixEQhXISX2b106x6lUy
pqoXdNej16F2G5y3WSNngM8CQjayT7efwjSyYwBeKUrJjXDHuztD0gUWDgz2gKQL
D+j2G8WUY8teRSEcy3IQ1Rffj8EWl+/JhJYTeiU7d/SnA7D++oEUkG1od9jQVKg3
al1ChVpxpNelZ+LJgsLtKyufO7hrlsI6Fx8RLhXQjAfVhVdVAsiEwZLkj5jk0JLt
D1k+z6nfhCbLZ8ktjXUPCYosjCA2EoF0L3VaWsJDh0jjLDE+vonAckRUaeNd6uTr
MIbb9wOHdNChaf2BBcZExNgStxz8XAVsDHtpCCvwuc24R9bGMkl0cT2R4gQSxCi8
ux1simKySH393ZiOJyNgkOFyXVlKfnxgmexqorgwOdIQpKa5oXzrkptySXYVlxxh
TSrY+aNfmN8j438LaoKydtvziciA8Jsqvn8/X9VfxMz8sY7Rz2vW9K575A7XyP6z
qh8ZZ97h3xTXFwvFvNw8aYOt0dyDKUxyi+5RRd9S4FJeNZc8YRP39ZgRiLR4vBx5
U5PDLKW0sUUd7az3UcBLB7nvXiyauEl+fXK06mQpte634rP9HbPQ7smp6luyZqrh
a/PpbvF2ItxvZ9adyUgWxS+t51QTDnvAdk2CsZt+j0nLt2HNm1PfkQv15exzjefF
2BV4544u2K7reuRQ3ExGJnxFepVkY+MYkpIhqJqsM9hP/ra7ILlLbXf8nzNx0Qy8
r+DWW0bz6+Yr6RejR23f0q4mTtwKBkID/Yoi+UR0Mogfc2bqnFUZFjm3LxDcuWK6
ZXXIoOClFzHt7pjqoOig2iTa9TTzd/Hbs0eJV9BAJ0aJ6GrOBeK8uXcAX7OByENQ
M15LB2f+5H3fHUIKHUPva1SvGtChijTgVLSCyBx2fzwV3w77a6ZvHNCnScDf4LXq
MMguNNeFS4vYFVnOr/ZT7eCMEN26yj+xjwBkWqhHF+vmPbVcZ7HOViwt6PZXb5Yn
HAxzY9fYaMYiRV4hxf70vIwmq5GMa56WzUHFvzMtdCTU5fK+O5Zs4jjjcVdG+6Sp
51rdGk0/K4J50aVxRyHTWTDtTXe8CrNS76YmV4rdRgitOIytP5boO/7/sEWc5bdF
3BNTO09f4R2TIgHPuEvLSUPFkz/qw0OC4HkvLB1G48V9auBqZG1dFFvLI/sWtoFK
NJVscId8ACpO1mmM5KzSGy/MvZK4Hk+yG9T+DNjP2YnBV8F9uqUBs2hZ4qYw2Ye/
e4pS1Imj9CkhtN4nSppgNTNyCObvSFvaSSnfCnXJREn9iBsZhP9CYAVu+61R+174
stD30l+/oqvF+oQ7AMq9yIqUHqkagFapp/oOejaPQ5GhLJC1o53nIUJM3sMs8vMv
3F45/o3IVHABkLURTiMa32+wBdQrTdwCrHMISh2N8HLwiyoGtQcZdjNj7YYt1EOz
8n0+b42Ne9cyPtR7+KfDdgxKz4dY3v+EeK5/rcGAaiPfNIo9rH+qqmZnXn7tVFNa
VLzEa19lB/GzAIuQIlYEXJZPDAq1M6IU6o1J7c481rb8YqjAPsrmNhH4DYQs9VaJ
E5HbdmdqzfgjlOfqYxfn+sos33nvwmuttLJlc6GqeVmMhWlf5ByOQpfqH4CyUY/1
kXeTBA0N6jfX8Pn9e4Z40pAvj6MytEC84+guhybRViDZH/dT/8sfOx1DeEuY5+Xt
ZFJsA4znpLM4WkzWiKwBTtIlBwnLeKXs7gj1mDwU35cL//AA34aAZjnOEOP3IZJq
T2ze1kAplb619j8IoP8ontgS6HzIm/bfXE9J+Sd/m6HQJqaXeXDQVOInKdJ/pHm3
Mfr/AISDBrL8PcYxohWlhbUXFT0H/JF1U9rruVhKL7UfuILmbIa0ounEnjI+AyGk
hIQSr/6OQqmwE5eAIouDn0iMjV1lzY9fI8m0YsFbZBiEqkfB0+0bFqmMQ8cLoh55
2FXfmHCC3gVLc2I9DHb7jWGxX9kqVgpgj3Tk+9C3bJScRFdwXgpdGt4O0CBrgWgm
8BpTAlcMBT4fK5zUufHJQ9dIaZ10SS3rhGQhgUV4dI2N3hr3Kv80wA91aoMaHhwj
vkHzaH1UJzwD84bAX/5fuL9XgIa39NpmJ6JNcaO0SUwwrqXHFp4t0BhNHccjZqtc
N0gQ+4X7J7lFcXX+ZAmZ6+VTdvqPW4+whPNLjUmXhNMTo3q7+Z/Lt9bxNdaHYdpn
oph99/RJLgai9IXfsC/p09l5vFrkVQ6v7d5/pffj6eeVabEabIlgP84V0dKl8Z6D
tOfCLPc5NcRCeePULpmIMSMgfGrgeUQOZX0nU17CCnNVoIElp332d7ahy41zGobu
s67lO9AinkqZmngIjfpnt5q8wEw4vVxS0K2u8WH9vQao3Y/xh+HKfCTHnSWLtETB
AUlYEurEVivliVTLfGF5vb8wD87mSwkxRkeiVKQAXI9BkQ+B5ADAKKoVSh+fYn0K
1wSkCMkqFguCdJY4AwURp2hXodoRK7zZQ+e9jFmxCKqbvUAfR1UR18lYUp0rWFKe
FzO5ceWT+TUmLoS7hhaAvnsHVB0e5MSNuS3pnZtyZvieeiTPSk9BuQoha0ei/Iq0
qRmrlQyMvsa9C80z968KH57QsrZCwrzrFJJ4Qi19qhVHoXyD7D8/xv0Nk1HdLCtF
gogEOG6PQEUNq2vDLlna2t2iSBSZTKyiIngyqefRmgxEeQsZ8dxwR6cLeTQpfr5D
JKhMCQ694kGXH7VHnks/1D/3+34ypGtMZEH0PbYkzaz3GhKzWGv/gns+If7/pjrm
I/xgRk4cssXB7TUNPW9sYB2N9Gi7wzogzdzRK1+jmpz7oe6ie6d/RJSRZrv1yX8P
pF9d157Ef9eHik5h9Z6zIVsjXhfgXJ/JE3zWlpJuoQ21oq3NJKX5e8ROhIyfaiHs
bgS58gQVasbWh5u4QPYP3ONcpDN5V4Mc3IurCm/9IKLXcJ1uvabdYjB8lu6+EFa2
O3ICJKbcNU6nKl/bSK8FNnmy/7I94eFGzUFsq4wKZWkf1rhiNYmjvYbFE+Y89b0g
ZtXnG1cWbi9bnFT5CCD4CYFDyl6DBCfpfEK0fnxO3Uyiria9RFeyHnRwrGTpE8L+
gGQHwaWB6UMu3msJHllFe6oMnXuwZ9lhOzrjXkyIPBkVxkb0umerCIQVOJ9Rk5Ki
dmBgraOeIdAMTyFsP4JCOS2DuhCtJ4TQl1snU6kPLt3HOzDzJLsG6uIbMYlNXmNC
OyZazKt2qnEBWObert94akiHZDdtqp4d6aFsWh7sozuIaGOfD4GpSiNpMc/x/7lJ
O2vNnfTtTJ2pv++eceASf/YX31FZ52+PbVhByBbWzqkOBZ339exau8hjQvyz/XYe
z9SY5lye9/zA8DurCxgNuj0V6ivpQNXBCBjVa4G71NO+BUqsJADFp5zVIUEuoyAE
yZmpsCS5PnA8yiGVxDL4k8nPbNIu0dN015Q9A5g12CgK93I9VfTrBe6fBfEHVKsn
m7RTVP0LDWp9pJQcryW+D1XVbTe3PYC53uVJwlZ2rAPqd2vxc7UZYE6tS6a9V6NG
eGbwyXZcVa75oQ+eBf+Rv9faXDheGZEQlviTcVDWyVWiT4VeCH0ovJB8aQRk/MmE
/nt5zWKw17igiH+xUva29OeIPeECmOkF2ptQwa6Plb3Ma3xqID438QABuv7BJ7fO
28Zwp9O9orAXDwiPTDauFgTjS7yKkBBvJduWhQKg8ECu+rRIZo8Vd40hkRqC1vNJ
Ve3Ybm3DagFWOL2Ml6d3euY4zbaUxzZBrgXhtiIo7k4lfgVZBJxp3kybXYSan0R4
fuTXtkjqJ51KLkUdrZT7RLnEmeheZVykwzRfbik+jA+yNHYmJmau5vmaukdcbDc+
6sKgMGJKXhnynXdKhj4ZPgX6epJI/v7IHKZ/h5TpTNjs5JjxQr/6gMsN6q0egA/W
CoOYK7Bljv9yVznJHj7Cu6P4hiYKW4ASAf3twgJ90mCsWgiT86cWofbKODS0a4ov
N3tN55BDf266TvcyJG5zjYY+32GClm8Ln1aDO4KsW5D6A5pF4cYI6oM1Cn/Z0NPZ
zrcs2CAoagjoKHdU2Vb+u3ZQ0/Y3XDXftUS6gIBdl859l1YDjv9XkfAeuQtOj6aB
l7AU7W0yUExyOtc23Rfe+YKpPpaCEGUwYfUQdoESknuaVKWK+JzQQYzf4if2B6Cf
ofwQoMJB4RLgcaaMgmAfJa6GKWmscASHzd1MhQEiwO+aac+tFV6mXQRY03cu5ciG
Vp5rjRn6TLFbNQtxB1PLTT7Wf/JFaNBGWqwNCyQIGajuCLCYkmxJ3oxp6EyFoODk
Mzl6YV5Tic7gpyyPGhWN6yiVokjNLySbm8C5nzdqmfma5IoRQEioDn0ZZdSZbyDR
ZsXhTWYy4+9lbSzsCYqAqobf2UONGKF50jt4AWt+lQ7QaFQuJ7K+962P6S+fjWA+
AczWVYrUvtKL7lyCY0suzZpJnPPDfH/JjhmWRlSgrO050xS2D3ZmVfzsTL/yxY65
X3pKgEfmiBvgJtlu/hmzciJlgKI7PahaRAE4FCJKZNNcL3lqiu+NxBmfzv892qG/
IXFBsG97yb3d9T8oHzHkqFeKunNrv46/0MBu9UZlt7REslENzqzG0LO0olnrbmnZ
z/gqYn8zo5uAbGrTomJNB0rgzPO7s3Tt9qB02ugHFTVMDd5tf/icpJohhTj7wTjZ
vFeN8WcnCVydcgVnr/MaOO/UOmUiXdp66Iq7NI5NDvmm2e61JVAzOW3HdzBmIys/
EJTD1ZK5Gc2iE02L3zwxIa5OPN7zIQkKE6qTWB4SUgYLdIfedk+H8OJu6NTskjwV
QUCmA2vjGTIIuLwlqKHl6QgN/Ma3C/YIVu+b1+tCcfmQv4z7QnZUTTrbpjH69Mzm
yxweaYvoIbu3/sWep9vPkWy59HsDcVNgaUr36hgRipLCzdjfgpz0fkEhl1Rd8wfQ
O5HuUN6KGjZx97bt5tjQzXXaLblNFeqMCzlC4mylFBkjOJTDjQXoxc7nFnohBNTL
S3TEbqbT3SBr1g8NSezL3sbDENlWUXEdRaPi6RfzC6LTII/kOBjwwWhUSvuSgyT6
pmDKVGCMZUde6hEcFTg6GvpyUwBzF9lPt19JUJAMQeOUzlA7KhWQPUme9TNx3fa6
2m3xPbE+zACEYC6Y7HwLxMUCqwRNo7zNnB6G/Sn04ZAdjNF7ZYkG5zM+uqyZr0Tx
JNlkVp+GnwiNEm20I5qHRj1ce9wGNsWXUTmFyeBxtQlnYhccyn5BCEjsKRdQkDFk
KayrRcYzWvuCkZC8jkDbD5fW8Ynk+ZYY0oKhCxtEn5cyrYSbTUPmB46Yf2qk2eVL
tTwkoBzu1FFhgJpf5IOFThEUdwXgs3NM3BoU+3RgszGqfBHK42pfdBciTRskH5b/
uxFHqEyPoy+iZIHy2OdtWigjCpgC8QtZ0FYJE63c3FDh3Y/ynGgpE4/C+sKELzbZ
zuKOM99rrXjM3WDknK3xKO4QbuJchqDMOBIA4ZYjjT1wfypIpXn4VrcJ8RGPM9oN
rsPYpbcaO4pEbJtNZZqFVPgCmeYw66UWmjttrJE2BljFYV257EiWSJYo2ns4yp0S
O2c8jRkTpneuyfSmnipG68+7ndAYkjC7dr6z52wuNSpJ9Q2SDUnnr3sSIDsV1S1E
Zaj7I82TPtg7BIhTuNwzdC6LV7mqB8AXU+0VvTkG8/P2QjXpvXmtf0cM2ATmsQSz
gmT3gIAkDTHwttuXaO6dOAHaUQUfh99yMTqtsr/8Ljb9CARXOqFMgVHatGAjHAsx
EFynDTb0QyWTlrzBQ3wvC8MasS6XRk+paKmAVLFjOvbD8OPyNhB/ZNvgWLYeWv1F
JJNw12glec9WTbZ2Tdb6LCRnprSBdppZonDPbS96Wq/ZpZUF4S1zI2OM+1wGEnAW
WvgDh9StGgblYwIn3oDrqJYAGixL5r3hY6pXDoUAy+xy/gGdED2+lKPtVAldMyKb
s03Hw2jrKlRsY0hzNeFoS0L8lsnqloHRqyIygp8YpHfb589cpezRqGkxgkOG4njY
upZangBcMuKAN2pQC+0T3QvOtamyHWZiH0vUow50OPzWZcozEwKDiCBj2KlQa/1d
x9Lbi69VVWBW3svMVuWZf5zchT5jD2XDwzs2lkQChbPUr6ZkaQyKNtcsrsfq0GCG
Iq9t7ApjWD+bxsUVqnM4pEvCdhxROeB6v/3l+U/mGO1cY2YOmN9bPuAJ28jVH58V
gC3sFv98rwefPzDDd5Xd3HgtV+Pmqd4AUrzDfWjEeoly7S7lhKBDa3z//JxkM3pG
W7h9vAiBBbg6i7bkeBo/F9WYMdMuI8vEC/1bHBJsAx+J1vjPMTIUOEHjAK4iPNm4
OYwBVbFqh/xRDiilamz6vrSTFXcDDoY09FXWpf0lXXhVJKjzh1mfsCP0lWtbg/ua
KPOj+n5H1rNm9tJULTkvuhno32KlfGPFcWNnzEY0B+t6CpzPacIPEtkqmfEyVLAL
BtrCBHq4CyRES3Jpp/nbEEcxvCU4mUQtD64a5JCyES1NxE2os1h/IyJFptMQRqxa
pEoKWMFnP/bBGDdEyHK/10itl32ftit11frLXceHtk+FoNRIRqIia91CTR6+9scX
oj/0e6jmePsC1G7kbfG9My5VHcafDxEQ9C6QdA1CSMtyWKJTqmkM8Xm+A3WarrYv
xDFCK5yfHwAyQAOUenqEBTan7BLls90iRVEVDaj3e20OY8avlLYSOYmRCe2U/Emw
x5dCpczAayjqphNidTrOEVM5xAtvoix0/WaMtFomT9ejZe/QXeBPxcGKZp/eCtV9
S9Rw09F6CX0lyhHAMo1aoyKD87gnTJDCiaYxO1d9uhZkTEskLEYCoqhrVA9P6F1z
RD4YjKy8pnAvoYMigL8IFmtVX8VcRrynFc+G/AKtEEccbV5A3Hqx+QC4qrckJrn5
ZWbdsPBj6Y2ku3aW1HP/qQGsL6xehDoIpHt/2ZiGbx5/O4mXH+oPqMrgKjJR14UE
ru4H5URfBdgxE+LjPE5PC0ND/FTdbpF2B3KyvR+WLVUenBcKSYfShH8Y5+nuzQ4/
Ni5nMfo8U427bHo0mFlYstKRbMWQ0exQMebALTzG+Cxdd3FuSJABz9l0d1GN8HVz
fsHcy9DsG3w+AtuS2T/+SAh0CiI47n6je7tOULwp/N7RTCksK7VBfnD8V28wc7ne
OW0tmUcuwTOADNwq19vH8xYPUyQ9GtfibVtTqnA3Bp/uijjYln5sbDyJ3lmehzAf
OgQLRqE8JwmfW6dsXmcsoDYKm5Zbgf8dUvXcce8PUcpdNbENydVatkZhIbxBm0Yk
bBPhJWB2o9vpXqx4y8sKJeCsnSFGp85tEOONsPaTQjVWvSM67k3qsAydVg+5rUJ4
Q0T5ql8qWfJ5J6tWI6J+ZedNeLOy9vH+7FNcIqiIUkc/VIEQHSpDyZpadZiVvgQi
9aafmX+138zTxwQtKIxAgeevU6YZOOKoJHIqm0nAEgS/YdhLWB1bG51MZKeHj1vF
0+tfkZL8vyYN2KKYr/HFmgEigAqnjy4P5z9szC9NoVdRJyyK9lN8EuQ+xhrQ1jIR
6w9WWnWcLSO0jDdkdN3HBPQtArLCGj+tQEKO3Xo/dXojyc0+QRNYfieXHuIIwblK
ldzXhyt8QBcPhh28KQ3GakY4biRHmQD5T4e3na+BM1VgyybOgTT2UYuQPcWvHhrO
PfOEwsvAarvt8A8u2JEp14UV1jy2sf95uL/yazu0ieNtkePQ1PZoKFVffowhdCMQ
mu3oSEBsXZg0+Ber1JYXVXYqPPTTJpLExZSR5TxwLyfEmCjg7io/UkxzwiXywC30
KY/MnJFPEEJp/7Ui+OuyFXEYHLPWxnh2YtgWO+MlXoSgOfMrLIll3Dygml0jmfqv
q8R+yILUoO857ols+2Zp6xZ7tLD2JSyHgrYDwGi57PioDW2SZ06JFUntwtWg8rv1
arRGT6Gil5OCE5+xarfS8rqFwgKnqLUy2FFNEKiOseAbCj8rly1GRo1T35Z2HBA2
FtYXkk/Crks0lTzMKycBxsZ2ii0Wvug6xmQBXh1RKe9vtlBLJqOHQ1wG7AQAP+OX
0lK0kK906a2x6RbEldWTuokwfbPo3RHJv6K6wdwMy+fX0FsA1UQK87JiwSldxhJH
5akQYfRYLYcBUWghnDuiIMNDUbD0/f7w0HtDJjEJdbF/u+dsGaQe6W36VENlhhTS
YmI4Q/tRlQG2CscycgX6TgS7Ok/3RXmLEJV7Lx/GBpYCD2n+SE/v0Y9T54RNvkpb
Jnarpg0pWDgTtYw+CEny7vPOWzAptUEO/EqfxX3Y9ep1iFIPgljOBfl6VmqwiIn/
ECC46AV4pdfiGhi/HjxPB+iR44nYxBK+SL4CNdEmCtfxCAKHWLn1+1OIQEXt9PxZ
cVAba150QZCxEjk3cjDgvOKDprHrPUPAITUHD0/wPS0V7g+KQnfoEsgTuDhpoALi
W1JQpernRc7e0K47UAZEL7fcWCu6qVMYKmtI7e/mg5S2hnBUAX/OYHGtusm95ewK
by7PBgREG4VJ4VEIw+hmvKNVlw9YwopkYhUfUomd581cB1eTW6f7N/xopkIOZUjN
UPmGhZrzWXbSLKpUPgPU/tGT7nYIbsdlFY/tKnF/9/xseJzdECzyYd2mQHew1nLj
OENQrd5h5gtvWnEudOoJAARiNH+nVRD3Kybh8xTJzFINZus5C2xrviuJQ6rmNKcJ
H3MlpBHKGF8g62OVkNdC/+SWBXN8qPT0B28eGZi7yjuG05fY6IAz4TN01/xrhR/i
yRo05GXIwIlS6k5eY2feDECdFSLZF7qzwor73olm423dYqDdl9S3VWBzwd1sLS+h
TZq+GFbAOywApUsOZ+tne0s0ZY8EObjvs6EnNQgMrQy1wjKNnICLQDjgjkQyMDmV
yNcwc3bshuPKYbcebwUvf/Sj5jBHlM4haQksPH7e9Pe3NubRYc5t+PLctxVSC7Ri
eXvMzGhwlkyKNtATAGcUtEiJKAedze+nRRkP0gZNg1y0v5ILsMXeY1Ms85Zy8vGm
36rbBxCoa/qG54ARAkzbWJ2Dp82gjsiXbGBfm10wYyFejQLPx1F7edQQzQjgCwlU
cg5HEqIfzp6PU8soXxBbp9q0fVOsJwUKR7WkYGn/crSI078rCWocuMV9oDf06IqQ
ca/Ci4vMcmQYBKd8EDEm0ACNSmo8DGDfCKmcCnllQF8qu56HTdk8MQ7EgwUO8CNs
xtxADv1Pz6IafihK2a00qCbQnbSOUhzC9wB/AKF/0fCxe1jtSm0JNAAP46yFfJ6l
oVzYKhYR8oBR75D9oo9WQtkff6vRWjjMa+lpT+dx/DfTwZ7M+w/ms0XdeJWDXzZj
blcWSNRuLHzXex4VHJ8NVGKTXhyIpBE4JMxnmNuRfbwSzxGTlOA4O55gg1eb0uq+
9UdtXcXkfxwV1TOy+/lScIYAaflEyM/4jsC4vMko8baKYjFczCyBJzUV8UbcX32C
htNgWDBKKN1zzu6nUDxBCAxDMxjqCTwUykKsF8kKkz9YGDdkH3vEB4lWztdDsWZL
NNxr88i2MpSetAlMXjRnKFHRCnZWD+i0FBkAbSogePd74MNtnrlD8Fn0Q71InYF5
N609W6K2/YDogggGKznXklyYNOaaujj1f7EbPA1ZnWI5aL9BGnOzPhXU2hPOiZPf
aQbTHK1A1WV3XWmstdoJJ6v3FuCrlk0fpwuzDWEVe4q4q5uxxF7Xno/OudNm7Dn6
tQH0zMLLEGNEkekuyGqWlEydAnH9RRbCwXSeNylNwhjwcdSnbvRrPIK1pWfBBRpW
7ir5QbRIcvE0Ut23qEC96CmePESHgk5NOZ9SRbtK+e8MD1He71xlrxICdJClQ9bn
wzR/Xsp+AB/mZhcx1nThnpjlVdO9OQM8SRpyip33EhIczda5UmPC7csLUsd8OJ3A
k/t3KzlFP6hay0MatrfIYJ+qfzCFuBZEkijoAl0SVvbgvX2cBXZAMh+a/fh4EFvD
WebrozaaOWEIDssbGN5mPeP3llme6BG5OBLaiDnI1ydZWQcjF/+n34AdaPKXRVaF
JDcY8iBgrFbWWJEgsAbzoP9voDNUu4NO4wn/fm69xu+rRDV93IIiWJHu8TF4uoIm
/lgrFpD4EBQ7agNQKoQjp7ZROkGpI23X6d9JMsI40pHzuqu+EYsL09Hn8CZ4Ve8O
GJLHejf7sO0dnuJ0FkAQxFYmBYE/+LWRLndYZ1DVZ6wvmRIbQOfvZpqWjyiCXsIf
5/c9kfdw8Esr5C/I5k39UevCL5vK7Fjir5vxMsge/llHTC1tVqutPWZtB8/bo1dV
eDFLjjmLFM1dRBTCKPyOht3aAZeCkZo6DO/+w95SOZ8DUW1dPtm1ssHZOMecZ3En
BVtNH8RCeEKgPofHWo3gS4P0bP4l6I8mmCDFv1QxIZk9Tjdb0Oo3SD19rK1S6pqg
Xr/3XR+wDZe2jTg2zFvd1DDYnAwDo8RkwzhUXU/1Omsy0tHHrzoVkfLf2A2QPDCh
IUHEr65lJDquEjuZNsXW+R/hCHpaqU9WEIwwh6Lg6jCipnY23l19xt3asIlm/h6k
9DuIvid6SQ1/H3ET5HOnLjDUKwMlF/ZE5a9JDbmbXP0LsBZg08m2ckDKm/xyR2CW
9sa59y2O8HA7Ch2BIcgFKxanKwCIQSY9bKY9erbgzjzaFG717E64KcSN9FB1MAh2
F5FP/MSfsn3WsxgDwfoFAUxsZBQy+WgSC/EsASFC1rl+MsaXpaRn/Rw+Fs2mw2aR
H4Z3p6IcFAPOdfabBps4W1/rW51i9mk3438uONEueEky6W99WUffMy+zuQknXpcd
dzEASlDa26F6J6HNxNMacFJ4BoCxwt3TiuI4gxi4ZDv64L6J69RPLeT5Y2Fq9pxW
Bc2OhajzvFkuGr+vjWxF7L/v0yQ2qnva7bF/RxEaFEKvZ8j3gexGgWCoKyJ9/QnV
22CXxYp087CSrGf4YUzNqsF+nm1z/s79cMHpfPPMWisSIFVkfGenJv74Gi4MhtfI
YOyoTXV0jHyU52m0/ANqwWhD1/G20MtXm0DcKMVs3zfr9BM1Fp7PaElFif0rxSrh
D7Um5VN5JRTyRgj3VSMg7jSIFongZRk9o8WuzkhTWygm5wvIgNLvQAaIMgK07kDh
HIbcTiGUGHO2fxNvL0bm6rquUo+x4+o6w4K6kTTJtxoFswm5ZWOGLCJhtSOmiTUi
fen1ztJhVGdhL6HiMq7q1p2fZNh8vWU0OfKu16jjHBjKHoKkYCZI8flWdB1xFjZ1
jzDML5l5Le2wTgXJ0Umi/6dJOrL2r1QUIYQCUkdYEdKG8S2rIv8+66J/RugaKlq8
zJDbb+Zgyg9q8GBsuVQz+GPlKqYPDOofAuafJxzGhT9jYFMB9p8FfzQk7wy1twOF
ENTXZDjHu5AtjT0uqZjx57UiDRfCZc/2qdosf49eGfM0r+6YAL7RVPHLf7gAJ84M
bspg4mcLCV8v/fALWhtLoFOtiRBxKHS91bWaUfGs9OX3Hzh5IwZaKE5An1nA5r1S
jMhhJbN+AOh88ROmyPgmJKGkl3cm4t/Lz79vuXJ2/PxtP5NcoThoHtM/HDofZmJV
e93rKQ7kmfaCRzrkAa85kAB8lfUtaFfDQ5APuat6IgZbtJfMubEKMNhVi7Lp2T3z
IW84NKyDnvkY7kdEC300xloSNSSnP97LOlCLJ2wL7Ua7So37keC3RNNy7fdPJdAV
nZ8NX4TXooLbRxHGrrhWyTgk1X3ni3Ulq9AjdoVNjJ5XnhXVmVJRrP3SlmGT1HaS
Sw7oAMpT9DuSa3M2yrXuyuJOOigKTaFeF1Wk07k/FAk46qBunXSRJmx+C1Oal8Su
+SwKzJUm2O0TNaLqoEAuQwuRo1/yTf247Zv8u3ifn3qvsqaQKKXYESSeNv386NLv
x+wP0qXn7CNzbsoXtbymKc0IgQPrC+0upXFnIF5eWoXRmGQYxspdmyVnNtO8MlkJ
S7Ar1ZnKYrYVOz+0Ianini2u0bZpOQHBtCbefTtVPoyLd2jFLbLOosi+eh7C16he
5auE5vAZfJVDap64TFDJyodo4ti/PR6G63RuO89sYi8mOBPC+uxzsPGKWBoC42Lb
socJAFiJUXc8xNJYJ/NA0GH3xtQ/mcx3im0VvG1vhqYjRudNXY3ymJ3iepBI/97j
nWCAE/1+yUVO3jXof4FBHfSm722mmmCm35w2hjCJ42gLkO0OK01pyWwjRpF+10Bg
xr1zVDeEiL/4aUohnKKNOEpJyxdJp9xuzxP7OmDfLZozIDoeoOcsmHZ8kWFa+lbY
2lgXR+KC9BgbNbIfd842irJc6m9NXKmeNYzgUhAsBm/YJVO0YiI5lvDczgWgldnB
I43XkCjg09G5Pd014rwTgC5D8ckmGqb7FXx4MQnQcHg8uF4A3fGwDVN0PDB6YIBa
GwHwdNhkPNTD4kSW9Ioq9szTLJm8/YHXagPPkJ8BUgD/NWfbq/t/Vr9jSH3GOM4z
0G5/WOsw++jEHiLLd5NsEWK2JVh3EorsJUJEfx4WXszIseIrNKZ8N12lUuDEtbMS
IwJ3UY5tG2oHvo4Ctw986NcDCYucKFJ0JRpzAGe09kfWRNmGRt5QAHKaN2mKfea6
WcqBUIZ0DXNijzJ6pGHQRuAmzQeNReb+XjpaVsRUGaR0Fsjw5ysa3upniZZoh3+M
zhGIi8lqkBELl/bq/WGbLTn1OZweYNtoZ6T36TijPunDrPlvoMY206fvdCo22k0L
madGv3Jnu/9cDe57eOUOe4bN6D9jnxMKV3XptCH6kME+d+NNUkwYAA7E8gLRAt1N
OegHqYoa1uHb8OPrLPJ6SOo0ybpNITNsqgGbADsENdECuicxaA7vLJUnPQ5fiJ+O
A7PPENLRgo36nkGU1c3hjS/2LfGtQF9yLq5AwJBFIiY6z7IpmGpi4E5p2e838pQ5
d5GAvGLfGnUPd2PG0+vVFuURp0Yn5ugSLXWYuOIAl5Vcb/EJipGdu4Cv409E5Gaj
qr0WllGmprniY1foAAlDnnJ87dadtb8mQ3eCZycUWdLTHLyi0bEeZM2R1UGLGTs0
uCxjxK8aW1oXGsKcSq/WPWsPIBcpO2+MAGXSasrWrTsOxQeepBFrSDLwvGOUKtDT
18ioGWcZrs2hbzO3/CfZI84+hkSvughCANkWWPtiOxkH2b3lvFo49mLnC213SFw6
lsl1yGWgJzPOoPJJggOfVl4KakPJBNuEJw9W4HWeMf5puQLKytgwX9rIaG/EKSIJ
gxJWrl4aZK3adWUdR3bv85WdYq2p97WvUManwTP+B+aDY3EhRAcuLIA9HNtBoVUg
WTFbE2sPfaUBShPBFGFG+UenyUm2G3SysXu6QUH/x8Wu9wkPCUzIl3ddSAOwZBZG
OyGEKtMHBvrDr9pA+Hf6tYMLw1ehiMPdYto3E2xeNvl/b8FCILkgRRpiNSFRFDfc
iZLa0vG0q9DhR2krFvkgH/Py1/St8YR1ncwLYTGrlogHBaHcgAsECNUNYyStIJZa
byobEoMeMfFPliHiFxxnKtgbR5DDvErnygKGZP9F7L210Csq/N+DlZyJYjtFAcPD
tK4ICkSWPN4juJrIuRvvy5DAS+QYFGX51T7CYjvFvwvnJGwCJpMxIybX4UUIWGt/
/hKdS4BF1mdU9Sd6BBwd1PsziJ1ZlHEy2gY7XvIhJnXFDwKKmGd4yDMp7EjE52Do
SYW97p0WiRnTa4Eh9/v3t3Wm0qGxUkdey5YjE2gnQD8TPRjSQd+rI4o5TFjGBhtq
/OjVZ89RfmwEg5khRzzJeXa3T0bbWkgjMwHDwoynuFyQGhkYY1XZk5UfJRlxJYTs
BlvMo7fFe6Swbtg5zpY7MGwGcqNKOKA8jNtM8nBA3rjqkdpomRmLGm0HD6LiReQF
fk8/iuSjCFmf6LKxinDxINktQ0IQ05D+AihDSOhk+0gmk6VH9JsRg1CPhSlpBvP9
kbztYN4GvFYjAgs8+MiQVV1gxBynbuvtwGUauKIuKt8s6ySxfDpwDL2OcOIIm4T5
AtyYRuTIkOJ2MDfNIgDjmvoAa7muvdN0W8JyGt0LiGbfMxjfYCgEGKWlskZPt1Lo
i7j8PWniuelBaGxtH+MSXBHyIpAB/Hl5iVyRERnjIq0EKIsl7GvbvcKIhUJgrecM
I/sk496c+ceBD9uEKkVs0R3LiDyklPFd8CjGFbkZ6nd8Ghw6Q007VQtPmiEeLfJJ
I80kHcFCY2zRNiXtp7ZvyweGRQzjBhwX3w1XQQiXgow2YJOXgVtS/ekwnMmQ1RJS
XtjxthR4I5csnncwerGhC+YPRns9TIrDM0sbEMXDwD3bOax+Plr5gyVI7WH2kWY4
L8LkaKY43JV3KyIv/A5yQi314ZA91W7x3IrwrAJwj6GYIvDCNLLOKx2n38ITlrN0
ilaYpsuGFJnImUpuLiza3ySyBmX1HY4afGsM9m+AXsMqV7VFqLTR0quIFPNX47+a
cdyI9aARnXRVXkHsJuKHt1B0Nrz2RzuEC/ampZYXQKHd1DWWiJMr4csz2GfUBEZY
ORaXUoJ86YTlDEpU9yhFKWuRqo82BATVZyCPevxrRvzrDh66P0fkkrZfPhMzxzY3
RFQLsydlVqWfJPI7pr1QclA0iIbQDMixrwRbdtavmLJcsz6UEwp0vwkNQhxcpvCy
St7NJ5I5df2mBbk31Hp95iq2zgi+ZRcweEFFgx+CPOxC+19SCi3unIfy/gpF1ZoD
YJk8rOfKRrGPit3vBR5NdzhXduMi0aKZuv0Vb37HwMrVEwMtSMkbubQeDkVB+LVv
dfzuCQxl4nTSanZGwt8H8JykeCmyeqyIHd3RfPzuPxvgORZPVTkhHSKsvwPHjhw1
Wd00mXd99nJ/r8dEAsN7LND1e3s7CR7uJ4eNM8uWyqA+LP0rhbNiMQD9DGkNU6ah
rB0/i3qwqxeUM3KjagzQopcctVt8bhYHnk9452LAf+d0dp4h3naCQLNFwMUZJil1
iPKIpLty61dnrpPs2/ExwSZLQ2dKQNq3Q//ExIluk7Sw9pdJtBTjgAd9wd4as6WH
12VGNccP9kzHm42XE8OOGNQM8L2ZGnilXT7RdaBFz0cA9BgvP525irh3pCF1WSXe
ZKoBicU7GypZ3yod1PSHZMSSS50AYEpVZydT4HCS3LD2fXiHBKTuT8M79qwt87eP
Sz4dFQWp/mb8W3x7TLjWrzoSvRjED1qTL2D1uSThP/xrn+ySn6yTw4L8M3bPRp9z
p5+xeK6Y/vt6vqMqINdE+jljtqTHLSts1Fs3SwAp8iqQ7Nv9Pw9jIdfHvh2yP7M8
EDVW5ajE+a5GyIXKb+zzbl2oX8EhR1sMDzrMBIPxMSiU6Lz2avDY6K46QeGYgCw8
Crr9zqONg31ZZmPuDMYxJ7rn9tMPHS6+eeuOaakBL9ifCFx21tGBLYkmeMD498Pd
g5XaoKzRWOIlQ8WAMZaI6ojibOSHAU3bc65n6s5cZ74YAm/9y+2YutQ6xnnwTP11
3RTlbCpajV42jN3qGrXSDn5FwIR77SUDIGj7rzvbZJ9NKeCGlQtDbx3ZdxnbgECP
7vV8dNarpwLRemDR9oYBS6Ywc5/RgMmKPSdshJTRzXNmpcc1d/K8LAGmnSNV5EEi
WTDX67bCS06h82Jm68FNzQg2D9GGMzM1eJOEU6QPAx1bewlwsUzHBw5w+Fg/UbEu
qmgib0ZxydSmE+k9EGjAPHqTX7zk6ivHa2Tpsew4r8z85J/qB2fJdGJTA/ryTMkT
ocOLDQmH+D0FnUh5ErJaMBX9jVIzf74bXKvqpp35syeVr2DgUH6afQgihAH63hRl
LUhZ7Nk93hItjWuwUova234DR40DdHq+aYgXDKKKAKBrXMmgSDIJ+ghdLCu9nqnN
lL9k7xQPVaY2HoQztIoHgUHoL0zpugiSTCcyza73i+2vMfdgMiTG/jtsxkNa5Zn/
SD9lC417c8yMjoBndmSz3BJq/VekhniHuCFfgSEBNOAqDfVTTpaWbdttjISnTk5U
/NluuITIHisY6a4uPKBHA0KBmeHSb7L0hiNm3hYOUs1ohB6IWVYoJ1O2wtKv2CB7
oW7vbz3U8c6+nl6MfEx3xzrEH9V43XEzsxJqKliOAYBhOU9ZGIT+hRhTdNA7GTSE
jHri3jPXmbLzRLMWB+1Edrx46BYcHD8EAHgVRTSFwe/g+b2jFKlw+9LrdOePVkQr
vjmW/dYPLNXYDyL9SZRlxkiu3+Hb1ZjvpcakEjtUOj6bQPzN8PjSLQLHHOgJfLS2
mftlu0aSJOK9YiHBjXPfETyamEPK+nOoxlNFXuV6qoCWrIKFKy+ogL4Lhx9aftkZ
eSCvOPWqjsNeybvwbsaMqYStY4Zvy5xuewMvmQEXS97k6wvj50uDv8Jr4V3RFkLp
hHLbp1BJasG/I5xDBw3MdmZ/Lgl84UPRn/ERAIn1h6LxyeYLwipU0cgSTcajuFjj
cIxjB1wngSTuQG143n1yqRPz659ru5IiGAYCIG1KHC03FCE/EnPfTxa3Fhuo40+/
Eyj4+zL9omhgOwbqExtqMnD3JFB7tOVfpkNOy3L+XYxdys84AeXB+ndnpix7Cuaw
yu7ctqsaoeGpmHgRYpWic4B8nF88dHMKDtyeTqWRKfrIbShKdkFBs0swh673oY/z
waGhWOchePXD4EboZFaiHoqwvcFtdtpNFkghGtOOOtn0vlPyduLhSjBH2Q/2HWWi
4BY4GSjfDnz8y5hemX8//8QEo4gsudMwJxr4A3PBLldeJWpTsBwcRqT2vvNX6Lss
WBhdigoZrkwTeCpyz3zLkBWi9E3KEPuShKe02bEOY4GL/Z1FjfVbeUyt41DUzH04
rvtgC85Uauk9q6gsLcgPSll5GvdE2doZSdnOHcqoKQTNCAYlsgIm+PhZZuweFIQ9
r3Fh1Dq1s4BqfsNnbTh8B/MIqnEeswM01rhSxl88gL864vSPbujanWXHuLDhFDyg
brr7tGfqkADDsVy16WFfaCEDnESQ4JbozwXDtZ+0NKrtw1yAxEtlW2DDdmCbh75w
EKnPmJgXZi+ghXY5OLuAw44vSBs8WHvGA6xZDPEaKBWrdc/mv3TJgOqEtttnEUif
lOLDh5PT5/avvfVEoqaSHjECZxr41VFKQ2AW8xWp/3beCw7KqSxPkFe0tGN1TO4r
9caIdrdLs7DLOBFQkRgATpUeNYPqskLEsIS2DkBXCh86tmAz8EzHK1dd8tA/2eT3
ogaE3GxucWAbjHNobWI+iqq9OG8ZP1rfejY0VlOpVu8+7ignSlkBqh2EF2OxFs6d
HeYWlqw18yr93k3h7xgqjKRAkTnk/G4QTbUKRsl313PehHBtWcJmdy1Id4gSNCyo
EbRK6PfHxadvozbqbWEC1b7vABSTqzcHiLX0lVws68uvw+Lb1EqA5wDNO1UTCk9D
GOeLr0NHA9S2iBVUboeOBXfFXcl5MDHXX1xTGkYlXeGzlzhb6xOPC7n1dgAtbOR9
xhyc73nb3iAv/u2skfgxfAIndNPcV1cmruGaD1/DDqTGy73iJbDKN0Gupc5M+IYn
eRnNZ4mBAqD1iLlAIDOIGmJT88EYW7yZLTzP5JnyCYPvXpFL3+w9HQ+ll4L9qCws
9IODITM4oeaqLSNsYcNgVvqe+POrKEyUNapCKBpM3IgPw+qokGj/gAZvNwnuKIwZ
8l2kcMC9od5Deng4HvKfOBtiBmjdGZSpzBpr/IhFcJ5jl58QVrmX4U5GqU5gEXti
8oyo9aDCSYXP2hn8GIdRDHhzlYEcO/7HOOxgnMNaiGlErbw5tQeg1gSf2WH16mFO
4A2rziXinUUdyih7PLdeVrkbS07j9d0XCuIALf1dhxoetePmhg5bOjvPzpX6x8Mr
lGmQGrtpRQZxfFZfyyasYhN4nyvd8iAZ4Rf0IfgaE8vn/+A4mw8K03F7V90NDgTe
gNo5VQREbyBRwXdxagtMAIkgulPGDmFoj14M/TDZCIbAgHK+sjTOtgYNfwYnV2RD
ADZGDfduzz8emQdEul7oLC7FQ7810LDyepmZNbR89N070y46aw85uFrSZNqSrop6
gekt47uqyoAdFbeGCG9Svo9VKlxCO7LdodZufvp7xWroiOvKVUQVKkRCnqrSi0bj
5ZEs613M31i5MIqJDUf5HNGZPzfTi1+ANYzEDgiIKC6lxm/vjh6ahVSedV+nWXYl
hwlWWH7oi6f2sfqWu1SsLTMGLcI/LGZkR212Xk931TQ8O13EvDixkjOcmCav2vHT
1Ey3D3+DXeaWoqw35cAyMZzIIFiiR+oxRWmN2PbF1YmwDia0l3amJnibu47JBv9P
AwlTJJvnwoF6VgTJjMKU7/gclqkt92G6nRrlRX5UCbanBGasBYs3j90uP1y2zUXC
LWZs8XdPmSStpJ4fTeyp1NL9nIMg/Nh00rs/Odrg1rEI0u1KLH79EXQnvdxN8jQe
hhu2GCnRfIfKJpiX7whxLjiAXbXXlekjpdnl0a313HmP0tUR6V6JMXpIYgv5qZIc
t5o/dL0Vqde8kr6TFMU85PRTGxuytZMk3h491+C0uwz0WzrCO1mfSGOc9M06sUnJ
I3K+vT/ElBLWu5/3+1iJtpcEsOqfk8hif3IAGewf6N88ITOyrAieLfbnzzhrpWR3
26mcNZwqpOahTsgH6Y3bojwepXAXAslah7oGCYLZxmVdxm2J8j3fPVKh0ts8ycoF
bEXCAJIj4ENyTqSOkfbCvktxIRmdnMCGQDvM03NVw2FIsXFAAf54klBDHQzZuqs3
fqThXOYCuEcguFzKTd7pVxRAiHdB7wPceb614Yn7BVflkX5wscnmXHuiq7O3K5ek
eDJsl0Zqu/5xSi75WMc+F3VNhqRhRAqSatWtVnY/RQMK+/+aipw8I2WHCeh3+Ihj
HC5ls2U1yzwbDD/an6ak0RlsIh1xqi+sHC9son6xHqzPC0lUdRVNRxYJe+lwUsrL
NUnUc9839y/3BrQDuXWJ4va/6YiZbQ2a0bA8EL+aF+IHaIyIQ7tox0J5+ooiKZiJ
tP/SEwkGvYR9ZXuCNhYJIbgDXIagnJUwKrDMGBs3u5G9+9bLgP0GVKrbPBCmEPS8
JPIHXwNPHMHyO8So5Qyp/sjSmqXfDB7cAh+vccZ60/L4fVuC7DuPEnY+MjYGYRSP
9VxuTBa1dwiasGxuarBPMvTPztS0/kGwrw2jyfN4qKdjcK98DuGgc7XWDhaxRJs6
kUOXdMlmRAp1eOJMtYHgFuWAw3SpWnRWN/VKHnRv5b7v5TN+fCT1CDy7ZzzLbOZj
2czdOAu+IR1dkLcLgPpvqtVcz8Vv161hWFLogh/EkK+hlZ7/cEmuHLt0W4NLnYmT
1YVRVwa7Y+rJMLAoaRLS9hdnUk54qiXvx9rfXpmXiJ4gbfPUIBKRk9ccfY4P4Uhy
u0VcR/vHLb5R22nrBsZ0sddtreDpQEqmaKyLn06bam9q1+5b/PMIa9vDdbSPumjv
FmTtB0OX+3k+mB9iNyKQMBH6fQ6DAFrzLyrua8ap+Ty7guGhgpepP3/JcNZ8cKHz
rTZ6X5q2o132rfh7L8V16jb0/sSR73ULsZWf7bXuBHfrtfjY/PWWETUuiG+mwLLz
5cZfIYrSBoiLZv7g7olfZ4YXBPb7ARDThIMKvphnbQe1q08+Tm98R8N0ZLB5b5Kj
PsbWYq+UDfx6Ou3Lj++sImWMQT5cgik8gNK8cEqF9ifELxc1LKsFZCHuFf18tIok
yGErUs9ubFluVrN59KZAlp5z+3nD/5XV2RvFR1tyPuyOaPkQDa8seoew7YcRjvWY
F7J00Os23PLT9ziMJeC3l6tBcR42ewXemWo/g4haqr0QF/klWz6djXMjkSoUJRZC
OViDforvOf6BV0EIGQeMXqiTNRJzY5auAmalQIZlnw3qn+mRtnbJXGYt/NoG1oOt
uMWcEO5yV79BUKKIHABM0mwVvU1oKuMpnS9QCBpl5RNAG6kavTsOgrsSQ8B/r+Vw
b83SSNqgeAA0lVUzF4lAaUu02vKfAzQa0iOdLt2zLR68QZjdwiYZduFjeH2Opsrr
27XahjeIP6F7PIZwyNi/DoepOrDKrv9o2zoHGeAOrgBYlqZC17FZXs4ufFST9yrl
/o1OSR/dlHwTlwUc8Tlu526GLlha0PBXCeYEGzoSel4llyvZskh4WDV9OgzG8ilg
vgGSSfYyUEvW+XXnKyJILDRo9OQidQwb5FvYwAcql1roCueV7H2CMAit8Cy/x3Xq
BXUVt+HTPARy6OWcP0NyopafgQZg/mLsv/frlQsKWTzNdpAenZp7NNpw17/9rvbp
RT4KPcXDk+hzEIvjgoKQqPxMoPWRRCJ51qDZwK8lDgD0pYY5BtUALDTVhSv8DLg6
Mi+FM4fEQZRRyAAA8e/9n6uJ3MxlXmfkNicyvofNQQRVsHiZuLL6SiGiXMrhNLGl
LDQicWfBjczwfyfHjo5VJo4V/wICr4ZqTADgRXuBMkqBfLjsBspqxQM4bkiEK9r0
MT+nanX9VqkQrtHGhDA7GxR8WnWnGGfU4YeavHUnVA6WLfYKiBAqD8JgrJJPqvBE
BqkKXfOvneMhEONKU03gWJRe3CsDZB78F9HnPwYqGeDE2oQ/YHyic32+Jq9T1tKA
MNR+8FbcLUz+qfLhve4BZodF3cvYXXJLHY/ONQkTQQj/i4/Lab+qphY7bKATHsva
+DpYJXltRNpCcmvqcRFrijZaWw0H940XAKeK18X/cyU1wRyxqXXtW1Pga+XMPIsv
/GEyee27xASYraFLFqaaS3X1JkzCAmlwL6ShwdTZ+jCPKvUeR843sc8lUmBhiOyq
SVBoYuN04XZUmxSMtXCw7X3MBRT6IdQHyLDpovlpUjacNN5/dPB35GLWqQWrEE2H
6xccV3e1zFVs5IOsGSeCIJWRgErdwNrkv4HiNKXARuYqcbq0GrLJO5hMQBb7Vy7i
59yYd8z6Yxf+T6kasS35YH/u0m5ip9zU59rBq1rffh4GqicigodhUPMmX0PrOQzc
PfEMV6HZfPjipek/UGCzfrhWSOB31Ppng14RCVqVdR3xoiUZJZT7BjnEmviW57NY
HGBeGkBYsemcl40qaeFoPo9mrDr2YCMWEah+yoi2FHpiosBdi28TFfvPZlYrmD2D
i9Q1YCRTmerToAxjg3lRv3lxJRAiI3COVV5GUmQIdJzNWKY39MJgAEgKMH6RBI5n
l6GUW9xWMJJbmByvC3hQJDYl0dYnH4cd255cZidhqBRhwXkPExeVE8E+QTnkt8yF
QmlYHNjzU2GOuREV7XlDW8A3d7zDfLaw7cDmGDR1MJSZr+s6JUMdtBGcoegFJiUq
Dzr1V39ynkO+iQCNT3nxcICEkNm+2LS1febxWX5brfoMWd+uC4671C90FCyv70iF
+LPNmSOmB1fLia0fkd+3D99EgWdtGY7kRd9H23QxcoS3oTnSAU/uSLU2youZlwxN
sHamARUfUr/hR2C56ppEmxiHvVB5uP9vCESsrakeloDSI72hmldKxjP1jWGpcaaW
Y8o8zueAonusew/wQX25JFrb+mV97VY+ChDL8UapYn1mSu3e3vI+EB9U0EK3WeGa
GPSrx0Q8qHP3a4RcmIqfEU9AAx/GuNT4C2G1NwiqnV9kshohV0QMIrmvKELb6HQW
Eo7F0FAcXLvIStyh36w+sR3qo5ivtHAdSHzCrSighQbycnJ/0Art9tpOHVp0t3gk
90hUU+JCCVVFwz6cRMuy+Ktef3KmKk7uzg4VWUOrUtF58f3EovZyG4I6QN12AiEK
OPiC0WiX1MIcJl6Jv1d1yQ9vutFDmnEwxvnWMoRHLNdlKKDkszyW4Ux/iTXCvGz3
im4T8mz/grBaNXlt0V2gopMuCEKAk+iz4ztUjNvibrNp1Aj/PCZSDqiC5S1Ohav2
MIwDuq0Xn5pQogX/kkXmghO+BthLLubcP4dybXC2Cd0hACSKVOVqeg88JKzn00tu
1SQpkk+MegVkdJYoLKYwWwcAW72VhpCAJdzvl7AAjQpkFS1Y0om+ZBrsGTJ6qAvG
/gAPlx2X9noJ7dVO8WBkWELYDp6/Uqx+JGgRcGK+ZY7rOn8QMmlFbZO4dg0gAqvl
cnSKjIuGsGp58RtlzXO6Jx7xj4zY10BPONkTBrCXCcL7MP24K3bAg+okje6t328l
tDrDRAJeT2hVvx/jOybNCUO05mW21HdVk7RIXDdfOVdQdc3dTlRGWdSlhlfzPlRa
F1UE5FNU6loWoCdIjhlh1GIh5qTdA56xEQZ83C36fZzHYQy1Sa0XlEn7gkAyow2R
/2yhTAtKEbahxCp5jv7YjMZmi1Tzj1jLkJUO1ahdlbF4guhARA8iIeS9fnvCh3VJ
rL+kMwBsrMUg/Wwkg1aMdnsXFg8S1bEGePQW1GsuKUhEyDLD5Xfdnqm7W0gXiZVJ
RSjpV6JQ+2IrFBuLAef3Ffa0gQQEy1ClPmubqU23YYK6hVxvWq9u9+DFqqtE988t
TbpVW9MPKEL8PltswdCr1T467r2IZLAoYHh2Y7QliNT53fi/RtLprpWBS9jkyrWL
BVkv1UEA+hVXkq6A8B9qNXBFt1nxSoZiIXQfkasL4wXjpcN9bwCFL7J6u0NXjXMY
mw0O6AeMAy+w2W0/HN38R0b05+sjVSKfsY4DM4KCoDueTleEzeeZvfSbSoTfFSDU
IvkklLp5/+dJi4zrtHvK7Ey/Mxjs3AdbJlQ5CTameEW3RspJ+f5COB4b0vcvqLrO
RlCbb5fwYW4L6hTm+YItfgGUTvKToVtyHfcvzTJn0tqexKXts4a0fmEUu/b7w/P8
3roLuBOqDIKD/b70fYB+Vunyqo3wLwxtlv1Brhi8jzAGvxPn3qrq2I9pL9Ada+tl
rzljtqL+mK2Sd7KHBbwXqChsmUYYEUV6/fEv6RPssPPXiDpvHOoCXsb9GEh9t3Yl
PEbAk6OV4/2Dmv112hsyVlvcc49b/L1PLVbjlgH2V0NAfgSBvvT39PEOSxAGSpl8
u62cnG35I+SnY5xkCkDKMRpz0d5ICAKf3gY7049V5bRqvmeD2xPcGwztAUZQ0axO
QEHRy1Pz0AwsjngiohB/MwXrS+gCWo7xusyr5dNfNf7k9jy/T/Udyfggqi4LiJsl
kJY1eFQjcw3nnDb8iELzE7rRd1hkkkZIl5VgiGKwsjSkGwFt7MrbK7/5a6EfZroN
DKNOA7cRwJ9Ibx60LOKYK2IlTppqWIwgGazLQbifrJXUHP36QRoW30ZmqIheBM47
cDnalaCHo0NmgW2QyXNbjoxj/dpVJWnLJyriU5r4qkHQRTts6HmDSkiLGTT/JonM
6mlrL6tjQqX5H5bsGgv2sLMzVZ3+FXdc08DAH+ADAgcLRMYhGwr1EuRVut2cl45C
Y0pjipZqUwqMXsYFrnNE6VkDWM4Twf8BjS5BzL+kc19kXWX/6n3Q3ZqFxQS5+jXi
9VEqOI/r5clv9+d50kGbLhnnLOCtAgxtR2rs+eXeMteKcLIvFvLpVFQDlzenEAWh
yVeSVUb+zWCeWeW3ZN13OI27pRmszo3jPs4bJq0iNJE+CpxZy63ph8LceoY2ZDLn
So1kfdoQkt6HnJDa1qz24KtNKLN6+kssbKqJX4v3tc2YPBEsfCmze7IlrS7ykBbv
rOlZuUOJ+kXW6pANemPVpRCRQ/smZnBzwcFojmfWE2+lkhS+E783R80/jXnCcmNx
d3PN2edO810it63aCHfIN9E2JQH8CSX1uBL8kiut824R+XqQypSVOK2/Ot2gunJ2
yQoEYc0MHMCe3s3KUDr3nT+t0Te8Kc08FKWPLQiH3V67tbpWN0QP06hvwkLhLMrr
0bxtWefUy8ZSkvu7MpDX2ciIV3ShLO2xYk5DVNsQxLISabUJ0eBAeUvGU6VoIVfl
t5jc7VlcFnOu8OOdr6qaVj/5ijmCkH9lQMpsbf4urlRYrEW7o3iIIXP0Y9flA6qg
eKfCI9aScnxDSQGOPSEZTelND1n+0pz3apEFO7c2CtxuHkthvjX3Td4b8z/jWs+z
nInwzubp/DE2RxppM1yyTAsGqDAFpFnsMe8dg8ZJCBXUQ174IUquMFg8TuTPQB9p
OXJz+1FvcGOizUdU5T/iXFlJdxqloe9VVLE6FAQ2yV7aVlgLLfHKWMB3d3A6O9BK
0NYMamXi2WZ8FuniUX/67myF2LLkXiroZu3yHo8xBaDhRCuo9Kz2FqpJlgDI1UiB
Owg4MtiUDAAGyySPKDVmz/21HjRT7vsxqNG4lnkiLwNhIpxlNnf8n75XhTrsYzvJ
F2g3kssvQ6/CxJEDPn9tP95GmlgA3NgRP+FnVtCnNGlSDD/R5vaxXyH89DCcuVFt
mSaCNUxzsOWSG8pYOR8gFRxhXUi6DiXTjXWTdAn2jT0kOgWH7K3lz7op3sjVIQ34
/Y4RLm+6jNrHlV0L3eWl475dP+nBVzQwlDRtSqqvFv7HBeusaWBz8QeNiUjtBLma
qHmI7JgPH7oH5KJ4B+pAkfhNiDdETrjN0PQIa1Ac/8dBmwclGKrxGfQqqJ8/C7zH
QRGPeZhfHjoJgkfpVProydo9HN/i+jolX0nw+a7MxpSwTTlBClAQFuYjEY7fBiIH
z4kj5FxDiZ4HEj+ctD4FTgiP2hPPNrf+T1LdoVXoOoZgLvLr7Tjww4/G68Z723kw
Csz+/QmVkvR1TGmRV1Thz9mfPG3ug3OtA6vFEbW+QXF3qRyIuy+7xdbTkbhnhiBn
/BTnZgp2Vddi2qZmmTFPSY8N5DXQf1DloNJN/xzqRd7yWINjPUaaG4PFVCqAjpaZ
HJJPrx16+nE5vmnpDelwPc1yu4NAXVpVJGhPuCkQtahAxk6JmKdoPVmYiiKgDn7M
psQ8zflHRIaxdnIE3nYc6xA160zoVZmv47BQ9U060QxECcIDvnaLh3Bo3jih7CUt
XiWyfHB9LFbZPg3Agl/9azX6xHQ7na0B3emGzqGbHpEZPfkHszh0fz7ruPC96T43
OWFrZkZOybrM4i9oETaPUhowb8yfwF/RaQd6SXbEeAt2th9ni5G3rKE3w8iE9r1y
kq26b+gVpJAqyczkVPT742f6tHs4GR9Am9tjN7A7j3vIM3eMQt51Qms0e4fgFQUE
128AX2Q51jpwAGxjvhsx+HywS5SGWM0Jt1PfGkuwmK6fSflrOVHAcLjM6Rw8/aKD
O59lGL7Vs12RDzQv0XIsb0LcveUbrejcY9cvltVmbLws7oj/U23QviGeHCqkDz3V
+3Ij1qx9e8yKOfVFY9jwrTD0H+V5Q78ITHvIKAbq6BnRsG3T+qh/H/DApTONRb+n
+Oc03a1dp8hvh61jllvOlIUj7BQ011kyM8KnN0lsr9jDCsFKfOGte2/eMKOkdRT+
ibxdeZ5VF3QnXUHKwjobRo9wgtSnicb5CQqHyqqH+/2IluWG8KOfy6e5xcruBoWS
3NVf5J0hfP030lm/JWCWN/K42ecYTQg99mxDJ/5AGz7E2SUqS1CfSRs3A25x1/Jh
/NpSyPg+Zfk85iGqvVaJ25KRnPPPU4WO3VitJ+hGdvqtz/rAgy/rJfT2cXO99Ou9
PpPknoAyf/ELAdCIgMENlnEepy5Uu2+nshpPFus/JE8WhR3G02841Rd2vtpQ0/Cp
QT/yZ0hBeb0+kgB2p+8+Mlqww+k3ZH01kXKLdujOITku8tA+9I7RQ1Tb2u6EWB1v
AoV/kNdrpJayvxa/ruQlFyRbdt741SGCpqKnnydoVY6Tp7zoZT4RJ0R1t+mvBKUt
3LI4ff3v3sFcmLX8amq3PlZKSBpnN6qElx7HcXQzlLe5FzIRAzPtH+P47a1tdUVl
Mo3NPv08gQMysZBFfEPKnyIa+u7iUfFM62wFeDAcb2055PUIh84HGq5vybHKd5/9
UFzSS3iHwGX2208sPxXCRQ6meZ1B/MGfYF4rz0xvQFdSmXN2/Psur4gewEX4gDWL
seZmuzdfYtSOj1+KDLCopi48PR5gx6QDit5yc9+kkdJdetABQWe1zIvSmPLIVfKn
wDElF7BXmWCzw55f2ICYJPE/uGDf2WYx/RzygBkQEuh/Ruttt+yp32WUW3pQQEjl
bJCiQInAXHAE2K+Aak9R9sb81YCWzENG6n8it9chuslCPklNz4nc9whsHxqM1ySH
Gusd9ECkGWUrfF6lIvuJLvYAIoGG50KWgbYHPBE+AtmRcAgD/+Hk2CMGIY5OibH8
0fMMddRPhExJdZ8CSykgLs7Kr2P06Mxup6QO9WsbWYuIj7YdxHfR9iWZtGIBD4WQ
F0f4/ShpKqo127FW12HXJF63WjlU//RMFgpbUMdnbqF4GZGDSDw2PigUqsL4OsTB
oNHLQT9pq1culHfB1pFtfV7e5+yVGumfbMzzB6tZuTwtKXR1/aSHDys3uPoIV7bV
v2LmeiA9fLLcaKIaOMnO7uY3/N9pK9scxgrjm2gGmP41ye/DCy1DWfuLKMFIDVwQ
qDWeTGj6jP+nWCuhLLxj2JxyLytVzucMvRfxh0/8djoDMgK/Ia+da6akaHLsq79S
nmUOvvX8ahjk/4Ic1wfHMa62ToJMy7qfK/Ht3QWdj7fhSheKOm9DymsthabThIQ3
u5Wq8UX2EYCKWGt0D1+jVGPfu7ro1bE/OCO1ULzeGIuX0rgd3qAQ71LfyPpHXDyf
gZrcjhDVhynqUWrf5TMEtLx7dN7UHnaEhPVAJoS7eeNCf3sie4MsDjWLJ0NLfcni
3pjMtMYuS54pw1L4JA11r5l2176wPcNH0ccVqAKxCHICwsPym4/cTwPo0tXs7itJ
fgNnRfLZFhNhorcfux35JKaHTgKUgrY0Bu9FDr7TF3Az4Xq2uf12uBD2UgbqW/D8
hkzZtWv5Ua/dUSQT4ZT1B18MhcDVZU1Qu4KcfPv39BEOR7cACygnkbOoyFMTWx4w
soOpK3+Riw38NHmmChqiC4dgsQ2gPLLOLSBfe69lelSvBMNPc0YxGVfr9V7tV+Ji
zDXKS1YkJhXChFYLwvxbeNuaXJVst+lgfCxBKOC7/WvseJkpbPSDBK+aO7mvpipu
4ym0cYsw1ffEyBE1rR/wDYqIkukbMAT1v7zUcpoquE6kftrAZc/kndy4ASyT3+Hy
Wh0P8V97VecsevxkUgq3BhEwDQsKQDf9Qb2SIaufUS8VW82cxSD6CKmHp0RzKuU4
S7WIJGJCK/vBmLsGLVk/unxkNnKyrFOYF9rU/bXsw//OdVTUyqI5v6loDYxlqLIU
X75DuMV3L1tIwKPcF/6N7c23E2msD5yQSmecU02VtdzeEWQ7BPvlqqukJvmawNwn
8vUwHuIDkulO7XVC5GURgzCdhyXkjbMJ1g3OIcyhbw6sxutV7e1PJKiyd+navrPs
YukEUcoGxR1p+cbqVbc6RHcvJpAuDjO76AKPocljXx020MLjkUk77uLjdvOL2zyZ
NnNTByP3V/rXonnV/NMj0GMb9UyFQDEm73+cr9zdeTtgKAJLvAOcBWwKUxk8FM6G
f9N0qV2rSFQjCZHfv42KGpux64fS4GfmSfdH1LcYdiTkNznOB//pNlFzkqJY4UiQ
O2BCMI/e3vsN9c8f8NmMR5SVstYTq9cEdtFIH5x7jNKryj1R0DEJg9/ONuk3BvDL
Z5FOW38szNZFOv9Su0CHNucnM+GYr87vH+N0fTT9X41qp8IonH2nRHnvR1b53D6k
fRPjA656OTY53Vg8T0PiWhnVSiICD0Jgwpem3g8WWFREloHCAV18a5FOtTbqGFh/
3RROycKz9MHpPft9Rn/EdvChcuc1JQ9Vh0zT7JICwdWhqFRCOI61U/4n/TjE48qx
tD1T25UPplYvOktOZ5XBSMEN0p3YPc6JZA6PGTBTo86JYYCMf3+94eUeGdi8BJRU
kiJeDFqeY3BuusALX0MAO9vgUw0z0WrT2b8bw0jGo8o2vw12Qd5r8SCd177dSedv
ist7kJEKA36o/g+q+O8Cq+DpvfY+yPgemlW7eP5Fmyexmo42KCLt74H8U0G8iiNX
Mvxqb4cmAzenPrFxTBTu5hbNA7NjTuyBtB7FkB7qFmWhrS4MRoF4cbm9CtixXYMy
zBfCQ/YUAQfBMX7EBs0hQ/Zlvv6vMhYFSSz7Q9+rqZ7YISynGyw5zkXmWZHnLHsg
7kzOuL4IP2UmXmp1b//BAA4a1P+EKaKmiTnJWL6IxdR6e/q+lc8ZWg9b24AgxuS9
Dp9i0WlyhsDfxyk5k8ElEsDfBasUB5kQszJbrYCYs5B1hXhQnDoA5UZMZ1qt+ai9
MrahtEoPFph4mpArWUwNZ7XMlIOYFXLal8d47o51aBO0nnpgfIgIu2g3qBrqpi/a
lYm8ws5jx2eWl7kZ6Hy6Yx19jTZ3WGSwzM7dUvmvC3Rw4qYZznh/0fOmOJdtSVNy
fH+0kR98Bn3faozX5Qo5uJdpU4Tha10GnEUGmtVsXI2AHEO3jI8ucSNmSlTQr5nG
0+wc2bpfF7TepfZXQZ/LcvorfujY2ZU7UcrrwcN95/XDlPEIYy8Ja2wMTGBubcde
Ehn2eh90srsN0ClpoLM82r6vFnNX+jlgbvDkS3Ma+/XKlUJH+3Mi0/ZyfeePsXbE
c/cF187dBkaWk3B6PNFivgxMRvT02g4TD3KDu24O9gbit+Q9Ud5AQoKKmudaIaHW
nj0MDMKGp3msKKDTOXl3KPN85eNTKaCUNMNDGKKjV0dLVCPdgx0Vdgu/4unC8Vmi
LaeSDdQJvAXOctK2e4EVq9Qd5ovmxb7iHgZUQkE2S9Y4qm6FrnL11s7OuRVEPBAj
k6IBQaZwN9PUcGstltO/uDf4JACnj6miedse77zfGfewZWFhwHu+Toog7GRv+lC8
vh85jDlcoqmrSjg/GzZ2lEHJVTRWPcMwnLQyPCqAxEzmZ5H0Gpgv27TNODbtze1X
idMkSYrA+FCbDl4OmEmDQZI4E6n7n9lg36VD8FgOtpbz57XeHTYYj1bZoIQaiKSE
pW5zbvCaOjPOh+4FM4KPQF5wyQZH56wz2gMRhX7yf5GzRL37OZpT932+dTJ8W4Pt
Kp/G+dkFPenX7stsJ5V3FHzQf3miTvSgrvPSn8GNbjwL2m2bYWLxQfUtcw2nh/7D
I2oDxwZdePmGReEEu6ULwrAWkDVhNkySQYopu8dvJ90bFLEQDqfAsG5cBWtO8FPH
voBvNoZvaKECI0ahTA+FDE5YOxr0hNg/EEDH6d83Bp7rPbDRhHTmD1crvwlMoAcq
XZagpd3SWQ+xe30f3XHI8fBHhqq3aM4fBJi6bCxrVuGQlVCHCxFVSGXPvoVSbNW7
2tWLha1+Sgfh9B4y2PRpx6tsXswj35hmUpAIwzfJNeY5zm4YgqCDcTLe9wjtZTx7
sJU81DfsRHFMsPKpH/WLkwz7/rZSfmfM7HPh9awrU6X4MSRS9ErO6b16VdxdATIS
/GPtSkw1U7oM4IwPhwtWIN6Ge015cg2cYYgRJsBSx9AVYidUd+srg8ZwECgH6cau
4W39v755eQpuW35yPJklHUyGiFy5I94G7zR3R51IbjoPvIj5CFMEDW9iAxaKTIGB
1eUJ1Ny7i0lgl6yJW99w6GxlpdP3zqUxqzcnCktAZiU39GJjVpLMBpUK9dzpJZ0W
jL+rLSpkndHP2LQjNe40qOOnDnGCmtEzNNB6/5QCPqFH/7Z1lZkmZ+LxKGD05JGf
kLV1dKG4sjSFE4QNVBCFYQcoZJ52bujUUtHEwuSOreYOlTB6wsAUlXwAa8jVKVvP
uGAyPvmMAB01tcNHicDwm5uT+D0cc//ww5B26RUAawwujvmibg8PkoJ7D9Obc1b0
TUAwSId3oK1vG0zq12gg9VwGyT9u6IMniSt+CZzbxuMiMlnG5tY2eT1LvcezHhmJ
JymvsvRjP3cz5uGIfyY2h/2yG+ZpaDyuhiQZWM9OXCIuLs+Q5McubLksSkcNPGw7
SZtXRBxwflYJI3Q4tpSLbbFjCdj1AAmCn8kYcSp90acIZu1fOI+ZwQk0OUNsy5Dn
MyCx5Mgyn534CdJGK03DTC/ObYUiDsElxVkJGRWKm2BLk7Ah14Vqxd8gHaham0nZ
N+zNUIqEXEWy9dKydYt/C0uzj/EaPTOw3bwCyhmCGMI2YSTMBoBubDNlq6GxOs/V
LaobZ5t0ytyUhCEpOvjKydeiTC2mGjeDqxQsebPuAagbXCzgNARDgXDGfsUTTHpE
bdlmgNfx133KmYDgU8KfaFsS00qpZJSVlYw6WErKhee0nkacIjfOxj1hiaa7fBbs
G+un4r0tP4c2AhnoIE0UnGM9itaY6q+S7XtUdxuCtNnvc6FCHqmlb6tOJ/jYSIBz
FnTczJeOhp7IWwnlzWxWCtn7rH/rpJMUvurzDp1IFxd2Jl14kQpbqJLPePjqJ/3Z
WEy4T8ZJ4f5yxTpN223yAzQLRdBU3LAQKKNA/nopqIhGcykxooZuLymJLS9LTTLS
yWNZ8jXNjvj3V6p5Ecab1s4kyfChzRVbrse9Y+9HGOk/wlPVQtumdp734D9khkhR
6Txhadxci0mMz8/6t1183U0gQTI0QkzlcKunoPRQrk29SCChaE2mguNScyxNPCda
Jo3E9NzoLpqyU8eHhpz1y9t0Od9E8yoPA+s4SLSB8FGhOwj8X8+rNOfDkoGFQABM
lloprNDhAC22whqhxuwNen9lb04ZBzOo9ussqADzheJgpbHj+wxTHazLtjkSvg2v
mZQYtlCC0VWMnUhwCeAY5f1EpdBX3SclF6MD/35QBf/NrqV9nqq00x+I4MlFK9yB
sIFW1GmvbFracrwAlp2cEeKTw3Qgo4ewlx7uru3vCeapTl+5gecezhgyqZmBHMlE
i7ZRuJYxpQwD0RPlJ+zvPZT5TcWWPa+TLzEQzmRJAKS4dhaHalwvQ/ULc07R2VLt
ROJH5mrr/AKkE+MEgmyeVpEnD7VPWbzbpAg8e7LycoV3KkCvrbx/drPEjsKehkOA
5s7uiEbMLR0SfICb3H3Un4SI8y/qC1zrRtiLAir2HHuRbWr2ii06hmZbIuk4M5cS
U3SgI927YsPq6ZqkBsXoLth5J8m/D7CpbOXVUUXfoPp9+H37oVFfQicvdQX95J1w
6Ow10XkKgM+kRvvux3hUDLVPf9enI0b3EeXWKmfetvsxra2r6jhVMe06N+IbTcQq
k9WoGVbiGSmBPCnW/mSNFftDP2fd/ZUVhFqMmFdvPegE8NSL/dt1PmL/LC6WQDSW
ZnMcjIfsAvA2uALYcc5QaQcy8OD/Ofe3Wa9TIXiyZPHJkecAKEHcsw3pnQq7zCUg
VtAlgpmwObpJf25Eyla4eoxveCVDMrE1Km7OfswxrRc6ZR3v6s2G7XZg+G7WwxMH
33nD4Qs0cTUfeSUAA+UF8fzx8I2O6LDhVlaROWoNcOkSw3A3XqYoe9nIEAJRFocq
6AHbKPj4FwHCA41K+AnDa17FwnB0GQP/yBwc1QWN/mO45z2BxwJ1CA4iE1yhKfLN
0l2adaXkpMUanWCbUVybDUpSWAiHjVZkF+PMD3gy4sH+XaCebexK0PFHMTv+i6kM
8HCG/vEqVa4vViA6XW393GFtyeYBKJ+DU+foxZoXZLFxn5bYAneLZW88ny99qHyu
xzjpQ2ParN1d7HtzPZNUAZtIBLf9Tex1PsGVnD9OaBYmBWKDTfzKgDHHPt16N53A
0YMmJRjM9rvEDf/bzC3DKmIXy0sjSx5lCVweXmL8RUm7AaHAZVzwVBgDqEoMQQQo
o+kaRIAquOQOI90p2SoseSHiqUsZwBZ0VgEyjQk5+IifoXYK5wEbnt+thDU+dBhP
WJsqoB3l/ktPIki0vv8uL8KJm1+CfDuTNIXcdvZsjsUnAENZbdO1ffvzh3trYV+G
Lnz76B+0O68UtvnmE+Q0xfVTWZOFIPjIilo81FvnpQLSEzmTqArVczgX4GkThXjb
bY2dVylFiU1Awdiii7l2bKRLbTu9i4+zapKdfff77K6pMIHnW5cYuOQb+BpEGiM9
0q3Al6g55exi3IdGBXwOYHjqtZ9JmrUbqwJ51dX11Z1h/7crihKhWW/yj3KK/mBf
Iw6SnD6girnHdubBNdGL/r9buAO5mPvNQ9BDysNN9ViAKs6lmlGvQTBP0xP4/n3v
1L/tCNpx9MI061VyzjP8aDLSEb5wYhDPbscq0TA77rJY39Q3WWwdTEqirD9OXL80
i0rkvIGMK3oAl7xmpKnx8uEVU5m6OoTAlUsuFkhEe4pHTkeRCXrQd3e3XnqZQr7O
2JrAwRIn6JftYZSI43+uxCnytHqgUJ+GJcTjXOdit7nanyDOyayY4MdVC7W9WmeA
FwiTO/fGqXGb+XIcwQIQIyHfTklZ87ZfWS/r2jHCHM6wmHyi4LfSY4AlVBRiBKSW
AhJjMYzt+xIplZSWsWv7/tfEUtW7rxcSr0/rPRT7V87n3XpgoEkA0RT+vULx+YNV
zzasCz+AxFnk+Yj48wzeHO4MQWoIPM+C4NJWTHYkoN26INzVOh2eAyFRWXRysFui
aCb6jIE/RStseOXIASMPAOMbrgREo4bnibTYqA1H503c6v36NCTK5EeY6Zq6kKwL
VyV2qtWdFBRidCbrnHmT8LunfbYJ03Bz4ufyc/zMiNvSNKY//Ek9NZYnVmnIaIMW
FO5/tKJ9JEy1+64GJaEWu0YpszzKQhrYlVLYG9GQoiQOa2ZKn67MrDuyWSCSir7g
td8dv2YVClTaDzQzQA/163pQsKHc1LAJUxvIYuNGeH9++Dz9giKWbIUkU3HPRbGT
FzTOyXokMh0YeMK9HpIooMMT1X01vABpYFAT3kE5uN5+c7SygnTEB9mj5n8eD+Hg
Pzo3IeUEAeX9PsjKRB9V9cRv/upRXmFMaqgzuoTexG/sQ0W17m0VUJWYKjICn56F
B7USidXUvpgjr5DBL86m/zwuQntXOWjhHP+PxZWvIBrE6+dotWbjjuIeG0krAJRm
lYaKSIsVcbJ6EXAV0SWE4rlrrk/VEeEREQHp5zm1KswaMUE26SZPu0ys654R4q34
y0snM/l4fK4p92NJakKoddBn/l0dvzR4FL4uXvagKFKLXsrCjbd2aHP4S5D+WXcq
z/DxWUQlEl7A+RySIwf0Xs+EiB4G5roAjKm6fEJRkcL77IoIBhbpgO9lv75Wo7T3
kgiQUfttUeQ5KG+oCRP7k0Ad8vUGbhGIBmCqFqKgyXtPI9C1CViYvYfSbjhrusR6
BA6K92IegQwQj+VJ3WJrDU4j5LYowVv+HbPSR1wTPXU5BGgaCmvBYPSAiKtCncnM
25ABrbUUTeC3QEJGGTsJMqxxz0FcrOCWLapeMIMwE+z2qUHm4cPWZHXelO8vH5vm
rnRi30x4i7ea6xME+aOqpZ+CqeJxkWCvEKuarfTj+ydXjvQHGUzq6fiMNeFt7XeD
8bGQy/hOT4af7c53nrFT7FucGbTISwqRh6TF7BDXsXqCVw43z9JGCtxx2hnlrNmy
uqZGnDEi3RIq3oXLi0rbM4n/DR7J/ZE1utXWKJfP+7/gtS6bT0RUUcTUCPf5vD6T
CzTL9FSHO7rvQphgNz/PnLPsD8qrtWzxLIhBbBVkjPJknuWrNUh+oGafqEaurKAN
vqfpeveIw2EadMsaM/jV6rIfWagLMDgXn0UYeNoi5hzloNDSPbPsS538GQ9KhCeA
4iS0dQN89uAjx5uQI+s8DX7XHV0vbZz0aqgCSr9sT2422fbQVl1jnaO+W+0mlgHp
Stoauyo1LBE1oB1S3NkKFQUaO8b/Tz4SWca9OT/VTNWwgQJy7+GQWJsycBQPx7nM
kVWWk95a7TUhvGGB8UF2aras2nUjWxyGVos0Duga9qJE+4nG+cjvfy/8mwFlpJ9q
jzZxNOtgwMPKRCtYoMb8vHLgGq9DAlelNFGdzV7VsVaeOSw0curzbpzD+exHy1MS
Sq70mJyRiKo3sr8zWXE4eswmFfQG1UphVR6jF0lFANVLzT+YSmWJkwJW3f15VC1l
Waou2H/sTOF/kIlme2jDLjcQLWq2jtbW8YOiVYU1xGdQxZA46VHVmQtrG/0k+QAz
VylDMyxdM8YpTfSUEvAFfAINCnpd4Sq8/6L7gGNvbDO+c2ISQNdSNwVusSj43/8M
V0tuq2vnWiqLyGrRYsfY6O1Uzt5A3sMkXXsxDQj/gD3C2KzzG/JKKy+9ztjn9B3C
tiMkJ79zTyfksXirwhtmgFNtMEhgZQwpUE75KaKg+WhRqgpqS/HuUg8qe9DAkybI
eQg5Owdt5kKhnnM+dB+ONpKkbllocY3uXSuHqfqe3p3KiAywB56AeH34s8wgnbFc
zPa39rDgh1DFI2h71LUvWQVVxW+GsulE6D8U+CK8gQZnWKJFLIYLseEsf864ESqr
Svlw+YhDc18arVUFGZe7uQrkCfh0Fn69Ok0OGuvo+9dGiWr8TQobcR1QVFUOTioZ
n6LBLUOLnJtjOf8jttt4M+oF2JQrY9Mc2q/da693/w8DRH76IgeAfeGdYtJ7sPjk
ua1zJZ0OEfh8LkiOuAWeylo4ef3BJHVwECNR5HfjtKR0GdrvtU++vvRSSCkhaJh2
WlGW6D9QQkVDNzrE6myW4q4Ft/0Vu6WQV8115jXyS2S/fmc1ZRNSja4wN4Xp2IpK
kR0xiMXNuXHHbhxMP5RV48eFckOZVnGbUdcynGM0s3Sn84m4Tf2tTGbG+dtuUKB6
QTJ1pMmwOjHcCYPRNLQUeRbJIIgdqypwFZfDrJ61KiJujUkU6fOrwwYZrC5hrW3Q
K9Evx9xzFV+fdCmAbdhmZDmzaBqZEFcdInHOar/0xy29Egi50YXyCszwN67nfoFk
8V47RxjLPDAAjAUUTNfTriU3FshmMD3dJLvGizft7ju0QXCpyRs+w3hr6gruh5RX
aaMIkJKOc+lTWrY1UMzxtxknhkP2QhZeRXNeS0yIm2eH6pljg5HFgpz6y+AHgldX
n0M0ejmPKz8VgPj0Cw6dlfWXgkUdj1GdnE3s28oqXayq/NrSodo1BJMPdLXliZd4
7YwSHyTMsnIiTXJlcu7w0U2J6b7zHz0ft1K2BtakYrIXBnXGvw/zfEqhdTUQQ8e1
lxqko1n7xDbiJyVjNsxFPj/1pDlafhGCdlzBQDzq3+NcHH+LCe25Jlqt01GQThxR
gPFH6oH/czAvz5oWk6MLhWi8umgvOsVNSUmP1C00U1GYX8HsMU+uHhrHm3twMA1k
NTLR9yuQZ6KyQ+P4JLMhl/H4hRCpFbJNtjK54S+4Wx3M9F9402w0wmmJmxRL7ORH
wJ79d0/GXYvjIJotyHQe2iGVqmcFbMWUMwiZfqD2fb3WiqTCmMqDTI7rt1gQKZ62
h1ILUVXQVafue7ODpvfoOjOwJ3sDQxGM/h22xeDlJlHf31k/oEqCuXigFSufRF3n
+bwrCjnHYycoZcWlQcxKUlSdr6Ngt5Jk37unyORO64kwKVPhB/BdcSj8cwh5rOKo
WfsU2zsJGcz8Q/BCqalhnZ1Yecas1weXo8lKZXrJOUUnIvnz2uFSR78Ck31TpZtO
xuOIzJCAyhHnC27dCefKEInAbXeyoar5bdQhmgkHfVAwotAVqYC/IyVzWoVqUYAf
BlV9jIy8LXWh6OYEMPy797+d+QOUpxOTu7gsBfvvx4uegEXrZHFQfeXnezdamL0g
1g8o/OvIRZoBEdxxh/PEo+pgdWA6MSOKS4GmksKL1P9/U0n65GWaeKH+yIVkYjS5
cscfVS4QK16+4oWWWssI80KBLvv3bSIkIAAH0HCh6dxxN37yMeYXtf9RIYh7C+tt
f1DrDk9YR7J7renEa6llxe74d057s4Z9d6j3YVjzWT0kkHS2rZw6uLogvVvr4WUn
E1myvvmSfidE3d7ZBHlTWLhL0ZWJWhW7SJScCUQrHSBSyvqczEZUj1DMQQZhOEgv
ueb8SNP5TO8cO6K7s9drBCODTi0OvznzPRVeczD3a/BFvjbcfyD7WTDPAHSQHEdN
Aej25xeJtdN+2CMidoauhS9m5LIZgT4hE1TtpJSVAu0Kdg+9wNyV/CovMsfas3aG
ceCHJePA3sVPec8ssPQBLYS1gIoatMOye7Gc8I4U2Iuge8Csbtw8Ota1M72Y1q3L
KGmKz1kUV+pM+GS0Fq3wpT3d9OWwZkwPOWNnBEo0RjupjyUpja1pqvqlTQ017Rrn
/7C010oZ/x7svffElCksCsMZLGlRzUyhWGXzifmAXqb8eVyOoCHRfGsa952niIn3
6aWXwPRNVkAQngE+RqDTfBpdkJFj4Zh4juZ/6NKZL6w/qJCKUNsnMVVZpHbcLrOg
csU1DlsIu+o4C5KUSYtCFf/awRdCm+DHV4PljgSG0AUsKEsn28Rz8+x3eS+hdfra
LVKUNiP9UU9H9Nd2J3B9EBiqEoZz2MIs5xVdwrvnEK0U6VuB76E4DGsPKgNKjQEY
OxRnhp2tZTRsatHs9yc5a/9JMGU17FYs8zvIlBrB6M2XRRMSsbJ9C8yihcrW3pX1
OKyfpiux7hPlYAD4ag9TD6Cf2xzCfxc8A3sDqIRQEroUmbjCMq0zuLJFnktdZiTI
7tIUzLqsdT8WMEcYFJjZAms9KAWGxMUUdPIONCRNwWy1OKVL4tgfxgAbG0WACgx7
kdIkJCZqjo9ui+6FPA8u+yhbN4Z39NJvJ+yAuyF8AGp4H/4iGAmBryJ4XqzBR0uw
XoiUYu3sRh483wnJbFoe281WKaO2Gsafa4KFdzsij9tHWBAsX6rL8OZnhvJiuqKX
GuAPRG3iyNDLV4qqJTqd1SmLyDMtOWwYEhXdBkR2RXV7NlI0/BT6eBRougFdZ79l
jc6aog6uK8fl9IRmcKsZLBKPCuuHfEjpTAvJj+E65cvAvKsvvEO+dZuMYOV+0g9U
u7U36iNasqBo3gW0uEo/T14F2ozoS4l0TkELoQ/1ED2ECVXnQCImzWYvZBf/G80n
SCCuUUwysLd9rFVHiIBu31Xl91c+bmxAC4uvdJe6gLhzgQNveRpoMVDZ4+8Rsc4A
LSrX/iAvzAv8OBSTeMISQ31JPzZyQWRWZrlSvFLYDJ+U4B7CpfYGG+GGQ4Z3xmG+
LYQCgKdhGkOE0c2EoMOFYqAanw1WzOpw4/Bof88uFUQDRxzin8rs/XWgHPlGne7J
dNkkthfEzMmIAR6sYoqSpQvL+bed27gqlnMD6JLv7e+x8hW238zb0BMbUbUowgGy
nLyLvcegDfMR6bvucW+K3xzIXAT3jfXNgIjVmKDKCtgm6PlBvaaxuKNLY/Y1bR3W
Y3mZAnYvAkZXhaX49P+UsQtqRDKBzHkYx/iVb0jaZ3pa0G+IEVDB++4Dy90hpIjq
rp+7sRRfRRQ7rO64/75kOFRn3OYsA0dhmyqQ9hOAkOcMlPsD8jLmYLOCq6J12Pob
mKg3rTcTU0OW0J/4/OS64Cr5QqBeKh3DfWO7f04CqN+xp3FycKmh8S2JVqhwBwzZ
qMEClNkqAOxIPv+PATAXSM7os5kZIhVYSgr+cRvKMjgFBPFEuwu0H29HlyybG5yo
rTaTtSHfUWyVe8JGxh+detbbljF2mcW5aANWF3+M6kz7ZZNdUI0cXIiza7NT3FlM
TrMvjsTC52BwyKbts2YD3DPSsx6jlFVNzRUCqUGwZ/K/5yrHPVqSYcUycLfAzJFD
MYcMN0xWVdl30H45Z9hpnCBRa95odrfHs7/WQhzub8FZ39UqnagqqzvXgpBu42AY
1z5asyQ0kWDuptFCk1mTkS2uS7BoL2c7ORW8faZKdL1WjKpzKD6QFFpX/IQYcQSU
cL/rxT267YbCpLIS9OoQvo5DaI7QSvApQjAXg41y9kcWRsjpYBbI0PddsOl2gELA
/VG3UmIOoc9XX4SBR/HnsyvWJfLWd5JBb4l4O5YBimXHvzjM0SQ9qwuLWw5/LktQ
aPDHmWrM6vjJa+DOW2pp81LPhUMkp67cSUQKjtJsvLm7LLzPo6kR5dYxWiIr7SHn
KveZhw3vQs4FLtqTHvP9SLgnZW9OqyNV1EyE3P8cjqhY2pnTA+ukJuyk0qEJFWGc
m2TyhgKVCW6l/1czcTmg8j2l16KgNcUuFY3cZP3/5IVH8morcvWiAm+3AYxMqJDF
jtmgviQMeuGsqB8xMA88SlFIPyKIXyEBAr/qBBthJ8qF94JnG6M1h5IJwMu8slW0
3/biZQ1oO1mnkdCr8B5c7GVBOFpYQuolXtNZ1c/lQwE6LcTLFSauWP6tDA4PTH4s
kSz4iB4ALIBAqH+WD1H+wgqO8qDdqJ/Jk7D5m/FtPe0QCoLD2n7DiCQCMz2Wxfh/
TZspPdHMvAygsEiufo+YMXASN75DE7J9OijD86aAx+OPWpG9KfSrUIDbw1ts2fSW
uzb8/q0FwOeAgxXiFk4fmuqwogyFxDdTFeGPP5xDXgBgtn6eYaf0IhwHsliT82Pa
/cgR+IljSrn/lD40br9VjZy7wbnN5YmayBlFSTT/tcKmuAAmr86AoUNpbW8gWZKZ
cj4fzjYKOnsMsCrX5EX/MVzJajp3dJ/+0kj3JfJHYDQlEHnXd7Q/+skoiqXqjYTN
lJKIHv4PR0pHFgOEnpACqeRggRzAs8e2GW9+ZauYQnV54J4vaoJuw+W+iX9D7OF0
i/f3ja1vDeMP8w+Rc/3+L/e3StrCLMVfX41MqiZ0N8zU5c/65+gYIiKSxsW/Uy97
Ng8I3Qq/9fT9g2SWi5mYXEQVRq82K6hGG/qik/eRE9D638lZACWTjDO3D/YTr26M
BEp0TqMYnyun3tE/a8O/hWMB+3M9o9f0bySsBSdCRR3XpOQjiH9LH87giN3forpT
9s6++vQB5Ujkw9Twp/AzKr8hEiUn2s/mvKDp5hkrHofJne8amyWkId1K0Bl1y2c/
zREd+gUyCkw/l6q91YfrSxYrwB3X5K/ert/3dG71GV7opvYNsEsYcE355oagF2eC
WwlndaYgYIE679O49p2zIu4UpA8qytcJkTpS44OQ8rMItVv0slKFg+81MOQb+adx
YYjHcbnWXiA0ZxAYIcjxchIGlT8E5CGptJNfAg6mFl/LDKn78+zsz7oZFOheLeao
en/J+Y6tN3QkC+l+KXHFrHKsZH7iWviLgEFLjfISqWWYfisJESObrJvTGt0hoywO
t7O+BQBNFArBcuRNmw7lmEb+G6iwZnP2bPW9J2obWTiryQB/6jFGitXvnNCTj9vV
jdU8VBJMG0K9flN5U7bQKYj+ucBz8wG1+M0BCt6pQqeKRAXqkael1BEyakVgdk1q
y/O0pvdNr3iFtdHolDv9tGfVLhd+lKUvjrmIVCtpXtXUBqYS2l4Z/OumHmLIN9hl
yKceN/PP6m+TmRueYEm7C0jd5KC66vlISm7OrPx9ta6zJhXs7tSOJRFODGNCEFqn
M3tdu+Nf2yOu7llF5K7WpwqskgBiyYygVez5BA+aATG+dpm8Ij2CIVY1PZBMUCc6
F1TnNx8WqJLISjoMMggHMTMbRtTdiBjuW/UhLr/QdQDkaYYGhX7Jik136ns/Zfuu
SvLWIRS3KGwbEka3htlJJe8iXKMItM566BtyfzhEjI7s5DBTOS5j2C8BaBoguWrY
ItEwep9x5XyuAqTltUrtTnBAZLuWLMoS0nRZ3FWYLJ6SrI5nqAuBtuQRUykHzgOM
s/+YyYmomqm1Nva0cxoUlBEyxVAQfwtRrGKARJ8AZyxTVp3p3BW7yA97/9OMKAfY
mr8FDHn1QuEfjcTx0PBl1+QBlGidfpDOIMU9W9XFRzH7tMo6em/OE3VDojfM//v3
b9iRr3OWT6V5GVfdRtyrWTehSEwRY47UAdwXVJD7R7W2RAAFCSNcLmREtdaitXkI
oHxAn3vTA1GHiofVn8phyYuRgCH/TTJRVNdH3LxcPBCDYGynsrLTMippy81vgVh0
lltO7MxwoWUoD2m79psE5Zji8kP87poKEtAPl7LIYE9AN6rK5f7svoSkg36MDB3V
qn56thbGLDTNz5GbPVxJvG0MKcojLCtP3kiAH31nlbXh0rd4sGnN5tk1QSZ8Rvns
GlWbFM0RAJE2LmlAXfvmGcVJda9UxNVnhjO09O2esk9AcqMMOuL7X4LC9pGaQebX
tvThLCHZvX+hHLKiZfcRTFng1rxJxM2ifGMkXvAxfgK/7ZnsHk7lqzDkXO8OS+O0
5IUq8divXIwXgMqRfXYe8pKaPtyqAos4PFvclCVUThUBsJEbVtKrIYx2BKqlHhMB
u2Kizlo7pb0BLkmS0Gzkl6GS+y+3Vrg3FneH9TlkbQGQAr2WwtHKyIRbTIP0E9gd
nAzy7W8Lqw8030CbS/e1tqGVkCubRvyYi5cE4/3bvV06toUAafkUtySgPlNJvNee
/bp8ejRTzSZ397kmd7a9H4QErlrO7iKPT2n0adjkG9vulVMdSjy/QJ9kxBYNoKEQ
a06fDWBEwvQdqx064KzN8+h4qSD85Id9t//vhfdjo2zO7DHT9ERvLe4qM6W/BjTe
Eaz6JYQYxAlkorCoVtCEzkva8r6HGx/6T/yZAtrPMOuv+D5d9degyigay2wPBCG6
t0J41TZM97PHPBgXFLx3+7ohUbyMy8ST43xCgtfdSM3M/5L2SYFtUOtiqZ9EAjrk
yNHqVcoP/agMPPNYW37NRW6Si/or/iwg1Ey9uzn+4q50QHYotBETp/DLxMfsh/2E
QCCJ5smyLvGRx2vllQZTcvzsmw1GVKeNCh0Q9Px8WeFFkYAWpe7TilEKnc2/hISt
G4AkbiDgzUDesq6K66OEVUgExc63K6+J5z1gnPfbFeL0zxV6kacYk/CEkjdqFh4N
QCFJKJL0AGzkg4sDNIg7hWV8sgZePiKvHD7OlZyqBHHENFN+BYEs4IOHYfV1yz7A
lXMWhbxFri+C92faaKg/apTwjHGfbdY8cglrddMG1kDRjr6E+Yh2HwNSyd6lU/wQ
6wGHMGul/Z5HH5dQQFUYEb5QubdX8N0Dn5UAJnauabVMiVlOUEzSr0Rn6DXaI2pJ
J3Zng9bDisu2ihpWNFQ3JkSf9wCfC0w7n5US4KB0Un7D4kcdRS73EyCwZCSr2/Yh
H0QcV7c9pG1Z9qXHIB7EHIeD0EDxhFmTDijd27tfDca18NNPZcCJOR8yGEAAzJW+
rG6hShtPapujq5HADXOvcYAGzaWBjukLUTe3tvPEXTqSHzyJQ2OQxcqvJX73khVf
BkJylSdE3I9KyokAC2bQp/hbjNPzkh0bYAndrrp2ZzOu20RIfQSgI3RBwxFUORKK
hdfd6rwhOO/ydAw0/bX0dmtDzsYHlvDD8zk2Lwip1fQExBSOp8P9hf0U3CE8filv
0Sf10y6NAqhzRAoCv6D4bU1r1epdqSrwl2B/GDtPkkXQ29YXSaLlUg0vA/zlRT7/
0oeJZkgVMP+qOPWhjvyC7nki/oAEucXHPKZM2Qtrj4EQJqr3k0V8H+zGKuAb6Ecg
LRJNgYKk6r+Lu4ArWHB1preh2mxVJ0Dpd1eeVRWy7uRCBZn/ChDr1corO6zNQwTI
U//TOokb4x9mPFNdLKROLVf9FQjWc2oLEwbs8pBRrC/MXTBh6YWsh6Hs3aqH66eb
cahmsZ8Yu2St+cU2l9B12r9PJjBw9WCTesdCPRfv40s0tMqbxzrBm1yYcVmMmEhu
sMmSCm780jjq/PEqyNJFe0kgyxNA0/K1XBF0G775UYLgmXwbW686dm0nIsH27Edi
/beDj4d0Ir6gTLGDB21CxOjU13vC4bobR1il+VS6O+iHIcM56B9Ddz/ykY7h9cbZ
BkGPiF7LykoqOIDFy+GeaFmnU85MtNqQy9XrxFkuI6ZJYKsouCX+23gewaaKQwyI
zSp48pY0n5DdoI3omxQm7CHO2jbmT/lsxN/zeuVj6t882jidJp8Yp5eHA930xu2N
1EH7k+9dCA5vODwQVgoP/Sm6y+UVXo2oeVPNeLUlXLHzlpAybR+v0sPkeurua1wo
xZBTtN9IPfp5ovFMm1/M4+Vu+84yxQqqeTcn1yQh2q7DCpoQSTGO8QJxzmdD63BP
IsZzUFGwY0Jr4ArO4MPLgfwB0U9hP/4FRKNhBp9olZe7uSbdlHVE5vgAqJEvpY3t
7PLbR/Bv7la9AdeBtO0n41jj0mMqzc3Fx4KTJEA92/Opjq44bPo35AXnroZZ7CDj
GcjDyVolUFoTnqdvUYb7D5prq0spSKSYh/vLjmE+iEG+EDm0jeungG4HGIUXO/ur
3M03f71zuzr0b/yLjfZxtu3r2E+BQfNM0r+686eIlTpH7tiYtEsNpZFaspnRxoeM
l//7eYfplkeGtj4JgVqcmh0EZSu+ug9Jq9fIUAPZzJiwHTSjshoMNKTst6/EBpfM
F2lZ8AoACPQNkT23I+29JK8o8viaPwY1PTS+oVJdZZazqCc4PuNhfGmJd+A9pCB9
HNWy8U7AVfOFvFlKGzWvDw5fEet3PWa8mzB06Zu/eUv5gu/e9JxTW6JkQMpSTYui
r8qlAAV9FnJ79EIO6ISH5hV6gY1ImDOuWvqy0fdAFQiXPgLbfmzfQ3szZcczTc8F
+gQLJqLXieQKHjvQk75dISGTZjUDccXgVoH5uxb9KRP+oplkEt+c/LVB1wuKqzN5
IoEAoTDbZ0IFc2vH9GZNt6UltEn53uqoShfo+alSJz+BjHARed016O14DOec0S2X
z2CPuAFUCtJTkEl/WIvICzL9z38lYUSCtPUsVVQFJ5Whw8BMbwM6+x7VE7OCTfjF
6qCBHpCrh89VxSEfLAn/7Cjn6IsnWOoC8nKT4yuFUBClxJtdgZ99gZZWrf+iFcLV
NVIuTb0hhOnXdeC3M5EOM/3nZClq6As89FbkTYdPsSMA6Y2cv5GPRJq26ECQcNLk
zkmmlW4DDbPUPRrqz3I1WHAoQc2imHIRwwdOW9E5RK4TstLV2uRp4kFzM60VSiCg
V3ekNzfAnSO96N+8Pds47tFXvVEsnZauj1UG5NiYNUkYYGWqyLN8SIF/611XcE7U
mMviXQmGhuYpGKNwj+4312+OaycoQC/m+YmPosoHJkUdWymekdYwMU7h+Xpn8+Ai
a+hAaj4pOkwiTFOyWXbAttXJ9LOJywMEbfdtAm/jbbeG+7fVyoQNn+bA8/TGbY/Y
lU2FSB4oOnhKz7xTBYLW7weq5J1m3GqGCRPXd1yiNcsrMaBmM8ssS/gLtULzuDkO
o3fITQVgm7jHHxQIWfQzz+aQtstEkTj3zynFWM25g1xKw6WSE9fHLOIDZ1t5Z8+3
cBIBEy/Mcydh0i6hy6MXJBkRnypuA9BpCeL7mSgfSIEp4r0Cr7U9B1Ex/XqzxdtQ
/vp8eBlCxW5QjOdJpFoS7r30EBPWef9muPxcGh78INsHNcdQEERzGYDmohDIYZjm
/R6PEb+HtATDC70wYT/muzxv0I+3iWoJn2lQ1hreTjEXKNASo85WzQZ30D9Q+9Ds
d33UhD4t9VKDfEm6cM1y3RwqpBELtwQ85rhvTqCjlViH5dc0DoXO71LAEf+xbpBz
acW9simUpBaG5aB9L9Qs0zvybw9Xdr64pX10s/2osnNRbnLNjYDJthFIwkGUtPJA
2D73l/hVl/344slwqZP/LGNqR0Q5SbFav/qOuAKVvNQj1tKKXuWpo4kleuemgD4s
wSRWRmQbhzLsx8qDgcZHJZfO8kKBF8jyPs9OxawokSN/QRycdb2YIkip7Xkcdk+U
ekg8o9mXgsTC/h25MAlqz9xbKazcjhgbLQQV7lA5xwc0VmhS36z2ZcSREoYUisFs
aj9ffXWPBGP1aaZVq0XUrAL38TvwWkkT/COYvBtYdH+N2QmfrgggCeswrsk8DY20
T1eixGXHdrDwsTLHhNQA1b2xGUNgaBVZuursjM2zRMseYbn+P2HIEn5PIAoZwXa0
vFi5/JfHTZin5co0aU4NJGMki2Uv6MsgCLlQ75r79sBkNC5kwn9mMAkJfJq/Toet
7Ui4VlJgvWOG7Nym4PqmFjdDShAsiWmZY2Yxp8PKn51Km38mG4w1QmIx6Dxn0o8w
SpDdvueecXn3aYaEIqNA74LGMGJJ+xq5XYYhKyV885ZR58yevuHDK9ij017v2hRg
KsLutSDElAlwIqD3yt9IeBApE97UEq9YxpwatcetLM40tOAXKVtUw8qD8OcpCXkp
p/JuYUIU6OcXm6KhVs+aM1zUH1Ia4jFe6p9w/+Q2f+R7DNxvbY//mZGy3LiTV4k5
7Aqta7Re5kW0BXcbgVLzls7RvTN+2BnNWG6BZ/W2M97YMuLZcR9MWnKU7mkdM+4I
7Aa5a+BcVatjYON6+zuNO+puU5Gcds4zyp0aI9Tf5Z19O3/6QRkKgycWWh1jjlla
WSZXcEziUA7Wg7VFm/WIth2LlePzOF0mrSNgThPat1ERZclX+TmcJI+qQqTyzBVe
I++bsXdHfRXqQzgFBeoTc8OZRN1G6becDsZN1hJC63WlVyCsSMQ089HJAg9cMNQu
b+plA+VUFG7lpTC6P6UxmVLO4mtjgLqxDz4dg/msW8lP8ROWZoi3RWRk5I/Hjyah
KBp+ovlB+iFm95Jxvfx/38Dj9s6YpFiAunC4/mdBZedZIpJCQO5e8Mq1xtyVWfZS
atALFamzHUI4G0ml46Ts1z1boZvlnQPKSSZCYi60DfyAZdFlcUw6R2Zk4ZZSxc5D
0Ry+p43G6qfw8LEhX81tFE0bl30pF0dawkQIabLsuLCtV7uEtJdCS+oQzjPWaV9+
QwpB+7cilAzsMwa2D+n+gPaOyyKR3u7juguApVOlEimf3nRnRV7hvj3Upk0Zg1+O
RItcyGAdiieRB2Qcrh2IFBVgIN+63eshlSUrv2jIQoZNOpZEdk9Rk/gXp6hg9hzN
TjlXtneqFEuHV9e+cXWsxNv3vR7HRCchRIVxn8cOVHQkdHUACYA7yY9JBxCh8ZOu
B7V3fDp5zFF2HvWfABwv2XNySSrklCXUA4x37mGAY4wyfKHE+a+Ik+wFRLKxG63A
Y+BFIiCa/DNctUN+0Ykwoj2r8PpCGCpFUDbxpuINeD6fWozs21oyMEGH+Mda48vU
TRsdjiKbaj3g2oDGKpLKrbhIldkGAFJsTILi35hQA3zYazB1bLf9Fmjjf/JPUkv6
IcwiUppsto8c6xr6hBuGsofLOPQS1R4b2LIe0koUgL+al2LvxU1/lTm2oI7MVp7c
4XSHMZTPjXKXecQtxJNB8lMdsngrwP0vGR+WqSyMjJtG1n/D5g0cZP23yLc5mhMr
Ce2Bh+JIviRCxCJvEPJu8o7Z78UVb7xot04L8eGX5p8GJK3Lshz6GkvpwaWxvUPa
DA8CGezoZrV8TpxJbgogfJMvwp+av3JYFLIe2Qz3pCZnL1W7rSw7i2VO5rzFL5+t
w5cgJOch1RH/CgXIj7d4Xue7w+rDETbIkACCEaXNIuwQI94trUNLWiRUMrvcKvs8
`pragma protect end_protected
