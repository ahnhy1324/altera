// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Ze5Q+BR9ChLoc5b3ooFOYIvj/OS3Sqc75EQ93a/76WwScZQ0WY2+VClDFFntOWlgKzwgJNrcrX9l
4uyeqAtPeqhg5vFg5oRzpW52KiyA5K4m5sSNY9ukCoJA1/uSlxCU6zYU7dhgbVb7WF9AtuVBlxNs
LlDQGAIXD708h2BjAJGKAIOG9tX4ijDrsz4iqFdTRdUBKuE6fLWjuVppBWNbDp5xCoz8ePm8cjAq
vhxx8sUmAp+oA52+z97gmzeTCfwRVVpy5B3AXHUDDpO0RmF1FUdYKSorJS687E3zm16HLqxgLoJK
DQlJSZOVldXpqg0YnCF6TPML2R8PwDyqgpJ84Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
AAIAQZTPR0c2MLBGwxOyDDkiPyz3eCYPfH991NPcVZ5qjNj5Y3pntk34Y2cGFtLWKDMMSGx/HEpo
ICfbh+tI439kCe8IO01yf4Sa8dX4fyKeYI4YYiktHpFuCWF4KaXR5/TIcfnEwl4iZU+Y+9V52mAU
UZ2m6JH8T+rZOz+yLH9LGY+oCDUoxD4dv7iq2OX4x89YBE0ifLkn7P2bNrlA9qEo6PJZGz49GJnL
caa4B6X/82OVzRA9TDnoDTYoWbkicTszc/yMoGyebAFRScX4ZVIRF68LhPF7uIQL9lpdkcn1KI+y
tjNaducjr2Q5+Fjbz7D645GdLkhKWOlBiYZo9yyYaRO3vorfVDAuhTgeDOI4R8uvIpHxVjoB9nwG
oYNjBVH6nsuYzV6ijhDXxMc+wJxCdROSD3ayXYSmNIZ293BtwhDdh57QhKIBAIeKTMDKs/nZc+lT
JpT1VIg6+UYc4lSGkM7O6h9T2RNNtOJWQLxJiDg5h9fdDmMlxuUctMJzXjA5xKMcJlp8EAjgonRx
yZxgu7lHJWAdNWTskr6ZxDLSVWzihgzQ5Haj29ej6PcTo336EFoTfaCiH4Pj2fS5AViNAklV1tF+
7f4uhR/ZtfMia2bHYnSsD9Sf+MMmenQRQ5iMsvE5fcU2y3q5O+xjAEgeYcdkwqzZfK8jRJgXpMuU
gBtyY+q1Ewos17Nt+tOlsdVXBVUm8tNLdX8A/fp6cqfZMsNcISbj+Gv68jCfg0iQAOTCBNU9umTs
bNZbKm1Fk+co6TW7CZ8GRMUbQrT+g7cz1Iz3ULMoIRMaugnYepG+cJbsBqsPLjCfAbcPsLaFchAQ
VhSnnJKptrcnPxhr7XQ34AEyNSr+ZIwSuKrOLt4DFY8BG4N09U5Ubom+EfhdSxJYpSHs7GWqqEhX
Pcw28hMU9SQbllMtg2VkBJ7cELBrZqy1Ph3od/rgHZ9o2eiOK0g+Yr039HVfzsFdJWGaI0VXa6Of
wTBLmfDkbi9IBimuLbWM1Lwb6wMnrQ0kFjpkkTaATbb/LLdLFOQjALlU7ZwyE2B87p7KjaqSzOkM
2SyM0IQVG1UEOakjs7dqzNMy+l2iNYcSIOdlCapTrUxuqhluw/jt6fenX1oREP1/vDoaObsrgRfA
e1LH2FqhUTwTBfcY4LBVdLtEDBALk1DOxWm8B+5z8qgyQcZA+4A/y/afZMYOmgY6InYIBn/ZaCsl
SkmckZShnSuXLTtdz7Ejq7/dQCmf3aYErOZ5L7X0ys2f+Yx4A7bygGd3EvDX9ZjP27/XtFN+FD6X
ui5q8YE8Pt37EvCsn2TduRI47iS/6a32B1TwweqfnOCIlyxlOgYwrOnwSudZ2smgGKlLxV9h33i3
Ksc2XXMOyRMz7L8El/dUY/xBwBbe9MwieIOmqANB2QLBgLQTcnUpYlIrBy5aITS0V1Pof2mJXo0R
AQnnof/oQ38KkKTF5hNgpuZ8/NbsdqK1Cu79j3rX7xxPWDP8C96K1IgWPbgsvjLRTTM/PHbdQLIW
/6O5WvL/Zj/9iqHAxE77NjKZPKd/0fF95beOd3DUIk+mKNzrwXOl8E2SFjixs/YeSl0wVSK0QD2R
1TbFAC195oBHWFAlMhSheORawGXptHkJJKyCSxkyQSlCgiwt7DuzR6Egq6OHMkkpkkFFZxH0Ze6q
IMrSDpt1g6GyqrgmoSWbmz+2NfGMCM6DU5ffEKL/Pn1rWM3LWlipE/RxVHyksJ1folmLGf/E1VVz
Y5Ze87lLGaIA/LJZsYIZXy1c0gHqnoiDBqGJrzt9Sbm1zsp+zxYxRokuF8bUozoiX6+ThZDxLPo6
jz4TLZYV/u1Lcq9Lww9rdtqPam0bdxUGa48tPAxNB8CJDN16/5DQqwTNNflQHtVWOF3FI6okFBJk
xoaHx4qxyQwOfgl3fEo3MY3h6oAivl/hQRbbswrpK6ydw96yXcwr+6XueRR0ywMYRToblIMNn6Rr
ZwY0Zljwiw5FBSgfYnJBcfaNAE9KmE4e0DtxlpJ1lScWbNZgJRTRFCtgltb+BYcxPDZXgS1zBu5t
VuIvkPYRN+bX47i6WfMzVsFHbfiG3aGkNzwr1C8KQVaZ8CBa1QtYrsJNSeCafP7oUjLQsp1K7b8/
JsLDLN2y5Tv8blJvn2I39G+xkTUwXotNYpNilewetYHTs3gAe8ExkLqQ/aBFQIjQSbEWjEZZAOqn
LRPBDpWFh3jOWYDWK/lSMPoCQ83Fvlvdi3D/Ob02VDwbZEWZjkpQxhjg3iLeBDU5T2YGHr7oYXyQ
PYvcCXvF+PEOOTFZaRAsU+OxU3AlwbXzncSSgfy0T/SNNPDVEhGZNONapuEFWXtHD4gsJ4vY/2k1
9ChU6pOg/eNnT4LQgE+kcjj+jU998o+p2Yv4iFGjHMOoh0NCj2E8GppTkXAitQLRXI4dCs+eH415
U/qMb2xeAl8mfupO4Gd8Lv1y0a1LRum5R4wDMeFJDGAbzXCo03BBk0tdojdmMySskZIQtUojjd1p
/J7EQHdpYlvmzVqwVYp3NLMzfdgoz+W7zm2VgEgTtYRoyRgpWNPJSzkpbngd4JODsgMkWZ2a20kL
45NpQOy3V/ez0ypB3+Bt6ZZlH8Yn4VnRdqFxGSjDP5YmeGwsVS5qX6mLIB4/enLpPXEXq9RnDd5N
zTuS/N/BLrtOHkhYD0tb+fzxvLSlcBPgeUp/T01wcIUeC6NNxPAbOD9qPIijk9HG4QMI0TTv3HFd
PeuQpHvYd33PDAR1ezmbA/stJzX1WIHmEesHT+6uBIWCsfemfP/gl/8/DCiTGVWJz2UXZzIE+SFa
i6H86BspvKy6R+O4DtxReie9UztI1kFjwazhRrfXD2rUfyO3aceisMocyyiJM+GZsgUmA9CQ7lNt
Pfez5oPzhkDMUOkBb9bwfmX0NFPysCVQ4sD6UJNLWNo1MfP4NxxVVQ7bESM0/4sY3JKAGDiEbfzn
u7dOcUek2naeK1AMWKeg8wzyKStB+sBlBQYnS9cWqX/R5MLi7I6tfO0rby0tIdsblN9zFC//Vsd0
lk9/Mj4uCtaAMpzyqtAsGQKEALxcVlMmgtgzXHud7blbi81WTJXUdoed7UP7B2/wYZx+Y5TdVBDl
NkEfkVVYDpGwNkXaqAXb7+Q964EHKm3aUKuWvDUQNAZajSjshtZHH5rX/NaXtLCqhYwjMu8hOSjN
DvQI2eqcBsQd0v8lG9J4STCRnGd8RNI0n262DMT/4JVQk4qvmBHLdJqMdzRPPIU2toFU5pl+EE5V
zmtbm+rZqIgVJDr/EqNPjLqsIqlt2J4eD2QAP7u70+28AIk4amv/BxxHG9EsIHAzHiZi2TgOQ4Nt
cXDpiu4h8uPB41Elxdxfl/CoCWH0RKJDDT3NKcRUyM1V9ZMiaW9uqfZMjU8TW6nKC7m8Ni9aWNQ8
fBgN5udkCoTAUfKshC59RhZ010CtkIDOj+Mg2jKBkk3oJ3d+5yrPdC7LrBkc+faVFdg72LYzf3O4
u9tH01WKDCSsSGBhfwDnEeWWaR54kMzN41JXYETM7gWR7PZsrDj2WBRBjOAAcDrrUWHV3Cq0edV0
6l/geNIuRlhzyHxoqpuFvmQki7JEEVcbG2OShGJDVsVi6x03u3XhBdcdGh4g3WkNQMSs8rPauMFu
xL31TiiqCweV+QpCuNMnMcRxvZmu+1tZl0NDNaZkR0bl+LyxLNyMtBc0JcGRHdA542qU/XEmusVA
pVLfEhJdP8GEmr8drNzr4b3hwGP338HcKnVDcQ1wXbIA7beDbDmTjr4n9bQmIlFfIt2CUOYpUX0k
0tROCNeyMaUiNOjYLjDguo1ss0sJPuo2g77uvlTY1kFoQc7Dkc7IeI1MRvO7F2HScmILKTKDEs8E
aqBRqeWLXCF1hia9IBUNwpZPC2qrIithvxyCVImPuZ4t/h92fWPyykQo04fGP4/RIhAT69mapokR
d9KxhiKnyVPm9LjY5srPu5d+bkxpsai21TIENryl880FU9AQvoNiogkiK/FcVUM82OeqCE+Bu9UX
8+dGGMVDd2BoiARcXmBrt8FX4EoFVLYkfFC9gGAZ/cr9++29Zrdy7ROs9X7ewfQFTPLPLlxdrszt
xerH+IZ9mGowPPLjEpbbj/eOIAc/qZvVz+CDhOhDHNcNgqVV9Fa0HEtsrGEWX/wwBkQS9Y/flxG5
+RwtDc+C8QWkXUJOz9m6qSMDvhPyPvveXbXuEEkqqRUjPZTcua03WyeaMfmjtkW1HU/YqwtR8CcJ
PLO4ou5HvbyncJa+XM0Y2loDBeIyJIXy0xhI0c2IHUR+ddYGpq3uWAFIyChM+ZeGDHOi7MNNMys1
tpUCFoAjjUu29kCNiHwgV9+1Mq6Mu+SXPcVuggy5sQ/cW39oNsD/Jrd2mIyEw2kKVHf7mhgMl0Jp
lpuC4M/wVq0pMMKD1k4qq+vic9plDQlvVHfuONb++kEavn6xJn7Q6rRXI+9AblIivV/j9WX27u9r
ZnghjYk/TN1d+FCz2QoHkP/txilYTlwcJ+OstKKZ6yo6qgRAte5hRZDOpMOf5XP7o/wWHz/doeHU
os+to/YirKArL+KAcs7PELqRkA99JXcOUzWi4ZNBAdVQauOeVvP7WJA/y0xywWMl9QUtxlGaejga
Lg70fuVzkeJnkpx18O3WMcetSm8EvVaOTOfnXelUAo5i1d5S2PIXpFm4893g8u235mKzWrJGK29k
o66czRVWPqNo1MnVZouY4dzsq/E3bYcnVriy/GWkCBUthFHYDJijrTT/NsGvVXHsmgIFWhk6F2h1
N59a56yY3EqgIXYApvq0/BKRJU2EA3//Gj51FUN4n/kJJI/B0Rs8l0QWsC6cfXo93XoK7QMDRaGd
n3SjQR+kKGMGL/jQz+mMBtkhqWfb/HOz3lLqmQPUw++6TcIeYGLZYXeu8H+5U34qbXGaWAGCSg39
rZACb1jtz6H5YxdbIWRSoDJKzI6ciDHr0rQ/4Icrd81DhOPLI7MTp2wnKPjyQWKPE56Xhctxs4In
8jOPndhPC084eGLy37EG+X4G/0LHg6UMFGhlGRV6ZkXXyk+Z55j4nTFtZwTDPI//VwPMtci3k6Qi
mJ1JhH7zDd7c6AHPHEOhDSaKQ9Rz5fJlQ6R78ht/thngBZrvG2k56+vwq+HNulk9lqEINUz9QRLa
920ILPlNGUqQSna5T0Dlc3wkdvyWVOsTPHengf4zOLAU8AT0ksqHyfl+xNnhSnALqtlBKOftpSO5
CNlxaE66D9bliXrU3acfvmNXK61Wq/ZWYXoGWo1d28Fi9lQXHDTNTVUKuFk7ZKMdBmoyRGXKxEBQ
FLEGQaJzQLPD4kIzkEFSwAk9Lwu1QBDZz8h/ZcQm4t0T39O9xayZmOmEf22J7zlE7+qhYKjjlY/Z
li08UJyWWe1OBisO5I+lZeJxdak8xr91p4CWPIrRC4bCk7z3gY7ArD1R+xjBfFpmL0zIyPw87fvp
UKZHpPXOMtrsRsbEz8egDY89eE0ffYJvSjswOEAKWHMLgjNNYQco5bC8Wf2jKAHUWnqfYaYfqmlT
7qDicdx58uFvJzTy8ilyk2QOV4ofAFAZBW9G+92uiXEXaSengfcD5TJi1fODAENRRaIhQiU2KKWX
HW/8CGZbjzVxEAkUYklLBDZtGqGCcgN6n7Q8UyLyqDwXC6Pb/pqonD7z1SD2RHzGU+QFuCWjrVQk
sjnQxngPpmviV9VVBepH/0tVkrQT3zFavuzdcazlnwQ5QO/Qx+5tCvP+fI4KmlxNcAU+S5oPcGov
ERemeKAy9OWXHt6OTdsSd98WAjPCZF9+EALncMJaYsKyv9cRrkYb8vWutLcFrTP0G2quNl5gWVfN
bj1XMMoQnL+FzcbolBl3RVihV4sJ6EwFPld9QDGkzAFw61aHA+w6m4VOXuDZRzMo8iHpqeEj0e9+
tW3Tv0lsT5e+b1QsCMxyTDSvc9A1CezrPbZdmnwcrK3ZOD3ZxTvXec+D/1sxfpKyAzh3r4n5u7Zw
li8qzseWiXtfC7Ud/HUDmEzHe9Pd54IWi6JTmepO2vm4nMLPq6qoO7UJuP5+bl+zzifQ3EA8tm3G
7i3nBn+kNqN2xsQy472+sSMGyxs2pNOSEJC+OGjfexXZweR+hABL/uGv9Tmhf83KsTnvkjvYEhwI
q5pcJkzNDzMVMOFBrafb/X4Gbg0/GrXy8Q4E2f59lmfGF3rgEpkyfbMWCDv1zO35z87j7Q9CEid+
GfVLznRy7SYg93itSRZCTvMravIvgjx51bLYInwO7gXWv5VhqW9kdldgB3C8VCKNAFJKjeWvw5kf
2E91dnLpwE4mwXeBLGORiB/GDIdWFdZpa+0Q86609lsIz88CVVXTk2YijPJ5XLaprN9L3QluRwL5
F7DpVClaGiZlxf11ttb8sZ3ZpmMC+f4DU4Oc7e7ae6a8N5kEbDVHGRf1+v0hrL4/7HEBIKV5deSO
xY1qulqJf9I/SijNVNiFtgepuZdVJO5hWKcPr/kfVMdZNgJY+P03l2O2LYNz8pLCQAdl6R1M3nqD
n1Ndf7/DSTaSDaQZ0dq2CzyCl72od/2yC5/aatkl4zBSAdRHEepe0YEPDAQq/6zZdTo8hE/Z6AaZ
KOlMe0bV3yfUlWP+gKhn/nK2Zf2Id30cAKVnlVQ4vl4FI/NSW/DL7mLHeKsM3qqQ5fHfvv43qFs8
HmZtw335EJESfF9EkSDlPgmtog3FtF5r0QrafmX8TcQoxh6s4XM1VFIAIqkuTTjkZ+DQJ1gdByGI
uBaqqG5X7cFe3TAe5oLUZ/6tTl4tuZAWPGApqrfwxkaRa4O7Ync68jiXDBa8YP9wJXE04AK0PA7+
GzdzWZ5uLWspa+lEgAB3OdLLVdheLs1PeSH1a87f+f+MmGDyBpFCkIY3/Ivthi7+06Y4T/ZHdMmK
H8x9qyWAMSrKhiqhmhcH+z3AkcWstjxNP2IOlYScNfrtYuE2vbZ7GwXVm3JbT5kb69yVAlq6iFqK
EowUzUzEpTO4KOkmtpQPiYTQJwguitwDQkV6/+Px4CoY46gXv+C8uokSIfZ1q+yqJnCpd9yNIpEx
VZgdf5g4ySve3i3cSn7dZEtArY7n2DGUm+JwpSVbzys3x+fagsXF/2mdUclx0/Yf3W6QXcn4+UnN
n7JnQozktcYnghLzOt1pXsjr8eqlyp7AAEWiAygbSsa0sccqV3dtwEF0XI+wN0ifdNTL5ZfcTYb2
CvTzDLI+QJVjjIP15pLP64TV21TmolDQwj/fGLfj9Ygf0qaZ+Z2KXJ/4VOF7ODcryqB3VhynPA+G
g5N2b9/cX656XoK9ddGlQyNKhxkc4H94+rcKyD4m0QBWZEbT8u3N0PS4EMuFQrlBy6qBMp1bA6CU
rpXlX/4P30/YbTAQPCd5vv3fhJYO8dsVrRSTy8Du1EYjsa0dfTf6+rdBuTG7Ul7A0+6XPL09sLla
feOIUUP8Er1Vfd/Lr8Qbj69CmjJRgiwzN7qnvPwn5TcIkyAyyP76Vk5apaeNTh976+5fQxAsr+iv
+ZzAIubFE3OES2LVTwin8GkwfxbQQ3LfwkRl4dmQMXlC5/q3xoLPVgRobSoSHTjpTkmIEYv2dFxC
vd/L9tBrBTkOJsMKLOYUqjaCZ9jJ/PrJAPV1p7vBrv3uya+2aH5stDhayXhzgUhRvin9qWzVFI+u
O41zx1X799DnbANGOE8wKDpez7PgHArqgSlTzn0MGUWEQNHg6gGM6MRXzs58vgJJ8P3tR+u+RR/q
vl4cs6Za+yia906oje31jzYInOpcTw34Iw8dGN12NL3od7S0Pa0a7iu7kiEhz1+xrpbygsjDfA84
ZFbrePB1Z+dxKoNBStPpktSZKuQTyandY7AI+3ORAtME/L1nQ/Be4gqtjcbGT79fxXSy/fydrs/f
M1uU23sqys/leQ3kDsFyFQMo8ThBpzZ9HgphTwp8xy+c2+hN2mM7NAfLTIdxHBJA/yylLA01j4r2
c/+qKQ4xuMYcF28T3rl9eMDGVYtMISho9JJEKD+s0rlNRSP7Oelqniu2vOKoU9YLv2SRg+2p1lDT
fPPYjOInklCNq2Zcy82Y2jofMqPPXQ2QzLjnwnnRPDMDytW8rZgkkJyJfH9Edz0zObAauYYhlzoi
u2Chtwd6yx1S5ruTkBfYRvJUch3/wOZ3jxmjp8uQ2uiVe8q8HlhirHj+5aboyNL4ybgrQTKGXhi0
DzhjWQauNYd/XVn6zk3/uCqPTQBqs9N+OZnoVJTMPR1JdLVmCez1qRMgvbu/pFYDqML2ycRLX1kW
Ufz2ym3+UEDLTpKyGEPYTXENu3HyhGz9qX8f10idtccbRzWxsj88YbiahllVqoRd6ZhHXX9HtRoL
kN0XmNowaE6hKtyshtbgM5yNQQ++HByOsPv/dZDepCmY7jE7e0sIfsS0FEILwS8F5XgOSFxW57of
CfMgTUYOAr8+WtYCmbjKebIigmt8gXdsXQL/WsMNE8zgG6P7t3lw3d0m0PYHb6YzHFyTMfz8u8lp
jf8+a98hnQqyKryUAQz7tUB+cElwDhQUVSHEcTh4BhKZ/0HrNUSlMxczWpWMfJ+oKNZ9IrJy6SLI
5Z/Eq6IHsw2X6NTdh0z9ya1tXbV/b4LHCOpC0P8PgejhDrrkCffMq/YCxlXXUpA/7Ak7RWhgUZFT
rCoz7Am20mOD6NaMC4psWkDcxGL5EhzByUK/MZmd6ItVfDFWTTlO/CGajn05zCfnf655GGyT8Ooz
ySxiDZweC/gD7ZJjKeifKB0MEDwaDsywQftvGR6keU6SeOqA+VKuyP6+4aWRyV0E0Cch24WTu3wN
fqwWb/R6CjB9aim8+NWsFA+I3Ygji9ZCuZSdkk6N4Qz7C0Yo0WN339OQE03POhhucrLXAoRA/ldl
1D5axzeeguGBr4PA9jgt1GssYklVZ2Wd7F2aKE14U7KKMxumgp/UtZs0NCbC1BOCyDYK6kgzt7g8
1Ro9GF4UHp6hm58qcf5icld2w0f3JRTWQGQ3SIIeCa+kcP3nvlRUk7q7ODhpftHR9I1fsvnvq4x6
2/Z80aEp+HbZHDx4JOoR9wMt39VbsSGUKl3aoIGXzag3R/zaRnlWDM2b2tSjF6YHVrjhoeaYmiKz
7+ahdMQnBJ+E+AI36wKBL7Z5IIvcLDw9eDgwPY2GszO6MNl3voG/1x6ROy3xpPWhQrdMclgsKblx
2eNnVFlLWvxwb4s12uHik3hRv1qjVwsgX4azl0+HivCdOMuFmfSMag/fY3O4CdZqDIIxAWgAYKl7
9ptKTo/7y6jy3zRZPCETHrOLUYaH+HVWE2vtcf/0aJtec82iFdKq90nuRTJg3ZRnHJUvTZ0+4Sie
kcQjL+7GhmDAPBkzDHodJvlsJLIii2Jnpy27OxQ5bq98owxWqOmk/0zGH3hMP608B0BK+4f4BL42
zGPPNkTpdhfSyCGkotVA5C2TpZqEekJf4i+O0Sn5qSRdeOhbOGnYsjOzD1pZAzCUy3Q+esQmolbJ
Pc9c9de3xohYNHsTEWwufLODR4VYNbFAUNjVkbaM6CfAWtf+sdSgON1gpvvQcetsWPPuB6Tqx4Fp
ok6BsDuzOHfI9bRi5iYV+3iDOVyEwsNyJ0sG6xoHXmCYAQYVZxCMtF/uRlLBr7T30ecu2psYc/Vs
4Q/tf/uTxol4SH3oki5HPu74IfTasMeWngS9S3itVIMwfBwJcpneFQwi/u1VR10LpvePDHXR7oVW
ZEGoHFxVcoviXFlF0uT9TzeO9cyTVJSkhv3p+ZXk55CWv/Dvt8CRLAe2A2uTla5OIer5COQ/cK+J
iz4dx1CBcAcXTMSuW+PRgZxTjVGFRuYxJH3dhxPHYY+rSO3AZUKuvBXl3LE1tYRHtZTfF9j8AIyd
5TER8KrD6d539444Nd8UzoTLU0V7O9dNma3KQqGcgA6kPUsCytkmnwKZZ+Sc3oymMxaQJtc/pTav
q1Dw7CkMujy+aG48RupCMP9BenaQJxQ5BUCp7DFbZmkB9SAg9YOyreYTBsvMHT5NLgDcdiwKhv5q
x4tzJIx21yYf9JUEP13htBSymRdXVUwYHFCEv8xUKZwzLlC+HLNZJIV4DdTH+tfzvpVUEeXtB5TS
pJ4SMG6gW636GHewVE/1GSUb/83wT4njbGiZK/ya/ObHb/YfygWfEqXZeu57fmM6bQIVeEqTHXmq
/192nh70ihpczQXOs4jkyc5pbwtkQzKQSzsd/YOewegx/UEDDMtkkTbna+MbtITZme/uxCRxKk4f
N60jLYy1DTvwIZYRjLhXM06oULfoliY54ya+1fSF6wJddjPdzSyerkCsJkVRxgnCjXSNzpW04EPG
Iiokr4WiDqTJS5fUj7P/DVScrQNOxi3NrJ65okjc7oAYRVeCVwxvBakBRYogg6TAninh78IA38Sf
hD7gAHDVy2BQNFzUxKBm5kglkZ0xJ3oV3mUZL61Mnie6LBfcftxTdT/EBLWBSkZ4zxD4L9S+8p9R
jNOmBMKb+aM5jk/pRQrpeDnGodth0TO/ghHt+2pv/kPVIFD76GAqu5qOGHMArxCnzkqdfiOQyR3i
V7iJ9q5ijlZaU0elxAyCrPHxNcYdHuUm0o8g26EY5TS/P3CDApzugV8ernRqhF4+ocGAOdU3z4mc
PtUz2zzm9JsnfIeIeDxyQGicQ/AScUVXpjiBkvLGTgZiB3QWPWrB3UkNdApUVt4+qFgADec1R5qg
BANgH9WfeMJTCsFpslTFGkO13PiyNYZsMIrPGr4p6hzZXYeTXX0yZHgrdIFCfB6WB0TupQqf3RBV
oaX6G969OPtGN5IV4L35qE+6GRjTbqiD3+o0G6dj8vZ1qZA35JyW8rYci+oEirRqHI5EgrJ5qfE9
J+Z1sIYGgdvIh/hWNN1/oV9NH0vp+6ewg9R7fKF5VDzvCcNdEqGY0WQOjxeBsPFJeqmrLIoMaN7o
qq3yq0rpZj3XHsRnSJjGLYcR3xr7aOUSLRNYlbDzcZ9sTvEZRAprgAXJjg0tvkUFfg1eROuIJ/dp
Vco/q6LM58swCmEXyXCoZPqKFl+Oi+q/verNCK7Hon1mspmGEkrSE7/3IbFInqM7JLJQ781xhx8o
Smtq6Pc1bsVu36M96JU=
`pragma protect end_protected
