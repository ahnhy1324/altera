// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:54 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Dx3+RSv9cSMa7S1Km+YP8sgmugnkU64JfFYUmyJ16+WDClV22aLuFWjxJxerr7qM
W8PmyqsosmjGfrxExYVAdGp39AhEBXMm+0MaYdD0HdxsaNKt2mMd4SwKBmvYWRL2
H4CapLLKB2HudRba8H90qW+Sqq2WIRWFtYL+OdOtj9k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4720)
Wu4eDRupy8kcjTFIv43f2XJUtgMZqKtp9am0CA04NL68H40OAKjH2yWNVd3T8NJo
MDjuevdpycQJRdEAdoAytpvD06SOY66IdSM77WHlNUiHEW01u26d0Yv1QoCClZtr
XOcUQo+aJREySs5WIyQ1DiXgtjWFt/MZRUln2Ns50xYQzU8lHcbWqdvFMBAcSNeI
OJTW9tBbOTgz1QvYrqr6TUfHFA9KNxq+cGOoCtxTwpaw1Y9sL69YHc1YES4RBNMJ
FPkNkWyHT+0Y7DS3SH4NsC3oCXvac5LYF88ZKeLK02L6mPIoFuF4X4QLS6rkhWug
y2Qh7BPY//lnHglN/sHvFzLHMv0TT5Gjlqu/zAtpFIylfv55DkDJf3hYJViUSjn7
T5vzS6kb7/53Xq4utP0okhq8j7dV7aUGR0ONB7n/IRwWKjX33a8beZ74quiaMTwt
4MXcAjpxo74vMfXoD9ckIfgG2C321IG6UjlBCak/ZFBRIOK3d/Ka/XVGJoLx56pu
pn5FtZkOqhqNS0k2AR4mKpnWzPcEiTOkHdgU4yvNhQwcYl6ea/Ui8KuMV8B+t/0s
zVBGUiqgANJA72OR9IUqXzjE9CcEeOIRl3Xf4Z4kmrphYOsL39Z9IxWJis3B0OeA
gHTQrBrrlynnDg1CNvDGRwrG4kTaPrnZpNketPkdj3GyZcne5qt3+4I+V6eI8orR
PeH8AaCtnGU8di7dGaukxzePcrcitsXChdPdlzsD3qu4d/jJoW4uc9fJMtVkqQq1
xSKeSznnTmDiPv8IPv/Z3weBGfvC6xRQa+yM9zeNgMJ5YRYzXJEEQOKzFYjSy3V4
lIt4QWW3ugjHSCEiDZ04LPGqDPH+UMxkDnCPho80JhNpzawYrDX0ryVPmTVVLoR8
cwixXGNGL8mwJvDkcazHUjuokqbu0DEpH1UmSdj7XKjz4T2aWib4q6d04Sxpz4Y/
/f4V9D6X1IRLKmJIYtnB7hNLifMJzaM/xJ/hm5pGajKSY0Vq7kydWp0gJ9sb1m44
8J1Tge+qbg8uRkOhm61YnUNmXHKGJ+d8EWkxlgGyzOFick+FBTQsxzWaNJ/n69xM
gQQkAneY8+uMHVeT5yKKCuKYz1YpD7mhksiezTit4iQxDBwnrCR9LJPzgK9FTaBc
NqUOhbXHxiHVcibCj2jz/F3JL1Vo0gaZYGSrp7ct6EO20CprEiZReitTHeEain0D
gURFMbYdhxTrcGosK5K6rq/jrnxiQQnptfycstf0EHhyUeqlxir3M0Ykluen4N2O
+6GkuzipE2pR2i5JB4AhfY3OTBt3QMgrTaVUZ1OpqxVKWXKEH1Vt4A17BeuP/c1h
aXNr8FCCagYwAMP+h6ixLAVVuWAm0P5T2HQ2yIRXN0wpXLQmWTitJi2+LAoY30wV
TLzBNCqg8G3misrrdjpKUsmN9OhtjRTKtZJVsTXZqWmPGjdfOlFZU1z0aKWKkKTL
JtumYUitkSxcF02HmcarGbgMuoDdq3KztgntjLc3yxi9wfpjwREqNTUU4gk82t9Y
qlWOZPOV+mgptYQRJMZUTv5si8lQuZOAs+eTVpV6dvwaauHnsUX4x92xBtOANsRg
5rNKOSz7yYqcgHV1Qw8IJQQcZ6Lr9BC/CTyO8PjUm6Psy7rTCl7JyN8Ds4wxtKuT
ZG3m9Xn3/h/IhjKGRhiOnpZn8i/e9HOYy1Jcru73/ER5OGZlE/WPzSXxP0FJ2rL9
+HIAe748uHgt9bEYQyyKR0MOy5yTwD3H7VWIrfiWgB+mpTkpLIgLw5phZUuKD+IA
BCPcTINaMlkB5jcxu2oRQPsu0hCG540flQ8/1DWMZDRM+Zyi1g3QUrwY853JEfYQ
JNevJtmjJ7C+C+4XVxgauEi4yRq1E7DV4l3aUy49a8yMzwGIXr+SExi6b3U90LoI
ARGS6QBTjzTsFEjTCXWbSHQ6qPTCgH+aU7DwcKhDBok48LY7z+dBzlXjnAiB+0hq
Cruhs9LVRjkrvBCofcGHOlQpgr6yVgJfZGIHme50LCJA2VzHUKX0QjfBdsuxMFsT
iDDJc1X7fzZut7pyJJ+fSiZUjCKEGoIZm3SENbysmsIYU7jdpM5aZ+E+tB/NKSAA
jXcIct+Sqv/XCNqDvu+gqSvrFg+68GTrPrasWSJkxsrq/km2u/u7x2kqFmrg5299
w1FlaUBAygMOiUSGk7HUoMjjCOePU4R2hlYZ0rbmUEGZJozHiAw/dD9YQk+lEyZ/
65uXTzDoVYSGey1CAXel09W+QRGtrlIX5+1OxfSLvyLNjfjhD5p8DwLg4FhvhEYq
PP17KOYXyiVJBsGVQUquwWZgzzwkyCkNHbZUlZwF5FGvAqSmxxQIl6RHkqXCwfOF
RjIXRipoNCI/dD36nbeDY6zMdD4F9bmjxjJmXeDkSNPGpVTG2FB8lK05y/p5eVXM
Sq12+IVcO8aYuOEAWNkqw9LT85SYZNl9JCL2qdYO2hCqHJTCpIST2DSZY4jyB79U
6A+VWwwEZg4XbczxyKUmWHmrtqbYjI/zwZk5BucYZCquhhIEXJ/OrS6jATstr8CH
AzSmWIw1d5VqHqhaTmY8nprK67rxNvegRnm24Us8H0HsrzhySfq2YrSLylwyVLIc
UCEfmloGSjJ0IGioV46nwtJpShusH+rACw6MpRzUanhwU9ebHHiXxG7tS3qITYDY
OVIEaFuH4HMux9XgHzfeiMFCguce8ZS5jHEQx1uuCeg8nTEsIyyTnSld25Fh5cky
USnZ/5QGtOIeY5mo1Ttdl/rtbG+6wuXT4Lv3LydMABcM+gDTKdhHBBZdqTZx/4NI
Lj/d6frbiPLH9jtbFFx2Ya3yv+EmtB3mieSKCpUY7xqHiHOaXzWwXmUcgh7/3x9x
XX35jL+xEQ/Ra70RkYi3eDVSz8tO6XEc/oewdMxARVWeGiUAps276SWIQaz6LKnv
DwkZK9U+dxRpE/LWhWjdGXaH6JTTcN5eBPUreZAAeieSywjEAFLz+ld3H1x5EHgo
irSGsX3L9iWHrxWRPSmswkXOao5uprKQw+Tbv6UGu4QOsequ5u/Z8QZ+mYVCKGft
oSksQkcHwF4OskwHkx/pB97pGTefX9fF0eo9LqZ+WJiDCm5Jg8eDswmG9fQa2soP
eKy+xog5xR2GhAQbVJ6odY+8iLoIL8EooL9mypxCi/x9X4POmV1Q7WizTlCgTjMS
kiIkCcwg32Q2F0SGUkXyH6M1PUls0d3huSd4PG00qbcoU/DwXDHss7EA1c4DtJIb
Rvz0gNGcq50HG2ayEeUTp7B8AQWxJU8ObxGQcFFTWcuSpFseLBprUvyJLvBZ1eLW
YZlBeT1elWUGjKDKFB5ZzXlcp+jdDfgZKt8ByLb5oNUu3cQwWHVTy/fJsnUR2xWS
e8MhKkK+O3iTM6NaNP/In9RiK6ABXjZmxPU4Yydb8TgY171Zo2n6grXlZf2xRKAr
3iAZuN448+Y5KU4zWY88qPNxH5K9rQYZMX7N06Y7nEHGgZLi3bsU1ADxt/X8OX2g
zcL2KFgALSw96U9W9L5vuEy51j8UrKaYCRjjibbL2MnV7c/LAkPjn8C687skMiES
THjBMZjDEvqa92rfNdFjTZ3xDKRDKWyp8xgy0RIZWN2AyL5mun29OT+wVV4l2XUH
ws2eQGL6nKG5R50tRLw4FlGiPyyKOxUCT4nBJoj4thnAlaCjiipJBIPsyV+2+6wf
xX3gL7D5QRwk163U5Visy44yFzx2+4+W6JXHH6HTk3+qOJkkMo9pWe3cAMWCbt15
W5p8KJYE297131fBhqvIeIZif0Pgr1/enFHmPMsiVzrUXyp4sDAC5cMSHtP/qrRS
+XqQPdjwLW/qsamcU48MR1lWj6MWVGikrH7TKtURUIFQqmCFi6mMyJayrjtG//VG
RfUgIVEsV22DXy1L5p3R1xRz19fGsc9n2o86TccxdMu3aPTSEiT41srq5QfO3Mfk
Uw3buNryjS5gYBbCc0vVXjsiinL1c0QB25zVUxJRGZ3N8PmUKrpdemVKRTzBmpIB
tF8fv13WC64YVRoBQ/UK3ojYs94s4MNrVRYflG+lHo6wAl9HjyQLymV21VzA2kFW
zYruftJxZbUlXAAHatuCsOt2AAyekgMt1z3hwQQEE48LFSz097jnFdA4JkbFAn7X
iIOqDYW9yk0cLBKQ0mUR4KoPUUv9fRPajxMvkimh8VadouqeSqdOQs3uTeq5Dh1h
79BBNrBD8rlVu7ap3b73KbwCvVPhsL9X68MU3y1hjzkK2IiSBuueETg59gC4uDl0
dAml1I/YgYrAWyskQzPvX/mlCcZk4GzxQ+sa+1Oxa950IzisotIaupDnkTHlUNaC
poBmgYr8KTw5fcpWP90gZ9TeUFETeqOHV12W5XmkeGNsSJ0Jq9yKAO7bTcIiuQjv
WqNBl5/jGc/abaya2eHDLztwNLTHvuHP4Sc/9xQw9OhKR0f+kqnjW9g9Cp5cI2un
TjCylTV4X7WPu+zBYei3y0qnO3k8qdY2acwAtQIGpi3Ah890h4m7BusDI4TiAYM9
m2OyYU3y4x2q3/6UqIsHOxN5JaX6ubzfE1uSkO+F+occuQKimefiKsWjQsPr1TOl
GTDLlDW7PVe5mlQBjILRwYGjqomucnoJHLiufmsPWKZPV7T5oxJmFcgvgkKB/DJ7
Uf0dx+xkvEPSWPSdnmsbNrXniKIJBQ7nGNglpAUdDm3EPus3ZB+MiFLgzlyzr1kc
7239GZgORJu/9j+gmcYzldQ95QwhsKrdA7YUr89X8arR+idTxxrwCVQ7iJchSGNH
FpywcjKi6ZN5ZdVVA2z20pqSr//Xzyh7AKh00CzBdjrCURxAGGQPdKtDg4MToryn
bq4dKZemGIt3Gt3XHJ1RrCdoWZSZGfvrpZIQJ6oKhXXrnGy/Z2+uQ+ka2TuYHAMf
3e1+H6vO4EOmwlKFszNovSkLK2Ug1y+XaYq2yjzHGir7XM3B8kUk6SQ3GWeyFtc5
LgyrFNn+FWzLRHgUA9jESqdSiyrsOIIMs0HlVPU8mTnxzqpTgiIr1qMxQEZPMh34
awnPM6mnIrffmmgTKt2B37KT2NmL7HKZ+IeEJpNgy1NBr07H5/yLEnxUulysh79T
72ap7y3Bx6Kt6gnurs4CBhTF4n/3SGUW2KX2+dCBmJrlCqty3FpkmVrB2FINiVs+
xy6Ml8ubENBWITQk+mdJeQFP7OYcsvpoEbsgDo53stNE7vheRFOqXSbWhQxYlcVI
VD9a701gu7FTRiJEWG2J+dfDE0u1h6zzkGc/B8b8/GkxLkHPuzhm8H91Onxw+2LD
UAPlc3nkviomA2VcR/wTn/el6gHmvEOupfTVzJ6B7v1KsmRKyvJdLDQbTmdfLcLq
KrxJNkPTqXfWp4hOfzZblPXi3d/Jgv1yW77Y47yNIaTL2U+FBJaN9kWTxHcAG+1K
50PuUotbynvkEq2IcVXfsXVp17oS1/kwdXuAhH9yhkzyGtUVQMbRQnJDJ/CvUBtn
F4N5q+yirRKwrIibqXLa5VaGk70Vd76JYo1KWsRr5xGAMA4vtyJc/GMWvCmXbPRJ
roY9hGHuMGehljZkOLH0ZypU7WZBJEVX4zzIJDvWdkMsYYvhfxF/AgyETsoqvMEU
4e6AuV6sVTJngHg+4AsfBPQimFgVve+07aC2f/rxc7Ka91ZveRF9cXX17u9dbrOP
UfJMj5e7BmPGwS6g4z7WRO0XlNPOHz3q9LZFp38puMN9/hhkTnQLeL2AfPnwff1Z
dIG1D2qJt4EMBrImlcSBXdzURWpOZtCOK6YjtG9oohM7iSncT3WGUZlaAtFJAA2l
m7vxWrdqyNvZ9A5qHo53GYNKWkSp1IK8i2MQNMbOSxBPsLHeliQPdLi66aNu6IM5
sQHuk5BiwpCBCo1myJpLSoBAVPpsXlZZLXGdR2rpV4wBmXqOqKHvNSgB78BjArI8
/sLZ82MchnL2M+QmqF0Ww1qNrdoPyddaVZUmwrOPXwYuBqo0ZrQMk7qXis8B+phQ
ItMJK6FuCLKzG4R9TP1goTcNV89mwiqHPA0PEONOg5FW1thEqE5fhQGWRyFAUiSK
YB05bLZMc5OUptGbftdQV7rkvNYKDlzpISyITT1isKRKsnIYm7dUPRPBdAiARfXq
VxFgsEcP9FM8ccePk1ckvUDvZtoPz7aFmeAslgMbl6KmT1lDyNWqCdiqeYaeD0CT
qQvyoKhrEYZX4/bbirq93U4fGkbzqLUCODzYX5WkyTjN4aXz9WCt/a6N3cwwEi3B
bC/9fnmsuWlM4cJFM6jETA==
`pragma protect end_protected
