// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oGtA08SLVbqYszUlm8EHxzlJfQ01OcdfuZV8bAqHu2NQID3JZJwDH3kWuCU4w0W3
QAx7armeppb93p6NtzEOO+TVe2zUGqw2Zr3jfUMyGEsKxHOjbqMPEm5rqOmDBOMJ
RbsVB6HsNEa4uk0DRnOZYSKs8m+0wovujgSEEEmJ2WU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 86208)
i5MwqFoVnmSteSO6jO4dA1iVSogYx2xu1VP4RgmhmtjSmzMFZ7VoITwDSyM5U2hk
uo1X+UXHjCIEUsJlAIWy9E+5KF1uCAIrOoDpvnoXzvQpJEtnA+uFZMMYmFrCH2SW
g3HchaRe/vRb/I4n6F0h1HaX2whsRBJrGKwq0sk9g1EVwotRy9hiUY9IF5paUCRD
XdvamO9ZElwJRr8bzihm8kqa7S6gcaqlb11BfJHraeKbz7ZZTdACpCfWSbdoxUFh
/Gmfiac4ncAxoXtVTBP2PkTGzO5xigwumhs54GrNelXpwa6bWHt94XjdDg1gONv9
Tzo+EhjpAvqyjXl6X2PSuO1YXBDts5VcfFtvqnwvXIPFTO9/+tCYWhyLxsKN+0Cc
+Ivb9JqtV1nojhcpH5C/rswnG1/n2zliOHr4jJOTQY7TrRkAg3QzwLFAMUTE7Pnl
wsK+ZEc+oiZqf5Hf5mqTSWRN2+/yj6G8RKiCmCtqD7l+0MDuoF1WczEBGFmdXbKU
HADQ2NZQtqC7WYZwhXbOAbEQqiJ05LTvoQQaewns6/AFnHOyKrilsyy+hPeHpZZ9
OPNEz56ixAVRQKoS4cct7VPWADCc1hfybQS1LDvNt73o7ZsM42QwAVhL2L12P907
sYh9JFOn4iS9v3aifoJe+hff+PQLcwHsZunRCuE1pSnU8Ps07A0EC48MnxL2k7Q4
ugqIQCXZ1VN3aOUHur2loRzDGLBZqTe0wEz4tskB+IDZK37yw32MWHHKR8FTu0/2
PQ10YX7Afgkp+DZiU9I+grEaHlPZ75cJH15xN91no6g2/Yj4e2AVizfGHVnplUUB
l7aMfoQBG1NAV6rEqQrK/mis/cQ0eG6w3MTJdrXe4Eox6w9/KBqaidFqXqINed8I
hg02Rp7YTkl1BPrgSMrvd+pI9N2Au4OCykfPlVemJ3npEGXDLfJW02H38wRoFgiy
pRDo5/zhtslbigx8/mpVhGRZ3B5lUF2jij7eOWzeKyGNwp4y2PMU2DZ8uuqEG6iN
utGD851OMhXR4tbzcpFqNCGn2vN1Td+ZscWNKGM9lcJssN6Bg/KCdKcooQjqAKiF
CY+vNPosYDbjQLZKReX+krqzq5Pixqv9z1484nOZw2wWcro9lRtbvWgIpMmeNE0I
NXjYN4x8qPPAlmaJQ1uxSJ9NFIvwu7+aYm1VdQudkXqgVUpxNawL1A/MqhQRky8Y
uXKI4nAf5Nilz4nQj6ldBqdhecrOuRmMomwyO8EvyOUKpOG+gzRD10zDYbovTZof
/rLvuUhZBTnODSNZU3HtF4AcxmeAwQ1Rec2cSyCzDBmDpA2QVX9ItH9AVDTIKLDX
BFEp5q++zZfrPZz2ug6NAn0lvJZkMg4/dokhVWac++tLHbCWS406spniUY/hN1VL
P5a1dWuEkDgbA4l72P0jQXRJq8kTBGDXCIXNCmrzQm+hp6SfPgnes4CO9dMkxhwN
EHWxsOzUbloVqHuxvQsz0BN4YUloYLPX0R/R3p8n8dk9PTc0VGSKsl7dnGGTCOY1
sQVokTKWew1obncb3gGYzV1YyD7O8NW7ISXz6LMVK203yIvohRRt689mNXg7Gg6G
OmUtNzHo0FkdON3jpWJxB3BEe8j+iLgq5J6RJmLUVbdyyKjGWW/ihnrreijoC/8G
BeCxGcIKJ07+MXLXlINYmsNsRhiKGRTzFsGK0C8PRfg7KMrMf5ZXwaDIpJnilbsH
J2CZY+VkpxqXLQSJyImLTZgngrF1nKonlz9GSBld39WDBPY0MDtADu8zqUT4j2AB
taNwHaag4s/lUG2cwUfmHcg3RftJHkch3yPijqsQPgfUKM7a3Donj0eC/+TaHl6m
l9JhImEVuAb3KpG6uIRjWnxFWPVm9imqev0BgzGbqV/kaKz0g2VDKro+3lssRtWi
TvdARtKGX/fcN8loDiJGZdzFqMN1KPzk3NPqhF5LOTgC9XlCxZXlN5xg2aRozT2X
d++JF7sG11hUMGoA9xKKnWKzzrf79bWb4p2CyUAeNUFvIvs9LsVrU6GpzxRjX+fk
Dm7sra3frZTJNxRt7TJKUexgkQdp0Jj8KbhhuwVAgpdSjI07+lXpZmFKxmSWFwHh
0cEVmsGzKMmSMZUrsRO1ZO4KCKY3n1zn9t6jLaXN7yWVmWfdLoQaGsRZPZox7YeF
m5HFKSD6erMQTFEy4VKjSY7wkS4fKBKI84tl4w7CMS794jBSwrJtvbP5d5QC5qFa
Z8rLsDTt7lhuJnc3Y0Bzfbn1tf7CeUfCQxQ+pafcl3CJDZ809ZkVN9H2QiyJa3P8
rmRYVgRXtRE+0F0eKzFOLk62FIdsrCXEbZZwIGL4I1qkFvLsK8A5AoEkOHrzPZYJ
7HJfvhOKLOpJC011fb0HmXia1vq+QJRfuZR+kEGnVi/XGvdNX6c/yF3Zq2BHThym
d76YJY5yFmJDwVPqcoEGI9xX/QdGYkzSdfn/nNXjsrI742aRPGnbdO9hCoPL5AAO
GJozhT/E+eumzSqeQ9czkXX0HQvnz6/VENpH5Iwvp4E1Gx+0BLgVC6HKl3E9oQ9V
B/xqSYB8RH9uUyERU8wfPw3AdW6ItNi0fk92qZ6xCVNjVHy4mH1zBGonmv3HBrf4
e3pzuqpu1Jh1OKWoCNnshMweZcNtF+D8vMvFGxMpnOEwL/y5mhR6AAVTDl0Ok7w9
1rLQvVkKxIH6x00U+wr1+iZ2WFn4i3pVsXA8qr38sE5qxKaIoYoNLDgGeHiGAb2W
jSJYzT0XUwTfnTZIgeUAeOyvPfKTsGyNkgnb/0Ahip1MaGsEziGsOiq8EkY8amCF
YXaSSsXqZF2FriQ+RtcyUOLsTmnG3kgMkOSF1qyC1Ooku3+agzDVxB+wfzRgMDrA
oo91cT7H1cJuhmnspGUM3kBy8N5pZOG6rTypfQDOK1vuCMKLcLf4dWzCE+PTLzTN
/vTnuIVx1EJq6vo7UQyFLmTEV+E1Q+49BFH7Z2Th8f0H17AErPs77J7i27rZKRnn
ikkzMMbgZ5FAHJHNLoD3/kcNhnniudSISM7jEhV2Pn+6JymhLlajZZuWKnnkZOKN
wCmbLYteoijVwq8/K474cqPIGM4Y4W+l0oHCd7Hxe3ZGHwE2a4TqrUV/jB1HhocI
bebHwIugNLzdSs6eHS2btUPcmseY5M9vk75JDvR4GqAHFIPJrRfH/Za2cHXHvzRE
lCPOe52cU5x28PJkE+PvUqLYjeu2/vA7psxCIIHjK6cGpmevAFekwikiG1GxmqPv
SmHOzGId8DcWxeVX19TcTCvCc1yqr36TvLImfreRlCb4DvufGz2kRsvJaduo6pUu
KBRdee0rvV8HREZyT6d98phKn4rgc9We5DjfFZjtfAmq5mWHrRTJFqRqiLXe5GFM
UAE7t1S7g8VmuLdzlIWfCsa+ksk8a6qMoKpD0WLeF93uSXPUb4wNrRdij2AYQZwa
MXe5ztUQohR7XGF53X/TtGwUVs+zen9URDsrdpkQQlwuhrshfy/T+xBdZWeERHM8
uI144xNX44RW4yFgDXUVkT+8hG4rwua8Bt7uWV/YJTGK41p3Q2Dt/1UIYAcjofBO
FKRsEzDCveyt/fPUNmGVT0pcDIilD1eaugnVWW7StDn5jFOq2eajBfbLcHyO2ljz
YgduMfJCg0G0HgwzUzyYj8/h7ih2msecrQalt5ILI6nTGmBHQB+VAcLuk307vkLq
e8Uwdh0G3KKPqhHsf7j+iR+vn1799n6sbf/WDYSesRjszuYSGf5lFmJF0pF4QXjb
RD87p0poLem432hLaM9YuL5RaQvZjcpMwiEurOj3F5Z4+Nr1CR13euNzuv+BzX8y
a4Tj0ao38ni6Y5ZorDpEY2yj9lot1XKxzBFclmYyrlpVXIbAIh6Q94T9SuK3iCuN
gZ9AyFPRjAGq0huJ8RGv/KYBAui3TC8b/icS/515co8NTyrghw5OlGn+ZSVSxXMM
g38idUq26myEj9HUx79hLQi3IwCrfLsDJE1F4tMKPvwdExMHEqShXcIU4DxJQkaA
KxOh2xfZtGh0UxnsAflokTaQXn2YRE2XSFE050bK/n7lDfD2ePsIJrdG0KxEJHIf
zfApxC3V1IgeWAm2xRWMBZNTpb03SyjY8Tx16MA6GTfYfe1Pe3/B8qEMZnjvyX3y
9FNJN95Gl588YuvJ01Zo0hdGV+TZbMUk5iKsSNJdGUNNZpDMAR/kn0gwMBPf0RoV
Kqa17F+Sy6j8m1x7MHK/0PgqPX0y9aAVMlsv9YeYFPzaw+kHu90sbk1BjpH1AWAw
aMEnt4hf2u1lKkrFuHipxkDFWY7Bzdul4aWEjuH9QT+lNid0VQOqmwAwcaR0IEdd
vg/eLa6pOCT6CgnzbW+FwIpFKjlgXKCrsihyZBCMX1hc7fLmRpu3EVMWZPVLJ86y
zrl24DTh6yCfk0cyY+pcnHN0vqldZ3TfwzG5f4L1XiN0i4zhu2mIAwml4Ce5g1jg
05EHIrb5XWVXQMcLpJolSyOjFwA+a+LAI2SbKcH8RBg72AfS0bG0I7w6ETsO77Cz
eGSFINZtd74HYG0E71LOn3MWQowj0aoV15sSrOklArDBXe3YDfUqMjE4PDSriRb7
fFw8kV9wdhWKsVZJZyMpS/e31DczWFCjsQu9y5AnU5Er7t3WdvwK8j8zZY6Is/6K
rEbaeaXbpCLFlDkQw+Bz1oQsahIACWss4L5DUlLO5Y0+ogb7+MGcI9MIpEn8GSwV
++Jh9jtY169iNQnh7ig0Ce2Oc7BqKNR8S0fZ0lNkLphoR/4a7BxqChqwyqnwRsao
4GM772uoqU2Ievo4JYjEyKuQ/u1/eGUnwia7qaggx7ljP9+Fu7wjBRsLY+/hbGz3
MEFFCgqdW1CYiVtNqZ6SRlIdB3QCe2Y8vM7UeEDVjlOVTwhmqNaKLQC3Om5qzG1Q
sv0roEdpSua+foKHWrSKkQZFYqqO3LZ/VY9guz/PZvGZGii8e0iN+lIta/uti1V2
BoNRMPmdRS+SMznHQVXl4E/nkCoyMfhSrduDOmwvilnycDA+d0ecsXOTg1ted4q9
5yZElqMEQ9iY1ljkMFgAlT6cP4NamrXQcrjX/u/Vp91bovsWlPpPWafhryIGnX2Z
kMaCLsoOynJGPFJYabHD0bUYU0oMfmXdfeuhkZRrSOm5oZ+Q+wHC64KxhMMro5kE
52CsNDPzR4lphEgLUJcdsPI8khriJEyk/J/RqynlV2CotA7EaK7fYiotCgZPICBy
T/5c3hSkYwQ8n0i+4AUR+9uidOks799+gG6I5AOHIi/2FQMZvKdu5Dupr8LrPCjH
+mSoZvnGISzuNMVX7un/KmxtBWbpstr87XlH7IRFsahWGFkAeZESZLZU+IKWrIC0
g1TQN3bOHmbqmC7t2cDAbNYjx5yUY6SqRD1SobJNJY/lLxeUZsPKP2owws48I4k+
elf45gorMdi8dPCmarHWx3lOWxagIo1f0a7oBiCPRxV00qcIz5VKFTANlLeRWPTZ
vk4z9YWU4oUc1J5G3FUdLQsllgUjbe4bCNfAdePls1xEE+vbg6FySpb2HkNil5pX
ddd6XumBOtsfx1yhOqWsypGR1ztcLlTYvHOQha1ZOUsYDWsGzb/Hc4y+5lsfhPWp
w76jVw1vsQqOUcRjJkwaLRQBLJBaEi0D8j3qL29Zufl86ZYLwGGgREzaX/mmD4ho
wl0zXtSUSHAO18dkcNhXP0r2EgqzUGrwwQqFuuFKhkvuY9f4hQ7SD5Y+lgo1NhxC
87O0GhlV42m/E7+YKi5XQ0UANLoA4Fkv8jhW9TkSiteypakrzwP8wtWieMc5eTE/
kjorTdTShayL0e6dPYzokJA399R2SEL3MClIrmQKNO5Fu3O+eUCfxAOPESjBbdx3
/friXMc8dOR5ipIQmWEE3Cwb7qlD3p2Rfi7C5WBdWilUl+6HRXyodL8pp/CEp4T9
fCmcjrWB8F8jrnN5Q/ZqTtQpwjek3ji/VJb0q6U1cvJTgaWNLnMp/TjLXoWaNZ2D
FuvXVj4s0rNIan3XftGaBYTpp/IQc6O/Y9uilswkntibUMIueLBpt7VSykCAIJI/
LmwSXDXYEstTxRLjO/SwLDpOKWcwKigWMixB3ouQnm2vsD18F1ZulxwBpPzP65se
Y+xlkvlUBCBAcb7rqD9awEqgWPKSVUXay629qM7QkImtg8KHpXk7IETL0b9p0I4i
cQSNJJqRRcL5OBnBJE8S88im8qh3p5RzLbGUL1e95HAIzm4GCxey20/pOXWP9R9+
iYJOpeM2Uxa3zFsOiYinQMIUmB4GK62E9NZ1IJMlrmPI32RWHWY58amz6B23qyl7
diqWwJzzQaU/q7xfl+cvFlGT1mn+P8z5ZPuStAXMUpWo5TFk1H2l0vxMwQNec7Z3
QgqD6jdMI/vBtcDGZe+0SXC6HPShGuzfEamMIQYM3Z3dOXff7XCCpLAlIeyyajXt
eH0GbYOKfZFI61p8JRD9SiaTS3WQWVcwPjptpHhMvv39I5jFMV//FLBh9CA+Chjz
vDNta1UhTwZYnxewEPLSh+hrtW11CBf9sFUnrtBtW5YyG4vL790Q6ioZ4l47eLNM
7aWUSFGsv0mRMn5IyhjauVEhYn4f13WpWFx6059YVKpebo4SFgt8KQbLIvJjaElg
BeJInVzONrK4XVDsmBVMmhw1eP2XX/OJy9+n9rR5R92K1oTyAvyYu3GT+yjcu6jb
goLIemHd19v87PD0yf1f3dzY5TCWZtXSF5jjUvG4DPMnIP9CRwALYlyJufMrtJ5u
+H29QVsPRte5T9xDjKzZoeQ0PS5RyJh08U+Ua6EZtffs+cU6cFcfPLPUA31ogbR9
/O/KMzV6r1XNRJlVFoKJ2D17HtAzmI9CqKq/s/f5kyegyh1Bl9dOBvBrS/fH2P+y
c/xMFbZ1AcK4VeD5BBR6HkVYA3wxA9rWwQE6cfxGlLC2WtZuVIkHz2Y1XCnyJGvC
0ghNo2nR0tyA2gvRGcHGpjG9hmtaObphMsLm1X10N/e9G+zBzGfR3zALpY+a8fAW
HZuGUXlG9KdYXYtFWBBhpOSBW5XtAywrIfyj8Eomh+b4+QVbsFmx4OWAxy6MvEnu
MkEhtnIcDq3LOPZsTE/Hp6rQGNvb8nZt2SaZLm/I6TnsnbLlWK28Y7mO6PFRQ4BP
htRhdpOsdy2hU2Jl1VO5GCuJ0ZpN9Y82xSYd8BQXg8WjzaLFgyuigqxyIkkL1nYW
jQ3S0AqN6ba8rjOj6AIFMupxM+d1S6Ut8JlVa2/g8p0PRyJ2H5pGls3pl/rRJNXd
IOhy1fIGTBaOLSO3WYSQYs/6qs1Spke4dZzKQl7Be0bIsSAI6CRgzdcjTYbGN2mJ
8Ggx9/5ZgUB2ajiGrLTv+OKLAh6Sv9f+WR8A+xGYlm7OM8WY8nrJR1DEQ7SV5Gjr
Yf/gI9MYiMUgVNX/Jk3nqx4M308FiRjYCMlQF/4bB5SDE/hZG/WM2a749s/xoM6q
9JUBsGyR+JxNYwzlMnxXF+31FoTO13VfYdJWZzCCCv6HGXjvGXiaz5gxYpVIiypC
ACyDF9np3D1GPVJ9eUxZr03k7GrzjqiitxisqtiTM0ytSts/Qp+FBTlmnj79w5wd
eBnA9W+Xe80OcLUlPMrwS6atLrTb2D5E1TJQpeTo9i8E6NeeTtQ/AEChnqWEhzeh
2iQU0A/NP9crT6kOJZIFDTtnuh6A2SG+X1Ny1lGMdy9Q19i9afji11ER5FEflznb
5Pc0W3uIGXCJuyCOJi9HAA+9MAkqczJ/vwyDrCtDosPcnpTnCjVlQusIGYQUDbey
+l99PobLPoq36OyKjhwmBQ1Fs3uM6qwiN22NZHs1uFhZ3Hh3W3tAx9b/NHj0mSIW
wxVeazJZgL6NYcCw6BzOIq0eiid6DltAd0C+n15REjZn7zsrKByHsq2XWVGN9NJC
Q1h+FCzQXfpAuxOrXad6WUyHrFYrefElUMyf8Vffk3GUqBagnkM6dp4R3LVHomxj
++LR7PSFtXnVYci8394//uBt4T7+4ylP2Vp0ajJmzQxU9QPFzvBwCtomURFJC7ys
EeAOkfwn0KoqYOAEFMZPzcU0zxYjBmn5R3DcRRBTfWdcuPr/EyzvB2WKZRrSDeYi
XMg2VW9DwLv/SvyVebjq5m3XFJ6qY7pkPz4QJwqWEpFNMcBau98QF0JC9lkn5CLx
d8tXQsyinC3n2XT9dKPCQJvt0VHInjfcbxuHoNGW4yjXC/XXRN/ZZDC78d0p6DhK
8ZkjzKsGUeDq00jlwOhaFZmimZ0CS1NumV5AHQjTxpR5UpKdvqKDhBNTTPhreoRk
SgMPPAcMHCtKuQTYOGcljO8Rd8qgMFdz+vwCe+ynHj0ae7lccgyrdQ+FdjIWqe/G
NUsa57u+DtmJmyPH7cHG51HqcOtsOj1M2HJHCLcw0OMBL+mnlQ0ERQGGxVeeUdKg
wLyvv+8V6XWxNo8za4bLXHEi257c3BmfcE1QmQUVRivlx8LyZ1SagL5EfjjiBfI+
sM65l/my0X7M9JF8rImIAGVdaOHpJcGH+zs/8LLJxWkrjcJBbQ+9SjSgeZbGpWzN
wk8benyE9i1nsCksa0IYCtBPFNNCXQRJ1a9Vx2Wsp8dWutViVNWaS+PgsoE3D58y
Hv9SS03QXrrV/0UE5dlfdgBcVSelllCV5QYm77F/+RmIYSD16WPyVi29+obA1YMF
6JLrHcpOznAHg69mlBu2adRr1e0gMiu9dFVmNNA+3Jr1R8z2swVlqAH0xYu4sWas
32rXdoz/H+h+T/mvS+JQOLn0VCBgjJF1FJYlPCvLPpuMu9d8bftyFzwfRus+Xtba
UE5up3xQk4brjjDOLwY5N13hRmEBUfcIr5RGyuhpbfAtCztv9K5r0++9Vie8N9dC
uHdg1oMTC35HrbnGBS1ZJ8/vPRWRvyjJjPCXbYRQZD78gjYUZ1tXrZsXy+yOqRvh
/GUpjLDBxYyvTsecfcW7lXAYZQ1UMBLg7uz4UemgZYRIIIQdNRMb+srLlWGmWr4C
KS14+nVHsuxd74jaAy6S2wMbcOAfaOJhoVlXoCxKzE+/0t2jxMpy2E+LAwvVIX1L
qryvCyxpRT/wZIpbNHt9P9unZUHiYfxahkDljOf51kg3PTeYGR36WV3aIIV+jPam
GYfaUoB5KXMEC1ESNd/D0OmBx1SAT0yzHkg9zOFmnG4n5hwv2FburJWkNBncugWM
7anYDYAC8/EWKrodLTEVGJurcQx7Int6H95gvvytHBTbNY1fzgioEfVjH9WGmeFF
ggXS6FINcuZgs7Gk71aFdQC6as2bDbcRZ894k7BtudOHyl8tRO3ZLXGTc5tkSmdc
lBZdNnmR0rimbs/nG77QPoo1LhCHSg5qOIOX3UTYbfTgA58sOeeCjS5i1uzNIlrb
cWj62RJyJKpHyxJqao4a+qMcj7eJa42t6UGhWrf/6zn1iPAWPB9q3B5IlQCzSXdM
RpGpmiV/URM10buF8SZ5APMaST15e8Cok03mkFd9PnnTsPxLZ1cb9kSncBx9lmba
lW7D64gg87HpH5QIfj7F1Fk0CUejzY2T1KVAhBZ1jUZfocHfMmueKFnaKtCiNSFd
pogLJTnjZgCv/0JJ439lmBhrZN6L1oiyKNh02VRlz0kQwXtNUtrXo7PENGGNy4W9
rN1BUD2uKYkgQVDzPRob3aoxeFui0inyKGF42zcpRS9HvZaP0GYbBgmYw13COuHo
PJuEJzuQHr52sLADuO6iqvqiGxp5zJak72zalG8VnfIcB28DIDbvvPcStV9Vlic5
5lJfLaDZkP/F6FSbp4d+8695E4kk+XT13ZPolGAQNX0sv4G+do62URYWb4FOSSTX
qL/HPg/EnYM6WZLMAKolRuxUf+6qyWmtWd5fQI07xnOCLQfVcKgCiz2nmKKombEi
CfiMLeJfIOlxOMLycoxVYR2uKWkZlxcuiqNgKNXv4CpihuMw65g6mLutrGC7iExf
m0IwwtHk4fdzjza+R0aPvkZLxStUwKvZC8cq2Z0axmZXY+FpgWU7xfEhjZzjJBRD
cNnsrK1n99/3f5KTgotckb6q9lqdI2+ffpaxCwZVC1oTFsCKN6/Cc87Who/FhQb3
RHnnHQqequoy2Ta922hU8h6IbfCr6aL/5A194eADLzdC4/6lsuB2d80Rdo51nAx2
7IX3rX/juqKhSqhBgTqkoMbJR8V6bs0+yo+x2ixZuAgqpJH1c20jy8wzHxTh0P/E
KiUOdWS9qE7mZ4GpM9i27tkWWBoVBntvJ/T5q3Vo1oaFk41LM7W0datAPyLiXhyO
UU5GWb4DpJw3y4xihuJHZa7tLN4mE+VOKb6S6VcDK3BR1+1x1caE3CaqytXQmnzy
EPTI0Wv9ALaZc/YiwAY4NPiHrO32CUGFhgOsW/rvGi8ifornsVay/ZUS7pKlJRq5
Ux0704P2wS+ZmKwszP0oA0/MuTD4ideCBMuBleegMTn8NtXBAGZR61TUgrzNoYcR
ALlzgfpgcnrmU5kUjWiWBOy/kelGuYqxUhLQBHXE+7MjSvd6pHk9vJfUKuhZ107F
sQxhQ5RZWHqCpOiGkWuonan9UV8qk5aiP1nMu9sFEA6G9mlIHEwsBHVrbfCZQGfL
VTQyAJlNWpWDu1DSvFZO27Pg8vu2Ap2139Xq5nxh/yn6FElI5o2oYq4KIUP9VLVn
9I2LsLUToIYRP7Xp5Mm1/pJEcxrTAtAZr5wUhJOLq4PWY9ISX9li7WRPXePHSdkY
azEH/llDb8yXVSuZwCOnce8jfalQoMAqbTo2h7OfIISWL2mDB9kbA+8stvaVUayL
XxGRyLfVWhED/6YjWBhHO2Maroj+R4UIfFQ4dCMDqVQ82sk3FTpvAnDizR74+KY6
8BeGB9Y+QGSAgv986znHx7ucMj/aaukRlyooqMRcypv+kfjZNZtMxiSO4Vo0A3F6
4QyKdBg5YmU+uMOMmg35ioEaxQKBWcjLsQ+BUebvqg5rO6GRrEHEh33QNFF8guXq
JkUSdbWq2T1KEJd8V7FrX9CMZgoKIugPrKpCiujwfU/NESv3pdn5mQvy2oOL/vOa
eKxmj0lci53GNiBZ0DKc86K7U7ZzoSQfQHzy8Kz/KDoUXrjua1PsEJxDg/QOJ46m
UV28TX7SMIl1VOTYzwYh82S1ZRcG6/Y4Z5wJJWYKitwT3LApdUFiqi6hzu4IslCb
aWLCyTT8sl80ZuG3GZ+hHWzKINATzOYhOqW3vtftja4KmoNd3B+sdkSOCbyzb7p5
wmXqGtzZ9CpKDMCdNKQdk5vx+zNfGQCfKs7aUL/X7CnhvMe3QGfWF6FCrxyg627H
uaKXv3BRyAGHuafXxTOmq5EhLSu1pC3lOg1EZ2o1/kfUayQGF/U2JNkfDnNpCYGr
HmQl0B8GAo28WG69jh0trswXi/a6QIRonDHLlKs4wtu/7jCg5oDYVZGverE1eIgM
S4sOpWyFwbavqEcNIry5KXr3zudsfmpRnkTbh5coQNNb0Y2toCEjaxlNeWWzwnbS
WoCGghtlajy/pQbozB2X3d1IXLpYP5mag2u3YUYxoEUAZzTjkVnP9SBeJBh23ZQx
N3ggN1wR+WYvBf1yU9ze7aI5UfOsqDvXBU7/vLA3agOfhXRDBDHsdvBcPd4+RvPs
f30Nf2qephUb4/QsJcsHK2fIzAQkV4NGlat8N3mrEy7jFOFNkMWPn65/FCTgfUBk
idQarkmMmzAD3fTwLOVh6pire3z4r3yipInhPwaKrKpiHlXx9QPLvJRbBP5pb/M/
IxH5TKwLpBG5KVsBVr6O9MSW+ClKFt6WGnKMmx3u2yCZn7/28uxtljxckEPTO4jB
nS8PKh6nSaftd0FCD31I0HTbR4GP+V2gFy+yecX5TiUpQCBnyFHcjArAKDyb7S4M
OCQJsMT3baiMY3hRKBT+sfRqzzPtGAvz7df+2M/lNZFmfDnLnj+l1kZPfDuqa43U
qrwnM7eqsZ5NRMu1v+8Bexy4cRYTbjNH4fM89/WHr+hgDc7Z2ho4rKRuCqkPMCB6
OYoIBYyGXgaL/NuF1YKySZb5knRIAjgkSuJYVwh9dR7wAR+oDztfgCE7JUPo65Ks
TZxpSiRZ3BosTzVfeUpOjHY0AYBQyPGMpmoeDk1qWauBsk2/ul0Aal71tSj/UUyr
obXnyK0QmTsQVlmQms37/LK/3nYPSLO3TR2NXEYgUbvP2CF8nZGg2S9VOJ6HzfbE
2LBNpuLoNopiCYxaqw79KFG6t8/xNjWI9un4yJ33FK2kBo7bHq21gN3+JbRE/oph
jt4x0CDnZ8TNwrnwO+QgvwQKTJuaeq6OVUyDLWV5Mucoh+8+QVz/H9SLi/5+/hy0
9SWgzTvRjuLjYJIY/u9ybJuZe9ir68ztixdPDneaPtaydCD73UF3rZRLcGTlnCM+
BG1PVLyTdIT7ynFSuCUn7wMK9KmBhAVIlLx1h0fTr4H83T7ADzv7WPX7RirzKOIY
voBTqHFC2kYTO78an9AINXa25dhThDJYK/4PpN0/dPLincx/7q2vo5i4pUWmr532
yE75ZT/Hn1cIpX1B/TWnuF89sNP4oB4TtjbOJ/EUTBlhcRTGxT6Y29GQHUX5FT2a
n4ikrmYO1uAuAkRCpksPm0K4b3z2BraTiv/Uy5fZcUsGBYKeEORbNygDPJAX+H53
g7ZXlMIkI62nu/zW8/v4cYKGRPeijc2TnWCMxMBNUwT3c0oNOJowYuRdkbBG6fX2
k6bwc9x6xxuN6FtYeNgbWd5gL4h1QA+P7rloUr0uCH2THN47kuTlMKmZkg+I/zGl
Wx8Zq8CW4YgZQRft0yYcoU856JVo/aiON4HoRjUTxcH/ODBm8uObG4xgLNMYl/nP
cJUqudz9j1FAKW0AQZe28MjpXtoG0tvG3v63UJjgsl9cyMZ97wZZyR2320bLZleN
Zyp0jxHiH1dgcaF3zAJghrBK/baUe6jl1jQGtVxRNkAb/KJMolCLZE3avytKLTmR
wf8XmfDu4cuPt+m4G50YPuR5mym9YguSC8CAvdvoISJQKGP92EQ+VZ5HOZIAzOSZ
Of5bTxQ0mJQLLh1a5e7w01i+Ilrgw7Hm87VYLB6KX9pbyNOonQNSoMkORAMAgzMb
2NOUoIO4rxC2wemDAiDuSEzU1uM4yTwdD5fZo22ZEqXheeK5Dv6o2csHspu3c3+k
hI0t8wzv08c21axVLU4hGRhxUw2ijbUM/Hq/h8E3YfzXbAlVyATGzG0v1CqMjqi6
0a+CzN4CEK2PI1RFVqVbvFrER1D28SyeQCWmGcVC+B43frqXJkH8vEfgyQ7rKtTU
mlpTMeIaroCnjc4hmxgmbgn4kpgDYdGSVTGOKj2ED0W3UkpZ9imY2v0iHkwFBohj
pmO12e6HM1/GZTZ6GXNROXHepfzc0QCt+GREBvsxosbjz1b2A1yvg+xxSpvQBnoJ
/5LB9azUvNdr1EsGvuHXF//oxC21kOCqFmP6xdsJ2XDo45EBJt5wTJzzUpVAEXNq
lzp8W30+C7NLxpfmKHcp8e8WJwgrlPaFwT6m5bVn0Kj/vF6FxIiCaH+oSIusqhDN
Q9I30KCZNMlQviC7nEY5FqUxSRDLTIoGx0HAlcPZmMALGVhgK4EFtXYWHfSZYFan
WcsIbQSUFl8ULcI8/c/tOgr3U5BXOhM6MiUV5k6sdPek/yNHIRn5mCImo/JmBgkc
WHMm2Orgfsw6605u2hVxf1wqHhsVn17BUVZ1UXMNGDX7zZUBAj2/2cVWrycEiGQC
clrrIDHXOuNp6BvkNieOFgfJDHa4fE9Pqc2ETCJ3biBiirL0hbmEHlY8WrIIvpYD
W77R80gut4wu0DH2X1dnjg08zryvSyqvXrRN2Boit7QAOGyfO8qH4eADFY60Wkiy
J8XXsohmalrQMA4jJ33WgsucenE1uvO276ALukHOhOwM3ZfckaHCEDDP4MAVTXaU
5Se8GtDprlB7VgJ57m6/hH4C1suln/wCokS0A7lDBflpky76HRr/PM9Ff3ZOp81n
3H6fI4VCbqsrWEswMs1tDINDR13qZB5zhqsICn6Xou+vMNybpbCdIQWI5acen99u
+Ix5TiVRGj+/0cDv1FyDFSFDRL2Z2NNgvjRoycs/jOLyVj7zMkKa3zec/0ufbS2r
zLHmKkQNJjzECJ+MVNOuF7TvuFk5XIj7FptOMveSfOp5yzDnfVnwJvO6oUn2D3iT
FC4qjjbWEl4n9rl+XwDrYnITTCs27BwTKERiaVjtX0ER/TYUHNTWUG+/n6hOLu1J
QU4HAhznahTqgaoqiBevyZexB1f5RXxUWw9hWAT8sSMtc486qnQlwb+94Cdu/EXL
lmT6H9T5Y6A1ZkaxcvjiCqKZKKtWIBssYTB4x1HXTlWxqgAzoG8TXUI48SCzVrcs
GpICT86zcivCNXbjkxdM5dDtAXLdQaoEm4ARr/xYBOci6e0liFvII9Bjfc55QHT7
BbZC2fWtZDI99tBOHP5RAeq4jEAjDkXy51QARwCVcwWqW/RPFipR36aBIDbr9xZs
fUH4G001CETB9BvUUZBCwqcM3jhg8+pBDZzjgMeQb8GbbvCpxV7qBe73SfaKgMBo
ozevUrm+zdvKDP8K0ORC/CqCFrK+eZtUqyX05VAocPGJwwhWB6/NBPACoU8JzZ3a
/AfB2+N5UW54b8KyXwB35iRlXqMxIGdCOD+jEPOK6kNmPy+R4tAQ4XyFhtK5zZZ5
TXltHt80Q31+9Xt4zavEvbMTibHegcI1tNNhHOuBtoph1h/ACBUdAQFB0iTVkNTq
Oka8HXsnJWFk3YhAAjdNJ9ir/3i204kqZ2HRe3mucuLbdUK+2KDY3TFsCE4Aiz1+
AcGfkYBQ0kDopVNxtZ0BjgV8sIRIdRaf4M7qLeHC7fZUpUU9wHGGsTKsBTkfxKer
r9XlU7oCXeqwj9UoKclt3oxjCqpC12YFwoNdMx82pNDxyDsS5e6ISlyWGkj22to8
7u90v1gMQ986JV1tBzO6EAfHqnlIcFSEJD90byK4M9jrwe0o5G+VN0rDbOWZV/db
5MVRU8irqMifniEuPPibZbfD39EKpfewUCHDACVHspys7mdUGyfPobczznd0/L4t
hMETd/gD6WatO/D//GWbLkajNSRVNoJu7HH84/Ky8LLa1VTOGYT8IA7AgTCfL5f3
ZsR9WSzK417nQpFYsdljB0HoJDWsL6WU6ZZiRMzGkfyr2qisjWKcsDWYnAr93ad+
00ClOcrWsAMrRdQeLKxnimRdgPYvu8eGlFlwLCq7RRVMTFSTjekClcoDdBeBKf+2
jIeXy6iUWM1MdEAkKzyu8pF1sgFnFcuk1IPgXwQBqtoLSJ6oLHmZ38aWh/yIwIth
CDnJwnSRP9hWUx25tNRGRS2l+rPzuW40zRx1tI5ozHqtOwOTCYuPzYzLZgktmiCX
EW8dUbJYPrD6Z9rxezyfB2YQHQGlQJfSrCOEz8UkdxqQPu+YziSzaHxHFhNgdqz5
5LIUO1f0eXGBdSNmsmGDS4/SDuq/oKgXSQsa4nrIibDsZeLNql4GGhfDlyheS/Ie
i/DNNLPq1+Uz5o+zWQ1cLIUpIK/if+7S+ABRr/h8rp9ZqWb0nDTwL6tULFdLKjPG
8wl7kUeRp6Hk7pboB0U3ESU+RbQ3taWqyN0+wLExXPMIGYgo96YiVQYYP2hsD0Aa
64hHse0mbe61H3UNDfTkZesqAzyXsBBmhv5bS1br0f36JmuyNBFBmHY4LHaKjJ/b
/GauKoxhqd+0E8Aw2f9E7/cH6j7/D6DJ0Ofm696q0BgyToPzdBb3+AUp4hXyM2Rz
YEC3n5QEDsBb14hSjNBriDHeysEEbc5guOI5H+7ByToQSTxiyFyMLCrQJ9mZBDj+
hBdA52YleEeQNNfAPsdU7eS+sW+ARsOqEO2mEJYqJR/T4njI9PWzaQ/Hrw3xeJ5S
jKCC1PK0K4lsKkQZszsfpamC/RlDJATTLO5tPpodCnCLEb36tRs6LSs5JT5GQ46D
JAhLwjU/0CwFzF66UtJRCSYoHBHV5LATp9IARWdpJrTHrolaOD9nufcHktJo+VF2
PIEMPDBxFb6UyR5Q59a9o7UcaB9/tcGEg7HdjTwo3hRQCkJHldyANqaMIgCmgGgf
mVyLA5Kyudo9jOaBe/bl68fGaCJnojZQ7b31XSutX1Nsi2ZJ0QBRNzbq6jDh4w9P
r8ET6f4wEblozC7WANHebN2RI3FcKrLm9SJjna2PTPJ0E0vKIFmtnqIXg/miQxO0
cF/tGVqT3WbNshycHercTgQg7JKkvONlU/Qp7ZwR40izVd3lCURjejQEEd8fDfgc
o0HzrG36mgMIH6k1hP9VDUsJKxe5asqE7SJw1l5YDL53iqn+xDisE+tpaVxY863h
zHhDJM/BT2UhiPNBCzq/KJyrfpADSnXo4cYKs5c22OvFAvGcNjpkAahVwcK9GzSD
LQpYE/I7xjqnm8JpOFm7WXdSaofqCd59t+dCt889M+huOo1Kw9JR4GWmXZq0ubAF
S7woXYbpwht3bVfwUKk0Jl6Yghea+7qceD1af9hK4SUY/c1CpbnMxm5/syeYAPxm
fKTdkNAOdnd+DIjdbBjiVv9dnFrrcT4K69gQkZPmLR/9cCbH2O4MRry+nxlSTZyQ
leWn0DOPg8vX9oCprrUKSzYyuXXDKqakyU194kxAzl79g0foo4zzG48lcAre6CRc
F7JDvQ6mhJWULaD1xo9mmmi2ZXruTCASRp7IiH4PoWl0rASyMrfFkXt1nv7RiUOl
/pK5IqsbuKrBSHomIpd+9itwoo7xB8CcajaEanAnF1U/oeOOcyDdiOQ1KI0VftrL
2p0Cy3DJAvUaXn16hztcyt79I87+u+egviPlfLLnGtWQyhAUBmgGLDI9AGG8+kSa
TiORQF3l7tvO1Dll+4wq9PnQ92xdj/2OCoRTxse5bi+ehS8M1RmS2VotFdXZeEaP
sVa8weFH1SCgnY2tQBBs9+JmFfRX5E2aPinVOjRPIglsjdB9g3PqYqHTGWrmB4KZ
QgNvy5kjxz3cv0tImCRDBznqjKgOzfIMUQHlxzSy0xPjGzC1ggKvWeUGKYpHYwzc
BsBsBBXFq6KkPHji4L8VMwSdZiYLACowE8fQquTdHb/7pARB1IK41d/4CsxZ9Zqj
gmy5nJYqbTXBD+DuwmRcjGjkcIbPA2kuAomfO9B6sGzQDWTjtv3TD+ZQzAD1eyUs
43LaGOZtEwlhwABU80dHG01KTXXMZUi4eY29gL3hd4r5o+D20kXRphJ1WPks+xsE
+Tg/KhEjMUZOjbkbROJm3XjCSxg+cBJBqn8ro2udGKIQUi6AoZXQa7ac/Wfaap8w
8BvWf0Xjr/3BU6OhgGL6m6+eW05g2H1T9YYLXpXI+zdrMUqcBF1asiACftS1qIr+
2PqvOZtQExKMVvJu/2taa2dcxyJtGj7iHMmvCY25pdP3bQ23m1zY5znhxahPtJX1
C21ZBN8BeRXYfWJc2T5tIpUjttMXSvU4SaUYLqRzPsmw5KVaYrSMxP3JYr+K2Hyv
tvH6ncFVVNdZelpac2re6Dbr6qtRyCWfk6TipwUNXZ06WE9ORe2tNB3j40TISLoR
A1Zc9TkWtHZx812r+PVwJYeYCHKiMp6ArOFVDnTKpk3NqTCzSXvasdDKZPCX1Lv9
3M44wrzm9QGHyDQ890L1mwzpS+Uwvc7zpFjh+crtOJeYGZFj1pPalPmdkK9ofXBp
dYHLNTDyl9Ept5H+w0pYDJyRnFlSXgoTzJREO1oO5kvN9a1vDbnPXaVGLIWASnJV
i9M3BsHENgapVyQtigrV6U61IEQdxgmTsVDxxN+cgWb7LvZiqg499MjL4tmuMU1C
SApZKO1NhZy5htjL+tdt9h4KdV5iFUTJFORYsbUAyOzu42tgsiR0yBm6cRA05VJv
fTyuzC84N5YJdjzmN2m9RQAxrYXihKV2sJLL74oYksP0LaEHTbqEgYcCQtqFczuM
AuXB95KlpN2lraPvGSCcbARjHTA5E9cqWKByUPXKHvC+fjOamkPi5ZfM59AMoyZG
7tCTzQZT/7uMFpWt8SoOPEtl3o/SAocHzxUv/xpsg99FncBYiFdbOsA9Rwbhvf6G
IYYOyC6VGt20cWWw0jkhHtG6wlI3Uz0EoOw0KCyzEwIWFST0nCZk8+UBf0SJMD2h
FvkyUMT/UoTvGN8mUr7/bPnvdiziHskeXbkIc+cXD0vGWFmtiZa+wNSig6kQAkVb
4d+rMHmFk28Ptf015B5UgYUAiLyYQDe288rqY2oCtV/bGEbfuo9p4EAa2SGLQt9A
LzJqny7mR76Buxl0CaPlocsPKXmL9spZS9k4mUISnrnKXhXFuGBPJbyqysrSVdK8
5lnGZAYlX+VFRK7+qe1xxszIIctrbvkuMtcsfXZHDov02LFSAAsGxI2OM7vGZvA7
DheOaKTz8mSs3Pxofxi7R6RwKHyf+WoislGSwMcEiAjUM2GdWJGI6ACIkTjNnsux
gWfYslxjt2OHgrI5/KwKXAILGdmbtO4puOyABOcQbVtpLJO2sCqpjlQVR8fJGvd7
ye/RG+3Cdn0enAgfzLKvd/3aq7Oc2tZNL7x5igWFLljjcPDId168ZCP1XJ/0MdlK
qCL//kXXTPGcLD4eenxhxjyUuJSolPmG/qLHCxHRQt0+fb+1Y9RYqeal/7ndhzbU
Uewoy0i1h/4S3yOU+2zFpdSiu5dQXCiam5/bNRGyxFuBmwEke22ByR2yBNJ+COAU
xXglWSxd+1Si5GCTCv+rSp+Qqt4Lyn1xCvq5Z+KhLlrnKtFZm47hSaFN8b8L8WUz
HIcyEYpNYooGT9fyMCMuo6prFh1CPdAhwYsombeifhr8DMEIuxH3xBaLrv6Allr0
P4AfMyikU1AQnUM8ZPtYCfz77Cu4Vn32RSciICyh87CrJM/GSQTfFJcZKa/OERJd
k/lYSSt7Mut40OIu3xVb3Gs40+4ndaYn71Na8S6HDBJw7TdLcWj03veVLJlnII3J
W4JDivMWFc6kut3v7bhy1KUoWSrS6Z6pOCV6gRE0Zk4lKIhOFvez0O/apEFSZFlL
LcW2z/ppbRZurAgRqe/x2fD6mahm4FiN1iXsXqTqDC7LxLGa0iYwhlrP1OGA1lqB
qU7eBcnqm2aUYrKpHWgKDXxgCQ6rNVcDiFkMGPIfdcrwZqsPZemX31NCaL5YRD/O
225aAC1Zu2k864qL/P5ZYLUNanIht0B7/kOlAzZ5ZsuBJYO+X8GDsh5zeN1EigVd
sFmdU5h0p8ao7m6rqNdl+yAthbaBqoRpDfN4lAfcsggYl8/dGYk2tdhLsOZvDZiQ
zojPiaxogHX9PEvI2xbUt5Z9kRLmEz+AxohXS5OSN69YJOPOq5TX7UgUPMjkOEuf
ODJ+ITPrEDjA8ldQG7mln5UYZbjP37wsban5dRAGZT0HkyKjhyCXAuPK/PETFusr
NPpLINXqvqs24shifdaVjIFkqGgLHLEtSzE6tEYobia4m/LgiKlXd0gvyzKKXjri
HTIuSidsYVrHhRtxzqjfCcuom40qYEwJoo8Ulh5X6oegqdiPN+XcqnxPE8BH0lNo
yy/laqPG7p7WzSwMnaTHRDP2KD6c3jq+7PKtG7t92F5+k9S2Juff0oBhxMIp7abs
L/yue20HPyxuX3ZEJpv6JZumLB+X8xylhjq6liXd53au0FHRtgFUugowBZG5vMOn
OIDJmQqGlvKo/jBpeu3+e1CKlB5H2/Ut14DLlG+f/Qhgg4auU06vcHx76uO7Nn+h
xinICWPqE0I9PehswXWN8ifNhECtEyGHUlomhoW3yqPrNyo5YapjOCzBxn3VJTw4
aBeguMwPOtHuoSxBrUNd+zrAoQODTkUoVH4UECLddcd/pobjiu1OjxmVkdKnrooZ
3q51ztcR28PZZxvbHMWbwJ4qHjlkERBIvIWuthghNG07iAJM8r/byLcrAKYKnmWt
mwSl78lwdtPIJQnwzgGZcMKYFAAKCQctRFYzMKK6RjqwQobydHK4CUR991nqQ1t7
y/hp0x7Vd1LAUIFnvIoZqJXUGtCf+G9eAMexthtW80SYun9antuUd64jYspjVSo9
LKu9o3yznamVWADbuOR8uXGHUn+dH/YyTjpH1/XM8zy+owzB77oupqE4UiK8Lq5q
2vMCt6d5zgV/r8NIM1vpgDvm1e9hD4L8rvs4wB5SYxT6fiOEEyU5WF7nhm57ZwcM
ZLHJDnk5tUfeKw2Kys8HmnXlXBD71DlTqd8tQ9UcRw4n+BIaJ/nNH8lGkUG0MFFt
2fnhFpF+3bn7RFHZJm4tsmjunnd6x5UtcP9uHQbCkcAN1EV3HF8OMpFmugognufC
jqRsjiLOG+e3Tamn+sxgblS9hHKiyi8ourKhIxu7VKf34FLtmwOLuprggZ6g/Zem
o7b4IJvKKHkSeZCh/mgDjJAeCweBC7WEay7TU/Liqfzi6k1rs2cQC1SxlfLBScOy
zxHWmU3/o+ewS67gI+KJM48flqFnmNZQlHpQjuBDSspJeNaaJoVps50pyQP7ZzAj
RDNU380cQM/DxKHzse21FCzzqEOMIOgh0LOQmnA07AeOZ6UBI7ip2co3OUKTRpGt
17GM5VM1sXsWqU68dYC5jVIuVsZL1csgdJ04IDbGXQZthZO29OPDjLQRXt1C5IPP
+v9jo01PWa1+pg4Ez5XOisl21a/dGqz2TdgZIuE5B9jCxNGC4Jhd4bQlbMXQAFx0
sOCWSwCqVDaNSw+LAZSWINQy+1CvluLmrAUquTE4g/KPT3UxJfrCVO080mIEdlqo
dlYZgnrAP1HUWC0EQ4HON1rziigToRrUz3VQdr5LWYJfrSKIro8rwUQRC+2vYbno
EoeHHCpRuvyZIfN2tzWJv/oEiz3OnhzrbFCLOq0z/kL5hyVbTdk2a2kIFoM+yY7d
FT1S/DWkBN7BEFwrG81x8fgjpQdX3APpGq55k3X1YkIr++zL4Lw7Ic9JnciwmCkF
rfQtlv4MNVNYGSat4oXGBq4cT15U0ZSLxUfOmsvZEIWwBCmLPXIwO6zdCFpNX+hZ
YXG20HlmI1YgOK1HtlZl+JHUEi5wraOY1mypNlzlK5aYLvd794cKEqgq2veuSREh
5/2adYohWyngbisP035nNrISHP6YLnYY2g/RwAi9KRicAz02Uj0FFg2MAoJynvJB
2hWO4ytJgQuKmIHGDYPyYLmiBcksVylUBmiFTM04e34ehfQBOd2Qm4tTUUJX27dW
a+rn/UUChFqLyamU0StiyEHnn+++y96HXMS0Qx4HY88rebt2mqyndeGYdRSy7y+1
OJKhSARvxjiO1zg4MRiQNhSPJsWjJP0FiQmPbGtNqpsolu88ts8QCNMAxY4SQVhF
Ktj58XOgH92wefiUgvqtwSyGv75MURuqiMy9rmMnNHg+P8NmZALZ74nZz+fGtQEM
UJbOI1XfM5sB++LT8qFDhbmM0HTkbgHk0U8g0Xrkh47WdFnCLLK3l+tbTeAUdoJo
bMIBzLS0xlYsF/L+hgaJBGnb001Wv5g4oAZoqrsK1YJqxEly0XbR10Qc19Decgnq
rurwzItFq6DUYatyfofvtKdPSEY9QzhkkLbQFygErAlOFJ0oUWgpGVg4df0jeVyL
QnyoLwDJSLz712gv1sMk7KiRn7GsRz0QakFOxRQHGHArqR3UMof/2kNU/i0nYwP4
u+7z597rTvU41gjViohZ1WlTRRYn5EwbgSZ/BShhBhOzpqOaxxd221sBclhXPyv5
f738Kar/mLYuJzr6SY5j51xmzW4IamFSVHGWS0DM01WCv7JsSk6N02UEVTGV0554
/dMalomKo1e+AjibFTfa7V7URNw6/qlDA3I2bIAKdf29Np1bEki//VZUgpHyfZmZ
N4mMug6c/eTqkvbkNKNcp944zfqoSxqoS0Z1PkEdSEZ399h+e5Z9/LqWHOhQ8Tji
YLxi9hZOkFkUEZdmu0KGFtW/cJOkov/2i3uvk3IsJCssmxU8a30zfWLhgtjaW7+H
1AvzW86lVtEEo8HG7re0riLC0t3ZTGvfUVWsF+iTTvEsJJOVWYhpQBxPNHNxzKkY
VFV6z7ki5YLr1fTAH4YMAfsTBaQ8MfViPgWINZmklsL056A5yFNs9fMM6S3F1D1x
VZ8cjhWptb6NHr2ixcR1i29TN05Y+fayYT2X2MP/0p0SPYMAioO3uEOc4rjSX+p9
3tvIi77DV4HVZ3TAKMnzNREl2bOX/SnF28iP9s4egZbpDDpUnZPOCg8FF1cKcaUt
Kc0c6+ZASc8wrmVwjce7oHnnUqzWUkuIlPvzhx7l/tvxi5+KOGi9Mu/WKyFVtAqL
VgIMOXnNn8RYGcZUt6+6bxxrpT7kOi5v6wR6XEnEU+25edqCRnhOyoyz8EZUi5uG
j8zkPv3GahNF98/VojwCHt1oZNUtbZs8/GLyMZvIlSPUYrE3RNojAe5xwtyjdL6b
lYBeY+AspPlWaXMx2vXZQ9kWSE5xQlNtoa6CzuPTRtjuivELqKl8CLJv5JlTSATC
BYG899EBa3XZbojVPa1rUv0qQY7BQEHiOQ3WzegGsmx3j84jggFrV3CcGYhfiueM
v14leBRzK3VG/Smyl5ARe0ipom4R0uSEx9kgotR712RdSKvSwypiASVhNo/XtuPH
d7Z/CNjloseyw0HP3uA+daANNZ05M0Fs4++T2Q5haR1Oge6L4A6RoIZor3SCcsgf
hYU3pR3dNPCs8p9tPIaDh5U4zWsDyNGNv0NXKm1qZ6evcu4cTi9LCDwfNmLLCZZ9
juYALacRnEzmu9zVKC5Q/TVohA+YvChJ+HuBmscLdo4UKyr3l9SxSaAj++xETm3H
dAvHNoUFbuH27/yZbExxyDBEGSLCdCrDJqlGS36Nc+ypWx5FaY1OsRJ4ChEL8idF
8aeZbSjgCvtyQoN4sdlEq1nivER0uY3nWWXPSPo/TWqJzpMufVZHmrJIqCJtjOpH
dZ0Ic4TE+I8XNIYlTCCQ0hwoO67D3dsr0lXDUHy6TMp3UVOaQ4pcVWZDBI3Mfgmi
b7/tWfezifBSFkGxYhfs/+s9hLwMvQw7VGmxOAjAAFFRTC2ufCIX81gRiyKV+8R2
i9wjzzQszGHCeEIVImrYTTul6aXe5+JdyUHYpRqkEdGGts1AeJ7x/zi7lC2qAJSK
XBciT48XlDazyT3EdRF9hN6tfESpKJKrOgmlQBiH6cK92THInHsH+na91TZB8H6I
8OwYGCyH0DkKUVxqnejGPLXWnT8nUAOW0WR9uJ9luOkT9PG/rDZ6e7/hrtrzKwSA
N/AV8cckSrXcofj1YnF/DB74NVL9+VYUoHZCuWC6BSg3o+s1H1/7KNpXX/Jyuxn6
ljuTPkH3clwvqJ2GaaQr1P1B8gEBvqPcJTchYnYtZQ8ZsJzm70ijJMheqdlzek6S
yi5NTOxPR8ctcX2j3EErmCEt3NMr10/QNcnfwl+wj83B6I5aOpLcobDdEjbdAkf8
dMfE/Nxz7jI+pRdhGqLE/z7IAvEkXj57HvNLfts8L89WwTOdaMfybip6foKTLOwU
Yuhe4pJuRoe+8Fff2g7iTWFkknJGpsKhodHCnzTDSJvtSWVePLVoSxOlVSeA02sv
Ka+BX4J5aCsU9Z9eLC/ad+iiSIjTw23v0boOys3MDZ2Wf3cY26Trvfi4Qiuk7OOS
dc14+8b/al0NqcirmJvIZEm3clWwxIVmD19E75Pp5W00Uy9iGnjbtJaYemsuI/A6
fUbLzDgH9BWQeanMDHGHkKwzcav7zE1Apmprx9ecaipMWtV+3Cj3YlJZklQWcYJ2
CIdwp5Der2MNOEHmMnz4iNtwvzOJ011pcPt9viXWew8o61JbS5sp5+cfBhNTmFXD
As2dcsPmyuXvWrSWucF978t4UXGH0csqc489++cvOFQ+z8U3hZbR8tZJipLNIrXF
nfTjGbWCUmx66jmvOujrqazAdFjvVwYcjQkRmjnDDy7kCVivmlEdj9yvkmsU41wj
hvJaM25VSlYeIuw9a1MH+dVzS/UKE5wRhudcOiBMqqZqVIODHe6ZS0vUEwfzGsL1
pfEhoEgqwaUHrJxcoNNuEIw+2UGJO8+Y7G8tlwSeJhPylxMF+EQc7nPcP0QOuLen
EEBYWkpWNRumapcHehJ1atq+unfAGk3ya/u6lDofZDl/U8jvXuomXptswiMRgcSJ
iem9BaYGZI3nm3KUDvRmCv+JYNb8T2EKkL2hclVo7Q/fJjYqUtY6LMumc+UoPiq4
8Sb31BrigJ5sGAKRYtUXxc4qvzY+GQltEDgM2MMS6anErpirRcjvM2Dp4hphJvn2
lhRb9EBZ/K84OK7zfB3uuozMDyKkTwQTYGFf1n1LfJJp2OXLv7AADC3RcCOrXchF
ApXk74XwoGuA3HTqCuuaNez6A+FOUxmQmU4lBfg89vdx21jj1BmRAQfx99FzqT3/
NhBtvULlOz8lHA6RvouHtSuk9zT0VxjPkoAQX6vfCK/wG+fpBzHz+5oSOeyHXB5n
8wqVow7rFpJ8irgjdBdiD40/E378opiZ52sF+qEUZIdnYGDeIRu0NufS+LL0I9Z2
HhdsfKPXfhTmpDZoQWs9jRzq5GJ5/xnQQGQueojG4mmI7iy7FLZ83bme0ahUmk/N
oewpZFei7MAFE+kmzR5krA3pM7CVEIEIK+UQJsUP6sacyoXy5HvlTGknK0oWf41J
7Rt4sMEC8F1+YDr5BRO680NNOxWVYI0J0nNzP2s+RP2Ku5tdIlAhFS0L3c7BC/nI
njgMSix0fElBAxAW4ihBEEO7WMzfYmOv2fezma4TI8mAnJBqUMJUOrgDdo23A+4E
e7soui4QLoRMMqOsR+w0wK0Kg8oVSAkNS6gxZxHo38V2H/gYBtn4B34yAxqpB0Cz
sYkdR1wb35pI3IQ7HeYicBCrYc4ZHPoQLwQVRAXzUS9BjG84AJidPayZtakQFtKt
6396C/VpKskLfeRfbhjPhBLvK1mxLtKBCIphVKUoa432IHc/pegY+V1YuBirZCPb
Vm2qU74MTOZwSQ5uthyP4TYaQkupfSnAJ9jSufx88cXoZezeErMEiIXPzF3d8wnK
4lwGoPn5CIChxqOV8E8/NpVlL+s1vNoeNtRO7pMbTFhVAilfTgXGqHYDy9oOIuWr
fXQpUe5YheTehHG/b6ofgK9x2oUcbwX1BK91y7upnwC3mO/qQba0m0eDDw3zRJb+
6MupYucidKKsHgiHTejuvsjnm0I8pekxygOTudP/73I1s+ARvV8OORJTN7fdvWOD
3RBoK2sAMYAyxA87IK4Og1Vt4LKna7Qxbf6nXPhHN9k/3VcU32Bw/RiMK+ZdcWCO
hOy0N6svgOHK/TIUo3nAqSSGSwTVkK+Obi+nQc2SEe58dodpjs0JTBjilyuj9JnL
5dtUPl0idpiskkZo0fTmT7M3Eq2YrB4PL4x5Si6ynPUnZfg/oZLIMevVo5BHeE0R
U6psnpc745JccVY0bhk7/EILd2hkpG2V6LlOMElHCZAizzXNqlLoRl3BKSCVyLqh
LxvU+n6EuQxvYieCp9p7EfSYyylLDBwhvOe6MJ0FXFgHdg3MJt5iflSUqGxcXhAj
DuKZ9lACkA4Voy09LQ+Rajti58KoV+idRcI9j8DN+8SbY8IuInb5Nasp0tivZIC/
J3h6u65bmHI92DyaU2ri5kgwT+/3hGDrWetdI4ikWf8Y4FeVU1jeaKFJ+dKNRG+N
r3boYUmVh7iyji0ieoXlmvC5ynoR7jag9BEBJw+X2Dcu01ne7xxg9yrKBZT99/Cs
eVhSMjMSjKW4Iq/Ex7nq+L8kMVaeCNBQudWkON8ml97EaCZotrd7oPclRX1ZiJ+k
J5efHiYAjxqBn0ZnMxv2yqsiuDcS43lkO8WjmMam5LOyOSLonSmP/NWzu3tyEC//
1p8TE5IauG1ylHBY401xH95AQ/fJu5MT9pYdApsm946NxsFX3rZw8ap0+X4r3kFB
38t7g1UL+o5G3WShobRtOPh3e4yE8+L0qM4SA5KWe3Z9i7mhW+kqg67vPKEiOw0J
flH+GrVNT+lBxe8kTwohVQyxTMn0BNEczOwyL65db/TKKhfc6aEFJ3rGOUtUmViv
u3VErUhPy1dyUmmduHlw/Mnuq0SojAj2fM6wfn2Sh72OT07i0HdDrT2TkFzoaTvN
uDM074CSLEeIDLyzxH+db1pfxItT8Jq0Nlz1qh5PsHOV6knm8SkT8z3qcZT+mJip
nz2YHUte/0Guj/0ZzDc4Zm1fW3lXgFqcNdAj8XgZm71UawOzJHCCnUVt5DfJTctE
S2L7u95+Esqhzomn0cAV73sTM7rfxzSXK2c69u8mj9D2BV12K0ctKta0oCI5AW6q
8x8oDCmVC/1Aiab/SFiAgH4xa36mF8UPxz2X0U8C621E04zJuV9xJ7MofwZdTrr7
9No+FnSkj/XlUehSKFJQhU+Ux8OUeQkQFKv/DdBAkxEn4fb9FxBF9pOUADPa7fOl
w+lW7FgecILd3z1qG/f+aU46VcGh/g+ZogVIHyKxsNk6oB93QQN/wbqv6SNbL0E6
iH8acGacECi86FzRzK7EG9LBgsgKvAoB+/PmnJTcCaAtlUNlSB+SXszU4B6PE+bS
jpWDbtMCmII7UOJ3S/gE6cnjVc1aOVmIXvstDTDsOGzpyaWdGZ/WerctFaLwyAQh
IxdnxD1WMAv3tA4D2+KkcLBRYFbBcRGWvADeYDENmduF12fTnu3pPXpU09WXXYBy
Lmc2rb/AYJQFdDLcYZNdpGSm00q7gXC1C2ePTRXzJmLo3z7THta0zahcIUKexMiH
mkSnhbePKzmB3XsV1NhsYfDQcL0P8utNXdCbwc1XfXMuQ3KiZBpg3QEA7Mt5REZm
wCuoKWat1AFOOMBbHr2SLaFAD3d1tGjuNV1wNdo98IFChDuE90kT+H4TjBz5aUIM
l2eA9TPZZ2uPBq2NIVxgwL87n7CpkCps8FIqOn34dGn/5uUPY1YbGwAnpznsiB2B
bBvQOPlSKnk5KMnSp4TZOYYoI+89uvv4/XbD4N1wr/uu25I69plpBmrXNEqhi0rk
InMlegQD0xIEqXjZ7U+mqe0QhcncuNKs34B1GnvsWJyH9T+2h34fyphMHsf3t1DZ
3oEWKsQT7umoWBrK/TIuKqpKG8JxNVgol2KEFh18EeWBMY5lmaD1mTbNGwFbogVT
G5b3smFHQFeeUicKjsCEI/bMLVnsrmpcXjV12NfvotaI+jrqXBcowYSFGz5pK6a8
mOjBXOAqZZrLIsJi5o/tlo1DNOIrOoKPJjaONLuvmesn9QFqpu/VHjs5eNQtI4VX
z1j8YU7Nr46s4Bl9aVlnEtzTEgqETZVSJsk6pk1BD7FJ4Fx3QAkRmhCyDUDXNFMJ
3vBJye48wh034hPpykDL71IX3tSXH9d3q0V41VejwR3hyQwYuEbd5udmAoNVKc2p
n+OXTnYDaUkoOlyb7Yti+e1BT1Ed1ecVlwqelGxcmNRivQLA3nGSn5jf5qFIK7Fj
hX7P4foTJpkTxUV9TYWXByyNMsHgptvzDva79JSWgyoQ+WNoIVfqZ4K6jo8WkhgJ
xapnkPCk93DjGpjL1+ye5hUvARY0BAOQttbdh1yojUHImVQjcQupAob23Mzz7FN4
j/aHzcRZ1DZJhJEwcbqpIBmo6J2UB1ZyadAKCu5Lvu3i6p8Dqlitinh87Xcyr60I
B/duIHZbsjJgS+HK2nIvGXx8ptfgg6r3X0+OClAupUxczisrW30I7YHcZstyYjSe
qZzOazo44ZqHMr+O18bag5ouCVhX3HtDpGqOPQuf/KYmzMlX+oQXsBDFj5D3TzeI
1yGvMpQ2XwacLV7yIIlJZsSQvS8hI0X/xZ9TN7ODOys/kVTY4tOtac3OecPzIfXG
2Eoj58EOPOaD/zBOAa5MeU2nYyHy9Fjm4YhI+xqaiINSt0wJ6xqd/EAazkUe14V4
2JjKY1P1ay84kHtAua6IMFenCWZBotPeOcF7bOW/kNMNNkqYXbhXsQtefA9ojwBb
8EsdmQ5udgkmSd3yNqK8CzF86zR9XbtPEUj0kJyT13HiLZFyFfFhqgYXCwFpZJF3
Kvo00DnT5v5oWPll1xQMcGCZYNx+0PgA3pGvZBUHP7isMhgydAbcCCOiOZVynO5T
cmXDQyUAZ/ld+kCnjFtAQs490IsguCK6htx6TE/kbLkDa5Kr4+TwIZQWYrSTG/YS
WpN25kVIFQ8pa7u92Gnz1P+Itb1Cot74otwho/E2mGdPDTNgXLU3AAnY2tZlnKyU
Jd9eNouOXb4DPkKP58OLhAfv8xFODbNd35CdIlNfx3Aqzkiog/JY29/X3CNsvVtn
jNHIwZ3O7V24YssDamedX2kdyLs9WcFosc4p+P6zuQc/24aYvI2AJX1ew0DbCtoU
iEEcwkPX2AnfEQp0QnpFn+dpkNRsu3F0alT/Nk4OhsiDx7YKpZ+/uWwwbKLr4U1O
mCS2ACfipWLWeMTliFe5826yTRd5QLiIqB+E/HnsgP3MjzBW6uZqG8C6NmpoSEGu
lL8GR0KDaXXG3SNXzdFBuxdhrXG9z4GEj54+K2TL6tribbzSwezKjfbXMxixkqQE
MAaLJ/n7Gb2ZzkeoBxSQTOJ3fvDdoruzRHLY7HgnjZz18wXu4nqnRhFYIK9FxgqT
jzKV28pUkugXPah8RIRj6YUj2spi8cyznlybXQ/QgvdjudfOmHYVF3qUusuV70f2
XVljcFBXMAN/XuGGnSHEfkxi4bRGYf68QrCb/yt+5bH2Nh/1Y6pDFPpSNj7IRfG7
OCQfrDpS214HAP1ZVCk7UOIgOumHmoTmnRMrF0/nTd+fq/gSlZw6t87a9ZapXgTT
LZSfM42dYGdiP38ohzD+gZjni54l6z9IjoBmCXnNYvMuKPh1WT6Dk2UvnR4ujOWs
G+K6sWz33Ap+HUyMvsXmfSQSNflEj2h2/oyg9YhmwB+iQXE6HG4RkeGNSsKXv3YT
unSdxM3Sw+XmOLU+2gjcKFSg5s4dEhBuGobKFg4dbdcVhc4STxg7o4rFiwzAN45C
n/ucOZbenwaWcdQxoSWHw+q1PyBsuxfPFF2iUA5pswx+ynYRcCcvgM/metwNHkjk
7ImOhRYraYVJ9UEfqfgdXdjlqLArY0zD5XEzJMnaFzh9L8FbJDVvJUMaKKa2tpD/
qlp625zgf4RMizplL8218RmTZ5fd2jyJCXwNndiOGaXchhHSzwPcSGYU6hbHd3Ny
hxcoExhzdpUq9mdzRde17K+owrp+9YKbB5ifzPk3myc9jGGTlGCutIA94RGZ4Dsk
qnr51C4wqKZ4J9gX9A1HXUWtJQI9mlcVGyAxN/nH4jy2komXAZr8T++8u1xn1hPc
OKidrI17cmIMwMZlsJ0lNiekV7GbvCTNLBJTHOi5b4rAG+ACH6ubssSSPZqK6NGD
LJGV9JT3cC1BBKgyfN5PjSYi0g/toJEB1n3kkjNVQ0Nvm6cI4Ir93LFv0k8oJsRg
ei/n7KIbaXoy/BCvYg5SaNzjXtHk7F+4EVX4nBvy2Mq/d9bRpOI4/QIldI2kr7gz
kyTgnBTrDB7HE+PhYZ/8P96faRV7jDaIvcL2NyypzjBM0UaDqadtd5Am/v7Q6im3
ItXCBVM1pjHQE2zmOnVNKdfAShXw3uj1nlbVDf9SmhDe70c/dNkd/kHyQQnlDou3
YunsDFwNLT9GjYQS5b3CH98cO/LmAoJoYMHdwdDyl0YNNcXDR864Z/jOT4oO9Csf
gcI7Lwohu5oESKO2Jjaqhmd8U/qEHW968ikQhuYmuKy9+O1r4ySNYA+yfnOPoVTz
TGwXtBa6ExaaNJOkZ6eGYveC9bzTZTe1WYthUA1M2I4z98vjl8K4+V+0/KX9b6GG
a4F3A20BO2WP127ZWSZ5NxjJyIyR9xDAx4gxlYCH3FMWAIP4mXMg9BBTfrUzL0iT
6YYw/sz/442HNTmEKF6/DnRe5Q/gem0U3wd4/yqsXJk5eOOQ198ZZ2Qx+mhJc4Ic
d51iBIN5kOZNK8NMIcV1m1rTEbnsDHkrDKVaBRWPQ5kOrxKp+slM5n9Rr9WRFh13
DH4BxwT7dLNct2Bp01p6Wh5QSEmC+ZpdimQ/6K4RtdDdFfJAGrttJyCWNAP4laKi
ziwX9sU4QfDx86aQt/X6mPFsXpUI+my1qgg0btoosRXw9ox4NzCJbrswFyaVJEkS
CrWM9/YVWx5iI1V5+9acdzAKGeLELi5eLpcntrqZRSY9gulz1Xm8N4kUxOeqq5OU
go/s0gQB76uZTfasH13EkqvgTT5wG3xg3C1Ny0eNrQ1vEfA6iGjekjHnAS/kw5b8
Olw+5zaVMZnMN9OrNBrp/MdbO1YYCVGgycwIrObpuloTd3hfaHSxmwNcodIXdkJF
+uxAzUEXW7acSMG/T518tiHReUdkpjr92MfhLw4PM1JM2zSkA+2yL0PJGbxCozQY
fx0+/4ZY8RkJWFDzxfOwFllGVWclV2SJqbxrdw8CjVm1a4Hkcq/8uLxre2Au1Qid
GJ4LFZYaHFu1yGS5pkRz2/qbrbConRLP1fP7/ZbCNa6C7c/oUDcKljdS88HUXKvY
RNAShxljiT3nxpbk8ihcJaadRWVox9SgpSLAz7Ct/PgYryvMAKphZZ76mW+jSoUh
2INmlxM06LnaPDmJkRuRSH7EyJgvJ7QGua4FRWGn/kRZgDGckHbm8YYvRiBKfaNf
t77Dt6OtsZgif38N2s3JxXapnLnnraa0rSm59P+njFSeZYb6FN4kB9vxTRrZQx9f
LyGcEAuDfJhIWaOGvx4OQA+fCQp1nRn1poBEG4R9fsA7hX2xg7tcKvyMx5UryShT
ArwmBHtAQot4OkvU5jDje7KGcRbAo2pMwXis5AknyXqqt4AIo9i7HnGO0r5IkWY6
ofiKYPkSxapoqpv2c7kRupo845gkTDQc38Ypape0ZLEeQfaWU/XxFyv8kmypgoIi
PvgqdDGlclf1mpu4Y/Mv4CGiwFANkmYtOfTmC4nDSWClu7pCpGr2qPinDebpATt/
uEaV1yyUJbpnOuk20lyLExvysD2yxJlHr+U+cHocWez+hFHCpglef+J3CC06xI6N
JJ0S2pKIGrP1LgiN83sWEw6uzx8HF70oqwXl8GAAEV+ed6II8O0+Vx6FixwPXoGk
CKL5BGJNcVeaqxtGsRlD2tHTl52Puc2tBj0h0UfPWnDl5tL86EJylTJykQUIXjrJ
6GQo85x0OWEYjqusLH1dNTYQHKtGvlMpdQD0nkSqCwmkdDp9u8M6gy55OwPYosY3
5k/j9RSeLwhNenwuZ11lF2KIfB/ZqKx8x+hCEfHNPkDlLYVSgHiLzCVPDXBWELK0
sOicAAHukk1ywZmpu83Wx2T8LG0qWLnfHBghfcDeI+TJkRO5jxTJu4+sHhO06mhu
S6a713fCrJ1XMDpRh0NTNgt9cfVzSFIse10vp/+yuErPRs6j1oGQlaYFr+ulENwA
GBLQ7MKMTlWpfbTxbTsl87fFL0GeH6x1LDCn7ysrmQnBYY1/6lnAqj9WP9vOCOg4
tv8sGziEfz9yeKphwJhNyRYbJtInTIrpmPqtZvE6XtN7GYPM3I6gthC76U87jANi
iu3c42LiqFgUMUW3cXeln4CFNz2DCiL1DpMas8pmloRYBna3RlKldmMYjVoHdAP1
wOTLYpOcGkOr0BeMVe97BWMDa2xT9h/p9WqR/Ka4clK4lxLi7d2+2YOxH5QYBrgL
lgdrRDl4E2H5APs+bfKhuvlmZqmp2vcZOuufQTCwxfjJrmAP7ahSU1EBj+wYwtx/
/gwW4IpZFy0BqcYNa9iGj9SHYUAvAXXdsK/jjv77PE+stGTzFAQ9/4/1UbcLI7jc
iUAogcfi8xJLtCXlMABUTIsRDrGkFD4mAn+0BWA3tQ9aCY8T90AgbuM/hNmc/tbK
hKNQnwpVuaFSFav3wsC/HcqSaoSsIsCbkk4RhQ/TyjLB0xlXk9eMiU22dB+yy53k
RJSrA74D/mUJYaLMHnCrREuBPvUQ61Lc/tzR7EHUsZQlAIgRg+drxc8NOyFSIQ3F
YeiGNESSzN3inj1twD6fOpKdwui7aCR/GfQF8ASmXCGX9qlp/9pYJknGCKrzfW7U
3OQ7bjuGj8iBp8Tr/GvidECrKigBqzhhrhxqKT9e5zEcvizoYN0usI83rAOKMDuj
gCp6l4ulzc5ICOjA5ELhfR2AdvXtCwTVhklh52AJFM2DyKqgikKE0uHLfmQzHYsr
qD/MLaMhDlzOhZ6PF+7bXFSxCXyLGlA70jaNT1510Fk+z7ReIilUtyQWk9JLkcXF
4aU/zoUHvaDwtHcNzLR1lPyjHRaTaS+TsqMPhAOewJMqTPyz5yhlCiZToScuAi0D
/5baBeAmraGSAHouqi5S8JcB5DCtLeRMDZsi1/C3QK4vwsAdTw31q99qT7+4GyEu
rxtlLXhCwMOIuntC+XY20tRD9xDZkbSdlF/5VcFS/sAHKx8Q3Wj9pofW/ZSKWVw5
YXrtSGa7lWN/j1iFwLj2NnIrvJzCX96CjnAgjEXirarK3kVuAgolK4+8vzzOexw7
YANr/OlUy/hNDE+/ELqdY6Y9jXaU/Ke29Q7dXHrpWJcqXWfOXatMMh+huh5Db1sM
WC7LCVMPPR9X7X63QwSjgefuP+kuAuvz9ESEno5mxW7XWWkT5pcYrqtFQP8hD1ZR
q5xXs6Ma1KjM3+TYKkHT0TCNc5JJKBn1EMQmImFhYpZaNN6dvBUIo2FedVDm/38F
xzwCtd8PpVSfbSMyACjFLQah0dI8KN17SU6/zg4StYvEx+tC8r0zYpjocSFpka1W
yKylpvAT8R8/loc9PwZe6KPEn1fR4HaZM8VV3sfq+JKYLiruxKqd6LxAIbFg0BQg
rRK+xg430eUR9akSUE2WbA9T+zZU3CGsnMFpTbJGjpQ5DMAwiMKPiTktgq3swk7u
Aw8GzvQdC/Dk0P8JNzAMT1dpGot8t77b+cTvUOSAFOBX6NhMJvi9UFpsUuRy0nFP
G3+PcwoX/fxoAWw7EZpDd2LBLavzhxkjDo9ulFrs3quP9qpwyy7jfDGRfHbJBDzn
Qw6ISQS4v2RFt3yeKcmlq50DL+EGJB47ppQ2UXKcv8NEx1Q6g3n0bTOcQ31PgrcU
mPNlsW1p5vmJpNdsEheyWRCc2o6upYPbSFpDo2fxnWnQ/8mwTtiBwNwmfBHy+zUp
7YbPd7vQDMU5wNqocQD5V9uwGc+OJg9PhyQ366YjExKi6pjUsqNrg2nJE74wF4i9
VbX10PHDZ+fsMEdN1dIv+kiPlMY99oePetAYO+kELgNIN//3+h0vk4XI59EA+JtM
RzdKsL2dP4xeQ7t/yb8kahyvTKysjaJQJ2A4uC+bkzyDwf1wa/xTwom+97eOHXsT
s8bCXe+PE9lhaRaE8m6ccC+isg0pYZjleK+2eWnBHmKysn3A+dhScx26g6drnpze
c6HJhrOMFFtO5oNeNfPvJlWJRNvACQrJxXU+OS4imSIfnS/8C9L+zWLZAf7MU0Q9
8D4/y2NtEZmsWOtIx287pLBDxYAuIv/1XYHjFtxGXRdMfxNNTaoD8mmZ2ntPzbdv
6e42/wArIcxYTTTCBgpuELbLj9LgQzolMweTWon0ZX9mLZeF9642oSXhyIWMfdDg
yziXbNFr5sZC7s8n7wMdXCCTU1ATQi74nhPw2i24atGyuobzTk+hLa+qzBSQl+4S
W4cSkO9gsnrXXz8jZplQAHEasyO5tZ+H07X/yRfPOGxHDwc42omIi9tC2tPOD2tB
S6SxufzYO75dKw5wLmlYfF6M8fsjq9YcLA2GZECn5JvwaSHL2tfurf1PCqU49H9F
MUNmGSb3NzXlUOmciBDOXZVsKdTlmE9m37DjrYg2zf+yg+86FVg7bEJktwvuKoet
4/NX8a+wcLYvzaBGpFhnech3Xtu/QcHZqMuE19caUth7G/YDepQi21MBOa0zIqJo
vLx2s+3RQmd3xb0Ll60F5MopMz5mRJ+aamhrOPuN3xQHecQC8v6ADCRRpni/yWG5
zDBfj6Rm5h534fyRgtryLEcUjg2Lt7B7rLwLEX5LQufY93qmqJGjVsdZBfwwSR1J
+DpV0PjLrcGyVi1DkpsZHjoLdx4utptQRPtyXXsBkemtwu6BtDAVQ2Bv3mZjayHz
h8xC8g5lVoNVuL9sYQ9vhmj3+Q1jHk4yH3Uq65fB4tri95a5lDcqGAD8PoftL0Yj
5spuOl0ncDxl5/s5txCPdlGW0g7Ks6qvLpi2V86xiLwu3pf15k71FYshethke1tl
jqzv0Qj4mtLvio4RuaD3sKHU+cPZr1+YLW7vR0vaBxh+M9jEDT089LsFgeyQhrzt
Ozq8z9J4WTX/gWTNH0KwmvhxYCypZYaQiDPU01Lk0o5KzTvo4wTlaWhBR25yM6Ss
wad20uO8MYt/gNBoYVTVm1mTLOQEurAj2YkXkz7auymcCUAtf1ejf2i8BmRVrN4V
EnQX26o5WIQ9MoH1NIa/cMasqQUCDeCE98gCmyjKUgiotyLycLVCen0I0utLpUv5
07BLHmkBbUgcNf8IEx4M2R1GQtz3CIvi7kuLLAIWHFnLD/NzxTsPXaT+0bHBdHvg
zDOTKkHoMmnB8BxdRGMZTWNwHVZq7ndQUCPXhLTMihPGIs74ZZhUr8nt0IhCEsFN
IaBCkPPiMCa+eWbU4kcr+ceKOqaIqZyEDA7cgGpP+yjcAUTyYLoKgwDxCUu3wuqC
Du0hYE/h4svmx3DWy+DRDM9vy5DTATIZHDlNp+o3yIYGvzRQeKvewG3+goOf2G4m
s28XwX91GLeY03pAFYFlZTrYUdBp8x10Y8/HlvmgsCMzqqULGTPAD6wUeFHmsAjS
hJ/U/Kr/SegvgSV9XTn6iGQBQn08srnqXEiIQuWpHXRf7i4VxMsEP0kEHBx0Y4Gk
rQcbObgH0f89ieNX1yOtxtwUbGIahEVZYXcI9sgj162SQ6GtQIxMAJT8YBeMhWK9
NOo/y/YnalIBEbooQ2sWxCXHHGJ3MLSGTIbqMfJt4ymAfqJdPV+1zScM8JVaNoP1
N4ydT+GPOuIyTlBAj/g6LIOkAEjrAVa6cz3voxM2cMlAmYRldIKaRtkghA3D96ug
hAa6ukasdKGtjwa4B/XsyByQ/783RajICzqZDzbdWxTnPp9ECyTxVgOVLVgiG2x8
IxsY/2pC/2gYMfEBo8fpu3j0q/7qgTI4TLJu/L3cEss3MRACZ/xKu/KH+Y/HWURU
CrjY55bYboaOYt3CwPL+9U/6b1gqbXL02tzyc40W/G9YBZuEoEpowdtBbXVAGlrv
Tfv/nc4u7ye7OZgD1lr8gQwYmzBJL+p6/j0xfqfHF7XOFdScvhDYOJWBw7jv7utO
MCgQSMb5g1Es1t5vwIg+XHuz4nNRT4grUHRfhI+yxyjSMPgxQl1zTthN96wGsdYO
Nx8iiu7BxpkLeUnv7YoHw4SMX7gZ8SSmvxOUvBUnmxTlCvNft279UtizFICVDApR
b/JQAIjTVs5zv+UEVHC3xVvmE6POsIj9IYa01mvqArotk8LhJjBEvXqB8Kgfd3W1
2JDl74LRMREKe3U/+ooliIMgTD1q61Kn1XyFfT0yaid8z7t46qoTjj2+/aB8J10f
iFAq1MbaIFudWx2FMWBJPJEUzE5cpCQPu7FG62Euk5HoOQN4J44df75mZQ7HuAZA
3pY2WOVSNqLLUPqhcRRGI9B5QP1CiBWUodFOThG6UO9uAyBlx9bAkh15YyLle+yl
Pr7po5Q3tPeIEwzCnM+YIxTc1xvrHgAVoCqSFhY5HZgG2YspMoTdb5XXfFI+o5DF
MDHJwaEpWDCqSl/ArlesBogtd2Mpt2dveXpmqihv0Zk3r2FozphWWKbrU769SDev
0Vfh4xh0lYDIzFSmW5dS53tTvax0T6Lt8wTWDARBC6i2VmDPEIT0WtfqXO0ZeE0d
/UbIoqabYU2I678qtgpW7Q7NRwhzxDlEeN5eKqQT+E7AnKQAwAcI8R3SjGG3vzl6
W9MHRs2/RDZtcu8dOAeM3mzLCe4Zz88b06R4wBEsAhUxoVhqz7aMwthGrVNrr2Mg
cxswtnaTcXriruu5AMYh+y3RiJL40mKeTSbWVV7lUKdmd/Eff6kQLtvtCEnoJv1f
as3CfFqNajH8O0kBze+51GrY5S5mosTm65ymifyh661km07wKXReg8L1h/sBiWIW
GqC186D1y1Tl/1nkbQB2qexEZv9JMpq7o09E0AAJSE17uVlQdBXGCFJ4/9aTJ8Ck
3/419oKd0ltr92DP7GJxZgGU86se99BECEjK9poSoyYq/J4o6cwuMd3Dfgn4+9Jq
gvDtW/BP8qL57IAi5lRDbZMWOBJcztUkqu2n208jNv7D5sEjKnEjila6QdKpAXmq
wOw+wplu0CIO4aEa6inDyQTPGafrjhmqdU33R4zUgwhcUIel2PSn0vmccu2fA9Az
Gay6UfHImcS7QG0RqpX6y2msf5QYgVKynqhFj6OP6fikiDdw+I7xm9dze3WaKbkM
QwIe42/enuybpFGmnuVsHrCuOQhNkz6NAS7PTU10MAkNNiPDjrF87pQMPL1LEC9x
Bu+cXkQtuJ4L7+b4JuQWMDAVWg5FL7T6IhAbBGBJHlc5XZum3eBGbRB5YsC+rX61
eoZworsT9EcsJPTzlbwwBMIfOZTetFJAl76oU81t9E+mtEhol+aam13eMRW6QznN
30T8kef9EyTwl2y27Df+4XlXqHiPQjCUN8yeubvCQh4yF0z56sWZgZc8mnweCla/
broiuHytTi3FfSIW8KDamu0s+lc/AqvH2hCxsqc8Oyhz+zaKasi6l9vdnmGTg+I1
7fCC7Acs/IOCmXMWrEdfGSzGi8/aT9cesE0H3zV7NeEWNKlW8KdcqJYN+GRGgw37
L4ayjylcRGeJdRewMUYxJgR3iaTIWqaMRjR7T0HuTkjaE338diF6z2nyswYXmEuU
VLErBrL9FwxVrjWEH1HSSttxHR1SAXFRkodFGxM9WSTaOIW4xM+v+eAhhRJUZtUM
dhP/uyQa+kFcNiIS0SyGOU6LxbUDkpFeoP9o++dnTz62ywqZhtoyMCZqWp20GMpI
gXdXPXnNfc/GJjUL8GPE3dx7A5GT1uvjt/EmNQCf9U6Z4KPm8PcS+Yp6bH+6JfQU
u7aQi95pusqhKtDVJ5Tk9DHRW41SOoNTnxWNqSqO3wsNpeEtmxke78C3BFl9kee8
LCEm/SoYvu97Q1zDWmWkHreMdnlFC/1RI0LOmzCT/AOndFrPYmST6aUsDCA6FwxX
FYLURYNln+FXcvEBYYiCS+eARtgAa9oPPsjpwEZavmt483HnE3UXoWAQpca/yJZR
mjQIBTBXka7ob8nkKnFhuxR/o5zyB+hLADxv3jkzOkB7KiFML6jto5EK+6nLLTiX
iWHAQjh1avvf7afyS0zOF6vgoQjN4nmYi3xwYGpP4RD4N+Y5qpZMcdoH+ja/md7w
1pRgkRHv0JWQeQ/2KSoAY4CJtqns4VimeItturd3hRQwR1Gr6kqscRLQXcgKt1F0
hsiSU24qwAdA0HoNJS+JgHobCNfB28Cjs3bQPIWc1BjbevZ1K2cOOsGDiJfTb3fs
5qduLmtXytQalUmWcZbO1OQYIAsAOpzWIZ4mjTCZ6RY5puc3RSdwf6sHzAVNSvrG
tVMj+P/YESVcgSBXN77wXjOHWW1jM7Ol+C9OGX/9xSdVN3PMfi3e2zoI2ON4fpO5
nvAwFlIe36zuKyegn2NPuu/Dfrozvmm//lTHxbGT4gEImBvdrW5G2xsYpN8/qH15
qsCmjeT7C0aPC9xn9oHTimRNxCsYB2iLYEXWBrGty1zkXUwW6Iz9L00IyPR5dhRD
wN6IkGrRS5q4wJCY7aUY7rhgYMUPrWWgGwfYfoMWSc5ZEua8i00CAavwmP8JCJ+T
e0r0LWQOQBby6AQMDjkSxQjoRvNnJKpMrtb1wP2W8uW2JwpymgJ3i7qRYgpi49vF
mT9YzKulLO9QgmH7gDZGVegrnbFSpT366+s+CI38slvJh2kzU6nbMfZcu9jwgbD9
QosiMmRSivWKxrszh2nid58wM58BBNen1AvvDbW45HTROQsNGvbaTJ40f1T4Uzo+
JgKyTb16xGilI/Lzm6188NTJCcXfVyfi8bgAFcsN7NNk37G0IZTPrV1VF8BTd0R+
eFuyuB9PeYFzwSViBnu4uMjM8FgltIacfKrZBm6DV4mU7ftPhiZAfadWDfeG/7oP
y++iWgdrzMjnGEoGuocBKGWFn+9Ng5Vjh+u7cGZl9bwbrtfAi8EFTb3bo3PRUGv5
qATN9S5rf10GLInaBJ64akybGTihq29ZVNthGFjBO4WGFv2P1/V3MJAA47x7Ep2q
bNlhSGo5ttKmPBD8a/9ctjgsxM0UlA4UAJp4J1kYyBKhRM6GQFOY2YL7k0iKJ20T
6XE6JtZ9wLCzLqYPaRohGbDIdbPasvkI3sCbXePxoAfP+IVXV54xK2mHb32iRgbR
va2CuGMlcr13DPpWlvibICikZmmtehVqALr5I9eVhT9sg1f6SE/AHMD16ds7CFCu
yUrAGZbmNS+S0N/UUxWppEDL7OsVx6Ve6HZqKNuHu0K2LoQL3sIluPtdo3Tk8zwd
dY5zsdC2T5Y38U3jA6836B+M2shFn24LT5nhrNucpaHakw8p5FXiC1rNZ2VN88mg
kbHKH8f05BDy9/5Z3rVhJEuWKSETRdMqkRiKzlGYvO83lEKgEf+NwlZQC8+PHg6S
9YvC0p8uR+2ZBGXSMH9n8w5QtFB+xc3Zl5AgiPNO5jrmM4aOV6SD1vlctmRXnOP/
rFpOxPu3Lu2OJuwdwUIJt+3DIwribsqqUFY9Txv+LzvvGH6tX9G7EdU7bV2iQJNc
J7ZUIXYntaNYuf+UErCyPIJ6mRToYRtu6wr5c8Y41+M1lXprp2IF+FOy+/JWNBoa
8mYYGLWWq9dMq5R726WdfhtDkXIdv52TQxlSuzeHpTf4N5ciZVwzqX22XD0UFhaI
ii6NcHgVNc0ywDpcoJ4L1ng34paZgerjVWqHjMzrfg4AEZIkBE1rNSamfV0WUT2Q
RamsVxqim7b02Y2s5lvhZkx46PUVZGIJ1ZNsK5FK36Z9vl8Eook9JRLqGaxJ0DYn
pdaZ1BetLuC3cSwVKBnEeKZ/+xWO0XGwNC0Z4/C77qrtJ0Rk35BKTc/fA6rL6Qz8
KWh1SbPw5g8Fl3X8J2bwFHNi3YVT20Bc8KvaAIgOn3DGy98UQVxa7oXWT+8YQPJy
GBzehcCfNTbjzwM+Q1htRXs2POk0974RchfYyUFbi9TkrjDf9cLWXnvpWDgWoTEp
/CpcISYeiUxK+ANby61maEg/Btv/YwKWwP4PTiuZnY7UVo+Kx8X3fxO0KM+TkiBh
FiIv1Nw7/A75kQJJKkUGTTyyK+PSEqeOEmRV1txYCbvO2aMcDAytVYE3FxmIuTg/
9pL0zgJ2TbVNuZHQjkV5PsfpsVTu7rcwGvHq+mpOQHcK2AOShMNcDngKeKZD5el7
NzWQEPjbtebj/M3BNNlZvqkFinWO4kp4l5QvWrJPvidH0MgANQD39RDvjEGx1rjQ
eF43J6p/KcoJQd8DZRu89dJAKn8MFJRem5+Iqa6dTmHsyZHcvhPvItyXW1oNPoJ2
DiJJ1D8p/Iu5cV3txvA0h4cLT3iNb96OcjxpXyeb0GlDkhYKo/Fx4LRz4pyI74qq
wcWQWpBZsvVBF/lOH5EbAC23b/KRUc7/eYKw6bK0hTqYiznZqqngAXNxEa6mgmtF
gvRHgfSGpMA5/7CCAFHs3ilQc47pmloV77foN1kUTCyihkMIAQ1VCGNi49awNweJ
ph2r247Ez+khhH6NwR/5aV2NNKlW1BR1/Jn6C3pe8K3y/R5PDOFf6LLyuXsAuQlV
RLppqqHtgkNfSsfBhEgWi9H6iCvSFBw+ahbwARuakmmG49+bx1dBkKQFW/W3or+B
QCYq+H+tWbaamE7hnxMmoSKDOsJg9QbaNqxyXBjnE62TNifAAxOy9MnQLHlRnmRo
U8LHDxyMQ4EtQCYquBc39RkDsavw56PYN+SHHUs4vtSmjBKoSHR3+Jhn21hPzWZw
NxatuG1EjULu41xLJhiEKi1chjvHOnKY9ZHOpxZAC5AuQ+3gvOZYDsIS3ao1nZcD
b78yQ1GRcajjw4Lp1zjS0fP2ynvP4k6sAHsGVpU9e38I/xLd9RU54tbNQZ0hb4iI
k3CbvsytOVcN+j6WXnx10TwMZSNKs7wDTR6iremxqfTkiAM/4DcR0fJAp3PdoBya
IghG2uTZ7FM7GGCXpjmRQGGhZyEhiphsKyeQoSjGHcz5iVZmYuQkVpXp9WMAVjia
MWq+bOYBKPt2I0r1B06QRxqaU/LevLVo/rZ7ZYAL9xAvQYgTAXlqYnYY6sCJCfYy
v4qB5Tm6GOVy3dF9A8fI/2+PAzMmsUUKulIqu3pr4YGTa/jGBRHlvIPZPdDWIQzb
/eiW0HQmDgtE3MiSaZR7g8mnq+wIl3Yj+xL0XKxvsQBRVSPzNHj+jy23ZcUm/aF4
q6zrZepDoJcr8ejLPUR9Pn0mT9CE07lV6Q2lITRXiOcsgjl6ENObuvH8BO1v6mBn
+wv2Er3+scFpduTgvB/h2wRVXMPD2Sus8EizplU5Jctyy2UMhsENZZmd3lIKM8rl
xzCf5TQWbaGszFSboGTmzAAvtOsxyNULxs3mHu28trdKA1yWiFxcqlr4tfZL2WLM
lDDQaKfCm/WvEkgiNCkPsrPnS+9LAtdI1YbOpOFpfxv1W9QtiTVHMBdctLkJhKRF
Nty8saRXqTLeFQn4OQPEnbfflVC5IqMJUB1frMyrohb490kFggZYq6pTL6Nj6KuK
K1LyTeNaDLsp9lZJYywVZAw1qrYOlXAc66QuR4S4P54wLyFn/k2bPVFJdju+FdJG
h7Vbk+p0kWUgLDxzuO+4pXiRPxI6Y9axTbwDQ2RaQfwZgBnK5H+gM6q6nX7wuCaw
Qj4r26YXW5rWBda5MtKCM4zKLiVtlHe1B/enlRy7xK+Z5C15uzdnRY2zTocyfLfm
WN1apLkDrAav5KtB7ml6CO1HGG1ZVMyro+cYds3dS5X9bQXTxd69JDZ+hVwEGGi1
SfUk3hSZVkybP4ozN1/kqUyGK/zPxZ8p3MedQkfHtNRepgOonRGa7e7Gi781STZu
Vq24jX57RgZzTVxWDsTN6wD0D0eTzqJOux5K+SSjiJNN4BZIVe42LPhcWF3v2PrL
WEZNZCgP7u6uPXhlDm/bIgv5hj/yecgYAlTwU/WZnKcw1XonQSdfKyeEkPOrbonI
7Ra+rHMnl5+3UnvQNo9M19FVCOORJU9JNQwiaamttq1FrtwVCIxrsvjq75/o6oQ2
CyO50KzexyeK+c5enUMZlU4j8KhgkM5Z5appcUMgIhDDL8mRijK/u9tpQWB31DjU
bfb4il7TYJ9yzxqYnHY9876X28wJjpBrhtUQqj4drBNq2QeC9ehIUr43qJcal34C
qep2nLcrBvyqkfuuxifmlc0OKyR31dUcls4pvkgaly44K+swb0Uqbn7I9/e05WOA
W4Ox304mvBvFTMeCbbMrpoVz9Rx3Lf8m0qJzYi3C3EYdSRCi8KyEQFVl+ru2Hh1H
0InIVLwj8mVHpWVqh/rUN8YgAsdroWWMZErbLlaowf32E1tzVrYJFOo3KDTu30k3
a6rzyg8YNUcNJtYR7mQdT1iLTxZtyyJcpq71VxVZNdwPHFhmmpcwWWp2UThtd2Ad
mhcTi/omYDprB8i5hVyWiroEVKHaUEKN2dH71YyJF3AzMjKnduDAmjuwIDfEIBvV
DSaDbaqHOJyTlTCg/13pPsQE7koPvg+ZbGnmQ8Kvl+3FB9SwkJ6PHJZUT8jH9Oxv
sGSM5wU6NDovTJL3b5GW1riO3P8sjnNkPJwdxvtuw61l2HdjGEVhc8LtHPHiZHtO
kJFIw/2qgf0E50pUVdHptaBnv27zLcS7zHJNVFBOpWHsHo+FhcxGAfYhKtXPq6gD
Go4TqFYngYYjy9/vsHMIY6W+T7nrbxZJmGb1RVE5uxMomSC5wB0fZbWsVAEpXNlh
kEcQxd85G3jXtD8ybQ+Wc23oORz6RnOADCLG9pGiK/hCeyXR1u7O5RJVnNVbBTyb
shJFR/M/U2v60Adnq1Hib2ncteyGjC8HBSKDDSV/2zdziyQ27VDxqZ/hnIIb8qtC
bRKb1uhhCtILSWDvDrWzJLrra7HvRtpfaWdIeaaQC/KBUWiu9qXkqxIAOO+CARw1
oGKoBsPzZEbeveYgbuiFjN5HRfS20v0l0S7AE9m1iB+uSokHF9aVjm1Qu35SHhky
UlNSlltTraRn2dmxGPIJyPDJ6uA3HfZ84QlxMxL1mQOPjDTeBjn7kWbNVrBe56gc
mrtkII2cPbgYk2HnQDwj4RVnoy7PzUpvYSPEXyP8RtX51DYFAwQteegQHHtp9pBZ
tOAo++Hev02b7mRv5TK9X2zQAxE+nE+cJ1YDTl1JRnPS6b3/pG+IJn+kUJTXFtsO
0BqF/AN2f/F4Nt+VmQtfBwJaoony/5iGz/3hNWeSuG+RYSa3fdADFhIv4x/fkBdk
p6DS/UWSTUUNSHaMF2epiPLJInjeUcYXYfv2quGSwaIXLO/EmkuWc6c+IwHNUZ3U
ta+K7D2wVrObaGph3NIkIhO75a3ufK1O6miB3GwwLc/KrwdbG9uN003uhWKXb7W5
p2RX5xtqwNSQ8yQKBJNcrXP/TnfFrhhE725ZwxgVhVIoIaWEgZ4Zhklze0Wg4Ibi
zImNc3h2kErn1GxVl2Xnk11oJzvAk+2JXjpNHZelsbpr/YOWAjBsdv9PMNftckbh
MVHghWqymReeQp/2BZ8FOvh8tBcG5VOtzhfe7hPDv2ni39iNqKVBXO6uMW0RXeR7
rZNQBjTBF1cgHwyf6i1dACxuc/Y/F10tHF5rb3YVRiZkCPmS4frZz9G88yXPLX9a
Kv026ypAjHv6yPdoQ/F6JG8pq092Vg0bTdP/POmTo44k5HVKcy0eGx8e1MMk3aMg
VJi5/+zHnhtBlGO6WxOvIOeKrcBhZyT0E1V2da/jCjL//DE3WV4pC9GQFjSpJCmE
LXy6BcS+KRtMOsaRMEBfrL97IENE2klaMJ8P1t4HRIQK8pksD4VkA7VCKt+tQPXs
3IZMQZtTTY9ce0aOUpj3vnyv/NZS5ayTg2qSCy6micgwWLmWbXZ9+tMD/Hc/PGvJ
KoHuDbcdughKPyabP6ZpNoE1AxD+JFat+VjjWpNB/Q8HUCIQWqyl894rP6uWOun/
7m2JhsqzulekXn1yUnpvqKgXy9oZLwGWVWoM8uX2z+4wcn/X9cCXunCMJjOx1tHq
EEKcl9ysD23zmoSru/PAdnLYJF2DrCNmUoADDpveXqHFZ7+dryHN0cTfBFYQ7nG+
EBM2vN5VSiTbp4FeSt1rjyvo9clyXG14g5dFgMKjU8NbFtAEJCHc0B/0i+f5Lrd4
X9Q7C4EPs/hNRWZ1TZhWjruHzSfGk9Ucc2dMr3XpBnbuSBeWSu0HyRyVpZ7awexK
yYLSfIaojr5BWFCbCnC6C3sZN0OKR6Yf1uPQX2XUZRYWghQ/LuAHTZtd/3+zVsS4
SwOEflljRHDKk+TQUI2NPKsAcV63HCCjOyfzj2GDZdChmvmo/8ct4O9rm1kyTYMA
mwi6uqmCgcJIIzY8+7ErRs+uRjKe4Lyq3h+JMGsDWLozv66SlNm16G59nPUEvAoh
ft59UG7SOka598k2MkrDfhimD9CttJB/GHyKjXH8eJS7HlNgnQvj18VxIMURlrBA
ydsxbr8NXLCP0SSXEuFiTkdxNqFi2ktzDaHkluAJvpPcI9NSG6HPGemcPLRulWve
JVSq0cS+rjv2R2o7G1DmBejhG4dksK2i+DpQZK8hLIft1WftGfcPxO6bafeRsuS5
MT5e1mrj9y5n7/DysKphB6kreysNMGJMrEDsKvosBxz5M96tpu7LpZlawcx4gGxG
19hlHu4c1wUFpd5aTDVkQw3eM6JpD8mINH0jYHJx8KWjB21AD5FsHqk14z9MQbL+
dHgf71sG2mH3bdNRnWhsLt6kwuie2L1n7Vjjrte1XyGSKuYrJcDnOdQ4HcSEd5y/
jQTrMXJAuEItVDEuqIK7j0g+akibkbt6xKVPXLQiLzCGsAZ3lPrWtIFd4u+uRF7b
XfdOp3dCDwbjGpk/NuQp1ERN5co8i+pRtjOl/fWHCAnvxRo6ah5w5XKQ63vma0Mn
1sWDH9Srng8pjimVNFEXBFXnQ7uDG1hyERO1kbYsIaP7Z1UtoCWkCe/Y4qGI+TSM
Sx/zN0NPpz2xiG9Qlf5Ha52z5vsCcEkYLqe71oKc5TuyFb07bauUH2MO1q+3Y/kj
aL+liYISy3xXdPiaaBpbPSjA3f5lMrU/KFlAmonhr62BAmcpdcB8FMZYzlUbOYmd
t0Zet20s1cZF+gVr48a01iWQzwXgbS8MiHGA/OAezpx0izjiYeam5Ooyh48POGeS
dgLcYYQO/LcUjfTq3FliXVK+SICTDjF+ebRZBBj5jXD6kKUzOqD2nP4uEAdH4JWJ
xE/IC6PIDdRD0X+hFKa0OMyTMh0x92CopBx8xkOzgSbfSao00yyYeQcnDP35jwYw
QAqATOenFu7Rv8n00YsSDbPI/s4IQUxxR2phLbHnxrLKYxHNZQWptfmkS8WbpZ1W
qV1lY0vaSdBPIevBH9ysvUKrx0Gwx2WImHY0PIfpgeBcCf+mg/hMgFjoyjIEz/b1
6RJB0NNrHarK3KbjmXxbav1pJinbmykNG2y2NQchSwHFea/B0lJrYgg5nb8+YGDr
rlYonPeQJDDGYGcQN23avSLEXjlDWHcJvsz19Z4AwjhhvB51gTP3PtTmUfH5Y0hA
X9ZPyonYiSPDj6lCQvEoE5xs/v9a5rGiKzOBmrAf/fe7raUZ+WI2Eviv5Ysd68Is
o55RdiSLdjfgjcmPNU4RIkUq1OVX/CrzVJw1U8rre7lIL0GxkQ1ujEsAiezuPxQB
j0QyEUq+0WtLb3JXOCm/jyNy4RAcDCELOh4bl2im8TowT51q3XoDHa8ZEGoLzWtX
tLlcuhywkIkU91qPpqrIUxKiPO+VCNqJbSJ7Fk6jGp6yyH7qIWjNzCUKXuihkUKN
U7Wo3Skp0mMeQmm/nN7SDdi286jFtAxOPxbRduL5noI1fvauW+Fygu0fOVhaXMVk
eMWkqZWhmnVPLxHWhg6dM/2AiGnCJ++cSreD/coIjQ2EPY6sKcKjyYj8U7jU/zx6
ErlPD5RioDTb0QFVccvXke25wfSulX4GXoVC03ue47rfGAa78FL0uTGZB2RPHOAk
a4QQ2WfhsZTN9k3B28z7ntU5VXhmjguV/VSKxv6fg/okx1G4yJNjbJOEhfytTGtI
XVNOI5ikU4PqOFaQVFP6mEwJPNY0e9ghfDs5yhRxYCTQHNQp13u/BxUMKEIbC7x/
H/JaEPCvqJg2EujPPDVEiMRZfa8v69X+CvQ+VNz069xIDOLqYrDP4QXh96Eg3rZZ
SSl99sNF9LtUjzPRvifsZxPn2LZz/sZOVZAx41LqrCd2iOEHFaVmr+fI3uNXOhH8
8yUp/curvpEyN4AX/ulpxcg+ido1nhmNJnvDhp896krNjD0+2KTOdTRIkVZxOXuE
seWbSwBuNDhq2F+Cys5ydda4xvraDfFdIOazIddLS9MdHw++w6jNeWk6waaGMnaa
VX+j9puFDmQmME3XZHHNd4iEDufUQV91GgAPlaYI96pfOThmiUaoLA7ZZ69sPcck
8eTCOmvCzNrimz9WZFpAN7Hax1ZDFOX8XxxavjwAKf8nTMdymrrLVLDU9nNnLw0J
UiHN5Lzwni8cgzGbR1MsLDHu2dH6Q0/2+uXAhM4bAaov5QkOp7NCckBG2C/e/pk+
/dOzGPx+qM9Qz2w9VrE4DA8XNC8LI/6FBuLX/HxXjXMDRX3m2jS5qBsnw2m9pgbO
2yFvWTozTGkWr8mPQARXJfXBw1mN/8rAZ5uMZy3lhJNagKOzoIt0HHKFE28HtfqF
HL3fNNDkd+FndnFQsqbMadSSE9nXhfIqUdt8zBKv68LptLqUmNvpx9P6oNkFxokq
nRqTMgWcIUmre6sTEElsJmIeUrjib31d7DmDcLSptJh6EL3WxL3yhiMTA8lpS9yz
9EMZsEA4ivIXtmjM7ofnfYdacb5M/f7kv184Lz0/6839roEv0M4820JQ9AbTvYhH
fUTOiQLrKdhz2jAvl7JV9VhROxHWbAX1/9hoQ9ybJbkB2zAyJ60WHQdQygGGh6x7
zAo9ErjREc3xDgCKjH5bx6NBLS5bxjwzV/ragjS9qSURAXW9E4S32ITknXt7342f
hIeMdE483BpyDWLOFTMysuch3ojybm1YDYhNDODI4MGvrOe8ZiO9LselaPrLX6xy
E9y9HCm15zRCaJTYlOj5kX4Kf+U8Fm8ENNX/uTNrF2fDJWcSHaPL8fcRxUohvx30
kSbSC19bGDb5sa8eglX67mp4cno/w64trUH+LfKY+BGyTwBpYZjrLMmvMtRYWVEi
/9CyUgHi7uEZRPbyajfOEjRL1ax0WZJIJaiM2l2WeieiPwXdnw+f3Q36yJ+i16MI
XZN7grI0/ZNN4AexfiG75ysPotsn0o/2p3ZfHbbxDZnYG1tokcG036nKeSE3BKHS
oEK6uGIf1mALX9NNv+aVmDdaevGhkXZh3B86VHGq+/uYKIo3w/4dFicy8caAasLq
RGkjj29HAUh30aA9HqbtbViNSrl941rwN+FaYH76kr34R9+ljplOHXZilIdiz93s
ppbf911itQfzjXd5S2qeafKGjJ28hEZ/Rb67UjZhneueQ6h1kBOcubZ6ox3EOVSh
GCUtX9Ryr1WTQadqRVdxieov3irEw5/dvijkEBwzW28cjsRy5jN6pVjjKH9rBJDW
WL3edrkJi6n4vVgphxNeXza+bBmOSe+bKd1WIwFZlWrwtP+8JGzcltoz5g0Ofryi
+7zM6weD2sXWZFBnWWFhnZTtC24i78cXbenCFCdjlVltTCXc541ndZx9dYmy6Hdk
SDZLWAQuSUsST0NII12CFGHYaExfpqlA27mrXR651V+01GmETMvvg+HEXdvIjXA9
Ld3nX5131AusVq0Q0KDRvcUxyeGxAQkOo/dcaj8cclCkUpcSYAUoqpZuFkOoXn/y
ihLK78p3Q0d4nvvZCzcEHu/jMpZFllBhU9ZI9Vqi/Ws9KHad8WPcFArZH5L/G8qF
gfVbukRfWw3jrea7jPosrg/mcM/apnhayoVTa5frXe1weYLeIGmxDQk77RQq2QzG
PlMdlRxqM+GRmb0ZCg/nkkhHzXhUylYGX1+Lc+GP0+BlfvZCX5MxlwzXg+1j/ZbT
sHh055xGLdq1IH0Wvjq4rJDo80v7iF917U79xBI04z3RIACMtITycFv6xl64M84j
qgiaVXDU4KAT/lPhBL2TZyW5zLXHIzjYaK5eEao/nM5U560n2GoH6C2JaDvTqNhR
VxaWB4Phn1izHKbEe6VH0sLWzFI8Wq1TcHZ5kSuHMxL8GmiKc/iz8OogHMIkl0uh
DLQYO/ov5Rx95yFWpHc0i2REf/++dXFo4P5Wo9VWeEjeu3YonVSSf/XEQGxT80GI
iM3XkRmnuYS0OMdZknpPw5YpySQTv1nH27FVPDEO4/K6NdObkAkAAw767dqjbAL2
T+vEAM5/F+uT8GN/VG5yQkUZZxrclE6Ooj1jBcRDg0OHnk9s87w9g7ofZ/D0E7GO
+9MzJIXWJxjTWZJhpjriREIkeRovGTVZUc/03MU0jifbxpJVodo6iWpu8X5B98QA
oJg4tlh+8TpBajSFugL060RydEA2qaaN6PCK1eKF15QANz7DOu0yq6UiAQq+OuZs
zs7CJM6/Noc8gX1s5WEKhla1qAgJPHTqxBKG2b593Str2o3NAH3JO008wTGp1Q9P
GGvTitpoSoK1lC5R5gTtK0FjdHRJHw+x9jyDQj2jT2+iB3pWIK3E8ZJUbCJjjQDI
ZbbxFtTw7t1FfXGf0kdz6FGexwWll8kYhupI7CtzjxqzFJIDVWo1jSBhBqyGQuuy
xfiRe+6Wzq2vVp7zMF/K4RSPraBFquFhocn4Ld/jLN7fM4etRgbw23rVCLfNU1yH
DJMyXkubF3yvG+eTZDZaSM52dq9APCcvQ+PfOR2ID5e8AUkX1lhBcSB8t+sQsiAe
Xb2J1mzQ4lAEI06at8nHFVBY+JkGdrEmrDe5yuAyH4JltStik8dWghQ2tQEUVT1A
vODBS+jk2hSjTca6LXOlzhN1lQjoevVRdChmm78ZqUF7N+ryHRUp2TvcdYsra30y
euWZu/yYyABtX+EQyd19vWaifKYyKuqTKegfGcSlBRObSO6G5F6e7waBrkRiVe29
HnAmMo+0Id0l2LEDGPYyu4mBbbKxP9LJR2hi6tuFW8Cwt0uR/ecDsSlQ4sD+fAzL
PFfNEYLXD/OeaPXM3VypjCV3dMCo42jxf/1mUyyi6bl9ltap7PbNo8990a/fyCdP
6SQDbHqWQj6levcrBpttTVZOIL/CMKg8u05lrjs/2rF2bL7EfBAaI6s7KQ2EbOnU
iBMfyv+Y8QMbLPZXNSwGu5jPKjJW81M5Rw4SD2poOdjDZKfhXnk8XhVq/MvqBSda
ajWIkgiXvQYjEOIGEPwsKuIuwTQpULsk1g2D0XCWh/B0um/YjGlO6smE6D06yDW1
zafM2he4tlV+nzm3Gs6Hy/dmZcRXXlM1UIkcA5TP2wwPr3Bv24BTYg1unssHyGLU
0FfBthNCxKFI/OPiPH8hAntXO6jm4zyAfQ5/O1FuPkd89ZjuhcRigUFVeu5PiwTx
OTbfzLVy6dumjPXVTj0xHeOJs70MxzG+01PdWlWFcR9w+D+Fe/TP354qWUEvU/GF
7dJznJ3C5j5lU9lz/+fUM6HU7i6k79eXzZroPUwvqVQ2CUiDWAs2I1V6gXYY/RwC
jKpH+FuyKbeFZhrnU9FRVXZq9xXOGJvt+N/3n+QvJV+PyEuW1HCnvQZVCVWnuEdD
KldTvznS/w+bsTr/oH+dDnpGbCs/dhsiwK8mJAucFNJTugg8KukDx01CAIdE9gvA
BClyeNUzW200xce6eeH41eqvS7krYE8VYXjzsDZrEGUqzdu2rF29hieXGy0psb9S
+wSrXZm/H7PUfV2NASCW7mGBEikzWyAufGxjctecOLWSlzPHyTK8KnzLN1H60YtM
kYasQvMTIo3PK5rwW9Zcq3i1EGXbc4KEZfc9iLiRhnl+lxsskpkr1FQhhumqrwx/
ERXmo58/Yk/GC8RTVs+8WApeHxsOBdr5QPEuarV8z01wc3KcxwZMn83/VHtcIzvG
vaqF8bFdUgMxMLF72nXtJYwT8nhZa7S19k6UYFqz/6dYsllhjILHkaV1DJbrX8Bn
FZy7LR2wauuqEAtd/TrhDi/omSECy57SWd/q+4dlWbKI92I7UX+ZAqdlarNCxtdk
ZSHVC0graoXS8+8DsnPbmomuIiQO4Rv1i6RL0x88/gqpi9kbYE7rF9ZokbxNjefq
AU0NPR6urPdcFiUpb5zX3mOo2oxWvFJJnKGOsNU5vfj+qQbmx6BeFwcyQFMwxskl
GrDZjKYHW2T+Q8iec0ylAL2kVRGBo7QJ0GCyRxFigF97eiolY0k/C133DZrB+pB4
/CPnxCLQJHfqdclQUMv/iDPlWbwswehN2NznqHCkYxsQbgZzhsPvCefeWK1wOkkO
IRKff+onU2b/qih6MMMB79O/MaJ7bkIoLuhZAMQca2nE7oAo9iqrdtAT8tdnAAyd
LJkdelgk+JgKktOri+lvcWkXErMcdiUCHFbpm8C1olBEDALHV/3FbUQgvm8bKUs6
R7/YKdmyeFBO1AObzWI7j3eG2xqWtCg6j+Yc4WiETjszfN/JiEd/T9XheXbNqw48
/0WAVe4H5v5/fox7t+QNg54CIBkN5zxFWrL71jQpnFkyYOH94h14gYP6HKstClDc
lkcWMsov3o9usloX3iyPuNyrBkfd5clz7s5bKBxlzI0XPJ7iLakG5tFErQ9lKhvQ
N0flaz1YDOfmz4hx060pO10G6ACJpV+CAzlDhUWE9hOT8JKSe3FZTkcnJzjEApVH
P6xf4P+XvrpL7yOZgiAx2bztTZ1pmXzkhBSmXmn4rqFU9xsPpruwQTsY/tveuVHH
FXVdKq9KUDFMwPTGOeb0lh+1gdlWl2oUYj1hmtvKUlcXOnPFlxWFDc0K4Vnsgiap
Wb38RtjrSKRvh+hi1jwRSQUwUYsLGYeVBI7scnRBkeE30m08uQCUdvfytGrftvAq
3Pvu3SWnWIDBMhKNqlTWnRYQQCQzaVy/k1iKsu/lT2haayxcVafxUGwCuPGneuXi
kMKyXANCWf1pcLShzZvxSn4FktHURJu2R3MSlpN697zep8sTa1q31A8PLjZ7uf7y
J8UBmcabsghFjq2cvxkhvJ5CsqLqSivWf/YyTN/5xRJUw9OsSMuGE6kpa5R5wRnV
XXk7Z91V/m3MljSac/3fierUcUstQ8V1kSS08hmdTloGjWAo2IMyYxvwj81uQZyE
gk1ZUBa+3JwYL5kMZAeygDHly3Q+u0Tm+Zm8u1G17xCchmuGICSSn84LSUH53uWV
lYm0VasunuU/+Iy0wAr1hWc3HYUWUb6dW74oFJw2RD0pjEynlmY5CIIDVrxK6Dhs
p87DlRONl+CCtBcoThVHfDPUix6KXlRg35czVD5OC2WEvkWgobSckuURbnMY4TvZ
eTntdlHYVc6/uVyoIddBGP1xzL/FSXlvBDkInYbGonBzgT7jbsZ1iiIPsIJkrKRo
VgFCmU7XC/VJO6M/+9SKaSWLFmiJl+gHtkOJ2EqERBpNZI2jbS4M6N1L4IjoFdp0
pa4tlVshDSaMIkdZ8CYYu9D8z/1xDdn50TKIgCHpWNzITMPWjioJflTxZXreQJUV
0rCrLfDcsz/y/5wZf8a+PQXDLi4soI1TIcb2L3QQxi7XkOzFfb5W0iSniXrVhfEn
+1BYikULLXnXYV8fyixzXhc08cJu0/KLJ8GODj2Lp6JAcPORbZD/9odm+foO6xq5
btt8gIznVubbaaOYhYMZ3jpL6NeSIqoskgqAWPOZTuGzsX3EVXEq8x1aUNGZ9n4i
YtqK5IvHeU1Ds8PB94SOCIVIbG9FZQZmyNi3p/Y65DnalzrfYtissRZTiDbNfwtZ
gjaap3yprJtkhEEeE3yVIbscRoGbfdHmQu1HFIaJYInXq8Bc6+Qdh8TMUIBGs/n6
65uI+0WOSXRkkn1+S35NhJQGtBkRYy/dVxLpfGHRpz1C8XxPMgbn+XrU73P4MPnG
13vFwOs9GVmJ5xQKIfipklAoj4ISzfPHt7WtlEOQWt1HUD+7X0uvnkFqgjtr1tAz
aHyJMVW+C4pk3iq1c8zPohsvBwE0e6gqx468R71yAQsS1Bo8+ZTpVYQAk2eOQ+fX
3rYzElurszwMdOAblQ5EtadFuEf1kKYC78bNgUii7BOu8XTzMOD1YDV5BgzS27t8
rPF3/W4X5SsCXCfMUTb9ILpdAB37yGQ2qXdyGlFA8N7HirpMe9dyCKwgNC2HdAcz
k/JKm7LhUEQ+9hYPYfwiWrBauShlGxhdOXpmGX3oAy1yEI7ajrsJDd6/ieOT2bv0
SfvjUcLWrFlZC7pGH4ZVQK/EQUCUeBALOM2UErIxH4Z6XD2ZGGw0gouyLXdl90RU
Gd5wjB2cfEMK4W/1x+3kYprl2NkAvuR8IpE41MAE473w+kXCUkwC7LWfRX+Fjn4N
qMV08Ixk66qgHt5LfvTqC3WM5xGl9Nb8EMbJkngq6ntANNlBNc0uPTgQd6Ndbuby
jAtCB98/1f7sKnX0lBhqHsRUpwdl/6K8xv2PBO/nIe9yNLXbO/3P6DTq8N7N+bx+
HGLkRcpf07rGzFE73mnqoHZCIme8Eww87x4jq0rgx8pksRE1TVtg4BLch7o3/MFV
ANHhGoxkriGD1HL8plgybgSXe6CklOJ6JRNPosE2NPlSJOJSVlLPgez0oE/3gn3w
jGi9hTKQ9ImO2Mhdza/i2Iiq5oLg/JaYcQeUQ1dSA/gvPOfzTa3OCf/D5SbYii6t
wyJ3OlhRlgDvx+d1HdTs/hOiJK4jLyvKBek+r/y8j0GP7tUULJb1MhjyPOaSAIxG
l4wA8yhyq3CQGFAq/d75qmas7GGODMI8tYF9r1arR7Io61p/9cuVBYnnF/w8IhZU
GoRDX3GuVnGD3RnNdInePJuxH/ntZTb/I22L3wfpe2lodfSp1uOcNrM3o55ylilm
0HtK5awwGYG0Zazp5YhUrDnn7ptlLd59ZdzIrVj3v5G1NH0MI5TfSRpy0RXhESn3
tw0LCwiiRha/b4DV/Rm0KVu1y93BRQbkmCy6dWSysTl8bBeKeSXI2Xo0O2YOS4a+
hTe0mZOQumB40rSU5rvUpuLk71/ENF+8eqPcvTkJX30NX4o+mOdrMaGVFEcPD2Gm
emn5dcuw/vJ3m0lF1UOqUHGhgR8m9JxNo+Dc61jiBCf/OXaUp1r0eM/9s1TaZgP3
/B2J530iFU7X1SisFAVPnWqppjfOkamIXUrbYGAO+ECstWk6nJwn5PQCJ+ODMT6e
H+OUZRxwSjv9rSzA21iZ2aRNrHk3i4SSm9kP4vqvTHj5TkPGEOsQC3LabYekNnUE
XiMcRgUqH0wrkY/TfE6nUr8hYLGLVA5fLzw5LaYDbQDI0fvkGa9hnvZTg6tV+q5n
Xer4ifOCLHxlOejsfCe/a0hmxXLvBLdbEftMjkb0EzI2xQX4pfi0UM43DZX1TLdB
Dykco7MLUOH7YuBQe3MMZiI/KZgf4Rl+NBo6f9Sg4XFi3Wmcs+clh2Lz/JP9SHPG
qzRYGYlw3NVcObVbiEmzZMg8CRRCTqCekYEpjxvgS5SLcNbBt4apTDKBLQO0l7MS
cy4lMY0S/pLL5x9Ey1S5EsOymS+wfjtiqeI30GnH4aPEg5jDG4ccDO9bgiwEa5G0
JhcyP+2Izf4uRMp7DoSVOR+MRdQ5cNb7ys+bHIsMY8DaUGDh8Z5MYCgyisvSsVkp
oJ6SXXoJs/oc9F4uFC/RzwzeP/r70BTTHCnbhaKZtoc0rHsL96lTnnxx+CvnS0r0
s/r55fZBOxnrP3SkhN6UfO6u6s2H3M3qq3AqvtnT7YX8QpffsN0dIvxLHuxMY+vy
6AaxculZEyJ9WGAaWFke+iAWahN26YAC7R/hlAA30XQlPLjFsT5Kt0bwIjqlmLrZ
Yc/B0IZxEV/lILwszaSVhN7Cai4YzzbNWLY0ChftrFItKJWxy821N+uZK5A1dVsK
L6K2tGSzJUAFuRXtQSouk9+0occuwoRsYkq4b+Hiqdm5QtbbfAMKzfD/XOE03BUh
rIi1OIoCYz3I34yJdi7/gvkQIwB6BhPKHZAQnDieItApWi9kJY2I1Am+V09pDpNI
LnxgDFxEbbkZlQV6PHGMgeJjWbhv8Ajr9gOPewb4KXLVjvOuht2H4z6C2Z3sRt2I
wNE75A5ShqUrJ7bOQfCc2Cq+4RpFaBk2vRvRtXKOyGflrjVlR6SJCy1SolLJXQ/8
krEZkEo421aH55I0OXfyMKwLlAQjpwbFjmcAzCIIF2dBQ0/NvTTBib8f0gl//IrM
ce6+QWYbCRQNrnDQ6la+tt/XcO+/6JytOWN/rD6rFihLv7Lbh9UpU0C8NAvaxIW5
mZ9Edc7JQWgEiVPjozHW8V01IgNUJc7LsmMlkOOTYtQqvcFprYgcY2k/NWFiVUMP
SKcALuEPQxb1m2lXguRGxM784yxfS2BDpG9Nt9DzcoXRRGlSmO1eJgEXjv70Dbeh
/1IOaRX0py5pdt/YUPMRXLvypYTLrtq3ymNHUgfnP9Zs17t1J8+eH3XvPjxOogkC
8L57F+HXOzdiPl8p7Kb/r7LfvKDeQvVuTOuD+E6q/RDtH6QknnSF9dczxknG1KSy
Upi7LOKqGma6SZWVNoKoJ03NiKywxEFWurT64AKH3qvVpqUkwpTnYFKil5SqLRpx
f1zh8ptXDmN/Iri3p1DF5+c09/aRMgDG62fl882yvBdVjf3msYEvdkPs5F9F6M3m
FUPhA76+mEy8b9TYDRBdZY8iJ93TvXZ2aXPyadbABzVrBn81FJFvSCeU2JwHiVuy
2H3/WBYFld3YAj6xFSnQCnNNxIM/26uvG/1N0gBfLWcPeSQ8nAKog1Umnx9HOgo9
0gcMglmMHQF328HAK3LWZKsmd65AgXouVnuMdqC9N5jCBSunEbEColdPOYrX6jFO
V1NVDh6BhpxWjWDHtN1LrNUMk3UFGMVFALghBQ9UfFEeirrTGUv/I2MWTRReHDnT
f2lzJXTQLKM0atH3kJD7tFvnnRxf/FZ8SQ0Ewwol6+UrUQLY+3b7VhqF54+G4SNC
yyvx+a6wt+vus9PYrJWqj9pmn19QuTD4RMdcskmafxExZblnwHcPMiXgSDJfma1w
kmLSh/+c5Vlym/+vVB5CBSqb8bY+HrKWvjyniE2nHB+/sSd0fuac/U75sMueD4rS
M29ZPJWFZQHhc3fiMdSxKZCjJbkYkMZAlbjodT7jyQN+YJtuPWyHuzhokseH70a9
Bo9656Ac437l6Ki+EYhP6Z7fAzyFPbyTFtRzSZz4pGqbO3PnGEgfndqp2qegIqXL
jK3RcviCFB/6BW+pSL5NOQDA+YpN8d6qjkbFZ8CSmG5Pz7OCQZguqyYohmsHsKr/
GZqauSJbxroQIzN2M9Atour2gIFxaXi4s4ruuU0rrkQ141KkrWqt/XDGNmzPysxT
SVa5sOaocmrjdmpZ/kFB1B9QFMMvaT7G1jYeA9VXyXXRf4ecxU3KP9mMNLIxEm0f
n3riio6aM0uZGE9m7jxBesR+SlurH+30rOl7iQ97mweIZLVekSy5vEQU7dw2zmlw
GfUYyu4PU/gyRIrBY0am7xhVNgaVDeU6s3a7BglRBe0EfPUJMAO+GJvBOAFN8+lF
h/zgArkoVEW6Omy7onbjx8LPZw6KVHj2NCd4xcuvQn1DRMv5pQpVRmpC7uwdpZ5X
pkPsHHrQ1xV3T2EwxVIdcXR5QJ96J12reOLnL+MPzeBy1TSK/wisoasp5eZ/eG5k
gFkM8Ury+sXoI90yZjc11/VbNWah5P74b7pcFmuwVgFnpLqLYbkgFybRdqwNV3wL
/cl0y/osKFkGZ24qugLl15N2+UNmmxCrP94tezejtHmupzKpb9VaNAHbH8r0NJyv
z29JgcpRlbgLsRq+q+c1PgDLVCY9EKexJzHRsWQW6V6bUiEKbN3VMcrWGUJUs0Nc
ioh5uhLIhReqrKrjxPYZL+4WkMmvYpOWF0p/U9afY+ZG5cch9EQtrPeXMC5vLUtV
k4T19heA+24w3Vsq43Fsxhtw4OVhfUgh0tzGP1IaVJyE7ID7tgpTaxUuD1sB7WTS
TGUsikH1a5sxIvr3qVE2eh1u6DKZ8Dm8zACdi0NyrdS79fT83QY4mwNbOHTe6M/+
/kyRp2Rn9bE3W+A+4Gir9XNE9znBk5ujwB/S8x0CKlPGUkQPxpsFwDizzo4M01U8
04xqUDsxAmsDp0x3odGhGSd27buB7wZ4B1MALHMpiNwCfPCvk/wIU1Xbhs0TTtpB
aAYWWC1zG1ufuV1LDxZnpecFv3AZMRmG6eKOEhPPGdM8OFSFQM46k6+rAmwtTFbC
TWeUcQjsXz6XS2nQv9nbvnLJB84/bLUX/GZeSaYaTHpI1A69vkJYmrwPL/Wa3Hhm
mFTRIKZq1nT5ETNiuFYxXfQ+zPf5RL3cjLjDcwWDcPX1Zo4c9b/UaaFWc7SWP28p
bkF3GPtg5r6RWY5ybO4LmuEMFUYrAztVF3uNTHVwFb4VidjOqtW3Jd2Iz52aSgYm
C3sBtgHPFiuIYptCy7BVFEXU8EtgvSNi9jMt3rAgnSwVE7t3GELLaek+0PEYYlNt
rLhGnU3ttHta0B54qIxg6V7DEJXYUAIiJF3qqnatVSVxog4TxHMpyqdtTTD1TJmZ
g7DvduYgYbNWu7RlhAWDCMImP2yP6ghNHeooMwAPYZXuk2XJrElZWYK13rWEyet5
Irdf0mEOLmjgvl7JBIOA0BA2aHG8cYaOUIChZUZUUDMBDVjwpGoLBifKf6AdfIIZ
qOoSWImK5UzYd3WRjRfHsSimOAh36qJDIyt3JJn4xixXk83NcqrKZ7eBl+8HPtU/
CgjpDeXtfX0t6BUmDZZdS40BSXDlgfV5Rnr0tylAfztlVX9TAbloDwN+a9T0VW5G
5qzFVVlpOp+OR+9BtHRs4MXM9d29XpaAaJ2C46M9OSjCw/3TR+V68n3NvZJl2n4r
oXfgXJ3fM2Ma6TDaNioPv4QNcirfXxOVKIQH05+a39BByOvL6ImSoVApFE9+Amii
z3MCtHFRq7zs0It2OCj294L6K5L/8IQSwbLo2dd5Ukxxxwyfth9ZpkjG7KdBCU3s
n7uH2TlgTnk6D+/xApjvo9arYsDEjcu5KCCry+2BJcwzsL41tAVzlBlMJN7Kbspc
Qblr5ZargEoa6u9UUHgI+9A9DiyiOJrXTdqvvtPf36obXha7ypogvrzUMzUT1HHd
x6b7o7hvw7kIlZrnOBowtRwdOVPcJjNMzOgHi3AhWmwpAIz60JKpnxCZ95mhgn8V
DN9Qyol3iEz9OruiG/AzIurUUyIv/1GR7k+1mHofMyBl9Sq9HfV4e8+MXMC6Rk3y
njaDQangsnIpJAvqyJbeCFfgn3ec0cu7tkGj9Vm97cQHjZqIJbwaej8Ti2Y0AJWj
zQGQDwMJJ6TkAiIX/6lg5/ZFOzEXPSc6sAwRTkHWqksOGlKfbd922//hPqe5lwf9
+Osm2qaAgGMbMwQeQFTTiYqtCoWDa9DeUzg6cA9wE42s9O/BcQhdZzWEs5raUTLC
gw7sq7RQULe9829kBHCFRhtAVz5qdtBk/fCAHA7mCqgJK/+zxcMfxcLn9uuFCS1j
u7fCfbpaqnFG8xMNhRRt98OQ/GoWNvCTQ384O7gB0HnGME9kPKJ7UHNWTyIRDcti
Y+OeK73PjoBm3qYmq3egyWNU5IgFqm0ac0hkX7Knidcx6B3IXC9MPyuEQtTHS6C/
bkcjAZ1ExbFqi/lUn5Wq26oWAoZILhfgdiIz9NKoUZRBmJQcMat/XjU8q2s9W6rX
3V0OG3yX6r31li3HTHUJgRfTrtCXfjoRk1gHDm9LSi5fbOQQYltnS9tyPUY3T8l5
NYO07Fp5i7ZPo5mL0IUxa8fhZR4Ry+o2g1I1/vYjw4WH0SCS4/NTxRmh6wtzWj6L
djCp1g/lVhqeJ9vRVgsHR0Vewc0Asb6UouZuavAVU/C5xCi0bKQ5RQ7ehiECwNoD
hJ8mcKM87gsVRey7rvxK9juZbWbqjrVaYHjdiAZrTv9hMkNV4abr/C6fzv6VNNDn
g9AihsaoK3opHrfLPzgFjlGOThjKBmkysgtK/DCBUVzX2LtYE+Rw6r7KZx3+isPs
SQFZdixoD69zW5c6U/lPXSYcN0WvDyd2mMtr5g3vhL6vRqMm+ErYLJ/DXhWLlN1k
DWl5PwJlw2Qk9YtDcErzJ+ALUpNrIMbFZYOvuOaqYoRuC7QESZGNfMJL7dTEEVIF
w+1e64KQ5ctsphTzSoacSua2b1z1Tjip3/O270Qc5GTTEzi3u2xlOABQUNzsbDFB
KpxHuq79pT53eC3R9kjJAwr6ePTgGyq//Te3mzj1VwWAfZ1owPZ728iWhSuiXlXQ
2Qt4gwy2ZHuFh4+X1UP7oj9DjUFEgLRRCvGHFkuyyrdPgVo8yPdTiTA2Gbz4ZXke
XxCQbLrUkNyB6Hg9PRCICrs7yDrTUI5KBIbk05a5BvFFCbHRzClO++hbPWIUrc8H
wkhw6N2LzMI5fs2ONvarikaK/pqU3gwvnqEDsBtoRBBeyRoaIKTh7wn0OIIoVdjK
iifK0tyZF/DcfjcefcXgVqM6Of9cNPuP3Y1jLsuQZoKy6c6VDpaul8FmJTtP8jqv
dyd8hRxhJM08cu0aq7RvOCpVq4aeZsN6pkJzPQcCgmSpeQl39Fvdi3lE4o7uUFKb
s0tv31p/QT6IcX2EqMPXJJapUiRSMWN7r4hNo5Tt20FR7coF5X6571DOqoDRp8dm
n6tyqOHi/+sAdmJyUbD5AmcJ+RIh+hqcR1w+6HgYX1jpDX9N5MbOAskrZQcWFsJK
HOaDuh3RJa9HlhHzfJZOfCubqg5fwOQ4s5b67FYRHU7o+9f93uhmO41fivwEZbHp
OmcGmJ8rMU2dIX9H6wKUYIonZai+aHHHKQ1hLRvS8HYAoKKZQzgrCpEwqCgBV2H0
GHjE+xjQAMf2CEiccoX2O5ukKNWFhVMQLyDfHOuTv5Li5Pjl10GpwRP5VdLwC/iT
n2xtFivqSQgEakS8vfjbBl4Vy22iwYxbacPFWw4ygcyguHt8S78lxQCZSd1XU2T3
BTfTBBrhFo3D12CdbBPhZ5laIfFNWXwAqpSuuuuA0a8DsQVs12eN15m/WaW0B0h3
bfVJ0d48rFes1w1vhLbKSAcUa+BAoZke1Az6JGBQ12VwgGT1CVxVJ/SV3BrZP/UR
DfWLIMRh6CeldHEbCXTMAOx4sX2Y0yYBK0vYR9YLu6esaJ9uOqMhseo4wYx9usdo
K0DecnVSEWZWGmlLTwotxE6ArtU6XNZlR+j4YGltN71yzds/Jf/p0m8AdPKJX7TE
9pkShgQoK8ISyxJRIobyCP7cqR8N79Vh1rbGIzP+XEBc3EXMM+rTKV84l407EaPe
j310vpwHx54gpcUxAHoNQEpfy2p+8bkBqC4bfw0ejlNsovJ+zFjjpxole/6YKqB7
zJxDsteRqTgGyq0YLrcjNj02c6LTNp+iaHVFSTX+igg1PRbOJFg+lXmMjRgWnlSv
wwSHn010BjreUZg9M2k5DJIphO0uaKj17BrMYofpr2VtjMTKMdTGabzU4wnonQ3V
E0M9GJpjCjlL3KYEH1sEiljlgH4Q03q+VcDVw7O9TvxO7IPONBPqFutdcWFxIbhN
I6sh/LrANtvhJYbkGb/ntTTpW+j5biMSiVcZa1x0lIkRc0Mvg3t3rzX5xtzzygdd
CkNv0vRG600ikR2U8tYf1SHsukBxeAOkOfRSTyJ2rVsLcRqd8dBAlm4vzcUsqD5l
5EZy0RTqHaa86Jjfgap4FCo3z1Bq+QCrlLRPx+L4Flr8RYOgNlVKcaEpRR05ja2/
AywQWOzCj1YtTX9/wJDBKchVo0cd08atP5TPEyspX8isGO077BLt8w1BbqYO7KDd
tmgYoKdGCIWT+yMogcu1ozytsmLBwLvi3lF4IAKG9zYfRZ/2JZ8EhKAhxYGc1ur0
BQXCXEq6RS5xLAKW7ve99pYIRlORN+V/Cycdb+z65qVolYOaSlHIp0aFmeAMvEvW
B7dt7y/x+Ga0RLimpW4P/GuqQhklmJa0+r00AncCU0ZwRUo40/Amd67dYYWo1IO/
RVJIPb0vxQ5tQf0TOx4hCBzzmp7t/tGNKm36aXsXCzqokD5KhektUmgNLrj+ESsz
4k6BBGICSsft7XC/yX5IUQljl8seyn+aDPSnco8zir8jNWXtdrotLbKzezkFa9+S
WMgavtfIaK+hO01dHGS0VC7Dsaif5xBV4s6GS/dOkyFuPcFQ9nOpSMN6Y6IdBV21
7ZHrSSeSyt+dLsW5s3t0pAx+F5wDbSpf4Mqq9yS5O0W5ItO6qXZIa5bX6P9bXPGF
ZsgvFSOdezZoreQEYnmhdtDJLcOkTwQMGC580cdo5z18w0ruyqF+xqMhvkkVSKZi
GQzOm76H6MxXMJvYsjPB+dlsrVB+aNhsGTf5+ilma167DGPEJlNYn0gkni8PuN30
A0AIQlFMhml2iwwh8Bn28mHNSZnDkA3Ys5TFeZ5SZcSRZyMnjGIObmRnKJ/t84LX
nRa0wN/ZVPxx021GCrZ+sOypwINA+HCqxixuokuh8D5pGi3gzw3MySoQzFbKeYJN
8VNlD8E+WBVm36RIEI5miWo+0VPvJzM1fk/Ny+ZRTlbq5xzqAY+talKHZ2WN9DIf
s9YQvLEoYymroz8Eg5JcFazpUHKJaUxhWAN9rmcOwPa74WJ0w5sKIv/+QAdQ0PGW
peOfkjveHHXDoC3YMr+0L6mht4rOgCrNN3HPomK1EkR17ZyOymFbQvCTJEvIGa+g
2gheFK2ZtLOGU2PPKvRYUtLjxe/uCiQWYkygJVHM8ZxB1qcCILRXjPyouliYXA/E
hnTqIw4RAmI1ZnDifClU2E9LS1zEzJfV0jT3vE+wp0uc2V1a5Qry2Uq5rzFkvn6c
GbiN4Wu5wlgc+W34F8eV+naqH0BQ23Gwnwgfkhp350lhdK5jxaBQ2pCd/rxSa/zq
YSGAYGfkv+nf8VrDNu6jEWItMLkbC+lnLimT8O/bMseGkHAgjzj9DEkVerTl8iNu
lFLuhyNN8+EJW5g7OJMgrY7uY+OA3Rc5V+Dz5+44oGPcbqRaxHLz2K4hX3PH6qFa
TJNkZRTm/2+9owt933d2/WnUgcxWroLp4mu7oHG4elSyhKBcDYJtsXL253PdN7qg
nJAfgmu9rRk0TPfhaAVufG7csoKd/ooQDWaV00iu7U8B+/kZdmGc0Wq9INcJwuJ5
jYV/eY2kwHmL4IfcXA4pYZueTJDvRiGOVVpLaecpX4CzBWvAM8UZedi6Nu9eC8Qx
3JQbpjvNlb8LQud6M4emX7EMnXfcVfZQRJyadLqJoQDzGR1YsYe3y4DEPaLhzM2h
lYjhupK/Nk77On+8oAE7pHfp3VCCkWRQsL+UYKd9asZ80j0Oyyi5WAGfqQs1NhPq
Sps1sno2Lg/2lM5I9CLV+dWgYojFKndTO3U73rL/2ebNxQJwBO/TgDBfmm13ZHsn
lj90OB1izxQLrpCAgsj7DcHjRXgsGRQ7q7LMDNC5lf6/EvME6vEamJOYLRSkAWJK
NSLW84gk8o9FN+ws1VV3f4F4EGHaJAnJNYio0ITfHKiy89DcMm3yzojbhRlXaaFf
T3Dq5xruokq7Tf7bJu5SxpNWfKTm9YBTLGBKStDbrd8ITynfJTAMhs+9q2IBMU7S
AxpQTgDei0Lnn9ldmmenfkLbtGzPuP5bj17zvxzPMWcUmIFWUoVO9VEXiS+OsGLT
AM4zr8ouj6QtwQZra1uI/AznkWxKqfEuBgmFYT00eg6eJhU8+qgI7bJ4A3pYwtOh
kDoXbiw/vdQuQMYG9+9UXFZ2+3B5WYHEqiKW4BdUyt0450cTbKUjd8DB7mgvk8SG
Y85LVGLzqh1l8atJgQ9dSbNFTQKYLMwXsnH3/SmWcOJlF7zSzbauBHkcXveFGUPl
IrNmN4K7GSbRiwlrpHAjBIcliA/icoFRV9YDsg4WTjdq8ycMkE5dvbbusOuPyo27
DHu072h7w9ddRc7fEtx01DsBb23m5ng+G8/c0mYzwIyyDr2k7cG80fXtUiCdeS17
ZLJce20OTC/MqVn/2yrjrJAY++fF9MCJYP19KxxJCmRZpE2kMSC1hckg9nw+eWhS
nEx4z1CJmqgM4kSPJ+FCe0WBpTSdj/D/OfXstkJpvzteDKK5ZwL2+O7MBa8dPlQR
MKzJUZ4yPbTCh3WrLAqPKSfEMFR8Gn/qzrRIOmWruCczDSU3XpC6AayjAdngbLLX
UwIG/reOMQ2muChab3soa9/fx6p5ZBzvz5N0N8Fxhb6hzSdPqhhHoqIjJcKLYUP0
e0CWVjvzBhZIUgyqHM0rcW1lqpN+VuGbeymoBzE5KiikxxLKEIH2bhCDGglMoxLD
fmCLmH4cSFSIwaGVctp+P24GP/DA/d43Lkv6zeIq16MARBu6NEF9ZXHIRoWfgnZA
26an0vs8aFNYYlAP+leihiC1h+aYrjcq0Z/IOWBsU7bdebuaB0z/lBuxYc7s0196
+odyK+4IjK0HrDbhL0WZwhHMa/HBHvgItoNeazn9BgvrVlKiqsItPADSvuoLpEW/
XBgM0bm31SII9Depv5+n+BFloQTUNE2q+doAKlalzsMPHpSQsEk0lOo4j3W/hnBM
p2XVTbSCUnGE5AdHj5/7iyc91SliFELZ86PAikpxh0qtxV0+S5mRXOZA/FFhz0Y+
5ZPGBVUse2NDToUlGK8dunQ5C9u71nPeCwrSChj0hvLZQ+MpwbkxayL3iGqqCVww
mZ5odd44KzLi+TZyojRkYK4LiBNAEhrrvlTy9nBz7KF7bCAXJViBTAggHQxRR5Ea
FHkFl/qg10mu5g4ty+M0WvNBpJdMjy07CtpRdg6JhDnHybMS8y/3DqKiC9cIdMZ3
ufcKWMssgVz+cak0N394FaZQTe3AU9qiC/XFZb2mddgJxVClhvxjUEV9LGggvWW6
jS/y4iOd4ltHZ7CRmOAARxj/f/tPrAHWKxI4qMnMJwuG2dOau3RRcQ/udREI4bEk
tgdst93jjNuxdj7S/87S5mN76AcNw0Es9zuFYbDZPqSdo8GZtUBrSjyjFOlk1EKh
FZ8QElw6QSWJ7fiSXycQyNNBv8c+IWUSCnVRJ8rxHyhomaZrFFe0Cy0UZ+uSdCJX
u70SSdWYtWl2XZESm6pA0DgGTGE5QTEpeuryCNWZJ/ZJyp0RZoAK7Kp0vUvl90lB
h8fj4/r+TdE1ekZQM3RQxLH7O3JhKkR1tVdH1qLJj9o1W3hdXHR2xHbhlzHXUAup
+m9M70lXFIDS4O35MjJR5iPbrcq5jIBxJdzuRSiMy4/YFcf9GvuawDIKvDTt9wZV
EQUL6Wxpltsy1YVHA43b0oG3NZr5zsmO6iNNfF/oYkpjJTLuEbqq1AI8cUwO9V+m
jSx4pIUlSuyyuaK3GU7jFLrTTK15/BUrjuBE/y8Egye8deWq0wR0V57vfuOW8uR1
JXxIV0amPcWTzgxYgMUlv4yJoS31Btjhy2yaicoY0e9FmlAwkmbEDG/5DuQUwfcG
bSHuD1RvmD9YL+1j/ufxmY4fMVrU5V8S2VqVoZNPA9BVOyMu6lzlh3PIYBc4U3YO
P5a3RhC5Er8Xlwb/vM5gOV71firzBA7MStRFHzRA3wKUcvcCNFwYMUJwLA8BI0K/
JjpdQsqRoen7q7JTqgJ2FfOlIcD+ze2MkKMS5mOF8QBfStsKGy6Nbcg3Zb4SCAGj
hnlU+szwqHqfcRwsoWykqOtErfxPTGgs3xLygQO5Q4xYFAnpjLBVVN80d4EDkOe4
Ffq7OY6rJiNRbVnBQXPLj8Dj1TSxFoyoLldEHoixhrkFmqJMWNOYxroFESJKBRz2
1XYISMuzOZOvVu0rozZJh1kbcYUoGDkWL/9Rb96ft1GklWvWeeKSpMPyOF4cFboG
kEtOUesc7otwH6OSUOyQVkR4RM5FRd6yISmfo4BapFLY9yH4fQGBOSCJD44vXyRb
X8AkoPksI9ig4fk7N48YqQz1uong++01DmG0x3qEbX75HBJMhRFl2h64wRd4Zeit
Qh+4/7usvXG5f+NAn7pojPRIwV+KaX9SmJHbMcXMp0Yim2dp58y8PAzMhdi9S/3G
7SQTBpzjKoh0OwZZAaJOD6a0pZzD+EMjJuGBIxlFG87h9C9ckRpQ0RSYailIo/8V
VsjG8Ea56rTjEyh/8pMFugiHfwW4jh0tvfdF8cQuaPVWWVTOripmLJEXJ6ihYXSQ
xTM6sOvNitPY8wIDPSKiuakZajHAiC8Zvr96rYmATDSEx6JdgeeNyJNPHwKJFFnO
hkcY/xPscoTl5Z0f3w7W+kVsw6nVvoZ4i0mxrJ0gM1CybrTeeS+NBhdU0ecs5vwp
SMnRjlkUK4NuIffJsvGYgvxexKPYrG3uQS3bQlXJPWcPmoQ99bd5T1hrUCqSq6R1
LQMULL3vmprUs0B9hCvum/WOPDv3uWev2SvuLqo8ahdTZpZGX10oEq3sDzWVggz5
VlEOZefTi8/WjWwtjvNBxNff0bchE5GOJG0YfeoKKQpwPc5H9skCqSh2YQp11fFr
0Ppbtp7LuMRPuLJ811qbsFCqMSH4yjufGXejtcOgvqKFsntpUCCXKUReEChpRxLp
Ml5Xrr1yMia2Z+//MAl1LCV+wFTHTJkxLIofUR1sSIPQfRmfM9lwD/nt4yehPeH2
EOTw8p1LFVcMF1Pxbh0j4mjeCOsqoGrcbWdbQv7S3qixBqOYkx0mZz1Jupb4UkBn
bSFyLUnbBoN/fEnhyL8gg3L1UhvRz0wTTE+QAlSpfnPiYhLlndEg5tRu21uUpyRF
Ort4amxbxUUEd4eyrJWq/DqJ6+dM/Tg0FpxdVwGpIOzXeJ8PJri9gXuxDfxjfO+o
VuPE6DFon9a6s1xw+RlVGnxGIEWEEf7yEfce57rUYRRhS1q7cr2YrtflLcXA0Mzu
auyCu3RZFIiptwn0DbgtXIiUEJqaueN+7FMzqqwmdFl6/J85Y2PbQb9gXvxb3amf
DdETg8chrewtY6Z0EJKLOyBByW14283kOuLuWVOyvDiYlzop25PMyrefHR2EBXPm
1GmSjxzrKg0TICbjWL3cnlydFS+LurjMZ2wNjawWIjkrfF3K3XKMAR64nyGTGzRo
S/bwzUge2itiChsYUstt/0Zmi1ucEhvFzs6G+Plvtocm0rxrRE93AqzWwxh0ILeO
WoIma8qJqh72EcGWWEkmmXWZzRGvuSGXqBm880gUkEOaUN101+chicSSlVBarJip
Ed80zlI5wBqsT7Cs1lz06FUYS6lsmle4ZX/Fy3e7wqmmYWOKKJ+qIWu9WYDYJWWw
JmyZRxQcs+O+DPd66D/qyxfKZ3ZahIpLPqgQJNrAl7DRvM9t8ldcyBkdfWpACqLD
RGNqILC1qb/NvcxVgizrMcxITVrd58WHMVrO4Co46Kv8Zz1+SkfI0lxxyI2jIMTg
Qy8e/bDVQZIt+cpcHBG8KI8vG7yBvpz7h+QFMWNv2a4X4jYwiWwg5BIl7HfIQHIq
ddEFv5NtxDgCwD/hDhG1VHO7vr1XSkD//Wf/MZE2L8vFU1mQdzdHKYI8hYYA2RZZ
/PeULeXqBsRxjGgYyuBByBMN7NMs6CwqHXWUNvbPdUb+fQWMDuc9dAwlwNGOBLi8
tUkaSKBmZs4BxRGhlsHSh1G23vFGpiEPT5+ZPL/Kva74vAmXwmXQMhs+eos6aDcx
UOy3obxVFqetsNOg4oI2QwLMViwMhozQyzbYsndQlhzPNjvbiYAfr7lbFWBMI34H
X/kwRF9FPrygGcGE7NBQaIU4xNWNYcOJzG+HHI3PDl+e+WBHpJ7do2s1sezXAjlP
l4uap5TnzsHI6rbG7thht435ta16DNpGrlfn0Ly9z0yAPOMhzdn2xel7/wGlffjL
tcgPDuV65uw0/6S7HHlCk73x4QrtTpiTCGGySUhDbvJh5laaxzP7P5GJMJBeWeXF
JVDkAeri+OGQtdJz76VJHnRgr9bKH4ZOrP03IjPHK/bp7DGm2zLbYKFCVcjQj6HQ
aiU1uB3tqffIJtJE8sqsra3mA9QR3xzVbUNxfzJp4iAdiT7p5HbKYSf9Jvr58Ay0
RCm4XXELENpR6fD2Z80/ohj0tDXbOMspSu0vLL9rK24jEAZcafZGGsuJZM8IqFaU
DJ58v0WU4ilqXJqlIFH3aYnrMB/6DRpMdn0QK6rqdNLrkMpLbQAnkUV6YUnqVK3v
AEabdX2fTWEJlYiTiMxDTbDQvhoZqB9+k11slaCHe2FCT8kYP9F9505fzSohi6Uo
CzsVezHJOIGUwxTf55iShYzTCp1nF43ZaMQHWewWo0LoOfYHuz/UKDoURotUt+0l
qiSsuiwrM09eM/MwFhxtVjo/ZkiiL4WjW5gZFPJdX8MDWnzZ6S0MahO7YLGrfPs3
qF6clmZTmTekXIVONwDUsaUrVcaTn8vIenWdHGLiuxz0+p5RL8hvl7yVe5SRyxaG
pcywzmRk+7ET1c1Dn4Vk3XPV1nWG3SvEvdPECXmdZhZ8Wh2J3Ko6DGJdTyPxReY0
MccAdcqfDRmBR38BF/KaA9iehVUOkUWTfQM5j5EsJY1efxlX/jitFzqesKGSzbf4
uTeyTZHpEu6XZKzznX5VSud1tQAnyb9oaf+NgLsgWSitJ828415w6La+YiAMannm
pf8lHItUP01irPYdtn20UoLFJ57QZN7CkhczI/3IDVMvKfx/whyrrZxIK3rmu2XT
bxX7Kdk5/sesTwS2xwWFYNKOTar+ZhkqwNKBmo9aQE8FQ5Kt10p1s0k+KOZrpWyU
brtRv5w4JJr1cp6iDcPCHQaj1ENUQvHq3TA+9H/3KgCXVSAV0ufwqUsby0VGOstw
jJ7hOKS/96rgWdimyDvjuJTJJwkL/7+he1FejO7TYdY/+gFJ0vyugOQXjYExWW9m
kToMICFtAf5pIWFiyfVu8T1k2jnhuxG7gLONEDcsKKOIwdXpAsd8EQP50ANU/LDK
LQS3nxTvHW9ER6ijC5QeTXnUzea353ALb0a7xDJN7fCiL+Ge9eF6FyHWk9lfbZ++
jzs6WESjxuZfYqTxnhdVuR2jJ4kILOLsfi3xuhIAg67VG7rSEMGTnuhHW17p7PQM
DjDWVnS0/7LGqVMrUFyjzwBRGri/UGGRvmOuydpDkhYCIDMCubi/mMzqlY/egSTC
qViox4UUpw+0x90wF2RWLaVrdhI6580aEcXn/TnznhUq86buNBCMo165UYSkOL6D
kWAYFUIOu5f7oQsKIh9ZuOi0bbV4PPrIJvnPMFbRthaiGpAnMw1IxOIFY1FUY3Bz
5FnnX2HtimCKCiqWDBkgeG7YCaYW/DmlOMRxa+pZ3frD1RSY/4mfBntdRorS7vEJ
1MR2g2ZFevHlPDeV108M9Hzh27dP9EbEYsWZUhQPiE5lmkmQhS6nELOk5oI5NiqX
IKaVpb8hJ6g4gc5Qf1viz74FEaVwWzNj696zhUWGRlUNd0VEhBgum2TyQ4FKdv1B
7LQTn581V7s8AkYnPpENGsPGtCnmVdYB/yG4jgq3mnvjKxo9fuore3PJmOyHNeSu
re7ZA3qQdWwLf7BVJrXtx652BM+01eiPnz7kZ/9TrLPIgBP/v+xFG0z4UITpzTzV
t8ni9DURgtuO9CEkrddXdcgeuZUtf7TVMk+R9ZOutyESUVCBsHLDXiSLuZKkXZQq
vwUML+hv5WTBjvMV8pNrUy9/R9HN9ApRMuJ43yMyHUZMVKyxQ8C+uv5QugNEpDHL
UK1ayy3XPAATkgPkFpP6cIWoZXc1U/xg4SP2aolo98Yhm9BV6Yfn5l+FXs2k2nJi
IpyllfmiyknEOTnATm+k7mRGUN5IUMHgGRRpkzMpjDXR/lCh6lyIdHSzP+9TBP0R
WRzGkd8xnkKxS96ew4Qv64G4fTqItJA0ICazpGVarueFSq+aoB+OV0XEpm4h2JhQ
onuhhZMvNJYXPBJ4WXC78mCK7zuO/TTmK9ecKBmm2ql3yhpRkEnELQLsRQEhCsCh
Fo478V7TM420MnsWKJ10qJlEPVjzBwxterMoTU4ZGs00478+CDqdkHd73HnRy2ax
nAGhFxmAoCg6NCEnYabEl4RzLySEJVmucEyFiXuM02O7hoeSvswxKSIoDe7oI7RE
9U8M/O5DMV0ca8GLngfHjlXIuTZHEIjwykQ2Had7FrNF8TkyaI5N4uc8o2c0ugYN
Lb+u+4irdf1D2oo8ePva8hDbCsXm5WQLT3mITU1guAe5JhOQ5og50/Px6FhtCRX8
mo6E/47jsO/OrrShjX7ZYd1g03P2DRnjfHaSncDuzHCxtml/UC7rebixnMnijZdJ
x7H5O840fdbwbsJkG4aX2OeiYp/FdeXpmho6gKTWkVojj+4t21j/YPdYC8BNllQz
e3ecPJp0tROGPDAO7zpeRecuOeAPonT39iGRtyczjNb+dHJgZX3RO2E6ihF24rRC
APn80uKzN4K+okfFK+rktkY+8dgVuusOGbIJLeacGJe/dBRtSAZdK798MMHpuRRq
pbWHd9GffnMroadcitfNbo/BIi8SvzcEG/IxkqE1LySfL+aAXRMwkb/wiZW9QVq3
fa/udatISUb7l4U6YAk9N8qrJt4xeQk6Da8PsM9G0Sg6/bUo0r2w/6QQwKv5DUHP
hHf2igVg3RwfUFNHb37Wx9OBVUwxVPC/OJ5hjV0RyQxgKZIhDrVB2cfW9inr5t/n
XmItQSSUfFiKh5puI7jFpyZR1k1mgGDx4xLZIqRPl41ACH6k0EsjQ1Ra89rabQB8
Oy+LrKIGICay0CvmcgP6LIKv93M2dEOJNV4aIwkMn8mjuZKmR8hfFwGTYTGDRIHe
DCjxATKxyST98gIryba8gPOxChhv8yjfhAkzFTHete1zIw9kWnfBazaaEIJtIke5
7Ivao0m3qA1AbTitxyTg7KIlIER92WFpO60rnOzW0UXm1KfFWewz0bBisGks1Tg0
Iu8WK1vJrxxRMQeI/TkrLV6VZCb56pGddm34oibMK6RfsDcotJg2ey4sbJnwzyK/
NrxY8LEb49EA4Z2nbAy0sMMMkYY7eGZkgHxA9t7N/zpeTfMGyEuQGmxmZ909qLiR
ISXN48mYc20+c7pPW+VXcKqBrRBpha3qU9zTdZ4kHoo4JBZGmV1KUqOEYQeMSUQ2
/qQSrsUm/PFkUzCC2pwKml1lTSJDh3bsBFs/Ylpo/qbcUn3T0c0VIWhJMZIW4MuF
XCX1Uk2PeVl2eRY+vUmYiyRxL5fVfs2CSNbZPHbklLtdxY2z2kg5zQkscoXRRSOA
6mWhGoW/MZ6clAYDxeuei5FTyAuMEv5sL3Dvcdx90QRFSPchlEC/b2cCAPCP6kUL
9PYqm5GCmDlIBBkecyXl00jYozy/5AMVcWmmv8lNr8q9494VXSzMWb5hkpgLTFGH
6aNmUCWpg+/051GNpM7B4AlaRidpvMKSLs9RI2jLK3jLMKKkpsc98Lr+JN3GcLof
6Pjxh5+MBtqZR3dTQ91Pvi6mvoj7Aw4Ce9/7Xk3pgln6tJKgLqg7rDPHWkLv+All
O0RAZcBGPUxpDU/k2f4AS2t+/V6qHCYIX8WxXkQ8xVsRpIoOrWKvld46I4t1U7jw
gEk5E3geseocaooAb8ZHXrX5JL2rNMDOfHHmvfACozXpRS2c1qFK8ywWDFOUX2uZ
wbp+LOe7p4y7loEkYuBV/Qe5+SwJi/0Czb5Un2fAxsKNWqJxHNoJx4IerBdRv6nP
vF4KcCAyPSD8T9OWPUCg1L6eEuI+qCINKH2oynL2LDfY/EuWFVE7y/htA7XX46ji
K8ZwSmcx06AXqflcvw6AOXL3nEM8P8jF4OyzBgGjU6CNMDB0gN4m6g4tNmr51Ptt
o+i86UUSDtr6zpLViC0HifcoIk0iZkJjR57Drran//AyBVfYiCAL2kypOeWvvwvw
TDVTxXxhN45oN9V90uTTZ8wk602E3AwEpkQW4SHOlBGMHf/7rC2tFHtmWANNRayU
wxF1N/NUyYm1pAF9VJ/7gP+jNGdhRmUJI82NQKKayltnsYNLJ6ARw9anzTnjRNAP
PwSs/Wb9EVKBVkfq2k+cw2XffA8Uo9qz7mEWl1DtXwcFNFo6mjiUYdTKrT0IFMaH
lUAWwlcGuXtjwAw2Ewf1qmbs2DkkJQDQq79+0kMuCPHb5uwUQcu0G6gs5agjnKIz
tYnE0wKk2e6IaEr1nV6rfXD31UN0KjjZlQX16ZTDYNdj9io+iuovigzOJ/mTDzuB
J2iLsXFoRQZwasbdY9jlk3QFQt5Ij28OohygKnb33BFCPHE2ivBsu02qFnYelGut
DcgsagHQJlqknivmkBPOSOaDWp5spHJWHg60+Op68SkEJYWVLOafOJqxto2Qfgte
shUH04+jacv9RJtIGpInSmxis908jnU8NThLqMTpKRWzSq0S9e1CViQk8Lo5M3Yy
9y9BJbUNUhjWNpnIC4kzhCYHoudKVA3r0u0gg6M6uBzaweUDjIcplmhDjuHRpWko
3lFvU5bPm0Q0iSg5XYTalVGJWImuz7LkIL0BDr3GIz2o0qf0DDWFiEY3hXWzZr6Z
LKLg1Q47ZPNhLONsnhXBbhGDIk7I3Ka0yCC7GgyCjl7ysdBt5qe6AMwRRN90N8Lv
Rxl9lBOoD3gvvm5PdXETJAKxbXcB20dFfWRXvyBwW6rPfP/ki/o1mvR8qRaLVwb8
Q0IkXsGg1V87+vkYFxYjDkT66Y/X8b8WLwH5w5QbeEMNl3tj2FVjkO+oZddqy72p
xMGc7SJQCbu9SxeHfj0fp/DgOEqJ4T6zI67/V7UeYzspxun2eQ67RMuQrTLqqmGu
TSIipdbKB5gyHbao0B8XZi4XI9jv2EGlbp4LZepzZc2n/e8xl1079PYy6WTKOV/8
7aGnWDDYg4ZDqe+jDwSnzXDYlVQpXS/vxhOFA+zCk1W3YkDzLAG4tvPBs/sM/mCL
BEU1XiCFrf1eg0CwxnJUEA1ITEnmgnsra8V5CuHFf9DeH5dk8GW54hrjswpZIAP8
AcCzJdTImynIOy3C2c2kxMVBHkbTHNQsP6awsL7p6SRvGqyEssweF1Ux7Uk7R03o
fABZm5YtWl9wCGgvEUMMoToy3s/wKJSYPAP/kpLkuWFw6BK2uAbiQDq5KANqAF2Z
Obvcz+RfFd/cNjVM9XkSPb5o8EPARHS+aCOuotqotj1/a+1z7vtpDzyU6hPd2aQr
g/gwBC4rQMaXE4YSlK/PDQEXsCfBeGsmaRsKGvcCPnS4dppRxTmYdFHL1KODjzkp
dBmSIeTMUMcmENed5W7lf63gs97Uz2Uj2U0as/yTtXp/WvgawBL1tLIH0n5eK90F
sahsHkjMN1I4inl5Hn6ENTk20oaynEsAoO9aol/ZAFaQxtJda4q3lJlzlKEX8I9x
pozKyozRMfyRFechBU0oGSaWYl7wbqtCIDpia8Il5fFGn2BrZ8drOaX9LXP1SPmd
SkvAWQlUxlrZW8uSjptyfHgcRUmCyhAmtMyRCBjnuq4h5h9e18wL+ut2W3woi7qj
BeiQolFgdJTNWgtR36CsuTy4Sk4emkZuBCMqDpMaVjOWDIZL0VepVxLh35cR735j
Lb7RutukH+nPAfAj+Dr5Kn1o7SlWYN7pvc5dsE7sv+eVpTmNUgh1jkPp8HR2S8yU
zOAbgOFV1WE0S4qwktJH0Ih+PJk5ffzEVfiXPL8/dgHeVRaA3pcJEdl1IVZttRdM
qgYSCabdesRXTVvC+jGl6nv3axfSLoLwuvYToLdD/3GcrmsSb/rO8tAeZ6klmGgS
I2KjabNNcPykBgb31bIml3VySLBySW9a0G+LKXjijES3tp2n339FqvpCg1z/KpEE
KMxZcomvM4Fn/ROC+U04+MNeUsTMTyKIymUWuabAQXwRDaA/4dm62IK10t2lGqW6
UX4JelsoCsjXFTFynmTdAuPJp+17Zeh4JhZh/AH/jxh6K2gmCPU2PFommqkIY8F3
QOZjDLW5Kni5HfwrZ+F30mBt6J6KH/cDy/kb6XEJDXvKI3wyHDEdh72t/24Jxye3
neIXYxnjk71nnl0jZQiJd6GPl1gYwe8OfEleUg3nFdOJAjJ0is/QlysvRuQiztaP
opbgzHl6btYWXEQb13IgKP5AAGe5O+kC1tFzfuH4x8Zdjb4XNHEUDRdgZH6ZpS84
LcbfWCAtrY5PAvEzWsL6ZlIejEI9woj5aPB2PcBngUiYxsqdD8yjd1j441A4sT4D
ZTtRttj0BYoC4EJOGVHZZF14UKAf37i4Ifxb7mfZOwc6Bb/uCfWorYFJOQCguuoF
LRmkYhseYM86vjwzolbHyryahMHSBvRUwKJPv1fpcO1ccfsZ2wb0uCbL0SapofMk
eBW8ohUUt4Ade2SmwWJI8dXZH4GP4NHfp182DKNSe/jYQAHQupcBrFce/l+YvRhK
QG4/f9gM06IyMrxLg6I9UOA5Wb2bF8Fpa29Yknbk93uLhvAXZtU8waGDTnSjZ4fj
XtozudX5ExXpuFl5ZI1EoKY7chWNjKVFOoBEtRtkaKK04ldVX/OMV0UnEOiRGQ9G
34iEyFjhv1fODs7Nn7Uib54Vl4zZa3VExjIc0q0BPcg0hGpUC/nu38ISSE0/imDW
HazkuyrnovabCKWiD/ugI8cC2igpDgcplGxq7pw6A2dtDIey4l+PVwPlWYvgfL34
lfBdzZ/HT+fMoS+Y/rnSQoqpHyujer7Iw6JNreuylM1kg/wFVw74EPfpfxs+EzPY
7V9rwS4j/nDT/lgAnioY+th+PA7ilQ/LVJzdHA5FG8iFmoz3gHluPEx8nUG9HnEv
1Drxw3NS/4olJo41JexB1qV7wVodIdtAwC9sQh1nvfjSs3cNiXdYydNq22syYo4M
TUJJpLZfE0wGyRIGY6rW6boK4bgsrElcKHm36YufNLiks8b/YnMNskIV2lRb/beL
yi8Spz5OpWlmwDqcafTaKo9E4rDI7kJWh6l+amfElUyuOBaGtm1Xy3l6uUl4vhgJ
aECQO4gdh7wijZ/mwVdVRREM837TF8R79/NkIb20QF+gbtkFDg29G+FAPTglrPdi
0D605ud/HctSL4OGU/h/smghaUkpVTIQvcdmf8Syut0aQwVW0dNMtAaC+QWz7EXn
OJsoSRI4FkSaJtq2nekY52DkcUSmxgnWZUw5NQOKC3frvDUH2AdiaF8qFcBSHgoq
qATNWl0pAPyVLJrp9lcDVuChDCyeN5W8oJNglsdq3jIpsr2fQg9gxaSsDy763B9P
nob5R6JfVH3SG/xCDEXv5qfDJ/aCezekRmCMYhxau2uVJPS/zbBe4IJ3UzQYLmVA
ENO/WNiUVDGaN6WhNDUO2I0g9QYR3rl+5IlEeWLMyPb2FhhWI2KDF3HLCvmlLne0
kJmjc/rqyverWn0P+/MU2PV7f+HQGUn++KO0S+LSyXOM4SI1SkjVtzxMDL+uQdFE
zXkC+R6lbALPoeiJPAKR4GnQTMeTEJIfMP4kTU3zvB+T5NUB3x++9tdUBCfWNb0T
/YJh1tZBQnivR8BAxciwENyCWkQlyPmJA762lUYCM6gAC3YNVn0UIdAuUwHW9FX8
HPrn9ahcJzNKdIEgRrt0r47lTXv3jk2Gd6SHIheoMSz7gusj2pi/263KPjPE6rgH
aW297Cl+ZbkDmGUqDgmdfnG99zwt61tqusDUjmJVEKaed9z3Dz7z2QKSSc4gtDy6
tRr74I2x8qUp3cJIoTCy363VLS8FsJ+lpwLHtyY0vaPpfdmK8M/IeVFUQXHHNPdL
OEEUpo20r1rjgI7ZlVnbiTP3010P/4nZQ+OkgZM5ZbHiiDk6s00C+PcNtHRC9The
MnECEDhojnzG7wMAZQL+CKALOtN+uoseckDGWYcW1I99QwKYlYO/WHWtXY8qWMQj
Le8uxvOSpBE4oAnEjQIJri6vw1kA/PjlwQqujq76MxEpfHAizTT/K8iVZ0DE336C
oFdSmTNKw0g0Cpx2+P8MI5orK6I4wZsIFQfJYDPD0oaDNQSv0ojNxSs02FWAmDGY
6pUlUBQCtaNvpVt6j+RZBIgtAL/verBzLIoyLWE4/6IvCQ+y8KuZsbR/zgmrvUQ6
Pioo8RrQvxyfXEK7Benz+aaH0pKqrjkRdpJe0ZVhnKJyuMuOJRX+t729En2YhGPk
SZQEaFPwkyYqKF1pqo0YsQqCfmE/tfGh2NSiDCLX5zfD2nxyLL0HZbLiyTZNICCG
SxBHMkpkGptkw82J4rIgs+43IuOGaoCvO9crO+uNA+MyOH2rchppOyC8bQaXeuAF
Hj3T/zaqXiY3k9zgdmrg8NM+jULW9CzK4CeJ9QChKtbosHQXJIhWlR5AkBmZadqA
5nsDSj/H6i++pN5G0I3+3SVmTlK4yvlfa1D37AwFPRdACl/muMekESdk5uCbVuix
p2xQ6sjuUgZtt+BVex6WQ5Ua2e3qLNVj5bhiF3jPFa3iuWDAIYTQYWFbIh0CI+w9
tmiiyVjELmqH5sLEWHG8a3aQPeL+y6X3cwD5eFjlnUc/wWd+RozhdHT746kEcttv
dOYHkIvDvzBn3O1viO1ADeMSoCRuRvtQbaqqnbcVRMHvvDmFRQVBw1xjXz42yGiq
s9ZEtJY+K9eQjkIkWGvHDJ2EhnIHVaCd5LsihgyvY04/ua1NCnw2DSBbuZINbRMH
pYoRsfSzo0tVhRLeZeOlIC2SUEu72rVz8cLNnZFLqmO1jBLjMyxbVTwz+wy9/5bP
HPwaqh218sa239cj030xjBVd+3pJFyvcblAZXAhZ+CPGXDkjrP+WgmEJVGKsTnaa
uCdOzrz6gisGBpi5STZuPaoYWFvXK5I+pEvh4+XCMvep0gICiVTitZy8ayfemMTW
tlCrLR7OollqaIQCJGCx+PZxNaOEjRIAQf1aGI87aMkbMK7c1d3FOMGBWWHHrRDR
XGPVrleEW6DlOtICZbogtI4nP1xjXXi6gwOMao26zPDZ1k57TSsWsL2KMgeIX2Ks
oQUNvhLFAielgHSoXaDG7y7YVSBH5r8SllZz5Xo2ckqcUjzMye9FazkTVdKr/VVp
hrBFilw6nVT4U9oNPw3cKO38kRm5uK4zHueY83NGggQTV8ztBH1cB3NrAg6JxNzp
JXH4JWwQUYW1PjplC0gLVz0TqORtRwjxh/TKIhF5uem6a4ErF4dmJ/SZnbN3vT+s
oTW1vRN8fXOiOtTLRS+dqKaPM4d2n0+XaYavocrDTkmbuXe7c9g2KxSX1cJRUbp3
8UtXt2pk3WS6QXhN/oKTaGyfLMME0Fqea12k6JBDpaMzAo/drmgBcy2r8PZ858sM
Mw3JycEZzk5R5DUyt2inNh5i/M6SY1ABka1A4ACPhvS4zJKjpEWKJmeQyFnmDIXn
KMqaD+bLNscFPGY85eAN9tGNLOJj8g0U1e0yh5EkGALbwGGwLcwgpFlfxeQ5v2Yo
9ZEy40kLMDokwGqOZ7QfTt+6dlMKwv/rRuW4askQ+C+qRt4VAFcXbRf6oq2j9QcQ
pFiP8RHTeyPpDbLDKs/UFrZhI+kZmVnJc0QrrxVW3oB+Lw3MSPW5iQra3VefSqGI
vF+BM5SC88oBAa8UQ+vcpo3+r5ApvdHlyH/pfffJR+QF3W90vKP4RFLmQwCVOinN
W9T6x48uRC3JAJK/+fmJsyKCav+/Md90sy7gqPAo3ExB7enlmYFKnGyMRG8ed3OG
p9Cqw7K2KQXcpK0l1hXTqwFxbfCsyT/URGLvkJpHhhyGvUbpefaLm7jjf9icosuo
DpB3JuVfPYr5SiovzJNqkxwg0BwvEj8ScN7pwq7nc/xdcIHs+kOrXr2CPErG+9mV
r3vGXrbPDcTco7kk9+MHK3qTRaL3hBPUnpCDFi3QfDpmAZ7wIXsPDtwzCb6ivhCd
dczwDE0PKx0el//Nh+Zo+wf+A0Tn6ujZ9rorIP5WTysWLUjLrIOhYdQEfnjL/fIz
3y8bmrfTrJsKLYBPJix7atHgdoQcKQOXKH0PlD0PDaPWdFTFe3YLyz0RiVQTrkEj
w3cyxdvrPzYbuZt9JZw0J1baXgE0Fml/+DfVJ4DkowBABGAVcuA/lxfu78dH39g6
EZaigkf+Efg+/mI/GrQcwHWGpXxmXaXcyfaRVa19pYLoTe565H/yabZg5L1f3Zho
TLdTg0wJcsnwliDdxNph+V4VF0NW1UAJHkd+47FwDJwAEnyEIuq/yH9bdZtzzFHH
kz5dpDio4d/XfLpgAdJbnScifrsOHkb/lkT0etAPMXuqHKGEhCqGnjfQdc58QetA
FT3XveLIPz8y4gnyLbAovCbs5IJH8366lU/p4qgIdwI2QGKdmoWIOrSpSxIt599v
uKPWoDdQyrTX49WengSO8EM0I2Iiw6yUdhoxLU9ZOBVryqhinpFCRZ13mJuLKQVM
WN+0NOTspjcNS3lVtPvYhdxeEQuKqpz2aAIKukp+y0MMPF72V0GIhE1jk1GhpMM4
ACubsoOETwibe6e6/3tDRroqB3ayzrPB3e85yOqNpCbde/3X154g9QPvfXXfoA3+
q91dhzbznT+Agpi4cVG7MnW++A7VlPTEuH+9Yj94p0fR4Pp7iZkqPZ6GBF1tHzoA
e17GGt+XSe/XHbWxNkRJbmb0WLvKvQMZL0+htUvo1SOf0RFi3nJc5Fx5Z13K8bqB
j21j3eotIDUbHDDY0CDufeCfoKgMXaRTE0LCSsKcI3vD48n1nNSI1Jc2jNqeM1xO
J0D6UwY5e4PWXZhK/PpAim7IL7nORzzB4nkYKANjtxEOG4l8RADPLgc5EbYyA42e
Vyk/Ciu4c+C1b4JkkjmPa1gkByT3NcYRAXlUzN+rfTVuheaf+7DF7hU9FqwEcZDh
ZFwe+eS16Eo5W90J4jnBPBT1EHnIpUUE+XMHj8QJ/nFdam+Nq328WydypLcD3g70
VFUNGo2Iul0Kool6l/f/+ObRsDKT+bG5PO70npp+0pZoZOerX7KdVBt3j0XEXfFr
h/YvYM9ufaLyL76STMd6aZuy/7tlRcYz9gVd16jLdb32IiK4+wUOQQJOi+ItaKn5
k/J7cY5NMYhfL0sFPuWHZsthSds1yk8QdejDkoPubCX+gIh34DFTc0h9TotafjbD
LJV4g4AVSQjSF8qAOhPdfbKBIz7M+ZASGEkZJ2bDDAMD2/uv9MuJY0euB8VHanhR
XmSCNOWYU2CGiErlTuAQShtEkjO7oDo0UGNaXWM02lpijD5dsBRvSdsfkFaNftj1
RS9M215q38BSE5dHLqe8cPCSdU5iuMgl4pB+nzbrbyHjfSja7yinjblP+ps+2zb7
Vz/8V5+ih0E+TWhy2jK+ANrUZbGFwSQDppO+OhcMeKP0nOid81HFQvNlqX+SM1TV
iJVtiVCBNCz4N6yKrdEcu5tpkV2vxJgSdKG/jqJ3Y258G51s+N0KsNdH14ya+d8q
my9VozuDtVIfQTf640Yf5Fs0STPS2KCZ4VSjs40XcVvoFGzVWJbvvpVY3fRZJfKI
Llsq5waRIhrJDJDbgCnORNcYY5gRJfkaBqux4GMN0Eh+Ilhxs5uEckVpOJSbJI9k
BT4Hb7zdDeJ0Q5afLiUlWDdB+WJ6M58Tm8W31MbNlb2XulSZ9a+ZgdBCu2QXqAMk
ZxjYwwlmRixpHCQu2XF18Qc79tz7b0VeZCes7nldDlvhA+2SH2pKd4/BYMg/JRa7
rIZUu3HWKWagyG0n0q758xfskkXfhDqBch4YybnLLzAsOUYCRqe7WMEjnbSCyXi9
Loz/v6pYhsB3e9DFYqJPZAf31E/9dXcJ4VVV0HM+F2rcP+sEbhxNphzJ5Cj8DuCO
HVOhi83sj/Kfud+CMaVp/h4kLNsrCSV4bWfYQB5eBG+u/dcWwYvuoL/4PKeUcqzu
Vt91w18Ea3tCFhPxOJhXa3/CyniGr5tCqyf56kf6Ii1Jz8dD8rya8PNRCbXuUJIk
My7qDyQixkeQ5ZWcqztLxc18Vr2YWC5K0/eIyFSsyqt5VT3a7Idcq/LeVLOQ5giD
H8DuXvwjOUPNBoy32Y4PVbW/yAQBbnzXN0wnj0S5Mh0qTPuZun+pQdkamjdcLwPK
aDz5X4+3mWHxwXvEAbJISG2jGpZlnGVcx5RjqOTqjtZUIVRZLgXvIXDpeO3Z51oQ
ireirQDMX7fRaq35wfQ7Qxel8uv9w41jY6a69CEwH2nPkyj48bUG35J4n6uKLlIN
UugQkdv+l9CpOuEJYjXXw5h6++cZgWTFc8MvWyTYrtYBGIoQls/NKXlqU6WP8Jp+
Em+ySqAF5G7VQ1IpAUDWpo/irlOOID5Q/+zsPDWAXIoARPbKocxacWPP0CLUfHyp
F4khoyKYR3Xc4eVQB/INkXaLREp3X3/tZb9hXScPCF56LCSfJ2Z41l42Xd1I/F9d
pabtX2eEQaGBJ3QzpSLmeD2d0QOQmWeZ8texGFVwQ7Nws7JdezyacJRfJF9w+icj
Ld7vTSkJ8XzQ76g1cnOmoWUTzge5GHiVzxd7c7PmZtWah4dUAPZd7sT49w5MX0EE
IMmCU6DTFls+iBeMylma9rW12pAqZRNrwXSFBUnfis1HLVo1jRE0YO+f5p1+enIA
vWatiPgXfa0JA0XkmxVgxv8gDCclDNOxXV9t2xRCgs5Hq0Ol/NMcU+iOwS8yWCK5
8Y6Qx6Bdi1DYWHltxLEJDBeZmd20VeDkFV4IungdTZdho1grh+DFYt16ntYm8caG
cvbuLXkSewqMhQSoyNnpn6ZEWbCK6TXPIOp1DypivsBxQVnzlu65qGWb0TFo1AB4
A9yO9RwHCB4up6wzCR2oGPtNOjBZeDfV20WRGpwD97FN/fq1g90ywoIVgT8DyXs/
oP4dC3YZlaxvYfS0GcDPVQXn5r0x/f4sVKzuRyRAOzIa75/aQQ6HD37ZUFo0ccng
FbyzCyO3Ll7tR0dJsa+TrzmEJKEtPMcq5TBPk1/DneoF2jUiGsEuylv/ze8cbsYr
t027FdqJ6vJWPq3u7snqlQoQY/ccXG5xu260zvdNrFxzg+iRC/R/L/lBSFSXsR8Q
7URKg1/Mp+QVsz5AkKLbOTnhLvmRPAQkSuLnnd2VNdrQvEYzCszbYe/CJ/Pp17MW
iCXKoBXHlmQuFCGBlm1n88gytwITQ7bwZQuza8XEqeNDxUK1y0zn8sw4K7pH4eeO
fgSpjOQUlHx8oBmtODioKSRsm/T2oWDEDywy9WLMbJ11PW4kGiu9RcLJ8ExGB7l1
UKAmDu351YNCOp7uIe9p4keIaotNKJu4PjLH2LejXddWDGC8iUai3EbOQW1B8+HZ
xYm9GVgW1e46y6gYkhtVuMrl5bFv/ek3PVz1cLHG4wOffdYznio5//YQwDbp/gdT
RcbF8roVr8XkciX9EHqJICUE5RM0tnhDYzENKY7eHjaCn/Bc2YmrsOKLQ0oYdZzQ
zmr9x5gv4BbU8voWR9daH4CgcDbF/5rmigiZ8yqrNEWwAaeXCHUdV4H9GU3hDdVr
Z6ZLEqCw8HaLXAQZZwhBNNEhM5iuCq/ofB76kofGt5KjreHeBbYd7URGo1tYgx1a
5l6+7IaftmVwdiMfKnkb46HqnqWwM2gvnToaxcXwHn73/c1nnB3gjBMXRcHdo3xK
RlEupeeeJdloat2/qm+ZUo/vOylGuD7L0aOtxugRWiHHbnzSrhcdrWhRGztXLbOG
Rvx8Y21eP/1hPplKBlSt+dlZS54En0iuINHXfiaJ+3qIYAu4P4nTwVLCm+S78d60
Iq3rbULQh8qdyYwZrXkCTdJdXYFv1u/DD/VRg1uo65t2QOQaDNsgkSJt5IcizFyw
vA+IXdjs485/M9twjEQDdc96sYFMQQIOtYv6azUWG+5Fiq/aoGmf7Aa+6NgDOgNd
7AmsmU92w9KQz7uJ/oCwTVU7KTigxXmOeJGSP1P6SdgbIidDQsn5bUPec7CVoAgq
QTsMDhbHKZYKZ6JEBSH3iuAarx+FF2dV2oFtxStPLV4VdQOO8JlToZm+c8iGlBJ0
dTJOJIzttf6GozydaJJfpEsGsW9YXh6k1jcHiv294JuIFphhHr345eQmYLUYpOSr
Pfkmln4H48+dzX7x4lLiM/QoCNO2uLiwV1TSAhW5bMiBRwLwsPikvrFDtK9p6tl2
baWCUZdcZP94EHUp91sr+8JUp9yApJaL/N22YYEHYhA2B1t9L0tQ9TLhQCy0N35P
FQOFSV4L+zvmzCFaOziweCzI/taQl56FrFe7mSoLYozMKyWBB2wIBZKJ0Apw5Cok
hA9KS2xMQotPl7D1dTYRysOE58XmQUwn9Tkuf9hwL3/o/faGQ/fSPNbQqrGdn7df
JnekR0P34KZOjx2LV1FX0cMjOeiPnrtSEKI6r3nRtDQZPB3U7OWxt/6KrZo2fAos
Co1qD7LWQfWWxnvvSB+mdI8jiEfvlzjJpmHaPTSscX9URf/sSaUoKNUeTaY/LFMx
FGdL3/UAdcqPY04iEHIyZQ0/9twAJe1sk0XpDpHjT4LA2c37rROYdPKycNj6fNr6
evMBelj+inylCCGPuvOtNuI3umseaK8RqYa2kX9k1TZ5fk1JWWbkLkuTVDnTjDTB
LYYaQhysxslOEBiU59SDxc5HvTyPxFjb0Nr0yYtFPxepauRXdqNB06Yu7+Y1EJO2
cB6RljfoYGWY3xc90ggMQtx54M2hgd/ywhIu/ggfrDiQAB8MXDmM8h1fmSmQ3Ydb
MeqMuJ2qkCcM5+uyoBYiRbjmauQtu9q/kPxADqKIfnJdv86nRSLuEznH8pyjrL7d
noOMdB4FgboDt79GW+nz0R7sbG+biGb24C4qmbxh0hwjUUh72JD1ezp0Ulfhyugq
oJPQ5gA4d5wioQwNygLyuf8HNm8of00S/uzxxwvF+wR5+NZcDhOkXjp37ZaEQI6w
RcuqqU9NlIdmp2XGn+LUwzXXRBZveMjByaOG+ST+OmcGbsBq9VieJyJsWr8x0xBN
3Kaawsj/9gqKV7KR4zKaQ10mlx6+7ng5VHL1BhzdsgUO2WlSCAyKtb6QYPUND8ps
FGWDW1r05Gh4eOffw2cjWwTfoH2iNkFzmWbZxdBKXLUO8kGI8gI08mFByaUFWJmX
gqhZgdi9G/azwnUNcIGVUZnHXvvPodfesIUhqBQ9cIx8SGxbhnq+nF1jYgUoYaaH
4Ymd0Oo9lrDc0RtGT9Wl18AmvVg/xpLQpilr6xeUU/G5MW9WqIHaNLY91PHQtzWR
2ZcLssG0RzMPsCfaY3wnzr36KV5XstF+iP5ijMLesfn2vzn9HMDNjq/Bgfs83Zh5
MQPAM2nPBBY+paiZb4vjd95CaKOi08SDSdFVovUmDONeYCNgbGL2gezjbwZysBea
G86iwEKtoE0AqJPycuPXPR3bhCuF/eVnb66zL2f8AOnrqJVNQNZTWKHbMRSfOKXL
Rek0OmzZ8K6p5wdyD/25lXQkWg2GRgSgMcY80HUlvxIVi/WQ/Tro7lLhEOeD7bvT
s57iTyQeN9L6eTE+M1prGsTwLfyWlyg/oGSlVXFKLYYggMsIJlELmeB1u5kijf2I
iaZLjwUjTKan2rWL/no7qRcMirzfwOcx4rMaCu6JLXN01YA+XineNJ/yRTmSjTgP
v5OwVk0CGb+E/nOeU/0B9dgBACkvNh9yg7FO/GQqt0JjJcwWOzz9vUWgSLL7zLC5
Q/TTGji1Cj2W7VbFXHHKtgkDoHcaBNWoZGJMMXNnRvCHMzM9iGcKcD6h0hWz6XRi
MAY1PpknRurigl/FBSKvXusl8AfoNWswr8VLAxKmaSZ1hLf1V8poj5Y2OnA7ntTL
lbvHJ0DPfo8YbD5OtjmQbV0H3grTiz3+p8suvSG0YDUZCJzPWqHxv9i61SfIsoaU
C9cgRoxNVjETG+yyqYLVfiK0vkOGYZH6Z/KoZvFZKcszYMdvFE/TXlCC0im8xwqn
GOyQ81KygUKRxmWYvJ3gdd99dNQ4FXOfOpyi5sdvYGthMnDuie6APeB+gFZPlezk
t/JSiOTDPRQJ5tmqELRWom4sl1kSNt8ww1HIC5xLim2O4ygU18qqL8Fvi0qW8eWD
x3tiXsWGznWPZscJdKoJMSmaAUcVjDXdNPFU9G7gA/DrnK4X1OeFJtAWuEbcK3YP
KIzOcNlB9ZDxUiKR1Af8zuEnzmlZvJvl/J6BNE9eG7sKcc/m78SRjbLvY3Wy1Zmz
H1h+eEqobgvMqPUFib5EnU3dmD+1YrBrPOlHwDAv7+L3GcFCnorZ/KHRtcJ4RvKt
6fPokIbk98UWqyL2p1tbrTGXF0kyqFPt2d55Dvxva5ByMbPFPzGjB1JwZbt9oQIm
Wb5xx5xQxYLiVIHS0KUD2O0Cdj0W6ZBugVNEj/fqYOtyTj4k5yaEpsnHyk/+Ynvd
sBU3vcB3gUCip/DwBhzQWDSO4nbresBpNUm5MDpw1XZvnWlIMRZDNgBXvgbbrYTW
9EUp/s1O4F4tkZGgYIgr4yL0BZZwOZ8tw8fENLZ+moQ9zJuWWaghspnRhjQnxBLX
zX5FWDixNrwxn/usNIK8VnCfGn58PZMsm51Zp+DUKe8nl0IJz6CEZ59hRW0Fh4iF
ArJNtaILd062yK9jiXAIfneumIfAaReMCQvnlcvwfzpm9yvSEpTyP9TlrVYJo25O
tr4Ra1m2jao1k9RoRh5HTROI2RLn6zO8f0Yw9afcGjDDUkFxN/ZIGgjaeeCFAe2y
EXS7qsNByLj53PSOMu6y3fSj6wc8YELYIl/YzQJAikekefPieNBTwNKHnd3NHlUg
GfTxJ+ueedB+9OkvmT75rtbXp72c1nyf/S48LH22PNbQzHAgibh1MaEaxaeC4BHg
ZVSezgVp69LmW2Ij+W965pnwHMT77/rk1uYkaJev2nTLwNGwc3PtC5Hj0/sHz9Yv
yHQhT3ojZLWV7+fVJZknsW8dqezqc4TlWli7nFaWdH59Ihs7ipVwtjDj4VSwz0nv
rsFykTwdZN1uYuQDgDBfbbQjIqUojx1JGYzuM9EiSeMKJ5VQSR2Ph+U6PI9jCutU
PWC2NvQa2ZfcIwp9AZ020/cw0rlfViG2qaZKpcBIQDgknCzyrBWVje03d0TFIq1e
/1U8nzDyvLGC8TslXYK8xkW9VH3eMKM5L7nIgVG0nV1dHJ/LIZgn84KbrQewq7n9
Qe48C2GWJNecPWr+7MMPGNoklu7kADE9x4nGUnUHfC5w0Dm3vBN3lR55jU5KiHmY
msCC+7KFDPDy7ShTebahupkxQOyKmT3/j4DAgvwMlhbEQSkM0a/wIhnTTR72mABw
8aGZY5r2QYketQi3kuAhAsZQAit0Ep505Ym9g3bONfEjVa0UUJSaI1khwkARFaBo
CA6wiY8gX98zMkTg92c2ByiLqGbUQtakyLWJyczeLQpc/Qnf+Sq/Ibl2O7656/b+
IR8bUDq63/hU/3QYkWuyO4rGcnCkxCcKhACSyIxVlrXiJO7MtX9FvfP6EZ6Y0bsV
SXaQ78tH5z0UGaS0cvTvnEwBglta4k0TTj2ho6RM9OYkAIwl4UZYEM+JUW5IPhIC
SVfbxCPFgWb8fcRPIne06qAOEn8nQAEaxvms4YimQssyEW+rpqWWEOKL+Lxj1ziM
UmdKJATwANGfSII6alVYoDzld6VZO26nf/aT6Uw+NglNrYmphfXiS2Kz5W3ZyOCA
E9UqLjl5CIksdNCXHQyZvY+SREUZrNUOqRxHMyynEi6kCR0mwkh9J+xSG20eVoTX
5lGgrxhhJvmLixwDPlPKpu8sY3w/AHLI4afA9TWB8fnD1cIyntRWctzCIjNc6ef1
N3Sok4qTq9tF8kFVPalQvpKtDAZPtYQ1GD4iKw2BZ0Tuql272OvMIDmiADkLEVUG
YmhMlTDp7w7HP2GWB4YK33uD2bZJQW27LlROMO6AMsTK13DRbFyOWH5kxKKq0rif
SXjJguBVDwFPoZGqy7/7VkyZIAGO/RI/UGR/slWyomxpigyINrr32KaAYzkap8HA
zB0NeeQTvGrYB8C7qLYJpVdQ/PReWvgc9qi/THwxC1qTIAs3mzJOCdTBX4PWwLFj
7ynGBUrQ1MsZ4k5YFnclFo6qxfk43cHuR7qw2UTF3xe6+fGxrUwJGFiDJ/jden18
viSx2ULzstetGiLKJVonj3Ve5UGZxH7zxxBpQJQXtYHhL1WQr0xgy4/9jq2GSG8K
63KF2knU9vF8rD8+myryhGJeV+wVj+yLWLzAqZrUK/hqx06K8B6XZEKUxIiW2gGU
zw6DkgwvPAAyeFxLYhHBtSSdwMjDemnjscas3OAowg4ONBYZ+Bu5ZZXQZej7iHvn
FbP9Rh5vnhoSdFTortJzEhCo7hQD5EEdA7NdvbG2qwOiDXTFJkln4I0FDir3pOCS
IbVu8CFowkjYari6W8pNTqOaGX+1jScm/QnJQwR6m7wrwe3I+Y+rSJfHeUJ/I9Go
4r+gAWb6XmacvL8Eegl64dgoRq547lLx66zUKJ9Gk7LZDlyGJBK7+WQ8A1oWwhFa
UMgXtxh5yVswSGQ4TjPWLsKyTt6mMq+CPay6kGv4QGvHDRakPfScZAq6dGhvT1Zy
aH0CT/gD10TTujAurtTGqgkN/HWpYubBWO0plw0NmiF66fWiyuVonNtT3Qwtq7JE
iUH2h8X58+IzlL22wO7Of+eEToqQu8am6sINlRZolEQxq0sV3iWKB3zwQ6wXOQ1O
BA8F7tlTWhEKClbR2U1hBuDk1jGkl709UYMjFTy8k+115BZu4EGBGeBoFsC9d/hy
G45pvvaNySAxy1bSS50o69fo3IfAHD0YvYfafP25QkVP3wNLzIgqk6gXm41wQ26U
v7Ng1oouvLqIxYttx79XUrnNUSXgpB65IsLVIOt7oeyQJlnoVdxIZeVmohPCtENe
uSvuX1JQpbEUE2BVd6o5st4A+xpx1Rq3MCC0zNT2DAUVAUbitPLvEhpDWv9J9mca
dt9EfyRs8OHb7m2dgyzRG4Dcbv7ziwsviMf9Y2QDBRZEc13Xfkk4ejVjf/DknhXJ
D9GPXhQGrYRo/Nu36zVjMnBGQRKWoTDmApngm7taMQHsoku0tUYYpaRVTWOkhC7Z
eASq9SDTKWssY/jKMu4iQRQrc3nsfD6qzjo2lSLDpA7Y9rQ38y3uabhx/6oViCf7
ThMD3h9ZoGqYbVWI+zWjTMPF6V6JgY6F5waGIk8CzN9GWn1gy+sgOcuJ1FUYbRij
+RUrbmtc/2CbN/+6zj4lpkqm4FHkC7aR1GEBsIlwo1vfsxLfz6zYnG0112S+xORI
vyaJ70qWQTfrA+vPl5Rbt7LxzoL42CHhtO7UDyMmaof8WquXdKM5P+dW4O49U+/W
pd8w/S9FDhP+UIie/FjXt6m675H1W5Nw+LaE22HDEKYrTjTRZIsGzduRBTymicWB
44Y7nt+4Dwr900w5JcfFaSwBhDfr6fTUpFIavWnUaVYDkVrdO8cF+M4TJpyWWV2/
2DjjnZVLag1TcwRHYPockqdtTZERbp3kcIIS8WqgXvx7XGA0hvBnaG8p/LMePd8W
UCAVJIoCbW2A8n9pebkVnlju1ebG4K0XAqmUbfAV0r7mEAIyJvwXGogCkl0+ipwY
kRmoTCFKLcfT9n0OpIOVIfbiuoz9MW8Fw8vCXtTdW4z37H5FW+zpSzkiyknGyEoJ
WyWQhjjENMCsLVSh//Pil+ItGQXVCs658vAuPaV7oRWxVvHwXt/IYCTIv3kbCp9c
Qe8yaKo9hCcRWNYlkjDXCzXAlB0FSYQeM2JeJRjrvKDx/glszzZrggk3e6FoaXng
XhNtsR7E206SJJlNo7r7XON4enrp2yJee71kYyuiFwTnkjj/v9HcBLAhdVZIaSqy
mVFSAetZJ+VYJ90SwskwF39gBp33r4iC0alaAAkYT0WD6yPZ1OQyvHcNY7PqePB2
5HeHe6YXVeuxOVIQ6mTdLLSuI/eC3E0C0M3MevP14M2wpxZjg/JxBUUEcMXMZXxv
B5CiQ1FYMa+rXXtJ7WBmBdIkGcQfmMWnweklW7JOZndGD3lrWNKzuBI3KpgcyHiD
P2l9Tm77peQZsdqdqe5i3ju+lqX+Ln1B3OgJgaZXg7Brnn3dX4RoYB1HPfwH8JVs
tKaGxpcKiayl8r+8B1D04lJ6Kcy4jKcBMs9k7pC0NHIVMuPtAeyrOi3DHzgYtiXO
NePbudLnpZgItoMEXPepgN0x29LqsjZHMjcWxqg/rt92y7E37Qi2n8q5fnonBKdp
SzosZjXosmSvvMFa0N1P9WsGIlCzO7WF6ysk5rxc3fqQFNq7gYVRlVw2N2H8Gx/2
VYci7HK35YzLwIBoSP7y9qKdA2TeJtxxc7tOCVTbML6hw8fiyzAeRmJT2PoaZgDA
jz7IPuyBt736WGzn30oykxx/jLZk5bRJaA0YTBa1719DZRQjNffN8YLtSLmgn3Ae
h+aNArUSPfpgs9bZG4mZKkctQXtI2AujvKVQYkgmqtNUIvoBpDICuLnHjM49GPrG
Mt8DXywlc5sOeIcElziSzuEkTJ5UjiFjIJaCl+5RtZz7n5Vyw8k+C1At/TlnlEbv
kqGkbpNiIFsk1qgGmw6M2L0ZssbAM7/RCNeD0Dcq/VKvGVrCI1LPNa/NjbRwwA08
oXawueuuNdRpzqpjz4wzd19pPP5bnwd5nwEDgqYM1bIDoJcjB6FPa5mEwk0O7MJn
suZJcKh5PyWWANX0JfLRnnQghfmZeM6q9upZhwIiALY0a7hFnGD8bnfrhspNVwn4
ihxZMFPhrgSAWyveJqXdUvq32uJfE34Jt1m7ZYUBkk7qO1msO+Pc1GK16tIsDKQN
TSbnQFCAtxBKavAzeO2sjSpR+PKgZO0XclfuPUoNIVq8X57w6ntdTPcZWHpXSZRz
5ByHg1NxEZ6pnLX42EA3m5q/Lcwkxsvtzn5HhkMI2fU/s/AnYFYVHsgEqlK5LI8S
3nolnhgSSw6Hp9lrfs9yAZgFexxKqvGrhKntagn5/a2LiOdhlY/zUfyEtard6jvJ
iDvn1B9lkWYu8UyHFw/pc4xY5PjJ2UOK1QyNqiymj5N9VQBOZw27WjVwh6dO1fUf
SWhNmU4KJwwQ5cxba+J+8gVJtmducC4Nqb+tAyZfy8OBiQW/Do5of/ihFlhogyoZ
yymNTLdz6wPFz8690PrxnHl7JBt8zAZynSDB1WQ8UiQv6QwxJRBuKm+WQoD7oIy6
lZwAz3NxtzduYMyIVG0a1kmUFdY+thInwKnqJjAhHJXYgef0AWO+yNSag7Pchbwz
i472XdbH6gldVRnVpD0YCOdxbzB1MLnqpmzzdQOhjQOewFIPgb6sLcNApPNxYqw+
sHcbystPohTmrnd+qiPJWZaP4u3XGYin4FwOyDPcjphUAbMQXjVdrPMi9Zey3OU5
3DZ4GJQLMNnEFSz6KXSLpL+tbQsfM+FuOnf0bSjXSinzYNSAAi0VhC0UJMRGZeeF
qLe/AMO069kntue4AzvdLWag7EFiwcsKFF/3doLD/z7el9f7kYUMsQEFuuCekLoH
/k8byytEekkZ6mcMKakkBR8uWDyhq8r95F6WTdXPdqaHq4ZPkahsRfwFgpkx2v1+
mjGOB1/KE0tsM5VBABtVhZT08wnVz7BEpbojXF6eki+h2LZ5eCqoj60IPk5tUBX4
tTf2ar1vzmO3lSRD3nSTsPYhNIReZOQda5TQsK0HcqQlOktfMW4t2fGK8bS3LF2n
+ALdPv56tKlfAfQOxsrrxivjSS7HojMpHpLJrWMqN3oXwGpCur2T8JIJErL4RB6M
R+of+gJEMFMg59cJAswVRcWSZVryB1sfSUrQ2VFW7qZ3IaLZ+w5NhVJP130LZJ00
1FWAlJoMkRKWtI8inXFPJ7kQ6B/9MT3sWpV9CMoqkNj5C5I19xu1ueZKMrfog8/j
7K5cytAXTzlmqEp2PsImMJ6AqglrbzkUmv+wgDglxmT2ccqy9U7gmZCn4fDXPKU+
fkZBmoD7zGaArCbSXQcBQcnAv+CxkfQ/pl2puuQX5z8R7QabSqeG5iT6JABNxHJw
SU3yQxxj1hw5DXUTTsiMmKoK/xS5roOqrQmbcnRsrtEBZyMn+6JCQ35tiUkI0k/n
KobniOaRQmmJXlwa2vfIFcZozzHAJwoCfsRnTb5LtI9n6YEJ6oPDVqHbYx7yOuxW
bvLCpWrKIileUhXzygDdwSW/MUmCeP+IkrgkB9kCPrUG0x3EzXpmbodq+C05ZxWP
hD0UtYyxUgGGUS2YuydAespu75ElPXQVvpMQljZwqowQoeaVnUvkNo71J5mPEU/Y
wZTdZT9zgrXLLsQgy3YGSSHDlqCP8Sx9fePgnaaqcblM8/jn5j2TfB+TTD2Ij5Ya
8WauGub67pGNQt9IMnORFr7xwNx9gkuTpn7KC8AjBmr/2C6q/UqIUDLOp7GCa8aA
EMwwYt8SyaLPJDwHqL0Hbg8TXiyq3uu3c8RiWFFOTJWVvo4hN26VOXzb/7kuPo/T
7kQteq2utHx16dxOhopUY0Wc5wdNzKC2ukQlpIjGVNwOqBVaGownyybMoRKXWsF7
GVqxtrCaHRgcRnKqqPMmD4TBZGrc/j//V4Q2x7bnSWMPmlt3CaIj5C/8rLKy0qy2
fr1E/D2a/pO+F3WFcy4bjydGqrvlsMAUG3bQ0aCiPI4PikoBi5pYyF6g2hzAHCP7
ZFgxAuDU7iTyNR+7BSq6hWsXLl3/mdbXkPfbhyIH8u71KU2FLovQc6PMqcTw2c1L
PlFEsysXWeSWn2Q0rPmfAhNlODe806cBGpR3mJURKCqXjaTmL2Ukdvl0lraB1ALd
Xg+O5Umgs9agTMMRANjKV5zDGa6VN9KGgsnF4MaMUU8KaJggyXt7lJF3Ctj7IBCP
yzJe3fFB7J72fULcUwcQxCHCi5Fi882k0AYRvEvbSYiUekCzeMd/VV0z4oBtloRo
UGibjwqjkq8Ci/HnFRl6d6Q7ZpynwNrP/1emzZVVEVNW8i4MQ/HCd7yqxJWCuR/7
DWJHLmH4uFPN9sC8CopR+h7xd4p3yACOPnG8pxAjKPMbEph2w0IucjzZhz8aZ8kj
+6ikAFMGoMRZvg3oAGzYOY8ygyI5vBDy7L5nlCmW8sM7tZQhmm6lo95RJ6rYxTAQ
UQEGWd4GYImtA6jPnHwI5Ps60jMehnCxwl93KAkrGb6PxotnlDYgpitDZtU92rHV
OPSALV609dky597QljXG6zzbAaawVj8k1r4gCT5i6gIyEj518BEZrzamHmJgalmn
UFg35kI8U7oQQJ0Wd2PG10JoRl9SX6E/Kqg8IKPWZfLb3Z3vc79jcGjtbTFksDWA
mBqz7r7YxhsTOFzb/YKaDYJUcCGyeZmepNh+bAEw5JvVrJ4JkAuEOb9jSy+Jr2+5
Me8u4P9/Rk88k5Z3mHnQ49ikyPfn+R7AJYmFNcohZtMsDVX1SlyeEZrjOp1uagTB
c1wE2S6lOzRLfWqngMhZziTV6voYitLH9QIN6cWd8gk6kBYeuTqeZZH957nI+XiU
P1ww3HiAUWFWm0lxhb3Sxp3wXYoD9tzawEFET50VyDEhKRSbFB+e+CCQ3QTyLzxN
sytdk+9DjjLN0jimTGVYEbxyxbf3muAVsm4RZoCTUZWtaK/mBeLnhDo80SDjdAVh
StIVzUuuQOzu0GJ+QCCYurfoZA4M7pHUsMjW/daYL3MCY7XhypErtK5Y0YvuMtfb
TlICE4JJAyLIs3++CR0zNakUDLROAh9t1AAasCtRxz87QKjSng/VNI+7dEA3NBG8
MKJSq0epXf1os3TBjZ0yZqhRDx8OGqVG6XbjWVL6/28hdXt8PVwm+BmHPIMyUboM
iY65tXUqnAEx0ly7/hg/HY0MBq1N6DoudcQmd4ORq7rY6pLOB6/3xDa9wLpN6vQ3
KUvJyeugG0/6RV5nqdu4qawPwlqLxRcy2RaR0Fv1VpfyZ0erWNlgLMAun3Qbci6U
A0+b1+gXC8iStTkUAV8lvr4hrin0RutaJzEjqWOnMCQQKqNe5YhdKwEnDsl22Z9p
RihhvRor7epxE66vsPyq5jx4QaG5TyCbMGaAPdPxY+5oZVkB+HWpq3Qrcdc7If7N
4IALtOooDKgj3W6pJueqUfbITKi5xU2ftnhBDHM+Hczi0AY3aAoLrwB76oSibnNy
JNi85R6riXYYEAXqgBP5CeY+vetLAzZP4kA8AA8/awcaOU6iU5Gwb1tgfOfWGPwl
IKp1GWL4AykGFODNbGKUbdrlsXK8w8QwqxRpvsWUDGKdS3e/k0q5/3GCFndOPf+6
RVjliSeerb8hrOjerxmLXodmYyRUAViwtIT/CKborIk30KpUWBiqc4DS36oWe8pG
aBbeJU1vfR8nxlZKwldXVoS962YXX2Uf1p+pbyDyPKJcPIqK2ygAAEkvhyWiXgdU
IhGmemED83asqXR/d3ihjkD+m8BV3OyjdTcVKrpwxIR2XnoWBuPeH4K1v7GgA7Z1
lgQhcq4UfqE9J7lyOOSETWb0S7rUshUAI7fsCl5meZTsA+9/syf/x7d7xKBtYr+d
clm5CHLwkbi1CDhmgzh689qBxzS2n20rjVcyPeggfHEotTPu9QDfIbOkFK57kcWd
uakZbcMjkWwZsTu5rBOb13+Mcxi9ekE/qaDOTHpKHKm9NM20yllxYYG1hYyKEEoF
DsqDcp7EpeaZohR+5bSRog363W7uY6U3L0S8IbNFJbGQJCIUdHb7O5HIAU35Yl7u
2GLBLrXcdHuhmR4ZNu9PJyqKg9SNjr5idSj4oBD7cdRfpzm7B6nvIN8WZFYctZ7N
9BLM1QMybuYtbnzJWSlp/aC1vvkKON8Q2clydZ/VdhCQaaJWrX4J309K1S2EqGFc
/JDNYZavYN2S38uBhOcOQprCoBzNTcTW7QcYvUu4eB9R8K7cl8BET4+jftEC4/Pd
LjUufaFoGsQucWtrrGaYo5FzmFJyg31Hs+vXo1i5Vvj6/GiDrG6+GBr5q7Bs0fq3
tyUwtOKc++KHjEVyFTKn6pG27aYH2U49PAu+RAi1PWJLmYV8gLFAfL7jeq+iAGuw
CwiE/rsPVTzujvItri+33rS/REpDBRYviEXKpV4S1DXkSm7p53TsgODz/H23JifL
4iaW7koXJgMUD8q1Dsz79duXOxA/XluWSXMDHxZRYDG9gGRGJmO3UzILF5l8DMEa
sVby/IiKgpYauBdBvLuj7ktstjLP7YKR5glT8BPiO6AGqnm2nBzDpvCAM7pD1d4Z
IGON6eZDXgprWdC0HFm9YduiXh7K+6pKbTwyGFQ0j36XRKN/1iNrfEZ0N6tCogWf
5vvUGbYx6er23bJsQ4sVMZwsjIxlYEdjE43yopAdxpVNRzbQVs9oLd5I8KLUNQp3
+THqjHeXj34tN85Sw5kfFUiqrdYxtFFXaFTtaHcmm5/WcDXSsV7ZetU0gzN/o01P
RkyBjN6HxGnbgVWU+eCy9F1k/FwRsJ2s0tKmqTxyuLvs3oAUiqxvouNlkBCyFhI/
ePMlxGbyCtDE8eIzo3xfg0x4Cvdhe8jrZ7ZK+vIBCjuOuBb9rEMNUKVtmd5sxBKc
7l7+fFblQLyh1BTxR+rysKhmL9M14EyGoEpW7BSl+krrkbGMPadLvLTCq5OuFUtx
UCD6CGMLpfq8iiA/eCrix0rOr2soGSY5qGxNL3Ly7YMTY3/hLYv6O5RJ9BWJptKi
9t4fa2D9F2xxmH3w31XdXfVbQXJalM42sTYO7G3AjByIWf9InzzBiTKtfN8hc931
ucRHXrmP6JnvPzYTJhLLgyX8ci3W99P+MVWVfJORH4JmCx71c7qbhB4g/wyz43CC
j4jydZukPDaXgtc3VTAV0bhPc7r15sKzXhAaNhtm5UKcfpKy9CGWI+0X5xfYz1jL
6bI/COfbtMci4a0kbcSSz68awCy89cwtstiF+ShaBHMcdu0sClNa1lEFw4IEtAaf
gGK0wM2S1tRfLYMxLCxlaXEiidJi2T5EO5yetzo8NXn19t3r50FdCny2jzDOZjTV
iYaEbAOQM8pyoLIAVxyBXEyOMnUNP+7IVGpKFzMcb8oHQ41rHWAJS81iv2yKFCdO
URtdZMoWDqE+E8jZGHh68cGglkawgZhIhICuHTr/74Y0T6SlqdlTD6yafPN5SLkc
hMKpue/n94ZMAClHir0kRvPV2yzH+gZbJaqmD0H8v9pSYJBUO9WfH/kAg/LPri/m
vdSNAUVy7x8Te+oiyKSqSs1W4h3w/w4nMExjeWThTtbfbRKU0LbpgWfIcLTwxohp
CaFJF5G6d3FNwIzz2ZFXV2Ig1lCU1Vv8/yoEjjPrzQyr3KEHMLEi1pmSsB7GO4/9
zHJ74M3uZMDI0qaDqm1fDKYx8iOf0/mFnEibyRPzerF6C7SG1TNrgCkJnVTzxop2
E8pY4RRVx6Cesp6Ys9cjyHI8EF564qjNtwgg07aA2f4QBvtGZVEytWb2JvZ0Bjak
mVeVVqQw6wB3lUiP4sDD/KiIhVy5OXDnA6ZQz8rMJmZbEchgMJniNrDtP+Ho9vGO
x2Y7xjUQ9kD0zd93aqth6+3cVbxO9Ki6SRzbEdgnw7UFKQDQVVAfkzr3JLIe48Ee
ptFQijrHnIoeS4mHWr4oFIYMSDgW3TDeMEOifKLGcILoi+CICqqUBzShqs9volmC
XyIXNAX1lb7TSmLSb8BXaCwNshh7+jaXKYEffG6EruIs7Enc/c+3oQpfrkHdnbk6
Sfxz6SsvS5eWmGHJ+Rg9xJXCeZJnlxEK1Ai+/EEyTkn9ZR4NisOOd4AD9J8KQwAn
Sd2aiAs2XshTwW3MUNUDKoPH4PdibHs6smcGvb8B4Zcle2X6Pj5qo4J+UT7PYk0w
7qgX0nBYvsxLpyuzlHSFhSmJcb7fLnm+WsqHwzLCYwuvmYX3kPEB7Sgi4sA18Aa3
29rA8EJcg8AvwHPqlH/OjfLb7org3SUXsCN4Grc+RnHwzV40LrwBuy5eoYxgS9hy
mKMBzOGiyABayC2RGUcEHqdaerpFvohfixm1tt/fdwTt0gXl2t5ELq6WeMvKO/Ey
2b1AZ4qy6LCN/qxAIBe1DEKEEFnngH2gHmCb+CWyugXZpke9cbO5czFTdHg82DYr
Eyfu+vAXv/8ts94hGu75yZJDN9RE3JwjuJaq9A/mp2sXQ9uaRRJyRtDX9z2nX+/c
s/ImjTTLNvNFS5LW7sq+GRIIsZwGVHROpazpPQ4x3/L8eKtRcGlncmw+TWhgTntc
Rfl5JP6NHCDmjGiRLdpsjXEgvkEDXmn0GxaXsGQgBL0N1FiBaBAHQu6wNz8A/1uA
4bCU2ZYfJN44l1pl7UJDfuYnDw3X/xkEGxKZGw/81U/6iVzrSh/mrB9Ab48jJavR
vElVTF9/srPsI2mQm5vZEcJK7zsSyeQSq5H8PB4YFeLshxrNR6ErGz12smo5+f3y
zEw2srKVuR7vZJ3Ln9LCgUCSvvOsVMDK3qQJaW6bh2sNPQ61J/2njjn6P1pTN792
P8cYBj5F6zfl2FYyoFjBQE21a36Clu+1FyAqM5K9Eyb4t2gMMki9XWn4qQAy+iEY
wclzlwt17LE6NjQ7qpt08HOb0p9/mUXZ9D9MrjiVhuB3aQN8YAXu39rXD00QvDWn
8pBqKpbc/lQgh/SJXOC9IL1s1sZMozcFkXcz0xll96wnKLOsOPil1rOHY+C4XAlQ
zVi9TBbTuXb2Lgvu9pyftzRRdf9WPvKecsbSUfrC3xMYoYEqhtXFdC8XTsNm2WqN
mXkwiGrOU1Mb4UQNDUA54VVkJcfVwDYdAftJ7xuTh9oeSRdHzFui2ZKCqEdQMd7m
eue5p5+xEwc1k3quwxRaF7ULE0CWN6cE5Nk3t1IxlPhhJd+IlAV5Wyiir1enk+vh
Al5GzxkD0Fge3hhRTBcLKKi63oFnD7FRRnaLMVppz5bfQJoSGVbZfrcCibuQObUN
SxlCk+I9x3axMisupI0/Di+jA6Bw5h3cBGOSm0ZdRGFgMd5fZDPVMxEzRuKvCEMA
hGmou0dsKZE8Zy6LM5Fy0wyGZiQ83rRsFhSF/BplmY6QJFtJt1KgVeoRPXbke5NO
n2UcjDF9Nj3BwW0WjOnAowgYqMblRguAD4DecbpGF4ZwyOFt3ddhaLf7GhDjLRtL
Qd38x2GncbYhH1tDUoI65HryEoULet8JRK9QyaK4jWmYlGBlBoOJq1AgjvTm+iZU
0JWEx+o7Jljfrto4fDGPyli0I1lJUsBS87RKEKAydh6Eu11ZYP0TiXJf6Wzm4OPU
FS+Hq5xbbONrfnOS0dBzeqQ2VrUIutid5s6tbNtl55i+vp0KN+ZDujsEczX4MSdI
2iHK8i0CV3yohcOHbH1sS8nDSFtlwGbIJ0H8B0C9mgi1XENR5DQwQW7n3yJtWcJk
Tev8UoRfIlAGjx4hjnm7A6C/dFnKNY1Mngtd23oHwLa9n44LBP9gCKEXjXg+37kR
V1zYw6CHk2KRFLGsY7slNNUQstGc5ez5B5oTwPqPRWmIKTM9WJKvG5zGbvcmtV2L
baR4CvktWvz3HA6T0GQpjBeL9FkloJgyD9P+W4f20H6IrwD0TssjZfMAtK0MoPSZ
+guq+wXMOZLdPJ8ZHXnXCGKigNaTY52U9Hp2yThqX02qrOolkyyIQh5aGXRvtVOL
99u0hImTxxXP5ZpymbYTvlxRMv+Rsc0bDlSHCpXKzyT5/iXNSXR/78JGaJwAxRW8
e9MO4IC7j2dxsk8/Qq+5IKPndCoeG+MiI+ez4mN5HuZXaHuMiW0ZoZicih5U9Hee
gccBU59M1xN4+NvHljc77lII1oySadgWoZ4I4ZvoNb4jDZ3dR2kJUWODU+ZnnLdb
SPJPGru59YnAzhbjmbhP/80US87rw/6z2m29ABohxvGqJsnO7LOYazGCpOPIIY5B
7ht53vbWYasy/rER6OIRENB3FMezZp7ed5b8ez1Te32+FgbyZEdqqPwB2Ogk7EWO
UGN/+cqPzsZM9EkC1rSK3hJeBa1r2/j8I9g5k5hgfF/rQPuv2N7HeA7jqs4p4wqP
8ngMjGNOeroI4by28/Rx0bU1uQSpN+46v9Us3raXKIEcwUvXibbOqggq3Sqfpdnn
yQN+htcWeiRyKaz8fVZlXKKBFA/nEWq7P8Nsey54LvgijBtfn0CzaDqk8oMa0lDC
bzUJ9/wOD9M+i41lGOAv87hvdPfz2fsRslh8TVjqEbyTnvMCwsT6LymN0dH/WLTY
Wst+jD0kk/duE0+300CxoFo3zlrL7EdlrA91rziCfbf+RhdblSit94vj3Ilxuxs8
CUSubcDFrLHDYgacOSUnvbuc41T7icgBx+Q6eWJoZV+jIfdinuT+aYvX2kf4XJmm
q6AynWH1vLIHOGdNI4gFGbf2WA3xSh5/gQ9lvkqJ8/Unn+gOvBOvd2DZB6teeYYv
0oNG+w1Ear8xO8FgUddS09prM0hVW4D043UGfxWYw457egDkjls8+itEcW7ZOW5l
J+SglwQ7lhA5pq6xg9rqFwIgZ5CUlpbTr3KwlqydvdlWlYatL3ktPqDTEOqV59Rv
HLT5vnhG385C5S+AyUUpUSFVc6A3mDjOLcMqiFyF0GnBwlK3LmpSGwOn0kTxJnzC
2VDRdcGZ3tKS339NQfkhGgE+n/mWtNFCYyeMLjZTw+yYX0XmwBx1/gRJGOqBqmQd
TJF8wxLJELsFH+Lyki0qK41GvqC68/OpUJfGYY2WCvcx1AsyXHM+TW6PNrtN2OdF
2t4P0/OEeEpt6b5BZIPKDtatPdANDY+9T1HZgtMzUYVdVrrBn3nPc17dV4bMXCN7
YCakUZfcn4RwYyv3IlyL229X6o2B+75jp/YLlPM3oLSK5RrDJ1NVQjxYkHn2RuAd
0A1db69yPZL81EejV/ExrVDqhwNYp2qYgqIcPvdtsrJ8yio9XX8POwq5wT7y54NG
zENxo7VfhZ+VRZiOOV1KrZmy4qr4ltgE4Q0mi8l+aYMe94qK5NiHB4wH3xLbetxO
ZdOZMhe0q9oP6WvIUpLSySxo14LBE+UEMiePHFG7xzszTG+2SXktvBDuRoDCEtSj
REjXzUNnyyQlJPLX6ugPIAhpx/slpdMinmJlm4ywRQXuf2nTDU5BF4Xj8/g6RWSF
U739iryXWoB2YQaOdIWoM9WLL9hzEnt1CADBnW4DKN9RJVE/IX93so/ug0OmZ1La
m6zZnHU+UNDct+8ZYr2Zf4MJHMujHEAXdiremfc6osZNw6E9fVRGx0h2e5xDrDu8
s5vjatvtchxCik09XUXJ5jYqZbwU5c/GdSn3BFfpBxR8cCRNALqAjLZ2CctRHLIO
9rMK0t6Qx7Lx2Qm26tn71vzBWhzAiwBpiEWp6y7iAu5vL2MQVY+SBP3HVLUrakWr
RT8ZIREWguUXXu5IzhsHV7SkHE4pJohpLyytZdAwCM3RcUmG+vBriPddiWtNONiA
MKHHGcVJ3++Lcd7L7mEGoYIk35ac84EpP8AS/9F08fZeydA+Ne/X+4JfJx7y/qXM
QJha5ZMJqjvPSBApzmIR4M9GraWCTzRqc5avjNfy7s3MofoDQ7bBLdYXx38GPYeP
Uh1BxWg+Y9JV1NhE9ilFl353YJMivoB77nbLBsw3ptCcZJe60CS849nil1enFK35
WMaqIUVTYSpqh/G5H6SJWHPYIeqj+6nqsbqUzkFn6qZSOnOcsfg9Z7AB8v6hOkux
5u5lW41l++szAwBVtmQ69OEBtyuJP9NZ+83aJhItFX9nONV2mLcy7/OPXxXg0fyJ
G5q3nmG3ovnu/69h8V7VoY7YcZSuPK0hC0owGfGFUqUHXTGLji/E0S0TszgBZ8Wt
53N2Wt9+7JTMKJaY3KMY5yZKPn8DzLVOuISzRb8ZDezm4DEt7tVsSs4+IjFHQF0K
M5mm57H4AiqJNkytTz3pqVjtdWISE99Ay3B7pwqb5NdO1Y3mamg+8fJ62UeqOeB7
2ycwUqjeSqQAKFk2AvPLbRtFwCABIl5yKz7Ylyn51piJ4uZTO/vzKFFx9OkCbbdI
TA7fWwv9WaeiVMqhtJtQ9K4iPNCxybd+Q2lIlWHrNJZBMWKPsdH4VoSHgmJKxNtI
oU4jbdw6ZBOtT+4+9CKackVAwuL3ha/+cc06zjd/K0HlqDvh7c2XMEr83/CkIZku
Jv+lEAGT/XdHysadZ0xl202dByy2uVU6WokFLDRcPeiiDqAtcpV+IfqVjx7H7FYA
uFk4Qe+U+QEE0FXhLpqABx0awjaNfnG6tJS94pRjvfUti12lvzUogIHjkw3YiF6/
QBbWZ+6ntTLmOF0Y72H56Hybavg1n03D4S2IUXgLp/iNbHIldoIYQUvFioEwuTGp
fmtFmuryz9WQuwJ3azPviB+uYTd70Kj/P1tHCOtNu2aGMxbdpFPoVtzoGF5GnoJZ
CBMLEnn+nEeO3ejkOOnE+c9dK1QvYkkceJUxC+TaUq2wvatvSah+SBzCERJUD4dB
vQFz9Ip27R8Zd8WO8jcOzRdCNs9HcOg9zzrhEHRqgJH/ntbUmrSRsmt7p9wVbhjR
+k4AXQECccyRANkkpzwK+5LSJQdK42p3ggTuVGI9v4u1Zmx4UxWMekPeexkeYw2v
Z42PtKIo9kzeHDbUkvIC00zzw/n9QUCb1zw599bcZrXUzBwIat5z43gA8/8EVG8F
QEmEYc455jeq+NgfDs1OtJpioRtvodq9Yzj+GmZ9OKqXgX+FcUYr+hBmapXaoHFh
I+31pmz2SncWMe2X9rTFGE8qF1lfueEsMDiTuwk2pms6DIRvPwlzmq/9v6wtZhev
TtD+/TFpUUrAZehU5vx3Ui/phfOKrGXzRRvvqsZmqgccxEozjL8JGp4OzsbEe1aW
tx/nwc3ay9ylkbYkYemobPp5w40m6Rf9ZNM6uGRA1mtYzwM7vCDCeXZ27RO6In4u
xccNIbGVNXo+2YnP59BkytBQTHZemjzkDU0IhLm0wYfc+V/zmr0hXswLRQnI/Uf6
BbTBvKNNgjyly5eOyRZSmPdvW2BSohGeYd5hY5LIfvYtX5CYQL+wWvsb6hE6boQY
ffMYO8FglQxR8B1EqsUYx48R9QY2GT0wuDfN+fzPdlMMc+dXlhm5DqItC8xCNUBt
jIYFvSOi9dkIbGfuuQwXvIiACu8eHZzAOSeKmKnYvewHPSsE+ip2qfoTOnphfk5u
m9yqGKIqKVBDBjNNkreQHRba1u0TCGA2YesEKPBpj2puEtw246ozARClqA5FlNbY
0Qu/3/lBrrDa8W03L1XopeJGZC/WBW+BKlU9THtW/zQUAKIkeKE0sSg9V6eob0aN
utlcQxPqV60aYfcnMcP/VXYYOfjW9/c6G4hVX6nKHO4Tw/uE+inL3eIdulPRqlQ5
Ri46VksSbQNGiJhiw5MPU8j7xWdsX1wupVMsbuh5QGmQV7wUjK68oLH2ZCaksf1M
60iJnsgvtAIWz8LbpiwyilM8ouMOiFXKcbEehxPwLU6fPPtOI/0rxROaMy7DY7rh
avYNkgAEG6ofS30XxIxVxYfUgY/ern3Ckr4LZeGRml/pDXm5zh6AIWqRL1tz6QDR
H3tJRvHL0DwcBwXkTF9NLB0G9X0zwLV8YUAO8KrMoJHXBhYUbIhZJ0LpCB4rmz7I
c7VqQHVcyGrA9FzUpNBaB2bw90Enk4Vgds8IslalypZWff9uCaUdMGYqpnEMwQc4
XvkWeEv9h5i7est373EtTDu/6AMQhlBTK4iTK0MNeA8Qx+TFGJH9MvfNHajTF7Q1
PdZU9F2+91/ogMduz9pgsULqO9Ef8dZ+foO3usUorsgFWZz3Xv1XWGiPLtSAu/tm
uAo1+d7p4tzJsydlaa/f5wIM1c5sGuyKk05aMYizlXc3NE2yTBZsBeUfbmUbCWZb
40CV8j06Ql/QQhbzEnbIQNrdZXHdLwpa2buhQuz0LlWoNGjGSTF2WJE/GlCgXzH3
l5Due0XPacFzoAuB4vYxqPD45zNqIyjsdb6riY4HR1ovEbYKUKjSW4kjEJWR/3jl
PxG8WGUf7y+3PikxlGmWGKoxHrdOj9OjKkotK1r5rPjzmLw9x2u4ialCw2lBUdzp
eD6yEJxKbuvJDOGxwFiVRfvHS+6dM5ry1PXzR6IhZd0ML+V+ECRdsSy4Sge4zagV
zViCW2qKtWKjcds8kJQT/Td7Vq/DXFafUxWSeKY++88OhvpEDpdgKShW/hulUmW2
LkWZVIBZcjBZwY8XVHJUB1VJdcEO0+/7bxBpX0SwIgeZqjqIypPhsKevT40R8SGm
l/6eCIZT/Z7cspi4HHk6MAspC53R+RNWH6JaGDR4e2aNSDMbHRVo2/pXNYt/FU/N
XD+suvOiZws12RUHuv4YryE0AZY/B8UikDj9275qGrHlA7JUQMabHq9APA275A84
DJLPg+hLavH9B+i6H3B9933fQrtspqr1SQZFwK3XBOSyY3wr2HOJ+ZQcjc5mWmpc
JVhZF23zK+IqQuZpH0HjLVDuonPIx0es6XePQ1XI4wswj7sl3WgpbK6y9HiXaCog
6uiVBQQp7AGWuldG6+kYg4YckjH73gN2TZh3XUmYFqsikg2NZ6RYHsxnK77WfN5t
oZzPj9fqwM4bhU1inZLxyv0w/hvc9HDhZeSpCC2S8WT7DpnxaZLgYwYPB424n9JK
j0gWw/GOkC7Br5bBauZAvFIdA/vNC+739si1sFGV/R3jM4+76Al3ZXSS9DQ12WLF
0wzMlrNXdAi83PsTOr+lLNLXfqNmoPPsByDJubAPynp5+nOtvR2rTEuyDCGGnE4B
jj4VOy8NroRRblixmAeWhao0CIK1MSjJhm6gVFPWHqxvqQQDEq+KqwsbkZfHMr9S
pV86RBC64kjtqmQx9t56oNt6f464tBHlBNwWfI4uomYNW8NS/K+MEH8Cyb3ED2Ze
Z5cTtTF5q2tT+VKQBvuvEcqp+aDJ8k1cGhdsFjJbnlX5lHJ7AspgzvCpeZSbvQF9
pADKkjvWOAQH4HGxHQCw6uzGCE06ztUP7D8A8GTc8lD+TJDZPln2E6VkkSsZojD1
wgkb0jeqXuaOB7mWXqV9HZZbZ0/9ANuNnjqf8Qbm1tUxT1XGeMUdj7AmwIJdH1UX
m2tWMlFxEKYDaDXDa7oa/B96axnJuQhNHD4tRaD6Tqswr0KYqkgxlJuQfxWhTb2S
Wgv/qcQMymUcnzPTgYUN0iq3e9AAERKWssAhN0anLTi9z12bV6GczoCffNPvBXFc
xHYxbMpIMcjV/tJfpG+Si2j58N34JM811yKVNcd3nmNmj3AN9h7E5wuhuu0GXuSp
G/a7HPuN7kQOMh77B6qzhx3oPPQK9Z93j3ZW6C3m5InGF4x5CLtraxX7NpzMh1c7
LEfjPNPgj6O/v1ld2Dhm1tGAkmWphYS7tjxnE3zJXVUGtwl0mNxMSnxRTCLiAAhl
QgfJCoanpuD04iw2JfLs3GP5wP7MhkWVlTdO6kzFBQcRYDPCUmCAJi9UxvY1XvG/
7lixO9kWoFlu62OfTI/r5JZRctMPSGFsZNCDIB8cNEfuRFFIZJzR1tDmc48wGBQo
711PXXsEBPng/YGBcKVlY/DsjTCfzp7kMO3x9UgLAR2U4JnJrK2/UwhovGutiMg6
sa8WlKpp+6+A7ytl95vFMWDNZZNCFBWh/foqWRNrw5V1VxRc4EJtryacUXPfJtSn
JdCujIerjGhlGO6xcyx4XCzjNj6oGCNi1WVA7RFu8Ncy+x8XIIE+98QGzMvPgwtg
1LTe6V1f0oPQDcr07uuoIkfGHFaqhUtcqyc/K+0fPJ/8Zpp6JOsk7/L1vnjw/PX8
OfCA5y38Zy9AdCRRMd43W2soAopjdD2+xaW3PZdAQx8jAVna3Z1DoHhCp796Pul9
dy7B+whpyPtQH4JP+Br+LreahO1Gyg4Rp2JyyeggKM7vwzTYPzMzJH3QQimeu95v
dUbsWRh90RQFXNLh7/aA97UpaW7WCcD8DzDUyLqXJAIdwYcNw0PRxWDJzAbrfwKh
BtG61WUFN3EKm4YOWFQWEFgIGbqulqTeoaVXkMIavoG5gQGyQAGVCJkm70oUzg5n
R+VtHg3zmUHJRz+ykqzKMQOH9unbPQw7RUPVyAC8SBDrtopnAW4pMhJoU2FREFYR
wW/m67DFO0idyE7guYBX6DrpqnFzfHIaf8Dk3Y7uYQqAMVJHAf10zemhzIjglUg5
SWv+kkbg3mK4IH3mq8RdQwzviSyKFl10aCVC6ki5+DIYgmlSety8X/iaWkfvkN9s
kFb9YvwfpzmFX9isijMTNZmhwn9wyNk0ZOq4DbMXectV2/eURf4UOaSkrTt/5zxn
jKSVPUQb/1mi9QI8civuDzLdf8UDyrKQb+NviF9qtVpeufAEyHG1mLnkiL4Baxfs
p2ipG1YrPyVcEQAdwLpOZ4srAb/8LNttuz8oy2N/c/JxOFs6pXxYsN7U6lduQ0+m
O8t6hWyHNDVnS9PAX4J/SJqtI4TymYJquka+blaRo2di6gqgtXC3sZQEgCX63tTS
QJSqiE+WW9P3i/fk8MKSBnCYsCyosDcbVyVQb/m3+tsmMtutUOZtpKPYEQqpM7IA
oDjBYsepeNKZSpJxzd2tLy4Z6pW+QYdlbC3qTn71EdV1ySBr8pFMTHQoNW3aaloe
mu/XuUOtYGzZMQ2dV+RdQ8Ch6/vc3iLDY1GN5gGZwB82KZnPzJaD8OHQsU0zA7Oz
5IVqMtFpE4X7DqgkLq+URvp52PIl/8RF6JYo+DeKKjWeB1+i4GclAwC3D0U1+o3/
9VvzLBdOtBqJlGwhC67nocWDN+YkMjAC6Qfm8o3j0VCslvt9FZMa3USiCFl6O5XN
agIJYUwAF/6nW+y5jxnQ/AGvsdsPVjNIPk+KI9nYYgylf9Tt25YNubx016DyV8SE
N2ftb4hTw2ZRx4S+nN1ureppCKuZ2grbGY5glVpYh6kaUYYMmVr+vVvdnPXELGOK
mGvXkMVEe2dyVfdjvMr06aQrPIjOTd3HrhWT2r3bIFPX0EOW+9Dngwxgm/08pYvE
/2HDtVgGC9+uip1iwMgrV20vyzrzLFe2OIq9b3msIT3TKsD9zU99YkAVPGHNiq3H
DHunkdV5lw/uLOPsWEjw2eqI3wMKNQwifpAofFRrwn/wh4hzOz3zuwvEJ8UoZEF1
aPV1peu8Fm7rUx3vmCmUDu32WSU1zs7muPMGc7p3T58hrgCa1PTGw/KMYhWMDr8b
EE19ZIBVcIDSmqHhaPA0XP3RrHG+JuguPe1pS9Ul1XO06CyZYd6tj40C9giiKFpH
1tI9Ecv0w6mN+GR8sTqsJOopEuBvSDySlpus1riTFEmcJY7/xiVXhSp53SaEp17j
WVvlFJBwMe/dRv+Sz1QU76gkkJB8LUTBP1atJCjPSuskcYIe4F6mvT0nyJrXtQS5
DINnTqE4TDyuoVTK2/r5FzZlqNqd0HRptSjgPmULGI9IvwLgroGhLKvyiy65rjK0
Xc6hEIWQLpYWSsztA7xuXbsmmVcZ0xdh61QxJN4+0yGOVFv0U+TTPiOPN0QjkBV6
B5BvyruqwAWw3v5/Tasa1JiO0JI/vwYwr9lFbKZaAik2Cm5PzCJj3vrGDaV30WA6
aZ43+kwqM7IsYlUiXnUdPd+drKUj5mL/KGjB9fA1bQFF9Er8GsGlFW/mhArn3kV3
b4siTq3+gK/HQ31LPxW07jneOBNnCPN+NqctR7erwk02E5PM6EFByY7D5Oyhv37U
WEHi8eDQNF9XOBE0NZm0GJ/XWrLZCx6AwXsG0y/3tewSxQ3Y4MdVHCNMvd+KKS7y
1ebYHwYYs81AjfHnALFapZnRjrJQnxMGo1uLKHKsuzwnLN4K6xD/5znc/zuo/5GB
1FKv77N55ct33spB8Tipd8Oz71B2nb4h3XuXy7QHveSFmdlaKe6AYmSvMqPP1Sul
yEYHIzE/o2icnd/P9HfSjn30k0Tv9kQf2g/23r/pqv5bBVAiA2nQ3uUUUElBV0EX
Xz79ZWtH8tu2Nh9JoWprKgwdS1c2kUW/Zk12OZkm+DzMltGRrhmmWersB7eu0gbX
qzl9NmJCKhvk8Y0PxeevD0SVzRxrKTzY84qWj71sMMBUmFhKQML6kVL25kEIs0NU
g4pLKH8sa8qGgYNOMBPxwTZ0AyYAccQk3Sj8vjEN1OsveX60REmJdS2QaSDv0cvm
WrcFKlZ74XSWAfusLw0jnWw+mhJK70H/voes51Qcb8qIXUAE6ElWmyDRzf3jGQUS
2LQME8ziKXTJOpPzc51QQ5vq14XaD6L6WhbdzA0lk2GCwMyTeu6vCGGGBrFrCTcY
WRUOPR0JPZMSjgbquNk/hOI3a3U/+9aXlGIXXLjmJSArcr6yy2Cgw8pr+WGi/dR2
U8yWRxf8bCFf7AnWGP8Uo6q7aGh1l4rRsECwcGasmZzvOkrGm9kWEa3tzjuzAGMf
5UQi6UFp1M/lljaEZJQ15GLI0jifuN3yz4oYCSjOa74GZTJHEdxxK1td1TALJWyR
kx5dMh4h6aoI1VyfMFb3xj9gBkuRls9HLWv8n7PGeH6y1RKu39CK7ZiQ6U0kNtwN
V0SxsjPwzlSKUm899cDdQwqFCCzwJ7sJ3V6L1XWaTsnZHdBHM48HOMBF3IRt4vGa
z+SNQGQ8/KLlPZza3Rs57dogco++OBV8/605X+bz27oI3gdOapSjqut7ZSEvBTDa
m1/xeVEzIUHnNYqdKN1qgEjwuQKTwyk4ynaWI8ERwDUEowXSvNxanwGnIoFgS3s9
+GAO0EVMUu6CPAJJhEa48TROwhWRGWJWcpuUmW9uFU8fFmrmykFP5m611/Z0Ic7G
ZePJVYhXzzYstD8zVyg35VKl/7+QTVuGakTIolqvSbU/G5fXACndk1S1GhEZbql1
tslanT3YvFAWHCbnqNZZl+esSzSFTkE54Vd4A6IbkAtrePB2T/ZGpS5knM9zisUT
YGb0d+ycciScQK0QbH+RQtwhAgNTniSlJLGJySZCUtjKEez4+M1elMmAcTvkk+td
TFplnVWrFq+PJrUDbk+N5SKFwAHsPQHnZNK+/iPzCt2mwREz2shzb6IifaVI0jo3
dA363Qus7mfR4vsUQsZL0QHDbxWUV5h49yO7TbV7Ev+1Yf1SWeDy7DY+ITNFRvJI
tpW7rI8SX3sghK0gXTOhrUW2QbCJU5NJahhFyHqfVl3qu8V0sRE5JcJ9OogQ4sYe
B6go22a2+2tGF0852PuT/Wy1J+8yAlKnUplqqZVv5fyKeaJAljYwfKoJzVZ2VZNy
xLL8EzgtavR2uwFW5gcBUqJ/AgQ2qU6wZMxhOi94k9ZFglTd3GKOCHrRaIjQStJJ
Q4B675Vw1sKQqdhLeNAAHW/UlF08ndS81sagHs5T6LjeEnbv0b6tP0N5+Fyg0KYQ
n1l8cpOU1fPXZpUN8o3TdZHAPUrvv0o0RRjNuLbqgw1VtfHtcp7Expgc/dPYe0cp
tDLuTSDiIJTAm6FtHKiLqoGCAGvXE5y8NIf/wuh5zLdT9dvIegpQYNhkNzvF3XVz
+X94MJZd/8S/AjSbjm3C4+q0Oi+pDdf/5O9Tniqr6j54xdzQ9QkkRreig6TcAK8w
HY05yq6nlm4mf6P4VtcLPyS5YkywuwJJY9TWxPqgRjrq/hCyV3uvq2NiLinAYRsh
2QlxTye0+rsfQk3LDpv/B1MQI+DioU6zcXFvyCN+NNeriVS9QsRb1eX4Jh1phv/i
zpL3Hw7kCB6hRXdekn6bG88rdc/AU0BQFA9s9aClvgnVr4uQgllXSOTBh2biA3qw
16zXQFNX8WQrAlzjy+WNptxQbLDC1c3295A29ltTXGQokZA7hhvycW1+thGzPu6B
ylD6lCHfAiwG1THazcdS9U81sNfaSX2U9yOOAXunonbjtEOFbB29K53ftCfPVQcU
k+vgFb5JtWeJ6+44q4ToklGnMKEYgkbwgJTu6zUriqYMZ01X1iyI7pJDAcA6nQRj
LHgDrj8HTP+kho69F6cUNA1TPyH4o7cTpCLS28pPOq24G5Wc7Fb5p/BdBNvzMdcj
2k4hd959ouD9ZXXTf/57sC2qtOQ8DQdhAMd38QtXFEEQDN3rS83b3HfbDPdfT+dJ
1/gRiGPRhDHKZ/6LBe+Ll+29Wro/qw7+uJD+RLL7TLbBRCovtkc1TcJzE47yWxat
yzec8mVPyEAVB9XKZl5xn7ty5RHcCfutq5zEAOFRXDvUoQ9OJvqTf7vR3Fjbx6U5
RGsKhfmnr35/WtV/7E0EDiqtNGAO7ofeMo/Rr7BZfM1CBTBNsTyFzeF516gimQRj
d/G4Jc3pnVJyhcY6Kq0xgDAst34k+AmKCaFBgyFGor3T6m5ehZh1JkvwVO6GNiCq
fIyzPmmzsUhOGCH4kU4MRTPfNfsYXNa++laptr0nF/iJqWCVov34LEnE0XT0eHoZ
HL0VnPAMVJeRaPxwSdKPUYrbV1A0IP0b2ktQK2xvlL6dWjAJYbCyvhL9AUa2E/Wx
N2xNnkVMddi/eugvbv7qJLO8EfAUf91BRNfnUoAjIS/sfoJcBc4DlEaJtbKqzoAt
eb/v+x/DBtSi8pCbC9JU4SWYMcSX1GGRhFE6aJwedIifjuM541F0lhu+zvshxXau
TQHEcY7md/mw6BVqkimGKnnyar8cE8lUxbJT7XDq1+jFvZQJyY7N0/dHWTg1WyMc
KHZRNXY8qB2OKDA5bOzYgcci9ewLUE/r08fqw22DsVX9u/Y8YatrbKBts1XdiyY4
G6GTL0b2Y831wRPpW7R3tzxdhqjZjsel0ruiKh+HXAFCz2fP+/48M3crYbsyLUHT
SRdw4jS24YL58todJ7rLjFPWqUPFrpjlLxVoXQSQzFRaIqOS1STYEgkDk9eKd6fD
EojAhkG7aaMAkRmL2rxsve4y0YyExiANSViN9tWjdaiDqC1hguMBeS4xgcDRfwAV
a6fuCNbrCTLdnia6acJiA/UqLKZxmVaEw1ycjxSmcXnpLE46OVAzm9nToLzUxlKk
wmIUnPiTOD37/L55qM+kbskaiepUyu61U8bcDOgi3ERXo5EV4rxl1vG8nVrslgeZ
LJhUl+2Jn6lPi6bxHM3xbIGXoW4Xljd1tzyOc6tUy/yBXElOgQ3D4yJlaf84paEG
55oCnIzwUBmFmavKrWBPkh2ElahkX28vyODT9mrtIPJ8RuZDFED3IeNB2rNgFDqh
r8hsgNVAKHzj+wRv5ly+8JKr+NJq9L7YwrdM6XsnuBTBmJVT3lvsfCP6FgGSwMIB
0dFLRwl0tzOHoss4LCX7QmFPdXDYjMdILOhgf5k1rLkwRSKhLlCYdb756ovi1uKs
4RgiA0J9Y2ltWQHrND9UeVfYA8DuC/HbWMuhQDNrmEsg/UQKGngrZ/iE0oVR2Gl8
LGr/e4+ajWFzTSoJvqb+CjOIjnmTpiIBtHv/OfSWxZk5JvVFGNVyF1Fc/z+7GJCs
Sae4P6pcykVGSo4WdJBCuERNCSl2zP5VIaoR68OcrrwPqEWeuioj3ZLhvdZi1LBW
4fksxywcVbrA4CWNhvybgSUmOr1pFLWR3lV8vGizktKcen+b/nBn2sksgeeMCTMK
lTpWDJU2ZLewyPqbLV03XJLr2WfmcvEMJIzC/2DlJRUzn4ntTRESiOsqOg3ccTAT
hXFG8fqKWc+rtwkoY57x7OhGhKJb+DVI73NbStev3S4A0Oa6iLb+dZrfpIoHRmpr
n/KLrM4dpzJ8InAIz/x6scTk0/ns8s1RG/HrTxXMUnLIfUJ7BVRz6eFnDSkubjJd
VMdv0zELRHF/NLXYkamAb+/jH4aorDoPHdGOcx+3vqHuNBIZWNigJri94NjpSKbC
vbjfjJg28yVhoLy9OJ8fhOK2MazMYjplUWjoUbqCbYKnOasBZ4zyY5kzf1RDDdz0
jnd327bocLqH906Dm86bDZHnVy1yNM3yo+rQG3ulL113QBV7dXCU74UXjDppDxBE
iCFFSgJ39LHXdN2a8zN9BxCzF0fcDUl6PeswuIASn+Ftrrbz5ll25jossm4hhBZr
EpQ7Wmo+hp9tDpvPjCB7WCGxO0DC8aGUSOA2Qlo+TA1qEhMFB9C8JJkOb/FzSUEu
ql0BEW+UfLacAQ35Q8IScA75kK81tU4FXyhYonYLVCG2L/0WG35CywNyI4sZl2Sc
K36ZcTXCTT+LXYOtwllkO9YXaJr3pkUnkXiuouSNjzBaJAODY+SwW4YNnmMh1X/C
nUPSaOXtBqMjksDV5IO8Dna6TYBnsUD17oVm5onllv/wKnOQjTCOwrU+ytrHbrvR
ZB6cEScw7DLPWfU9FdcFhL8b0AbCs0VEuNDlB7zUT1gljlbnUXSeGbLUgQcEFcEl
l5NNIWaA8hu+hWsPlhiYRrN08leDYJ2X1kghDsD/KxdnNTV+omJKV1jBAtmfCx1V
FdQNrxGbjwA97U0L/fhkUJLTDDim7IC42roY+01EXacQn2yoKLL4ud67jZFvoOBL
bfYHpBwYnJpspbMQ44qE6ZQ9TtDqa0wcHykllGdNd/ugx81qg5lbmQnLAUgvY68q
6LklHOyZWIWMxkPcsqmiAZWYANq8UmbVVol/35IAPYmv9E5LAbHOohPcEwrDQrd8
qZaNA6M7kX2JFYWKtbAjHCjNXDD6grWXzgNF+PTZw/rJ16KslR/xcFm2vthJcMT2
DZcRM2jgoqzitxMrn9gMSe2NI3UcCTQn+4NY4goC7IVVNb8DmU8WjFYVruRXv4bW
kZVK3c8R417E6IewR/ShMH15CQo5gNpXFTGmmogvTdsXugnyjgGisd5Xqo83+G1E
XgPSGZlJKNA9FeHrgk38LlfDDM6wm4re5S45NCq5XgIMQLJm2zMewizmcwQXrb+f
bWyMgKhHiTlmBxcvTR+OrptNcFlJgXXo2kgVIf/V9nS8AMDkkSHqkFrjOjj+h0UN
AP3NwAZolMO1Vmoegaqd0qAzzlUheNHdwbo7iCFnkpP7nPLqn3AE44mzO+nkJkI5
fC+H7YGjFRHT3PLsS7Su8YTSNN+vnXjf2o4oXD5a0oNO0GRNM7HlPS4llXoLJmz7
ZylvM7Gipft+uSaWJ1EcEK3z9ZFt5bqT2bLOC4b2/u4iM1D/KP4QU2OA7byWgmnQ
vxEvBOjy+uggZE0uU1ksqrGXchAdx2BtgPQ5Ujg2McqMNGsHrXVgX9kYkjtsSNYr
7EPLKyK0e7KaCfFla3GXS4mfkcSDEjY1Eh61PSMjLiIrrd660Tt/Go4sRy7PCyv0
vCIwod8kT4n99L/U8bnF10AvxaURwiNLTzuD4K4HAVAuYukv6wDOKJ1LtznPwY15
o0tzMpzr2hDTeOnlWYSg47jYY6ObPtinWn/LMV99B2afB0rPCQHnm9CIQmVS2XMa
zD0ETYEJOI0VfO7maNUB12mVF0Ob2NarlUVcIWPW9MXFrdYY374I4Q6gJTMkLc+h
JAFeBDoUClf2UMhwpOWFWffJY+VliLHL75jPyr1COCoBiftBs4WyAD065Zx+wjKo
eJBmY5GEiluoWAf10EAvMgBe8TQRGenVvHELLI9BR8f4fjC6HuOv5QnRAEmyVAGS
fL4+ljFSMOzw2cULqJs64xrt7iR2Be4HlLyVBSqxFH4FmSFF8LjbPfJYPv70N02H
Wmx7EG/RXxZCZqWEUzdsTM58llAjUNtqvuLbNE7VBoPIdDnoZn9LqSL2Dbz2Tk58
DHWfbFJ6IBotcNj4bgymW5wYQp+zQSzV0BogaBLOsSV2Nl7CfZRTNGk3L9LDqOx0
RKYxi3yKle9wrcm9keUOUrVr2OX1lLLyB8U0jp1jTIL5pncwauOVcC5qcIQiCvKJ
gp3ENNqrMmRr2TivaX02OpTXFSjdjZ9OykrVn5dBuI2kmUGhbJTst/M4WK6Ust7S
U05ijAUlqMAOsVj4tBuos8fZGfywOtxiLRTJNRbqygm29YpuKIZhPR8doI+pdfTG
Icd476whX4SYmBEdDOK134uetmFyxPy7vmI5y39tgVecHhw1LIUYqLMT3U9JWZCN
LTA+EY4kTHGrXY8m4c/prW77lQbPUvdiATmEtX8fE8hMIU0nxPu9ZLqwwagPQYAE
xPhNS7jqG8mhDz3EtskBTnza2k5A3vmDPLH7kO6tccHgdizs0DxTCUTe3Rw8yjYT
So0nyUXfiy2Xu/Mti8nIL2Lo7MNnhhprbhalbNyQ83OxWLFXH1NJZkeWj14URxxh
yA1w/IZBDGdJcTrqggRD81XdsR46SMDTFoyqHvqg8a4iMCG7ewWHLQ8MBtIDbTxb
3KpglyRVAx1HaCS/QBTjJuhQ260P2kH6RHDiwOinXp601VCJhb/mjlUNmURBis3z
LxXAd8FCnWT+mEDeXB2uGYTcW40LtnM7EODp9hXzhGvc98jCBTIRrbJ3HMgR50Qm
XpJQ4NT+ydR2by0/vUqvGoG8Uag3I696b452LWhV2NIKPj8YYlLNAePSNDCJ2BRz
gzvsS2OXKdWLifh9PWMhUx7HC8nf59PlOOcal0mIifvX2c7VxiHqL0pZPFfLUEnD
pMVIJvEXjibOwkl6v8WIHMLDT0Luo4XwZ5Ts9NhkFQi1cv7/be0QTucG5JQKaRQ9
gSQHIlIKQHWlF2vBnMhtiHD6mQhRI6nGhT/4qGfrAzEGL7jZzSelGvmwzH5l8ClF
tmePW4662tXD+QfoyhlQnr0kR9zKVLY7T2+dhc1lOIhNMshhbBTYfi19oMxY8Leq
LdFbLSNFM4Lv4oiH3wSzXGb0J2ybfYekyLHCbZECHq69Vquc7X+CMZa+OyaokRj6
3b+BqSNw20db0scwZlAtXDgMSSTWW6t439+JOR/IbS5a+1LpIueRcbnvBvleDAnS
Usf5Ubnh7QWj7chIhUwHQuHGom7Qaq4FLLyInWg/EI+EDzI4XNld6CDSl3XoeBsb
0lFxmOEd9voNNLTf8bupiVRlD9Z1D30K2ljxpzWMutLcCypmxdptQ/c2mtw63mU9
BwDcjF3GXlJo/c+24uBG9n+IXfJsK4DGIGoMoFhYzpOXrpCbNItetLa+GIU7IUtx
bQgp6rgzvk/nv3JV+uXVpHN7X7FMpb3Av0dnY+Sh+bn4pgTJEQ0VA+6o6pFobqBe
7RqFsatCuUaAUtFeKgQB63cvioFsnCzSsJ3nLfHywxAmqc6yaANuBe8QEgLvBIoh
zcrr/1n7u0EXNqWw+cKFBnujZlC2k+zh7riJDw+JeNLPkvy7n788BGq+OR4BBVGx
jBY5Gfc536SfLph1Ohp11bYNTzwtbvCQKSJrzrvliJCFHRFN7XvBqCGX5fQbnlTk
eHUJrliy9cqj7jymxtWwbeVVsTohac71WA5PlrnY5d6IOjhBoJAgTrnMNcqee6dP
JTSrG6Dzis2meztMC8f0BpzIhFjzjMonTrQt/weMjaRIpTuI1X9e8T5GATMscOZo
nBrh68JUt9y4KL2wlO76NFYa8WH2+cPG1iBA72MDWYtpmdXrtfnFEC5TvL+X9/xS
8iykQwr9oE3XdKqLDqCyq29pjTMBk+t6ukzFohSMacSVJgMtmsj6J0r3485pf9FV
8ijDZlUpTWdNGscxuPUeB0vXhBYx6tKnYd6r1tOqm5xYHQfJcemurNkYL/kpvyGL
skjqHRCKb9mw0agDdAqYuLyDxdeA7wRhh9BIT9zq3nqFpD0BpibQXlh1c98zNm92
k1OomgaJoqpC0e719z47/jBzyxm6Ltv5B7IkWzhHu96IBxdcLLEhAQPamjUPx0JY
o4Ql6+o3OUOCQE9WEz84o6KwHRPfxFHs7vrz5qyBlS6Rd2KmKCGgCvXXZ4ljVUB9
4+JNB9JlF4frbb/vTcbxrs3T9nWZYsBlNntDn8ag3WiE9J04LW7PsFmyau1tKNry
zYNjHXKPRYtxCVqYyOcsELxz4b49lxoM7n/Pli5VgQh4qs9L9LgU0AS2xQUt4U08
bl/ZFsMcvUB7GJsMnVDisOUIM5OJ3KH7BTjywAJRfUDS+amMTxym67ucZuEdmx7b
coIPJAJdtEjIfTs4yH5QxEZ2ri6NaLij81XcFvE2aCVshmIhiEsYfWISe8ohQoto
G4J/EL1G4AzKS91QFWNVtUBBKQ23sSFRMXdEZbNU6por4jORQKvcNDQ/TuDEdKHR
IXPBpmzBsw1Ms/XfVHuole32Dl4dw6bjisBUmipTA/D64Y0gXI7Qp1EEbLU1aaFV
JEOJQ1rnKPnrccZdWv1470kYXi+urgW4lDCWBh4H2x8gH2qnOFx0VN7W1SuJ6aie
0zRyc97fYqvdWGMBwYMFZqBkqYYM7WCmPB1w2V/0cuUNsJjZrCopsBxpcudSs3Od
qs88Ns+IwKi1wp/p+ms9w6FVHR7p9BuNR13Y1CkFQFj6gb9zyULl+apauUi/3lFQ
aI6s8L87goqZkOT3H83PGb103KiN59hQP0Os7evfLHfZ0h99Ir4blbHeMDZnDE0H
+xhUJ4kI0X5RUeOmsqvUdKg7Y8o3s3rtx9JS/DKNhJXIBP5/Bkr5T//t1+oUqbbR
cRmLT0x/V5PddvNlKePVKmMNWtqBj5W4cnzJbEFXkKVGM3pGZgjmrPxsJQUZDd9L
yB5ENpvt8gyewqSYrEiPzxKVTJUO6YsQ2/MQPADsht/N0MmIy/BoA/7tRwWjC1OH
bt+XHliedB6L+PzlvSEVCiQo9gLVaXzdwiInf0tlkdAh6iUCDVsoqzyFPKqb3jhM
ZL0uxaQYdQG75ABJiWIUs1J0WB7RFFvA5C76pkHxRI9FxrvEO6JwJqbisrd5+RZw
Tz5mqctWH8VGq922QldUum6xSpeEU+Cz3CqrRR6OlbTvzTIuu+bqXeI3/5558YcG
U21KHFxj4HGLODqvDs+89VKymWb8l16PaGiNBkqJkziBPxeYDnTHv1mVEkgahueH
A4eHLwEuOO9qmcaX3VNyKTd11+4ILDYkHar0Ht2m9UmBGCU1P4AKrlnEkld02+/X
XD8Chek4STLnETwNYZP1YaHQaGizfnB47uymlrNBO2K9dqlszNimufst6eY32tTI
4UlPBYyCWLTODeet7Jkt/0wv/FdHQoLZnz+clgOXyv1VYLGR+1AO4kDWunqPHmnv
L8Sr4vUvbGOudhf2viJ1wWNI3ZrZGiTGeOYD8ZBs2qQaEu/odfABIt7Dy640XqrV
CGUec6wb0pq/ASqx7a5lG9OjEteLw1WmSEyPn7jNIEB+pk8F34eCGp0jTuHEqFa/
L7kSfSofcpan1FmBSbFbDW9zdG/PLO6iXDDBNn38LxlDe44ZpwTq+stCMSs2dOGx
ELLTEOxEzPuGSExcaH55YCnm/tpY69oKujTPENOEZmeKq9PZBTkiRcrFrV7pPh3m
j0DXQJFECGP3sAlD62PE9MDCTaAJVTDx6HQld1sVYgQKwFmEfkaIkTtUkS2tVF7n
SAW8kN1xOgj/QRzdOsgatqafON9pxtPJ9rXyfwpvK1o9dCyTXW92/jMTcrnfvbQl
6pGZoPq54db37OV4uIgTnS3lSO0BLSHnNiINkmkvrnPCfQACVTLU9CvjqE//HHZ8
95J3Ni1/bA1xRiKvcO/f0Xhts9l3wC5baELlaQiCLgNQBHbQbVsrpoa9SUx50xdI
on7b5/+qUNHrYJZpKMkkOp/ee81/PS0XvXA/KG+xdg5cixJUqWFeo414Grutqozp
LZ+KScW4rH13dgO1etzXN1ZENHh8mMBZq37eaXRiRYBC3uf+dsIuC5jVokzLj5V3
j7Nr6KzVP90pQDHYiz0IJXk9rv5awFxSfhn0R3XTc/NZxmxKW3lof7dx77SKCkEw
ocSY4Bv8+gZft1kOZNCZSgCtqi5vcC7yMHKihAYmZ6Kz9WMBe1EEBZErAa5FvlOk
rPELSqcv8d72cjgxg8eRwAbMXL868ybCAeahMWesfWl2GD2ocUlD1YkNXq3nsti/
C9b1pZNscqYGYkwJJWUX+m3q9JfN1Q8LrSapKDjFWI3SXbLOHFtLwTcOm4aK8wY5
hc0DB1DXZgbL0HVap++oZFrK2AM7YNOdPGXeV+mJ2S9ev7vTtfHkEzw4QZuQAPfL
N0yx2sdnyan+5MnzXZ1ckY6xJwUOsJiAdvYbMCpaDo5mT9WF03Jar+whvH3OAgwN
mpKA+VHBZugl465B+epB1y5Hc6PVhRkr6NI8e54SABzW5RstYGUu3uukL8QqSAY6
3xHdUy7TxbayPToDzTtzzlgXkQ2sFdxXkRle4qct3Mop2tEq9SN41fMGtm9XWXTL
7VHewIiKUm0/1a4Lcn2XVSCqN1K8YNrqEEd89hCRm1VEmqPGpznznZtC1I6w9evR
HWMQreSf7yTDmp+Ks1/ndU9Ama1wn2RavSY05Drp03IANt4CKAK2ot20ISySs8Hd
ryQUpqLjpG+I/ECihM5ue1znva0gDYkMa5jyhn0lO3e7FgPWw0D3SDcn1A/RCkNX
3MS2pxL78IHC+aW3jUE3MLswkLA26PM+qkP66wDE095VeZoiPmA/m9O/T53GICJ/
GP7Ov1RcVBeKfL9Y5xVW4Iz1gzHQ/KihvJMMc1RiOfj0sLm7NC9GymkOOGt5JOzc
SZNYXm84PqVx94jIG8hZVldgDB/n2Ol+c7lKpw51D27j1xx4FTKdvfRVbAyxzMWX
0rpwVSnG1BIy88VEVQtU3XeSYY1aYg90MnyR7KwUGrbmniq+bMRzIqxq0bGiWgox
6puGgybumP9dBw8v7GHJEVkOp4IxRlsZGH8r+NHsf2XycNo90FAEaxS4nq5NGxNr
r3eoAFcQAOqjVdb7MScF/o8J/4ZCY/q4dLbZ4f/6bht+zat6rmxE1YuZeW375KFx
cKbVW861lXSGV0IZmMY9OTIGjHrpJuWmOplk8meQ/oaioIHIE/SNj6VFQG1Aq0Ej
ZgbbtQAuB4WBRer1QDAPlE+iTbPuw0fBA0BGwh1//6va/B8yav1krHNKELkYJH7v
2AdOcNpDE89D+Ukv7DWzihy7R+47LJXbGSU2t4/0xXcobJNCxjhtV+kIsJyRtBlH
IFnmSMmJVz++QHEtq8pssbTZ5L5kg6dfr7CmStCRrKcTEdlbu9F7iStYBZE++SzS
0ihW9hQu/7KRaGpzgvvMp5hFygt/IbHmBYqiypfv9xgTWfnURWxqX5stAZ/MpH3l
GFmQj5zDQj35Lwh8uIQEnSAQtDE3McmjYYp8HJl3+c8D5Z9DX7NXR4CqwVrB4LQC
CPcB1tndL0UgqdlpRzfA5DvxOd9ci+6pMI9fOlFGHGJovvN14/ZXjZdCiLhx2nUz
/Yq1tuB8cLAoSwQepyen2VBw6mb0Fmfg8mHZ4fQcr74ICswNpkjyqc73Vq9gB56X
4DGKC1SlkQECtcft2tsKLW7chRo4sLNnCWj1fNJm8PqGtP2qQVOiMB4aodyZXvwv
kDVnveas5qf/B3VzFX3BsxKiB9DPRe/5/O0RG8ufGNkrhzpDCOE5RaNCAIEUnHbK
PwKAw2fz8qczh39MO0F4MzA1R7d1FcKSfjGDQT+eth5Na450qtpMsZJ30x0PDCNf
b8T1Qj+kroo00oydzUyOcBa/A/VzB2QCK6oNYjhllQ++izfNGmRRUsr6DB9BB1Os
4Ssa3T053OLG3uJmxEKW2Q3hbysVQM8UD0GBVXNSXGs5yGkvvnzTnt9PT6MhLLJe
fJssz50Ub7hIzlheAlEm64Nl+o/3sAuXNSVSbxS9cInN7l7bZa5+WXLjv2nQBoI6
MtNdsMwZa6M7QB0aZuMoB8p7LK9gC4DZrpigKaHzN4qo9KIQqAtzTKU6J1/7yR3F
CSiH/qt6oa61kbSqNcM8xxjUViZFgB4xTSykB3T7bftqFVAhbwMERZfQ9sbL4HJ4
Z2RUSATZnyd9a1FpF2vfk4du7KvAu4NgyxttD+mK6yaR+ByOfsgMtSM08M+9eBRl
8xXVdau955n1S64L8uK7RrjEIoGND0CqnIVNDOhvZOpmNItd3ZecKpMfN+5J2UDm
N+C9lUcKKb8ulx3zhR+eUUISYsKxVOzBCjz46Tg87PQllHSXKvb64nFrUHAjMxot
W/2pJ1cI9dcd7nDkCexUKIoQRrXXhxZ9O0Mn1QvtOJIHGDnAKAkNTfw0Np2BAzn9
Lse8qfdB9a1pRsPvib+2NJbX36K9/DkB522MkNMUBWDyHmyhrlRKkc3FHeaDLJY/
gul5UXWEbFyA4Mv9ER4i3tUQazqzxlsdj/ifGoRj526eFg/eSZ11mIXrrqbtE5+P
ezg6BjbrSRyhHXjZhRyTfVdVSgqsUGPcMo1Mq18/6+yfETaBY83VmGO7fYnGU+wV
k+iT1G1JyNhk1HaS6z6XHejvaeR2C+qUDDwjXiHJwdPg3w0W7QaJrO4AnbHO/7FN
INrZ1dsw9bDA6HoS1PEr+fUw8hnNTEZAqpkmpZkWhnrnfSis9PEUmRMm6dIZQlfz
F1MUEkBAxL9glT7vbzWbkUQNho24xO3uczYuMM9F5OwpbwbTWtdQZFZ8AkZJ5dH8
YE0YM2e4yWpIFwFviSs22zph+6vNeGsloZGbxSNa2GMRuhD+xq0PnPDNbpUaeJb0
lzRp9TNTZBsowObilXk10TM9FXumrWGSGPO472KvMwj21mdG+pqL1kvySxAGDsR7
`pragma protect end_protected
