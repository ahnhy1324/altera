// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lPd7YHo26yAcUfvuiLgLdwQepyPWVn9SpjvYMbyUiGAd8VFhgKhfAgmN9JS1SIpR
xEXOJfVE4lfdlhCaQiFr0P72dzU7fga1KSZjmPu3WzsDJvz4es2zrKhdLk1fKI5p
UIfLQ0etuo/YOtTqXJuoxlv1CJwG/Abzb7oram4Y6is=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 63680)
yc0SSM9YjKSrEQ5Wtb/OLHr34KMMqZdhaE/SPUH9IVJ82KDHRgaAZi28g1SSVK/l
MvXGDwt7BpO7kOji0iC+iIPVKUwJzTZEcDaKHkxNXjU8jwWC73Ce9JGfcmvvZJEt
DdaGGnqELC/GXg1ykoyt3Wviv0hLQN+SRr9FNZR8P72nMpZulhTVhx9veeorbvCt
z6QGNv0fDas3NKZn999MLMfa+JnSYlEY+2zPQTv5tCReNIPpUk5rFu6Np073zulA
Qn6wL4DkMV/X5MPLSR67phk/FkI4sVAohSl/j/IVsgWfJBcb3z1dU3Jg8qAxcR4N
e3Da/f2QgJGDVvMiR9J8txGt2hPXveVfakfOF7lxSG5R1AkJZ3TTL+Jb2NrzxXmL
S1RMVWRbVyyKIT55UBLFpkL3YkPcJoGqL/UHBkex92uUdSmYcOC8XLiXaopmeFy2
kk8OjNa1TM+sKKT1HjSDIWbUMYUQcni4xS1hIS17V+8yJaKblNoLYGCLnXPmFKgq
AHaEPXWGERWnDvULCfFIyBqb90JsqzcYziyZipc0IhfIpBIlWzFICdh79O/uvUbI
mTpmC5lCaCojyOUHbCSG/LHEh5FWsdkEAJ+P6ZaqGrAaHAOFygYxVJdtlAM/x5tl
+TpxE6fo4NqTvFazLwFBolOkmYBlgaj6ICgX1r318hSV5S5JUTXvSMYIc0EGzwG+
hpviBt8G/HyXVh5FjT1VaOUCXWG2y68yCm2bcCqKqUTunHuJW0/V4eh22+3D4XRx
zJE/bVDEkSNW2tfXkR5l1qK3bf9hllbdiEDn6b13ULV7XVOBQGne7z8S/dJaQfDH
yw1q3a6Q++2xXOcdYrvlnsO/ShnO7J9bXKkNuxNMa10f2QQkMJ3QTk5aMDQT1zJa
Cxexf2kd0eAK8Mio5DDOAQCR70PvWy04bqX7WsBaIb/njJwOdbcRHiMGOPJasswM
QDBPqLn8ElrxL7QsYsgQ9Tl64g38g7Hg7t/6xYQt06y2GrWBSNt+NRdcmH20tDFj
pOWTEYY2BmJVvdw2rtbGn+ba/x00ZAbmmoytY6gG+VwMTgJOdCmui35kmdod98J9
1ybtIHLDuCB9YuxQWYbZ4tTnj5b6FBw8UHvzA4Y/LFzJYEuqHzSe+0qm919aLpk0
A9hoLmQUfZsBdeDaIgGW6hBKjYgaGTX+nG6hDkFHdmLL1WHy3FFX9KC0VwZGgMGi
8J+lmlYf4PMY03MTFDiKsykLczsJzfPirNr3dQaiX0lYsH6B5AL27QWMe8Wm1wMn
fuiZwoNcYtdLhrRtLnBx/tSSbEbIDz4TWrRYV+PbSYytbE3WT1q13XsqQlQHErrH
ZZqx/zajzVwGb29WfJPZsBhNKS//RHqxShxYpz77Lj29roR4XJ0lWSJrDXjWnWm7
Zr+rbWYqkDyBUIGS9/94IYZwUbYspkQQKi5O1jOL+SkeWUKu4Jcpm5llnFPtUape
E9JFdga2Bcf8v8+Bwc0GiAsSiGhJHtxtl0klETIBDQ5sHnoI7wUqgiPNaiNcWqhI
Dw4/2a7zasIojE9fE4QMU3b9cUdlTDIinAdIbYiVWPudVH8Pbk0cmWpt/rOsZ5i9
IdamUxFgF41JmBn4IGKs4jBwFzBQrZWWKjThi4/7kjg+70aPhRENwHWTR7nZMqbt
auP0biYUVY/WLpO3jAzzEc4G2w3TCJExQ4okKLBG1izaHWYIYax9eX68+FVdAh2k
P/EmE4Ve/wAviPIVwqadpv+gfmEU0b2w+JOXe/cc/gI8yGA9UX/63tEjbXO0p7Gg
bHc/XfApHMB9QiUN9wk6uILUDm8NB4Fk17/wwMlQa50f/jFF9BWnhkGmSGiZlO3w
FgPDls/Bs38clf6T1LiaymV0mDDXb9Jg9gFqrYFg5bNvHNUE+as/LHjvNAeNvNde
elZaHzTHqqST2Uy0hO4FCGhyq+1qXP32YdYQ6kCUT1zMYUDT+s/Vo0wJzS8HOZoY
CderCkMG7JRhWwtZk22DYUw6eaQTCJSCf8hRkezuzBQwseAzlcVr9HdO7g/rpKae
48Cflwqv0amiPYxP0/k2j7ccXR9YTjKenSTUMA9saP1WW6dY2G9tqHctGkKpVAs3
rMAxlHyIxPFzTqEyeMcuZOYAqTk0lPnGdm+LjNu++I+evbpEvfKlAE54zExE9QSB
FL7FVwqSqtLqJzUheVvpwEK60nJN/ssQNjRCYzQQQ/x6rJyO9Iw0oLt50fzozfuH
K24HqwV48BMxRaCmYwMi0U3SHNNlxrW53ZhvDxDHt/I1oHF64QNBrLgRfNHPoh4v
gbh0x+djCGbTOfJnDOoxrwFBS8i9I2uBc+Q1yEVW4brObyD9IOYvqDcSjIHyFKRH
1IcP0CCbEdOHvazSQ7sYZ3VA7uzNc80Lh6CJAawVCSUARxD1Q1/q0AVBf4FTTBmJ
3YTtSu5C+1vkC2VAbR2+T+EgebM0Ip+o+zSjn/nl/YUgS7vOc0gfdZEAfqdRaJFj
hYTqZe8IGqGmshyQ5/xOIcQkhJin26FnWyNG7/DfwbWbBggqBrDg7WB/Xxrep7nd
BMocykfAPSvfiy0rXebTC+MN+pRXzr6K7h9rAEqIFPHD3rbdIZVKJTitrQwQ5WJN
N2Tyb8TDuXR1aHiU29hucsvxT9XuILGhv7H7GCanZvz1z+ZALbf+5gLwT8BtJdSZ
lkU/lhfiGYvUcA/5ybfg+JIJJa15ANI6w4mVoPqtD6lXil7QlAJDVbgnz+s/0EyA
GHOj80gIt7J5eftt8RfgDOBHWq+MUah0Ydheh5F43sO+6uqnDfO3+HKkJIlXyAN1
P4szp3+sLyPXpWQPYJjZzAF8uBf4fXaYi6P+fyapUIRPrjcvbngoeI4oAE9X2FyK
3Y9hyto6SQPDZJX4a2twtVfo/5HpruEednNMQ1f965Ys9rAPeC7L6sJ4led1wkeN
4sI9CD8jysiLinhoHEW7/imOf2OYlCdAhEY3pqqnv3qG9pxdrSMzk3aDkSAgxoiR
r3BIBuzNpGBceVge7GdQ9doanmDeNjueZdyty1IMDk3snTHVOnSTpFVHvci/pT5u
j4LoYpdYFz9Mi8gpp/SoL365A4N8oT1K2mrovNXUKF4n2WZIHZQqTXypWx1fhwgt
C7rYXwRDhV+H/UTXWW02SZMgxz6oS0l7+L1YtVXO9bVZHqgzkiOJZLSCNaZyjhCQ
TmL4iozxyCWXC/N/gpeygvt1Mn1uv29HieO1Zz+wnFWs0wUZ20hmpVkQkpnSwNDV
vvi0jWkAG9NMbWdBgQV6VbgCNKNop14J0S4XgmfGe76hhJoktRlxQsSw586FzWiB
/oI7gouCffiG/9Kafe3goCzMNHgx78fADwzxYBSfJPfiB6Ab8XjwxSFz6tAMe2Y0
o11fHYBhkCTOpl6tZ9u2HuLFX3Gp8zD9ueqXLrWZ1912yvOqwyvRJMd5iKANAiPj
BuMCGK5f7OcaEyGo/H9ER66d2+5VjUS1tu1WHfq6jUzpjfLjx+InM1lpCkvOzQoD
qJ9ZW3JpbAeX7+OKCov+XNBsevjVVgq2B1JafOGpoQe4y/+zKm637+cfFmil/zq/
SUfaNh5aQIxlBKT9f6dg+HDS84N2CwMh+jSZYOunG2oQ+uZqbFKMmPc7Ht/L9Ykb
DDFYyB34X4pjtJ4Y/JP8hLuy2/VHvAfvjE7h9fjjB0rZ6d65ki5Kv+CQovUPzFkZ
cueJo9sdLlW6HPR3H2uad5QDpwjNkhVNu2Y3xFPaL0VKEsGe+Xy4DhAOpi3V8nvI
kEb/JnxrjPnEwiWQ6f9APW/lAJgTVsOAa2auW8s8pLxog/tw0wQyzZtVaSXf10Sw
kmmJpp6q6ush8c8vnEnoYuRgH0Vo5tc62h4VjsDWObJ2ZvCAIKuKbaXdgdlxJNM2
XaMVl5D7uuCIN+pLs4hdtYuVf4cxS8nTuiz1+XX07ZWk5JITSlhIK2yN7nVoZFnr
zYieKjwEjahCqnTQrehG22p7q2fp9R16qwfvESp6FWqyfBykGD76XIxFoHYLKuJ1
t3doEsyUzfubu/BXsxvFciwCbUDxUd45YY2vAEtnjGokTNc8xcUt71LlhNuEho25
ot0DTRN5+8Zc148vATOgHwHK0Grj3XYHWBuBblh13K3I/IgvjubMLXio2Zg3RImp
xksUn6NJY+gMfHcIHgSajDw67u8IliqjqN/JiyNyLzqb338/4WMlm1MN2TDX+Y4R
V0h1yXjYQX0IqoL8/0Wd439mYNKcBiXJylv4E1JTJNgC4EQKEawxDRzmbe1rA8xv
5cEoBwfLGRvqQEOgExz0aTa8bRhB0Fai2VE8KQpVmmGE9KWOB4TUF4Ydz7oQX6Z7
eC5Xh4ORCLq4nAJJvIYzHtOPrediAIdmQ2VQjAHU8zD5WpWDb6fa735YoPcMG5jH
JS/JI6586gPDnaHckP6PfNZDeaZO5Dso4LJ8jyRYUPtH7/jlgb1b8wKWrqh/1rmf
LsGMG/Igwkc1vYaU50ndv0ZPza9CFBOHBSw89Ii5w76vqsp/phm46tJ8IfCFU7qn
tZNgUNIpTLfnGcqh0a1jOsUkRPneT4RYV5KElf4G5EPFG2mhV41oCZLCoGLvooyi
V7wnSQLanB3ulybD/rDCK1hocdGTF4YkVKTFvGhMKsdflXu904q2LzxYGt7Lbd0g
iOYUo1NBcqqjVbK5pG01NCfiXFPKG81qeGndegtB42P7sHf3HMfJxduifpCNd7c2
ex28vPSlfGZu+2aOtUSLQ7laGH+jKgmAafoRc3yhanSHdg3HKPxynr1NApSENeZF
mhEgoI+8k/Uior9gwwjX0mGLixJt0uK0LvxRTt0OyejtVM++SOnlXxfQF/Gp7YjW
PS7j5q4SDdpThbpdrJmWAUBih7IejozyTKIu39E5mNRT0f4XFb7Ftttpd8gTJ4Sq
oVyvy+mC7Qk/xSeF26Wtc/JFlLlTzaac4j+4mU8F+2h/BLw2iiv1Ue2puWKndkhI
0AVJJw8pYIZh5yoDj1YPpebD5oRik38IJG/EeIWjlC6U+36Casx0zc+uPWNCM082
QulRaCG7XUmW83VYlWrhDZzQ1wWOuuiRRqTcpid6Om5Yxey8M3AeK94IJYwTK7yH
brSIMbWhAvM7Eo47vTQMPi1ET/Mt34lqPma+RzGjgIDjYCjwLy27LL3bBNeX4gqI
8vI5K9chnFKEduMurufs/0gE0WoEd/lknc57ljYoJv1PYw2L7reZgcSm8W9jSws0
A9MbVwkogjU+MK5jNQO2kwX7VjufR+RrN0t6rvO83VN2cGzhKWobWoWVRbhHi0Uz
btChuHCUT3GzbsCQoHOuMPvSnAmkw1+594vUvWU6PeK6dahtLkpvqthU1Y4ri5Ay
VghgI/GKAZQSUoAcV9K58R6cJy98jeN9OS11evXQEQEF/YBJ3GlxXmVmQiw52URD
HO/mywkP9kif4IfoWieI6DJGT8gaTSY69PPJ8rhBJ+rs/NplfAlaWYQL/H6oNu1f
1CTlsUhEYHcxtd1hvk8aXbfXsbh2LeERs1wvGMCNo9Oc2d4A09iweAt9o3guA/zc
kfGTt2zWHWpzbP9RskEVbETTTgbxW8e4bBORTBQ5S4wqm6E0Yv6hUnGG+Pcb/3mS
JtLLrWToiB1FCx4hUF2womhMnOE14uZPQewnwJS9Rw7+QdabIs+CgcqFvPlLA4k9
PCiYGruoO8nNHH9MgDiuJI1N9NHXV88a6YQJBk36pSk5fILi51tC9GJM/9WfiqC7
XYEPDavFasSjkhc9PYJc8rGweB0uYkZNROxELWjneo0vQDuJH/fWkDCzfu8UNEH6
Up2w7qfNnX6QUZgh2xuUov04jm3PBVV1D4CDwqQ1F3cBrU73q+MLQMDA+wz0Qpuq
zjZL/RhcVXOhCV2BJ481lmMS3ChGmkp9azE9xTgt256ku9m+P0m8ZLA4brwr6qcA
UkBfPQw1bTAo45AHdt4Gk19pRyWhA/LCfKaNg4/Vf+bpOIRpSBphBzr9Ab84i4xE
xMNqrb/+DEfP/XXTTvCLl+yIL7onwv9Zf3Km3aaZG6tazHldHUyHLA6RLeMpRVuV
iah9eKPagrbohvYIKM35BVYJcTzW0j5MFwO0PIwEVj9CG42CCZzpU4WXyUzNwb8H
Vyyy4pOwZhU1kOV+712wEYT3bsraLcUycyRAJysrsxtINbByJNLBEhy2RQlsqGxa
1c3twXQr7FRDd7RLMOFnl0ojy7oPddiicplm28W7bbpiu6sFeZlh3L6Wrl/tzlQa
X5kG9FLxxazak+Ai/GLRB1wDgUUspQth4X2EtkhngwQoAsHlN80y3biB1aMPSKmc
9SKiV1YqOMPMGYOn+KoJeTBp0SuO6nYW3K+qhTNx93PyOkuh9l7vApcP6MhoRe5Z
2kkpP4U0hkSctBvrH+5LkSAL+b62SOEaQFTs97dCqE0OrK4kL5HdWRiX4ofMqovn
nP7FJzQoRgsZZFDhPewJtzuObRY4fR7/AxLeMeS640SIMl0UVJqBADMCAexswvNr
r+uf6/GpAbz8hYFTWmeA/nd+JTn8hv5biKipBnJJVFVYv3PEw559m6haJgGnN1MD
SFtFV8ypw9PEvU1PX81BJSYNzrqDJCFrPlfHuO8h1o0DkdolVRv/5Tw5A5VxMU7P
bN4GGFCRkVRJWNw5qVuc4S2B946s6e8PJwlWXvKymbFSUP5YkG0u5mfjucr38d+W
lfvCI3ArqhWwOwtQIMGzshGERSe0vRQONynSnINuXBzjkMsxZ4YoxA2pYCdcyM5F
0APe+S3C13XZYeZKyF1h0u6LhY1qnegzDwlb+TP8MP3xpUSlHHqbQTj0bFfyiz5R
BHv5iBi1vND0TA+hqH7lUkfymKmkZ/tlficLZPKPA9T8vTWjbM2qFmUeq/kZUUzo
nKNpiLFq+mun9M6HyEDv+xVcDQdMuwIT1qpoTwwpQJknmAnK9XFuQY15T8tbetMP
l643un6QViPIzocqGcccQEbwB27X8VM80KZad9k2TytLll/KoC32tVEZEJXltYG1
cnfbgQuqpRFmvNdObV4lMbV5eNEaZ44wGJZROaxcAbWXKZf2fUUpnkOPxY9PuCrd
6kxiSMwWdv+hcQT9ZqFJrtkSjKIjjFV6yfp6xEQusl14P5LuSQw+SlvBvn4LYp4x
VGn7XGXijwsIMrGh/sTk+7o7xOD523orGpxz/JiR5eAnP6Uxv7EskuMWx6qaXlHd
LB83W0dpiNfT40KlfQpj7BlCH0peYfv6Lsg/sRbAhGFFbj/32NWv/tZ+2fWfnkpd
PK2e2kPaXde2IJAoQqBTM9T/ZHBKjx/hpaHSnjen04uaE/xdmtIFZqjXmUz9uky2
nHR1XPSts4aEGb8D1CeN9aU49C3LZLLT1XeEf6hnC3WsgmUdq5wvdDB6YzDKxLaz
x+Bd9Eu/duEWRZ0fweEyGqZkmAsobUdNmk67HBFfEDl0l5f54uc+U7afELSVRENl
Nb/wLiOMKPFe7elrfQxV47vkEA8lwTgYP77i1kSVM2RnKV0XohCBjhy2P8QCnXKs
i0CX47k05qC0pprP1Tj5nMHbvUVRwXU+SpMb80QWcTXGvHdn+P/Ps3IVvTztVVUu
I1OqADbstuy/qyW2nR3rJImLRNPJ5rpbSTm5ELo/RLSSrBxYGcV0ICTaJwe83BBv
4Oxyw/Mrp7TPm+wdm+dkZwvKGbF3MAtxaQX+6+bUTifLttOV8nhfzuj0bMhAbkJW
LEvz0rOXUF1dEI6bl3ubKzw6bYE1NqMbvrlFjD95SoI9aqZvdjZsWc0yOtNBXC1u
RLLJs6lvoOOrEGlv8/9JozRht0cmT/5VilPz7mpSHsiQTDFt8EqyGfDZxyXPn++l
tXREDYyG6wvqTx3znqqjFaG6qigUOSxw2XFe+IoibHS7C9B4ypDZozK7Ife34UpQ
LxCN8xqGek6l5vj5qo41o5W8A3Ki0/FhYNWcjba1XipUA+SeYO+tqQCllLOj6d2r
0DruoK/TlKY1g7CBt5dI/lTLZecG3dIsp4Lgdb5MX/pzlElzdQRjOHmdkQKTsuTw
QMmI8Rm6qkkk61kj7CpZCDvzYAcctB1KZf83CGzuf9gLe+V48yUDnGRTeSsynkqc
rWrMJ1fgU+mQK7qA42gbXa7dByBCrOPJy98tdEK7uo+W43DJu6/bcbr0oCfakgDW
A2t3N6SGNEJoXZehROQx/8MvNCZIu+92shHIdx3bPrRSbM96fnB4bCcQNdpNlb0b
H0/GHtWzDKh99NCnu904WUGyLbWpLbb210aQnjbNsdO/c+Mj2iBzI2XfQKhqUIK4
YmTZqa+BWPXb/VCfWKLEO3nzdHRwUhZDRXRPZQZ9hNjT8/yqWzg6ornx01wHf8L9
7zjscQTsUdejPzOGRQVe7kCxKBDCz6I6CrlMa27Y5gQq1+wKQOQiT3k8YLKu9OId
8YDqfHloxKbuXEf0Ht14WHs2/CiwA4cfLhl52LXwVc3PbZ5XIKRjmXKsurerJye7
xvyLjb/2ZK9XlKfB6WoWKRDxH01SHBNlKlMexjsVbXQP2bquvGItiG1russj/KLP
s7Qh79pMceO+gRwVUR3ICrwA4rXkDf+v08Tje7mpaFzLPdXf/4u3517ZBujRW7bQ
xlExn+ysVPFICKGHkKrVesH54UTUijICX4vyox3bjzbn6d5VgTaxzINjfINUtIvc
rVu4uFAg6dD7aaD94H0IO2MWJze+7/YfWVC0NKXcmmzVYGvEPrIFCvstusuUmguN
6OskWx+3BLHyZMEbie/W0kYSpqknSQCF932Uc/IGlxKQ3bEeQzvDwyaFaDK96bhu
rZSQdoyMcvvTSW7602du88by/K0LXRq2PHf/+haICN/NwrQf7v8nX2z4b8u/L2W5
t12EKJtibP+RW8ckKbK1RTI0+kErQ66Wa/mVmDVuyX2G8oonTNh1zcGhnCc5t8yO
ACx6A9XnQrKPPwthiqolPtetM91U/tFwV7GYwntb0OXcl+6WfqUQndDaK0Rr5yHH
wOGsPg4BHz3JvGS49BcoYdnU/h0NLnM2LOufhe4SWyU8tO+2gzTBnIYF2iLE0LAS
eyylR6SkgFW31pUCSRJv4cez9KD1uTei4ePR9oLhl+QwYbNXheroC73WSFXSKngb
qkQwg96alClPWUOrhOK3wwpQ5dmwCsETogoQbvI+YND38p0+EkPR8z2zE7OCHWfg
zdUlqU5JCQb3VGK3qH4/N4lxkEY0Yh/hgB1Bbg4b//vNCzwQGenMWjH7ZTEmbwax
JvcbPPFLx74GyXuYF4TsjHbXCoI1p0HScjl1Yy59zXGNXfwXwsApbskq+TTzobst
LPYbxU5PTBUR3z0YnRgt7Ud50zqGcXlcXCm9Gtswn0Ou6ycI1opok8pCQAcSV/nY
drbR3ARFcASmRnuXRDCAMqsDI/QWUZVOZDvOf1p3H/qtPHiQmYA9Sr3htPSHvHp5
dQ50WGqlIqGGS+0EsDg9T+uS2Ao5LellwDskjtPIKSN1JXVnsqopkQas62ZgIUWB
SsN00P0kokBS3hxt+4sjXv18y36OZjegLM52otJKm0Ti1mlVKH7rbkgQi/+1ItJq
NYI6p5hoo8fjoHy9uqBIAgpeOcM+q1xNrSY6BgO+U6D06Du5T7Mag/xll6aY32fL
vZhtodFklZuteDXIdXo2dKGApX2e90bVYRb/vJ09YSxyPQvApGaQvMAF5YpAJ42i
xsiy0zJG4XArEXfwzDbF4eutVPYQ0oZrHLsg+MaIbtB9KDBC28+B+cisPbg57m7/
Cn/mzayWQbwWy4Tni5thq7SgbDKpw1ErzTKgUBad8lt7x6fSRmjKTHtcc65zPMVv
ZnyJDX+KxsdhawGZ6g38OmLQxHWaaYoOLtUDw0DNrBud+kvDFmEMzy1ggaP8vAdw
6Psu03vSwkQvyCyQFp7s1lsGJn//uEK6Tkev4pgD51LXNo5M2gOhdN+vFPHJbLHO
JqP9lfpO5WUUdW+6b4OcaHJEqU1cJjqu0lkWtuSmdGBmyrk+HTrnjElU+rCrI1GJ
LjT57jHwlbacOudYYNwHzYdo9vufwQ4yiQ1/VM4Ypklcq8L9BMDkoOuMF2wgviej
wObuIiLoEYcn9rYego/NGHuNoSbGwb0vNLS5GniE3AAZLVsRuHSLCqqVqrXiqdb1
mH9Q2wzvkVHNFJ9+CURaWTorr42+AUxOWsNca9k3KnOKyGuZ8EWPKnXq5EfD8buK
PKaDOyFe5egB/PK7vSJu5fvuXh3bnjZCPI7DgV0m3bRJ0rT7cOq9ix8Qp79S2tPR
blOm2bFd0o7o6eSwH/hpRlFaT0qDOngJgGgxDKm9kUsVI3G3s5RydUKxFbDT8xYx
3nzRcjsGEkLcmbCCpe5H+WHO+NJyrIualOgc8FPyafNyIcxl36v5t46lxm/JO++w
6cZQZE8vTVp2fIECPCvNlfV9MXIuNGuD3u2nhLxRG6K3TDS5wbHE0iGJ7wSqrX4x
7l2zxzDgnCXPwtgaen7iKsjSCVBJ81dMaKb+zNo/cvWjQHDAsDisRrRT+st/HjCW
qqxr50f/aAs02L8N5mdJM0psr89/9J2kReABJ8CjKWL7dDLSZjBabm9JW0zndVEs
uqiy8kAURB5M0+/17zzV/XP7cLmmpyg9br0cuHBpy0E5bK+AQWHESbWzmZSH+IQI
MjYO/YXiSeioFA4kcgEjo5dMLlA6wBsaL9g6YGye0xZVyIB/XxjtgIvs+pqL5oPG
YgY8Vcg3m2ODAXozqwMkfE3B5Q6kAtG4ie5cDIZSx0G130kIL61a/EYnvBRyDMke
fNSfyJITYfo9GGc7OfJUMEVqSVIdYQyEPgDdSxDqGUpZ3jVzuMEJsL/lkki8NxRc
+QVwifAMiOzFhf9A0KB95wIOAjpMUO/4U1fzjNwkHewPw02C14MJ2JwupRcD2ANv
G/nvOoDZTM9xbuNHyc40QrQE0Ciq/WONDS/t6NnfYNtveZ5RRnNwNkZTxB18fFIO
OfmHUKqkZhNTG/ybLrmvW5Q0+/KeJNgN+SaNKwxQOFdJJ50whvqE20gmXDl4Sbe1
RAZLWRXgkG2pDKiSB2wRFSQjzDpJ6w7NbnbNu2XuCYnRoyRFeEGnDIsHFwVqYbq8
Bu+/ZTzg5ccs+01qKG6hcJmqyadgdhHbEZrGcX/ug9JHbwmgoRNZdSxt/hBQXsTc
qgrTuzeLbtqUV75sV9jpiZRAFF7B+0TMkmJCDxGc/XEYaC4zAbtpiD8mZNmbWmQR
7zEUJDQ/wuiwTqzKt/PBzjCU8xVBlN7TzZQTFYVbJ4Vwf+PFWoOY0y6B6zxd5MKH
ML0UbmWrJfZQt8EANQcYCk939chVuqTvmw6fA7DtFT82mDNiObXKYW20K1fzfQuq
ih1fBl8a+UUC8UmdxhTIIwzeyiN+LiiSZ4ZGanIyMQoxVneBD2DbRLgzEWk2BS4w
Mzqzy24wH9Cm67V8tIbEkuqRShxAmRS1ned5GlOQFm+Ed+prU+jzXzJZC0UGsTXK
8XT7HsPVP+PDaCG2KaA9Dot2vNRu29G+UrcgDbiW99LEUGFn9fI3gh6PEKMSzRo8
jWCQ8oF0uoUf0ZMscTOja51dKR42fMIUAC5y1d+0ExTtXvId6y8SFlnHoukb71g8
CCeBuw2XHzoXeM4JJIYOYsEzSBJVXQXDZm+doKn7y244nvEQ4feMyghabGBeIBQA
wZNRZT4sRnfVhtricxAz+cijzdV1iKLaLa1wDjT6lchhv28U+9xmTGo9qfSY+HuO
dysqrDnty26cU6P3cytpXsaGH4De+y0svyM48Bh6vbp/laETD9Skf2KiH5QfAQLj
A3c/9dBPldEmj0KNB2SWMGjBFzG1KvdJdQql70vyBgf75DQnxVffL7X95289VtNX
MJgL21T6kfB39Uw3RMwcmxM98q8xnc92z3hnjqV8g8l5tHt8anUgs5DVeAnvmthU
xLgm+yyV6spN0XXpYMCYiykWWBb0jjcJz9LlikCsuJIw2MS7BC53k83iIRGTkzG2
eQAD4/MPCvKqH7J4BVvDpKTYchSrXanUJ1XDGASDHnRSXHsH9fiyir+VqORs5USV
2dKCdp71inhP/3/mWYywNY8bokIREBdN2Q3i8CaSntXJS51XwYWIzBOFKxVqaHnc
ZWnXOE3xXhDw4IWIhMuTJSNdsgcOeB8VnQoT+uVMllQTGwrsNmZ5/o9aDoC+d4bZ
U762LoEZd+hsa9GHAflI5QuRgp6bcqrKt1/PiSVRimmYnHDI3DU0o7/P7zACbz6k
hbCCycS54upStFK8BcX2eRP/awLHQurDXkyEC+zL0mimp8n/mvaBekudnxsYsDIn
vnQpNzregUert6nM3lIrtwP+7Pe0YQ9cjIYycsK/Ojem51iMq/J8cK4ONcR4j/5Y
y7/xfA/HH5FM/WZYZhzgXts2LE+FT5rtJIHBZeRpSVgN0WCKw99Jx1WRzJG49/zZ
vVT0FcXBGnhLp7R3p1o6FLL7aixT7TPI9M8i94nzr8ApDAmXRjaGjeP8jHiXCVD5
bhNEuXKcOd8cLdurFFvVdQy1f1HcKs0MlOR3yofCGba01Ty3kXz46Btw0uCe/K4J
9mrPYaOF0q9goNk1ORhaQrhTjoIOCj728TPqyEaL33B1taPvh5xF/iq86kN74MZa
zl7WvzQi6ZGEqhVxk3KvZKimRrlwO+ghfYZ+DPxjjFsBSOnKJebWp6U94V0++EW2
Xx0is/NzeHuLYZnzQBHjX2RAYdFOZTIOAZYqu6TWg4y+AG+9wBlY4ga8SI8qQFis
moZzEwDGaD2IYZjvF100Gc6/wXmm2BjVVQosSYlpA0lmeSkxXp8/iE3uU1539aha
mFFbj5GQ7U5P5LLmX7/QhracBoGyMbT5DOxiWPYm31dJXoGdqAKGTfevWKUoUNuX
M2ufeINUFCP3g8yPktLBSpDIJQ/8nGNI++5zpI1Mlef/dZUo9tqsXEqZzLs5NN+F
PgfIlFOiASEog3FwGx4gCiDUouomV2kwOvF3fEChwIEkTBWPu/UsvDjHvnjSAwqh
+PSj+gich1p6poMvSWCrfn+niHRNbkAskOQyW5/FbbksBdOHg2Ny2dOiJnYx7Q3O
2D9kz4+C55eEl24XiW+imA4Scxqg0Cur8XTlnUmQqxAvDen6s+eR2hPxhA+LBHUQ
Kmr2+1l++yjbUCq6ddw+vJmWH3VjfTYAnmbrMgIVhLkzGbqalRBzOy2zVwAYlWUP
Xy3EOnhdeTCmfkOosoQ+4K+PpdZ3lLrqeI0QC8lgy9lSUPSrbWpB4pbGSfk5/OcZ
sV+bDuOjz/nFUuioZncazrVFc32skoXwzJnOHfEr6tMBGv/Kb492QG1s9Jp+apK/
+/7Qu1DVESszTiaKl3QkPH/rarMe4ijQr8A1Q6gihLARX7zpHg6bmzkP53w2Kic+
Txgjz4sF2ZPJPmsxSvpLSSwI6pCWkJgMrVoI27lGLKDMwplgFVA7QWbYDGpD1z0d
Sho/iZw22iBUxs0kdKHVONzV+g5dx9W2DlS2GIaVG3S1oOhm4Wbm1LVtEF2RtfyG
zUEOCrQSIoTWm7y2A47x8QCxLJGWY2EitSkfNNmBvPYWEFvB43QOyKQqIG9yzdaP
v+m/gOhSJMBappFTEp+SMSofPGvX7L85gU78vkIpaOT+1pl3snT7CLCKLmuxgO/w
XbNVHGk2IZ38FtgWGY8I7ysRSffSt1MHVXdgx1dFLLZ8m/nd+vxuitOGIQoiOGRF
9Ex9XLNzxoGCjHBv+vtDnDk6VX9YcQG1IC7PJ79CMUdKGUbtfsPbhzxD7p5ZPeBc
b19Oq9h1sEpJWRW2VYm4MkI/d8YNvi/F3FFhSOcnRXVsi3I1tiQkx9tMGAp4YIyO
G8RUv8L/aRFR+1pyyDLwHJlEvnHMoOrP5TeXQ3VkOT8I5sL3ZBe75dY4pCAZZnUv
z+LRtVNiOLiE4z66tJhM6yh0DZlLwHyrIl3kDsGgIrM+yCGzHLD92fFB1vv42g8+
aa0+iIRzv2d7E/eIpHH6Gw/1fSAXbOtikjOGOsYzkVvoiyV9VYm2iPiYyODYeVrR
1tB0gZrN3Nzh0Fc6eXnQfqikcVwiCKOhuQokJLDhcVFLz3GuwMTwPzNUKxOcuG9V
DAd39seEKGNMt8vY5sal1A2BQ9f+/FVURha6GDb0/ntJ/MaZ09XouqMpow+sZTdF
gYKtKg5aA6sXLcgYG5dAHiAxsiRiLlqLCBaCkv248sy34B9MSio609FknFkBI6Hn
hu7sDgN/j/ibqoRm340IloLBbYRhDWzZBzPzbwHCABz7W5X9QdMpR2L4DEBsuIP9
nWivnZmDf+RnzOfGuvjlnyx5oG+l/5dgzKxYp52rmhdW5/mq65Y8+F45hYbq0IcI
pkvVxGUXcvrykdfiSmdHRWkKyEym2VCdWVaw7PU1MDlAZ/VpFTybtsr0CSGWisNT
tIlNEzEdZrE+2nBff+BPH8906r2QEcuI/XJacCeRL6F5gmRDeQH0RhQeJo6j9U82
HRDdmXEHSadWtCYLL9k343vyH4Gxdw1VxOqYWdIm/IXZWsqZ/jV54OjJIDmFZnaK
mEUHOg36Xm3okF7eA1R8fHDYExj7cHEbD/8z+YCNSIbaxn8s/oduEFmH+3OmmOcV
8OnoZz0PM3MWxmJNHn0/l6M/+fEg9qWGlCtuHssAdBiGGEuZjXSv4ry8u0EEuDlT
pbbZI5RfXv+lfQm5okGPQst8nmIsLZGkalPF2m4V1cVo/RxfV1m4g68RCNe+O9qV
D6EXBDQFSQPZ0BTDXJf1uHCIiXnjLoHmAYdvSbVUcayEDn5r2pbfnEg61uToL3LP
qomAD8YqBq6oCsBln2k5atvalRm77Gz0w2nn6dPLrDbLqz9e7J6DxrOFU2LQeXLU
DIQX/7qnIqc4iBYhSgaQbN8TVu5HvwEZUJD3ucz0h0LCUvr9TFg0zVsD1GROIssa
UKLIU8poUyaCKNJ4A+4QX0/oxsPzeC7h/G6givMhyPa5k9z93eW4uQFYtSRzwOX7
XeVZtjKwfwjQvK4twAmpVUhhmjtuGi8Su44V3c0ZoqC4vPPmj1+4E0zK4lqFgxY6
5dk7oyYAIE5mjfAZCMsuAh9kJL9GQBOogOMJCw7DEXCuJYdf/TmUH8U4CjOTZ9QK
S1SoQ7MBY8u6bc8KuGEKWqbxZXym9HO2I8ptQtdBGaCjIxH7HHapVKI9KjMqrOGf
mdgeb5tHPKPO8MNdOQhj7ZKOQ8VEkiVvcrZdaKH0qsCd3LyAd8yqHDX91SMcUSd3
aXwnOYLk+0Kwd2Oj5jB4Rt0Oxwfpt/yp+JGkdQjHPKbVrFYb0Hg0A9bN0rpn1j9X
9glPcPPnpH0oa60omE2TbftP0zf6TUwxprN/UJMxiacJlp77kUizjguMYhhUq4zd
sVyV8ClgS3vbaFK3zclyb/kzVUFAPMR2h6PNasg5Cteu8vzkLaGXjKdtU5yA2iYP
Zhyjt2fvmIaYCuGFFNwbv2Sw/ay19KwRWa5IqqzMu2Dlb2/t0x3UUCPiW/iHGwEI
wczkGjoGz1/Gd9rY6obtzawifX5mnCpAHMmexVuxLp1gyDtKjBpfZa18609MKmzd
KU0GWfkWiBChZOr60hSTovbQlg9ljl7WhpwBL2tHfEkp9KvU+mrhA3X6tH0V/X+9
ZxFZ2YA3R66+y9xmWzSF/tFDGMAHAMn8mof8ssPcNUEK3dVkClUHNIKYMJHhroMF
3oy+O6gCgYjwJdHkrExVE4yTukrpAA1RT06Ir8kwBo8c/fwG83Xm7XJERjEVLFG2
Jso+wrOSBbfVtYXT0vgr0wfqDzxnq6V3Yf8D96kFKSPUxHw5sVOAvUJfaD2Y6crr
dB1yZDK5+L77LR2FNAzA6yXSLiXtevMTeVojGEMbB+V3DZeVAWvD19HFvWmQAI23
wgu1QwD5PGn+VhClaCPovm+1uC+ZKl2s9gLYguB98gwx8Az3cK5NOfh43Ameds88
sb9F6OUS7H183JisiFBafmk4iVkvyAI3s7INIdRC+mixYzeKqg+MoTvSxWf7N6/S
RVbXDQ8jIhNeBhXsuUlwALTptE3uF3iUxb135HhWiqSyWbjnjz7rAsbmrGlbOH6j
N/Ff7A3pFKjwYDq8g4DHGySPx3sSfB8qVPFN+QvOORjGO1vNBqJ5xt4+qTlay81H
0GbJtCqrSmVZY4JHqdF1Ah+9juk05ulz/f9FMvNxi1eHOFC0C4uSWv7S098wq+ta
K3xLD2BK86FPGn/kUziey96KJFUCjGqzkSpUoTL1drJ4MmOqNzttZSLqWpQCUjRj
hQldQjAHouKmcpjU9g9zcNs2Q3sHydVqpf47oH9WE2XIVvJ2WP8DDymL6nfv0KWn
N++gSWLGk7ZzCtJbfvWYvc5aqeS36aVaNGaHTG0c5xdtMd24tyjDeRl85nm36ncW
R+OvcYGzNUkDf4HkvYNix23uhcHUUbnvGBRjUodTefNTrPTWa64KLMNmUZ4VEpQ8
6YKbPi0WGq3umV3Fr/+meiT3Mv3zihyixY7F9YVAeZbnq/lhWHGSDKBoE2P022Sb
nF7b7Y+OjwVdHhKmN4eBfXSiSce8irmuoiE85/kj20Xi1GiT352qAtTDZw5YtaAm
n38CrTfW8P4YEYeKTnxHEkCnEw0tk4qBPiYfIxxY9sPK5R9fVu8pJVvqmMMpUtj6
XK8oEzx5exnO7Km2BliIwqd2Ehz+QR/020sEZozLky/ZwgM6Oe7lDgUJ/+icLh2S
Nqj926kn1dCB7lvYiJ4xvtAdGi+MsmE+LuEWWR69WstCIQGbiG6qQEzw+MevuL6v
LBbe6VAYBTcMs4jVgx14FwUE+wWH5jfVdFc5hWc9uHj7JUoAcX5nrWSaWMMG7q55
JUgKMGSph0m17SIRT75F/4h3no9zTeWVBmViCj1os84kSsiUmYT03EUsnXqMLAFf
av0hgjFR29L8zk4T6I0JVwIuENCch/P1RAuRKanCoasqWubys1gnDv7jxmFZ5Og2
JsVftsRzLji9rLrhdRxonGLJ3KmNwR7If1E+/CSKBC0amzqpjio7ybs10YhNyFey
/AT9R/3rFtFIdOB7C1mrAY5vkM2at9lv73ocDjN3DCdMdPdi+slA5wrJh00R8HP9
bBGDE8He9MfZUF0FKlFEyCgFQZptbbOJaSAsh4cOGi9CoMZnW2iWdyTCjFe74yfF
UN1CKQqt7aSe9u3AerZNUz2dE9U6CrbOAK/+IgkGgy4I8VlO4RVS9UxwCUTg7g0W
bnlDuYqNDs7l/Kj9+9kEtKoJ9fQPHIr1RG5lE9H+c6gCDMEv9EPEpHOhfcbohgN0
yJoga/5LmyI3Rt2OKmPNzzbacoYHKDUwi5+pSJyndHaAuzfpa0cncRx26OWa03GF
H276n67cfCOaSVBvz44bgYEuba3+bNVudnp5eKnF3LwF+iWKJ7iwtTS6pV0pnJov
U/RAEZplSlO1+1WgK0gBssxRDAUcDU8yoTaAAXga6nhudcajhLi8JIC1C4zmoeRc
XxRF/WUtOt006lnc0KFSZwQyzpBN57+fCFpvOhhMg0x0WyrQ4STL4Uj0QU2FBh0w
WJdZi5pkqKwahQ+lQPiSxqFc2aCT+V2w/vmzgQkW6Ky8XCxbSNC7tv37oYDC2mQS
3xhR6R52Z6AxB8WuCQlm46F0gj1f6lDF4rCjJLj9fHW53IXV1vmZ/2qFvp4bQxxe
HbBzcJzNvNlV/CJucT3MUoEcCNqxv3VcAfI5LCAhBLUeS7v7xldVtjRDp8wvTjav
UT+cwKY4qfta82cZAloUUGpyzY7rZICEEs5UN2ldcCM+LcFHXMeVPS74DFN6RST/
TdAxFgRA1yx0+S4iBKnmQIMZrXto/pNonNsVQ8mG/XdTpsBdumeW22H9IgJ5VB0u
+Bn13sHriAgIXSuj5jLhGxsfRdAKclZRo1PqlrzIfhpo+eVrxM9v24Bl4he0bl+3
1HCi+yGEfJrl6NN4+9VEPoYldquWYy9pdJyCpO9ZR2NnFIzb7doO7g5W4ztXtGFm
AzDBkRGAilx0ZnA7o3tnOViOsiC4I9C6bW0kJo6NLBak/2HEwMB1aoWQp3u7Emte
7grHrRjNTlDvFBlV+nF4ohUXhcKbiP+Nhc9QM+x0QeKjPKFqkIb3+4R+IT2eorCI
CKll9xKVeEH04c5EHstXW/zAXjQ53dPpR2NOnssZIg1VcpdDN63hET0Ynt/IbKH3
uAGlHmPFmO0Ga1+ZwHgVFWz3yKqbL/AW8sh4MnlkYCj4lMwz0EQRLSVxgDmDbC97
jOi3/yTJor3Nbquykzb81IJ5tIVkvtNXR/RrJvqAKUDdwPt0euJD/gCS/Y5fA/5f
EUgRCaTOxO4alHEzHhP3hPbJ0EaQFm+77mQEIxFGUowrsu+GXIlHpUP2N3wXB0if
ig+LSARitlyNAxehzz/73Db368FsjSazUBM4AcfNkOTlJr8AJoYTAFUvZZ+9LH4A
Ln45RkJoUUEZt2qSo4ilVGs8cuQEKo11C1ejm7fXSIeWfk3iy5DQfBAZAV/ObLvW
2SIYEX6NZrGcRGxT9HKQSgJY+OIJ594OLpDdwZPdaduxOE/5CqUfmdnEX9OxSqEa
FeNUwvSZPV5At3SlIuxJrfS+jy1lm2wGXEHfvLMvvcrDb+2rdqtD2fSRMI1QuEuD
ti1ZfdumKA/Uemzr5sROjVJvEsjsaiCT3UxxYvPAYlWa2yzEOOFK4EUM4UpkIAJ3
+0ceWspe+ztYA6eeCHp0VkmgTyDK1kcGQ8WMTI74/YFOfxVFhSAmEQCcyIhof6ch
mHDZx/GHSHPsSQKszJRZz5UBZXPpE/rCfn2UVGQUwfP9cdYUdI2EvY0oiHZrWOT4
XzQl5NQuVKcbjjOmYB9op6u1TtEpAo+v6wWDoi/y2mn7cJ7zFkS+43ECgKhqp9mR
D301i5gKX9JoUw/pbu294K25s5JA8vBlRDe+okJWGJg42QDChEQb1zzwqahltYKu
oh550AM02y61VhOeJ+96hmRJgF/Yat0JFnfQi4eQfj79+oWsbFIO23VsAW9q3UtB
KbIDUW6OWtdLZHniHqTXo7jZkxWQZpLztzoMmpz9o4tdsY/c90Pl72BMFJvxR4dl
LP9yxAMYeFxqXI3qTgOcVSlsPVC5xOnaxNTmTq55RayCRR2mEjGMyINw4O/qrsxG
7kPgcLIAzt5GGTdm7W8sT5sdovkSYIhTjuagsdbp3DOLRqzMO8l7LqMHw8+oWi0E
44N6gA9jf3R2miAi/aop9X8cpSBeahFRLBwdowbcqs+9Gqbc3BXt8UlZqZ6weTwx
4NlYiT/t7NMohQVr9YyvUL7meTgu4LOzB7h5wFjLhwYjqlRU9tHs5cdEvg6uPMkV
ibfkte6uDWvwyU0e744fi+PRG0uhbaHQFndEZIAoB86RLJclJ7Q0mRTwgSX17ZZl
Pmv9EALIuhsARUS0j7jz/LvEJ9lTD9B1XqSQW0oNiTmvmSRbTVLiVGiPjku2DBzq
unB7sNutQsI1gxs/CfQr+RhSWfI/jP8uPeYrk/xxiH4YuJvoodRwKEvaYuv6lqgi
RYA1rMLDX9OGf9gqXeqgtPb9PVP1/CnOjHAlH8CSqt0MGUQz46yZI4gITSpmHPxh
RJpXUgWu1BbAnWXPJd1/y9Qam2b8aozKe8gCGWMCV9LTpPpgW4RoRi7JRDlfib/x
t/vTkcSztAT0JQK3Vw60ig3KKzGSzy3e4W6DPXN6N36L9vNgS9NMbrhX6ZTbxeEw
CLF1B9vtedGBRsEo0F1s3YznHvc4h4ShMf1i2xeGMy8WI+vArB1GPccCj44WdKuy
V7V0bpPWAAGzgb3qD/oe6+k/NPIFKXaooYJRsUKfB/3uAhjkD77+upLI1p2CVBmj
ZCBVCNoOvJ/trMQ36lw/P0d5WiCLalupZiyQV2NtyCLBP3VkJC6o23sNuwEjkJ33
AIcWrXXjnghFo7hy4VY/uGykJ/2UH2io+xzAx3vKpLqKyVxxIICpHBZgrU7RoUn5
tqSz+QeshEfWVa+cCVSF1fEpzWs9vX9Vr2UjFhUjcEMh0caZy521MHSTvzThND/A
zdDTjU/h8v5FVjJXz4x5chbxR9OesMABIVYzmd+gbCd7UfHitD/ptex8H/IqXfUa
T+qvd5b34Mf8G86kFv6Y/gPTAK2qVgWFnI6P/4jRI64RYCl/Of6Q1+tXLriqJhSo
DyRNI0nZuPi5sHpunK0+Pbp4zhDRWZgW8jQtkoNW/yK+S8Ms6XeDRigenUsZwVaG
k2xog6jwWJoifp559JDpCS9Sgiwy69f0LiyEmrU6X5vSeJZGOJ6b16C0enJmGFPI
Mm+REJ37koTE+8DreCN8x0pf5iYIPMAiJ+DhcVWnCxuAf/kHBIhgUimsvOzEu3XN
QdHMaczrhxDzSYLqJd3AM/Su0Aa88UG5JNhBdkOTTbPJI1jgKLlh6MPOkSFtT9W+
RcKDUdrZ8Doe94DSsvw99NEl8nR1bvp+wYdboyBZOODF9NBOVzcik+8uRrcCH0bg
bE38/9hbwSXjI+ZGLpV+NsAmwCqLMLpMpo32JdsZcnN/GPggtKYIWa6Zj0l02Afz
NUlDMWA5y3y2zpSUq7iiFlbrQPBGs2/SLJcq8UO9R+wwbV41N3W7u15cHrOvfWPP
D1bz6IUV7Y0Wvi/XsIz1+ppnDppEgIFde8DSU/d6qpVS7Yo4SCadxbbZG3+wjbW9
f1V+je4aNJJQ8JuY9o0jNbxvqASfoJALqsz0Tzz1LezC+nYksgMQeGnoZQrq2QuZ
ksjPvJttQf7zDOOe80OCmqrpGJTTdIHaGqfXeCQ0nwVDsAkXrA6ARzi8mnqLhKed
t2iCcMNoJ/Qmytm3YpmUkjC3MjAnWlsyRPxpVmR+wTXbB5e1/lfNBmBgMGnlg4Jl
alLa5D/QUsfxu4qrlNq5n+HVGMEw8CQAL8oSpyBGgigElFfJVxX6iGwpy3+EUaAQ
EwM2Elka/lTNU/NYAYTX52DqP3atAGqbeWGrwU2cq2ndjd5hKXQwGqj0AcltjSFN
tssdUDHdKB/1xPndGwTSQ4z97dKWa2BETAoQsmjrcp8/fiIqB7QySdMFSg4vfDgT
8Sz4GK2thuwwnUpkGN4zxOOm8JaUNTJifm6Tom8BLb6iYQAtQtKt7xcZHmAFWERL
PIVjRNM1pwiFhywmEQk10LOBdhnx8RwZy7jI0x9HrnAhGQ5FCNYc9tABUiVEBgXG
+1XoalLNll6+ORzc6x+JbnoSsTU/o8diCj9AyGWg1q0UwG/rz8dKG70bAd1qtIUV
RZ4ZV5C0BD9Px8cG7/SNn2LxrnQWBz/ljma7LaGtgaFdDJwN3L69aYs43qkNBKHx
IaY4v7cOUT5m4HDQO8fJQUJiXbezZE6UbEVRN2x7WPzGgNm3jB9K8maVexXbGkUN
Gmj+SHK2HBdVC9hJBMd10dipXnFNj2f8EbyNBjHQW8q4p0Szvxg8GGrW5Z6C+7jW
Ca+qVYhWYtJrelKed5epfXGYEGQ1AtDOwA9/tS6m0Ygl9a7RYfr+e79DPcY0By9j
zQvMAYIbPCgs+va+cHErtbS15t7DTke2X8KFkc97zjDY/c/AKJthW+zCDjbBzxBd
bsi9skcWy0T3T/kRkj0jABtCiNd0ekxN6Iet2NK5u9UNBoLYoH7QKzhMV5UJAcm+
Ie0uG7X7pdJRZFugJn17tQqEyocr3XfDvpk4fTzjgiaLaVLQVkVSvVxNQROl558D
5DGG4Pn1dLicdu1U7BRRvaUpbqH3Gs+Ijszoebp5UtqxKl2wkHX3ed3uPxEnhdNL
BU+iQx6imG8fVHVBSk837O22Fj2jHUN21llKGoGxl0mb73X71ssoTxDydR8cROKk
p1chS54hQ83volUQVQV9NBeoQPRYD5C8Z05Nd9uomIZ2r8uP5rGv7OZLgutp1rZZ
AOVC8p/owNGNJLnVVIVj6olILITT7WWqknvHF5uHpycXxAd852OwHqVat7n1A9lH
9RAqG4zqJ28z/+wbH6kZ3lX7F5HqHi4z21bDYUWzt3q56DXZoDZUbm4gB47t6Fqy
9lGverGqP8AmDGJXXdZgTYLeusq2FjszDuuIozhBSYXMkWsYEtQ06jTZJIWM1O5/
jEUfNn6N7aOkK0BL/aaIit1MsCovVekmp7x6jk86vFvAocQC9b6d+jBKHjEQHMeG
sLLXg3sXHQf6/1pAvAdIzYM5RWsHwDnB6sEzNDDxLz8Uto9FhkR+cQvCMLcjcIQp
OkZsGK5X2SBWbglA4NznZCXMhQIZkLvm2gJn6b5ONSSkTZThlDIc6hnXMvbNshsL
PDPKqv7mG4CSIzLWduo0MJUHm8aHw9nMuLgh2VvI0QdXMNpANCUCJ90wEfqrbcAh
HLUChuwr92gaKM0j1tTmaAOOmREoiX6H1r5kw4EyyN7QLjGKq77Zz+Zt9SFNeZGz
MJnjzW8pcgWZbGrTYtAGfB4fB5LlZaOXxXdbszMdiYATB9QaBwDQM+MGjeLWqB/A
zEoovrefIzijP2CwJ8QRLE95nL0a5elquv8cCbhW4pZaLSbF8JVwOZFZbSlhRSht
6AyADULRVWLs1uCZwdua7ER99OmyPlIhg5xP4/p88thjvqxCjc2qg1+k3IdYkXxQ
Sa8kzSzSiU7yWqc4BFwZegqGtEV37EF96InBVYHTTLn751Y+QFJzLfZr79iV5x32
TJgJK3yJkmDHiN/xfg8R20Swkw/NWin78NW3iDY8G0uU7mJqfL/YZgcik3OaJeir
XQzA8yJeDYTFDx4oYLg8/xVUackBFR1RlYqRhcXjGIs6f9bAmx+j7QSwgM40mB3H
f13cH7GuezRHwJM69LzA1JmKXGkWbilZYkcno/GDjPFn/cYbjbN7CMHmE5kOOjQv
yJMqQu6soJ0q8c+3Qpr3s1QAejJwnt6vso5BvwIchwvTtKQUjuSimt7wKbdn5NE6
dBzpbZiK2J+t+GpN4U4yXEKfzxaac2chf745hgSMhH0O37mgNcHc38srg5ekC1pY
K5HRUts3/79DxsZ0qb0u8FiJe176GxmWky6jyjWFqKHcXpqoLin9HZT+dFsswSa5
YARWyx89p1yV310VYBO9jVsHjQ6P1fisMHNoIxb9z/1GvatnF6UFXSLMltso2XOq
MUKwwMOqIbHjwkvS9f9eWg1xRYBNh4dp0bzlc1BjUBsGoef/hKhZK6Uha8HDsgnx
TzEjQ9g3Fbr2ZBPQmqK1KbaQSVMLYwMTelRNSRJv3Khh3VT5nYErbu/UQxKBcT4f
ZfcfzG5MLdvWKOjzvWv5uqBN7iTdYGb/Bnnsefv34zy6+7tP4357TRfWZ4Jy7Zs+
UMLeKEnrHarCBBVbOBFxxFs2MHagMeU0aYE3racezWjJn9MWlXdUwmKYZW6HtAYZ
tmFsvofSk4woVkTuLUDNrljuPYYMXv1Ce99QGfNmmrvV4jgJA7JxtKRfX8eLlwnB
/YLK5zcfnpIrlKwe8SxkfooIH/XkeJMydko4/7Y7UOo5hktkrldMSk65qnnM+BA9
UdALaaDvLiwCHjKtMPCHCyGo/cSqEGhTr+n+mIsh++Lg1qLOCbsNC/iMAbQmsKlb
aW7LDEeQrqeHtc70kLgnNVEA5BXd7p0t/QhlK9hSihJyChK9NcTslLrt+B4DGt8/
LuRfUmYHKGMnDIwu5gCP5ea3Wj3EjWFnsGQ/SnDtoGrt5xXUaVQP65GQSEYCOhUl
yjw8EKUnco41vUe845EY67/gKfjFc4Gw1Z7L918yFXUa8BWqN/qzcEq2rbyg7nFP
akKXCe1IYYPtpm8HchFraZ9BA736q+RQQFaypzJdYiS3iv9vx4wwI8hTPCktr+4j
JVc/Mb5BrgF6q/OwzXUVVXi3x6doNHbp7JhcAMwG6vasq4QXqs5WSPsN0Q4nDD/g
xdBUgNWICAhUM0nKsCL7xEl1EAZYO5ZSHV90zFecuPdrQ2CoxjekQJEPFUXVxb21
0Lpl3qDvL7d/nAzqIHKZqHGdKysD8AOoJVca2YTJYc420J0JPL5dcu4M2r1Uk+9l
LE8ibkaz3CkMQtU1MVmiwx+iPt56VR+vyIjcfpYhddq0GRQ3/xtzuQ9nkuWp77GZ
9wztjNcpeaAHMvYKX5WQBD3lQGeA8L8qWGMfKrRYkAx+KMdpQS9Cz4oMcv4GHi+v
ynPftstMk1BjIQ+aOgpJypCP9YpFTcnmA7IH9wYHyp2sPHcfE4ULyxq3RP8V6TbS
jHfbJbQ8WIMmRQQXE2w9OfFBdeFXzZ1/u2YBYSX0YcwWUT/lLIk/fEwTuN0Xon3l
iNg3DvMwRcZgpTPDIOLL39J/FhNT4rXlq7RNJ0UhmafSGsoRAXdkJmObWS6Np2kt
q4ih7MVrLyk/Fz8nfXzJmB0tnEeVoonMUZjbmEWbMdMWx46e6Etq+pByvdimxl1D
PKQjj+jPeF+f0LlVnn2ytG+MlFbubKHXY8h+/hheTTPfLJQKw7m1bJQUzUlwcJKX
UR0n3KIZyyzvyl6Ewx5GGmmXk9r2QcBarSI8xZYQHrw/zRhzvUn4Z0WeJQnYRXRl
utTS+s0NOqXXbPG6j9SCAh67IBcru3ac7O1lAJ41Ep5mmjPUXJJg9H9UK5JrpYTf
5W2XrlQG0w/U1AHqxJn81NwOFF9LZR2Sc2Vjcv9jYrOD63JThaS9nejefMqhPQzM
a3mExmbE17sLJAWl8DIUpqHv4y9se5FMFqsdusbuCfJgrYeh8pluWGNgQ/65Jn8y
OZjjQgVQVGcCowBddsaBSdGyNwKuyrmg57dLVssj/wRM97AJE5hxx+YDYBYM+u2U
j2F528zFxequprCJZnyBV47FEyF3qyQGh7X4vF5rGRnyNTiug8WgTOZfdCSEnagw
5rIXQ07q1ddn8I95NU4fxTqqVzQo3rnf7pebBXvLKgwGpt5qYPSFC5Jo4KZiCzuK
Mv4EhIiUPOvWj9fjxefbZmkzncpqrOjtxQclpNyZgoXirDbS5hNbWoErMw8VLF/d
Pa0HWUy8+CEAF+MzsXlu/7JbTYBFJkTQlv3++nKhOJ3ZpnDZBUcyGx/zN0VL5SmG
XE2pgAo5vbPMddj7EZWz7VfyFwFxtLengw3dFnNiysE07FehRLRfraTvJgRvs4Jc
PtlpWvR+WjDoQ5NxwEkibZTxgq+uEFAZuXeER1w3q4wyE+v+hop0brOBBGZh2/sC
7xgySAqatjshVmY1GuFvVmAlzBu8xtVtL+SnkXhszifqGF6qq0/H70rSKDvDoFXy
trjQugIlDlAcPb7XIibhURAllz9Tr+eyffGSX6Ksd9qjp2+CwfWT6lSqCyFNcj/4
iqj13u5e8keqASlwemIiZVqY3fY0eVo1dAZzpfyPaImT44f6/tzrjz/TUqj9x+mZ
CdQXX0YbhWSh9tX6uKAOdWbfm4NMfXM9J5fvx2CqV56qj6mfdA1ujYAAfn37wCr0
1GFkPC8QbqW74FJpCm5k7pLmje6HceO3IYhrela5u49goyVNeQqP77NDBZDZXqea
1OYsjo8V/GXysdSDXu6sfYdU5JtwQfVSJeglYkAkATX+Bnw2XnpTlu9CCHsJZi4P
QU3NftMGo48PBoC6gFrnTn2GpZM1QVIsPBxPIpd7FiKmklyq+npNfRb/1DcqPLYx
hsjdXWu4mzkTkj4Vvg0lxam5hVl3wrrBtNDFsLsm7kKYMxnPsSyujtNfC2oNiZ4U
uU0Fojnsbre3JcOaEOepgcylNz6cEeW44/JBPVatL9BGSJIjFd12cNaCWwUZk/ll
V9q3Y4lPZPSym+UXPsKjCK0HeN73MPRpUvRNReaAw+ow5UctUebqINxCBQEm3cPI
aVu2rAkntwQLPDsaxIM6ZhynspnrKoHc7xgNcyx3KQAVWMGc73BtkLeWJwOht4/N
BbUmvqRIaU6HpD0EyL3WwAYagmyJVuBy3X4OoabMZQ3iWpjzxcixuPXeC/keF0x2
y/SqgSF71RLVvwJUHASGu64AIUKkI1HTNDDDa2PG3lwOAoY8WpS7zOln9whnfXMr
bVKPlbU9O1VRclyHGu6L392ZdDXBUz4cZu98XnHvDqGk8/SqngI00DaOkrW+clXu
Wlu10ky97pMVXA4c77lfugM99SKT3cCrTlyibpBU+k2Vely9fouTFBUQM7haICT2
E1PBU1xAdFsto1rQofrK84eD7iG9y412u5T7+U6uERG31/lRuIz++aoktaT/kMzn
+kvr7fafTw5fh6kabfvSRpAyTPFW+EHXzSxv0zAmKLlleGZZg2DYuJyN2ja6ADHw
lCeQBIrQvwBhV7MuAqRUARCxI91JIOz+IY1OgWPQ5iQF/xrKs6edqZ3UPjsS10jM
29FgPBtw0UJkef/yli/oYGH+w9z0KMLeCXz9vu40+7e+iJlevvNTLpX1JsiZrrDP
GCT2Zrqp0mugrU9iB57j8OKtwQqShsBs9cR8n4fAOQnmuuOdw14R3pBxpdIq/6oF
03mpd+IrEM2/+QVGK74cCVwtgblGaKMY8klnu4gy/4KRMoED9Zji3TTnAz+q3fo6
MBrXHWUrw11kXmqob2w4V8/0iLyKRQqpCWz5gFsBT3REqmQAwyEmZkUukVyO49X/
JFdZBrWMDm5GNgoArRAtC007VhDgKUg3plkCIVJwXGv2i8cmneNTPBS+B7pcWmAx
b9q7ydXj2I2r1U9IubmmieacuseuE0Ei9AvvX83oA2SHuElb1Crb4lLj1nHOY64B
N0HP9AXddl4pKUsB0YbcgKxXAIbuToeAYWzDB87XBAGnkzu+triNuBeuhUfAlCKm
2UaPjgKZS9mxoTL2i5UMGENSm4qL5pT/dJqEF5pepHpMQA3pc5icumie9VebCXKM
eFrFWYI5Csyz7W17WV++Gii9ny4x+KRwjqIaAOmuCGUYZZRuB6PUaqb+hnY8sibw
PcBdCAbQikR4cfVc4vJ+nm9Flx9t4YJo9O+CaJvsz0SdtxmYAMG4Je+Hoq6+fq89
0HUmdgxcGNGulI7AyG9hv7xoMVQhn3aQAqyR0k22dtfzyVsn/WAPbKzlhCKRxagI
JPTOCxkQLTlvDR9d//JEh3gEsqgT2q0jp79jK+Mym/e3PiWEtWiatKs7scV8DFYu
QXFJieeN7ObxG85228AXSzYwzdeJecmD2yjIblqxYqIdR/IAZifkRv0XqzmYnQAk
6l8pH1YxzTu+lADOMY6YbRIPWA7pWM0NAxE9wcyApOddlEkqfB+j8LSeEXHknQzO
7hRa+anvSrJ0tDMRv1X8w7behSsOZpXC6Hs39uR+Gw813XApMepNMPjY9VoSD2tI
rGE2366nceKXpkTVacikv9OaKCUljZg/4WyYTfCC6y7kZe9B0V7NizUMr7YyXEd2
VCQvtdTE0HTTq8CHhDappe+/ot1bfSc27hGKTPvsXyPLk67GRsRdMhElDgNinuA3
rnfndj90udrenKZA0ILPBhrQQIHin/5trGN+d3T9LSWjGYZSA5jenCfz08UrN+XR
Mo5xiWb6/1LYbJsuwsqchzioB7Ln2rn1Occ8qScFNGLfBmOvxPAvwVopevEViVmz
VG5OQcnpKo/y713YY8rNYU+lwYpnaBsSTcxWkLJLOd5PqhtWcPF/0EQ5xdmzmzzO
mOJqISag209Xz6uWxXpNXZ2ISvw8+OIifUcLt7mNavcPTfuBmpT0DMD0ke3Mq0s1
pgzddyoDMWV6Jz66Uo15ZOByhMXS1vklFkbEKpujdK7gFzwTTNDvX9ZNfjRWyaK9
+pfFqWr/VQue3S9Nt0eTGSgV49YEramaFU8tmsiJMaDCYauFnAd49qORiyxHdc5b
+clY0H2VKtgSRuOCy6p/YWrU9aWTkexGT3ntXoSQ+TVWfq2jf0YxzZ1pMA/OlIOo
aDvvoFysRiBU6Z5ipqlgdc/Aw+pq9N0Al0Baz4N1e3bNSqTA94U2YT3RwXDP+yKJ
e/CcOzm/b3Q5+kqQpClGFQq+ec7BCKNN1d8yKI6hOm2fcRNKtH/HEDpkS7NY64pM
hIXMYxECmCgQdOFjK1mLZjjGmJsi5LHomJ50wf1ul/PZFCvwpmucM0qUNhv7AYys
6PXWif6R99maMsXWhS/I8hzXRFRxazqYdQNIJqMh/lOVRehHCOi+Xr08L8WxXd+7
l0wbLAf1wQLi3nMvGKoqPALwLYidRPxAVsmzaKUr4WZjATBPXQBDXag/tNMQWAFD
u43upmOXmr6IxYPOxb92GfoWroR34PW7WsEHRf8duCsYBdo+qeoPKIn6ubADt3Eg
D8CdOQLOztgQ9Xi+orXl4l9cw/gcl5CQj+6pxSLwX9yCQRzsiENNypdlnTqyiT4I
KJHrCJxmi64Dz8YuNnOIfU9WiKSQNH+IB+9yWFKK23rQKespyvP95zOn3Yilf+gg
G+ET+7DjrsSc16nq62M59rT5QgOIK4E14KGVRVqglCPZ14ilxoIBwfACGoFTIZKk
+2sZB2BesKpgW/N/T44Ra21qPwbD3Axnsmepb2azULoIKCvmg2lHyMIlIwjwopFt
1b9nhY1LtFpD83zrlnTmW1dUDIIY8peJRiRe/l1NIGthmvyFk8C5NUq3E5LCPT8s
JAfOk0Gk6L9mgv4XtCrU/mvMW4qcB3qt/7GCTBDwkTZyM0P/E1G7u4wn28eaIkIt
Ku0sMnsOs11oB4+XJiTNewQ8uJrFgOy6JoIFECITTum/vH4BctWF0QYO95sigV2P
IKMTFxW33GLf+TiwyQIABaYhwhf4EmwrxeAyJ/ROPfGMdhKtVJ3h1LD/oEk+PaYJ
h1tFvx3IF0UHAlGjg4qaGPCRdbO+h3akdqHre7rUKkNQPKzpenM8Oyk3XZAHyUHu
nSgDUHeLuXx6kzWzTnM/bZZoVz2/zrFi0h2oaHEqgMG+W4NxlT3hyMAD03u6BCKY
3TAYbj8d+NAmsU4b3CqN0XR8uhUz740sVY3NK1sPa0OWVSbddOGBd/hB4CyuQegD
JcvZ+FTI+i05+wNY7gPZhIroCDg9eT5oGyfO5Z682gX4QwLzbWOG5W1W5cphtEsB
VJZK/SBrl2tGkIe9lnXqDQGUl5nvO+xr103SiwjLhHBsuKhIN5T1lz6oTXp5OwKw
ndTYuDtUwmg77IdKITSmZXMZAQEdIOskss+E/3FE8AHtaz125D/yuoozrG0VkEy/
IMViw1dsT4RwFTOCESnghsJWxpSb8ocevG5tApXaiFF/vZtjFfvC9B41SK9ezmxQ
ySXnxAJw59N7WSgrKCtKr8Xcw5GJX5qW7pXvSqg+40KD1szGDyYLk9VUCfdJiK/c
tcDAjdaqr6gpfd1xRlVUaYMSBQvh9jtOQmH7+vyXxNucOrq4VdpVeWhPOjwnnrdH
360myo/rdViotHiHKyamoEUEwNev0ppMYNFSp8nE/P+91M1R/nuzkdT5NR9EiBIp
rsw9xNYPXUYMLC/LsSNdwUs92Swr1+RRejmrHTTH1ZbZrQzZHnVc6sUOvOdMT8uP
VzjtqZ+8zoPjKrnfB/q/qhpjagBVRlc+DdGAZBtg8cE3ysoe/nAt53Z01AKezRGT
+qwgiBHVd1ckXi6MEIlgtI0qDRpfI18pbUR0GAdMIsMwJxypMhHZoUpeT3Z266PA
8rnNKzb5pw1ndX+Iin2rVgSSfMKkHVlmPi0elvwge6LtU4lIj0Xoy8tcfmV7t75i
iJ9ukPu0mtVRcpLv4kQtCVK90nGdFDVyNhPc61fMRjuUfYxQGAXd/ocq1XgP/0bI
nShkCzGtbM1Da/9CX4lJMpoHdShNgEAwrLsbLKi7qQu48ijbV7Qtc8Bt/S0vlGax
g9xBdVuQkgIdeF3dERKbPa3i/A2lX8rye7+YP7eFcdB6pZismWG1B7iCVIsFfJF2
7QQ/SmViG2DH9a7nyBFum4jQPcr3EhABgKJzOn360ejfhOlhrABup6IpqVKboZle
q23CIuv+83VqoB+HbB4brG6aYaDqz+Gq7GP0a22Yv0M+VoUw1YRZS+uodzfDSxjv
6F7TXzGsJqheK797y/IApWUrdyR1g6cC6rxylHuoOYWClPI6Gyr2mxnkOQloHPRh
XQlGoLs/pK4ZBSkOld+XTSTXcpyLn+dYa5AEqNQ9PHwa68l/bzx9IrhWHX40TyX9
bPr8OjTex+rkgnpfkzMmS8ttTRWY00i1jmGhRKi++guNN3qXTfEHshMXslhme43F
c91Sm5zbGWkUNq0A8OdbDS62nh/UrU2AvgDkkmonvJuGjJQehj7jeknrYCqorjlH
3l/4ld97MXv5/0hgry2ChrnINzhicDnGeqFujtANlYRA9sHWgVqiS5Nk0Zx6TFkH
stFEKfpT7zaFgxsuWj122CnhukEda6s4aq9xqurNvFbqeYygrH2EbhqgjqqSkhbw
xr2nB2O4p+EU3PZbOPQsybVkKjwmAg3Gf0dKgbGN2LyEN14JU+z6Ep97sj+DnjXf
0Wx/in1ohPfLl5c+L9E+4RYx3A0H79owDiz9T6Ov2UPJrBi0ryvFc6gj28MOoHyd
WL1mKMDiqF28va+CJ1Sgwkb1MG9Wd+bP9ifNwb2EI7ED4B5dBaTGtbbBMB20VUtw
TvT29u1fNy1tHP7ALNMelpuaNBd04yFQLWZDc7x3QRU8hP2KbjSUXF1FnkLOpHGo
UNfvPrAV9plxCgqibL6zpDUW+enBpAnkcafIcdtFEqDyPLlFPwlsDdu8qrR00Nz6
puvONtyJq2uUGNGj4UJufSOcL7GMJchWqy6ySOGJu2PlReHMT/xScCtGNMT3h6up
1ijcIIP9I0bWbkQKEk/zTDRap870T4V8FV1AICBcigy5sf+R8Un8nfPWCMpzbrd2
AfsnDPzZbd30iK9q42G/5xzEyE2Z6msdU9ByHcoph/kU9YhmBKzmZUAl4ZSZ3/pV
4RFQ78JJFxGjv35NQwOg+uiGKgqX8TO9WYunbEH0QOb6q9vT+HsFggOlSl4TOZsq
Bwn9Mw9PwC4LuLcl94dJa38khaHcdJ5jZcS/PaWfVGsMtiQdGfj2jtzfGJaNWJG1
wceHSGBJcAz6iCrn+7IBLdV8yXrerMaFrsuPs+RMJV+TdDsk7Rb6L7gB5D1xVlf9
uQHU9PsO1Qe4XzRPXMwtXFG6MCS6bMtR2OgkI4ZHWe+o37wAB7EfriAPUIkTUMB1
cv9Ws5vy0UuEkVHG7TbR7eI65uSfRubT2JgGHwsYX6b4YAsXOSkO3H94lHELcuW1
S71ESjozBOrfzhCZE1luxUaRfaNLEIM5TyxqbsLZE8Q5mBlOVKCCvo7YDvDzjuJq
FOtoJBtWLP93Xfu40l3/LpxqbcUZt+VDjonmRmqIXijsqDuH7yPUzYEqtwVIV4di
IaYxe8vYg4nershK0ZMs0/jGEVPt5sUDCXOMDL832eoDULqkTtfgAa1ntTHSoftb
c8Mdcel355p7vB5UevnRTwWXdN6rHtBN/Sp9DhaI3R4gxdb8plEybyEl+m4ZjAVV
FFDmpx16kj6wrnucHtiL0/o974Ln2FGkIpp9ogsrjhWzYxTp92zKyEf0H3lGQJzk
VqaOala0Ajp0+STGXCOaj6BQ/9quUZCYI6ubZpx1iLLwnOkeHVyPFI6Xbtfju1GI
8/e6Ck+g2cbufxWlmrifIYQb1pj/2Pdn1JUI0IBRg4XcVE+NCVd7wqfFRRXZAmgU
kVvSljBntHmRPdpjf8QR/J06UGqMlh1qQpLRuGbWSLg6zaLgSFXfvvZnttHBQyIt
F10gutMd5p2V4tmQzduQ87KIIuPk2xOCYl9yRzI8LMZt9MJXkA1UT8GcuDNlkuq0
wwlp6Tddy+M8xAR1vnlFixUzofdPDy8B2HF2F7+dc48921dG6OOFBnicgCJIjXsO
/vdHYbwkm92LO1qrLz2GsHapc7cTP8/YuhBcBkPyba5zzefKuI8nuPVa9RVvpG7d
LTTPpFHDTU6VEiFj+cDFrXhL06O87XlG0CktmrXFsmImXGbrGAhdwKWgLelUn0Rv
6sQOC575xN+ka0b31fs3u/8ffD6Cdq0aBRpDGM8DT/M3P+5TcM6o5jDTU2sX0hoH
10cX06OsxzNFSrCzql0XGM7bRnVSIy7W5DguyALR76PLLUVA10II08WBIXIxFs8T
Y3X/eCQ4hJ6KeFHRa4SaddKiYVa0rBU1JfPGaBOb3PoEDnaIHIhRNPgh8zWsDwXY
j1BdJu3MR6Hql5i0kMJiYqRo2qtFhs3eQSIKh1aATVkjfw5+6wyYw+xOdnaerIlD
7XsTITnxLqXeIvd26qy8hutkouxLM78VfdbtrcanOyt3ZG9Un3KsGrno6WzX5pD/
OunaXvQS/8A1MnISbhsA6XnBVBtpo6EsGjlXb3eqi2OOlH23hbhbsTCeLRawQR6x
NbpxIx8Es53mfcxKaLlWrS2PqM2cI9zDt+cKzuiiczTSVCt9RuXvUXD4dum7sdZE
+YSZRRoSwtJOhH3DfL6e+TR6oFHZnMq43TV3dCsoUH+4SCof0cWB/DiZjJthmB5w
itAuyzwiw+itKjohFBcqS0iSapMbB9wjmL2w3/649wvhN2/cbRSmA5Lw9qyUiYJW
2SzHaPa1VGSULouCO7dWEF8RHf4VsvE5p8YE0mK/6BD62kH1c4wGnLTZUhsYI2TN
dVoPRfHxi5R+LhFvnfvSDBwGxXi+RJP8DDHmYUevFQMgGluOzcdhh+kEPfQpms9n
WgIN8o7Amh18UOdl8ol8trxVajJYMW0H2/BKAACXKHAWBxrXwoOfNBIL3x9yIlaG
c5FC3/R6jxjL9ri8IouMs3v0s2R5ZVV2OXaCi9iRbHBJwS2rYxwqwOD0fEfBOv3z
2lw/HESnp3oaCk7n8JFNJCP3waXAVClvLiXamyuvW4D31xNI7dfNSNeEMhxIDTcb
oHDSRY28dVhu8jJ7oDkGfWl9aPk7zve73cdo+YPppZYy+vZIBk+QefPEO0OxpvKH
A8XfcUOr+6MXYmDCAOaNpzMWOUpEqoxDFQ0cNGflj/2H1hZ97SNVqXw0ZIeJG1Oi
ZdFh9kCDGOdD9jK709Q/4kHu2/fjh5p3dDbNxaIQppcL1BrQOaZpi/vuJ5Lv3znE
if/UDMlS9YodbXom7B6L4+R6lzmCl3QX3ayyZh3uGAe1dDbgNIa2YF2js3rrH0wz
IocB8jHbUOunl12Pz24Ohu6iHUL9yHljPyE8lM0PMgiGcV1QsM5WyWd+NY/+Hezc
tIV5hDUekMtJSWG7JApY5PRDFQwio5kPXCESQKr3D89ATVZuw/6mgMca1d0aPQtg
nREfKMcfNlPc3vpo+rdVPTW/lot8lo0tYsoB0U90iDrJAMThDRi82rvL9Eag9/Ck
VMT0xL7TxSCW3oGOsraGtQw0fk48iC7kUR3E3JGSUmICmVuXT1z1Dnz6GQSrksau
hAoUgNwgcu5tqZ/WIpn8b0o7E3NkFsYoITufz72GM46ZnpjdFBPq6Sitq4YUvVWK
reCbmBt4AvZeoD1F4oyLDwbEuuPRmk+jNhW9l2pUuJT/8vGW89pSvtLObamYGweY
ZIcqAMm9V9X0k878cS8siiRSzFAyGQ0960Cg42WBrsztaiLft/AK6S+WGm0p6HMp
HC1AIJhjuMb11Ay+6Pf096EpIbMAUM6nErykY9EFZV6bhv2zgYs/pY1xs6NfjK3X
LnBcJn+6Gj0m3BDRWZMHIR+smALTrmWabW33kaaThzLeBg34sR2c8boKHOd/JhOa
sMjoLLD1lKSITmi5leZlIYyOqXeF+ynvpHQ9ShlfEJRHYljamgVW/IS1ZcDacW+H
obzi4tsingSpqaC58krkfUnLF3cP6y2UaiPk9JFOobbPL9LaT1zOA8IrQFy2eRIC
4OG9yKHKJeY5g7DUfTZ89qsjMJhTiCt6Utc9T/+FqglHUrjWDwSMm6vDuo7/x/0R
LibVHboTLrWe4cKcdTbavYQ01stx8kLyW5Tymv1F76PcLVg2u24hhQHkS7tKhv1j
nbfgsmHk04ZbcCMVRF2fRHK2qJ4s4hGMhjZV19vYGnzTIOfJvDUs9yWmAiBtSyua
dbe4IwdiRsby2dJMObf2a/C+LwRvXq9mH4p7r6xy+oZv5rhEC5tTlGH1p5+YeLEK
iLB63Yc5F3+j+gIejUQt1RRAOWsQNp2w72Q+5QOuVFyLJTHECJa5vp66xlkBfkfp
PYc+Y6WC8Kp/yyClEb9imspucQJf/jOYPPj6FHRPmMGLHMUH1nvS/dL9HXthjThP
SvC0KLpTD+Kpwf98Z8Qit7lqCf7ecBynJvrHNyWEG5Xo8x25mBJE4yUoABoYuo9b
7RrtOsDe3JhQ8X9DaB5RMQz4sqgrsQv9/HqKWhJnF1lhstGfUWJAGI9pzsBmBIZ4
/P/ZG9MQtpB/lEEWYRBkRLj12pl5Yi9t6I/WUoVh01eSYSlcUUstsmrgvji0ykWX
t8dkhzwR5pcEtOgQh+WCjiNSsit2r6k8c1IulAsHoqP5aIXGauvWXvVVvCYtfaxo
+VRdE5/2Ts3mY2dI4kgtL73haM0JpXOnLESw7GqVsMlKxeNPpUCAnLNdSWYlXZdK
hn0xGp7/GiVWXCKZPnCgw1Xo/cU8kWs4jsGzqdh4mueF0zCdtREIAznFFj3NWvR0
yGa0WKUGuVSi31I4m7Asw+sTBLY+jFNdsN62lu62ZaSE2zfZK/t5rVjNGb8ZR2tu
4ZSUWHKmUoaCf/mYTpuJoF1kDlFqDsH0XFcLgajpZF7Rdl8ziCYRvRAP2A8kZgoj
f5WMua9h0XZUJs5hEwcGIC6Sg+TyhfDFF4JZUrQTjjc9M2KuM3UjjYD0YFYAX2Ti
urLcYZpzAQCGbaz308Y3UH5pvkqYxiY7T/xqQbsAvAMO2GrKn/QcQyAdS0QD+zRh
b7itYHm9dUCDIToZW1CXm/P09ADCyNZC2NDSzENaB5kqP/TvOr2qVdXIknr9dYk6
vnkTbCQ4ydvan0bRQH6mmxDoTHMzg3U8R5hv4qz8xibioNBfKHc8zB1JPt7/Nc5x
3nHygXiJvCrxaKINdQ8Fh/cXnYBZyaZYWeuYsib6xb3HUMi7SRmbXB9TiRDG3OdH
61dhgKlZSAQNusrB8zH98qaH63AA5MYERn/jpZjIXt7kvInRSPK91Adt0lvbWkVT
JEo+g70Gnkq2mSPzIi4ye9HOocXE6Jlcisdy3HpPobMSD5spbjKJN/e7/A3US3Av
ZlMvqj6lsQG6Y1IvV/n1q2fUCEozD0TEjktisHQ9YPfXvvYE6yzZCueXyMQ+uMx+
aRBUz16kX5UlvqoCQCB5BkOlRSZw6BMiQRC2yasTsv9SRg1aKpci+OF3J6Unj2Fs
p9PoKv7RNoZth8tlcLjIIPERG+OLaaqGK1WsllbHFrRkGyAIzDFUzo99O+F7nHC3
SO1uOSO06PG5vlMjxclSVY6ptQ4WoSpah1bSTsMskvMPl4T4XQQa1K691DBBgFZU
l1ytQZAshUSE+uVI2bvMhxRMDRsEZg8q/VCFcZsOf/KOFPuggFGIwTsYUyP08RKl
aZzSg9brjdziWMxIHFYrVp4RkPnnpAxo7V7I91i8bYRID2b9VsnkcosqZpmslzCC
ouhJKOHq0UE6FmJ+DXkpC+mIHINVPYOLkQEBPhbmBm/X1N5pftTCsrCzSvMCBN6q
pRp7cTxA09gZBCd8QZC0ujRlS0K0IVIX50lmQPGVxeZve+t4Jtt+g0skMSbsao4z
BnXR+N4YSkm/ChMtNoThpVrtMZiGjklmG9Vx1klPJoXRXk85NRIgAcHi+S6jgqkt
FmksN5oLJ3iezj+dKx+t3ZsHE2M+GWN4bjGchU72FcpgngKnpnVoTsZ1yQcKQQgE
8+QAGeE1TiitoHMkPcWSSbb9HxFZWnWi+YhkjeQXRXaUT61MowiKWdV5M3suM97g
x8ce5RspJVjUfJQpqBhpNY04KqkDeeH8vjZoXecEu6vtGO4f1bfeShybUJSEMrR3
UlarjW8waqT4YFBokIUxJsakKQ+TnMWXjuLV7CdMY1txjX/SrGvm1oFJKVx3LaFl
xOAVThhjsV9FQfiOU3XDwbzahf0DXe/ojBmDujF1Xz7B4/jHLpfTQbk4pLcaMd91
J9BaPPnwUTXtsDlKAJMBKfuhz55o43Onlkm+xlPHmn96mVaVKdHXyVwEp7Wdb+Y0
ZQgUaqJxn3y0NhAJ0xyfPmL31/QNqRmlSOpUqFpRR9qJNJv+G/c1ewIVS6FpeccJ
BFQxmVNqUjF3Ub2HsyQPEdhXfolffy+au15rB9E+RJAaFcsk5V6aDX90nCSghsC1
0oBtLSvCwyrYmZ3GvQBCe35y1wNj29K/j2Jki7qf9yogG72lLELOZgF7dG9yeAGf
VGOJPub+JJyAav6yXWJoQ0N33Rci3Fp6Za8gUOT+3yOiBqLfEEYvnZoxNE73uRS5
D8Az48Fe7nySF99w/FPzKGfxAuv/yRhODcjodt+b4sNtaWgeYxIY2Z49o0EVZQaK
ZBYrCu1gAlGecKzbJ2x7w04/6/FgegtC2PkuvBJPFvPurI2jL3IsqQwguLe7vjvW
yzJy0zvOcCWZ/t9ikQXtSei+/MBJYwyti1FcgrTmt/RIoeOGhyjXF7xwwxS3qhbF
0wEEgYw/9qIOlZhXIZpEGLaJUQm6EUEIBF0TH5rVGQGGiHXR16BzXt3c4rzchB1n
jrv44rqqe1ajsjK1Eq2UA8g5K3195VwHqK345loNZhJpcl8rlceg5JM1XYeXOXAH
evksGZmgiH7prBdZtzAuTGuSy+EGHGI1//sWQTxTcF+uO5uDzG5QURJiVOWYhk1Y
NGaBFZJrp0X7ZLNtCIcO+kXz9nOzJCVDEJPN4lMEZXDQ7ZlA8lXVwdvAjnCZ/4UJ
wo+vTUoFrvAwjTSJ65rWKLKT41K85Qk6pB93pyok9M80yN3azUqibUPml7EC65FP
tyL6LFgN34rgCCFn9egv8MEKmxeywOwsBVeWiGOT6pq7iDg+yJ+jJ0j5xR0zUKjG
PLc/8BNjlea/Yc4XrqhMultyAuyR4C8+XxpQg+mxrs2FBJpOQtUD+SI/pnzFk1AI
RPwWuFdypA7FfXz/m8pRQz2CeodUVvAvzuVyediXcXlOLVKI9S1eI73WQQ3HE7VS
yMc08/QYNFrb18Vg1ck5dB5R8eqBfNY1k1pWjiCdBYmaB4YTiDysvbyRpBR/IeHe
k8+HOpQWMT6MCqPgLirOdd5INXiV1Lg/GwkEcSSK6FP6a+AChsZwYi9+d218cFLQ
wEB/bDwszRHOMqWOue48gq9t4dpiKjRjR6twb5Xd6pb4W9Hx786l19h3FK7SKeNc
whUquWodL6r4Vn2D8Pn/2B83HWqGlgoS7LdRuMTQuVbCc58G5aVwiWvyfMgGPLuM
VxDFapNf37cML7vRM/9mEc6ktC0ajHqdti9RKqOozFZyDIShIj77Jh+CWGnHE7eT
ngWVzf0pyFgILsdcwatmxHJnSsgTZm5vhocv6gM2+J+mdBBYIL76OY6ZCyvnC3Ni
KOhDO/hNvsgpts6JodgnVko4aopLe0zg+a6WejEcioogdDvnCFe3GpVAOqtzAdiB
wEPYc+/ifafsLSkAU6mcpCOW8saaAgLIOz1549lcsq81/TBv8NJBUXKPiVaoN1Tp
cX7dgTJb6TWRV3YAVKYZ21BVOcGpSoh2oDdQT0R0wdrkx9pLhK0ecpxAUlGxRl95
CnYPhjvXAuBICXmaVd0TW9FEGxtdcAC57W0CY71dvMS7ASMB1aDF1acTI2TnWwvX
Dl+XjRUSpHfFkKx9WVnTOqUHSngERjnRctM2H9XMwBQwYkXG7yiZFGHY7AnlkvZG
5S400jAsieQwV9FgO9sArUqMw+XQEW/FxnHE0KX22kzMA3HnbULIJuhM3Jq9vOVv
siz4oJibqvY/YOmsLImgyz9cOedN+9z986E2i/jutWnYBb1u8S3bywtZ5t26Ny0S
n2zSost4MZIwg2IFLXdZYuh2sX9T0AGfeLbqZC3a5MBIjD6IdX/p2sxBjAgf1xie
klrXzPt45Xu1cr//GCCxxWuAtlosIHGSK4ljeyNaxQEG9b2TiG9agwFj8BI4XbRd
CkaWe++Gwz14Gug1//9kBPBbbzUW6xwTiXXHuYWvY0+qDueGiUq1tSBQhSiKpACS
YZYwlaTg/MHYcSHFXUsDutfcH5FYpzlg/X2vc2jJmdKt3BmI+rKMpUW2QuDsAM4M
S/ocmTjdyiItTJj5GUxRx4f3l1vCh26nR8r0xlcUmcbxIBZx/+CM2ayDCCPM/W3U
CWsPx1l8g8gPjr1jUiy6cp9ddfOhvce42nJ1lgP1sHfqeXIA4WntHMvqGUF/AM/2
xH/JhCbBSZUmNmMbqFBVkPMioyDcdk3bP5WWSSE9+h9F67kJIcdkLOu5+FmTScUY
N859ird0PVJ5jpi/9vjvfjeU+zYdaB4oHe9V1isG/LTTxWLDZDrm9qY0Ec7u3BDt
tq1EHafotuN6RI3SUkWq7t3KF4ZyyzgMT3ESVRQ2II3VOhgJSZfdtas8yapYFHWu
14/JoEJQY7uQWoxE6VEmacw0FiGWCWHRv+amxud63Q0LOM9q6gXACDcD6WJdQN9q
ZNbROOrXhFZSkeS36JBC4UtK0ghAJEQ8KEyGxfkriK3KZkwKFhN1cKq4yovrQZy3
eYDuGpo+NU4iUYwOr3fN09lgjQzgFuyoHj1Kif8jW62bSKnKGq1Piy0adKSJJaFP
GuyiNeCEYLSuI7xELNtTHM+SuCnBKjSlgAH3BXbCW5shXMv8xnF4t/SFShnxvJtB
3pST7F5/ZZknBLqELDhtvPLwyFnqv4c0L1me6GCMDSkMUNmdQf+W2UPNvcpgDKpH
05cCBRhvnhfR2O2tWayUlEaYWYdaSU/gepPW338tQrX172GKf5rDt2pKtwfZR99K
DJH5XQQROcYZk6Xxxpu7I9oMo4J9uLhDVCq3xQXOW4AJPys93vA+KNnkWPGHQfMW
QVIlecqe6udkrVsgePh8BmXQesSk47XhPnfvAiKSz6AWSPFZ3NkMvuQ8sKTLZQBm
jT3aZFrd7LHfkdqnSommXg2ibfDHcxhpgpIgXPQMKOLAm5Z2Cn80HzM+t2t2iGP9
7Tap7Uzy2hj7igvWBlwQ8GrBdIuJ0SKo4OZmjo+0sAaAFn2/JOL4BshTik9WzzdB
w1cvZYQzUo7ci69iNJL7442x076/qn786l/+ELzypEVZItlYttPLiTVnCoNR4j50
v2kb8oWE2xINizfoAEwtTf3x38aEBpYC28GPBo6M3NuLEmaQYvXlLSliFbsf4bc1
TOw5pNYV91Zs7yBv06iu8lmIHOTiPABoipFtnxXnAVmq5ZY09UZA50q9IEqjR0Jz
yHdZC+5kePmWjWnys2547DTYi5/zaZuT7+83LWS7gDcSlAuzUywrGgexHUu3ZgZF
2bnATwKUAfoGb1SYqvKsABwRJzPb0mhZvJbGxqWC0v5XqnW9gRELRuxyNf1ELG5m
ycyS2DvKtLs6vUOJEfVIUFmrvtGjx3GqZbCpWm879O+XFo7YdUyjByCQ5Vd6hYbs
PngVmZCctbAPkrVcqtepBnBTyuYHCnk5Oe1s6HyCxpYlC14HWOSbPzHhGmguODGk
CM92MHEwYHDhE5ccnacmrsMteWiaY+qOW9pqfn43d9npXpfSHeNPN92HfwlYN5yz
mMEb+30QO+LmPcZdKskc0Wawqkt3pyY24jWk2390pvDSHWui5dgAWbRJKG+nOIjU
WH8OH8DGydQjWRUM6Fxz+DnJ6zDd/nUnr7k9u9m/LhD4OS+kTEgs+gfJcJGRJVVt
cSI8n/YGL1reGMg2AZpICbFdFW4dS3BT1LkaYf8PGCGlYwYlF1YBANsaUlc2eevY
kb710l3lnLI9u/gCZ1mVfk9Sxomu02iN6w5+p/Kb0P16MpAOXoHDbPCzIPIVTnzw
3W4t+Erxunrge+0eI3SOFEI+O8Gd1ril4RBBENqMxjzSF6JXR+LyoEqEm4CfqUrg
+9dH6PA/HM/somnu3Oibcrdxi5Y9QoEQrGUSpaW90x7yDnPmMo8pqX5DMQIaULhv
uQbkdO20Cn4IN0S079KpCwe+0t5OrDe4umWaYcvPwQHBUTsMULlPYYDmcMySIS6M
cAD551k0GjMOIY4ZiZJxQLgGpOx7CqtbVHTiXYFeo8iAKCz3V/3qTH997su3FFIV
6oM/4f2ubUM49b9ckYN6kGWuxDhK8gESQddSkX4fMXIu6Xp5LrTAdrVhnTzk45pc
U5+my6gGaJrawr2JU6/HQZLf4i9zVjJaO+RaHnqp3kaEZ6PtZLeR3otYOBsL+eeN
HWXJ9UWiMgM1Be0z0s1KWxrufqLO0a689Zq6AOiwaS4ltdNtgqDfcEXYSq6/CBj4
au/DRjkhYFm5YnfnXe/bzNHYEcvks0Q+CT9hFr5FhMYfffGz/zTTIevsLgHMLfGl
4p7sT7cCnG7L/hkmaJBzcIo6EZbY6YBO3v9cRcfXeDK+v2u5/nhUTgHCo5vdW0lo
QFgdo3i7E7Xf5aNNzkKYHYySNrL6xCazSka+0Up6hKav5XRowvhmR7OfT5DKQo7T
yVSjbYkiHHcEqRQheP99wQKqnMz427h/lnhXZMlM77BgiGqZvm5F2W1y0eK++5fA
jRgc/vIEMDbU8N0edFRYRgMeY99lJzuB92JkUv+QQYa+BPFKHPjPXzxCSP4zL8DI
zl06516kp+bQ861eGoaPMc3jFUAYh5BHnJoC6n57Dew6ycvSPzFPJQLJKlcFOhHc
Nto62yrp8eL22Gm48M2k8t6wOTB4/Yf/y1F+P+s5awYMiPWwM0p3farqpcwKLo4o
s70veXTSs0ygjiNVQ2D0j/Fh6ocmVQhvV6JbBJN0ub6toriQ+AbWW/HDC24V5hOM
Ge1A5rsV9/dV+/UehtRPm0WYOY30QrOkkF5aNpwOhKUEalmO5kB42jNwRKTc+2yT
YbzR5Im04sF7U2ipjBFh6oMUdk/xw75JPn9KdTQVg8ospM/CAOFv/ZhtMncEQbED
KeYjHE9KnjarsJ/QuSRqEDmY5mcWczuFz54PF/fBxg+CxmTmGlslLIkGRyriMljY
jepra4TJXUX8NTa0ppVEyjfMXgHiAzXjDWX+WxmKZBr/j9fQXN9zMgTFuQ+P2FKC
r2FVEHbsg2yPntNkKL6IJ4SHPzyKZs+iLBjnNsX5DnN2i/lW3+BdwhL7buMzD9tK
dq8HQZTD9iuPyzbirZUCvaZ9vbTlnVROSffpQiz36BDIJd3X0Euh0vzJwrSk206M
HHLEwmXYehrjBAeKBGS+8KlprRl79Xsf+kh5UxoOin2XNc7rQgIoaapfj8ePbWUF
Tkl0wo2jGA5AhYLO0c/5UmpD4Rkvz4oAFr55JCergcyNFbh43PFRJUKhzeNwn7xW
bmMAMLbsf0CUhSQETr/k7cFNf4PXlkH+2QHEiFRL7+PvnYSNjFOyK/aVZ2JFVW78
rjD7sUJWVpBY+Zz4PFmbE0l+PGs/UAn9pbHZ0ftkDtW//rAQwD+BkfuMfrpKiBwa
KjS5b+s/6bYvVxM6Y0TqsAg3fDkZf7Oc1LgRltBMA0OZd/27oVwDVwarQ1VDmgr0
FqUjgdxVl/cEDVTYysNdDqbYMc9MHNXNTilNtmMcHOBZBOfrTx6ICNxd5+yfWxMo
BhZtj9oWJATRY8ZWeYqspLF8l7EKZ2yav+U/hO/rEf0UMDYXGezH2Mw4OUnLH79M
Bd+/V0j2+ObYn/3a8DBawjbutuK9N7gb1vY1z7FafWrtUKugmWqFioshkderZh1L
H2UrfPxpu+NWTDoJkgUdQn/ZlGMHtle3r9UwIC2nW2T6eNGsAJLuxyzi6a0Vy6C0
DfCFlbk4xWGVJdDW3gyaqfiuzkYcM+Jo2LlK/rs3NjYYbultBTBe/Roav+mtVh38
utOpIaaoWlvrwBmatVbq2XcEdJ+gXXtLIivpZH3k8YqEKEy+r2SgaPQpPjo0Ob3Q
Hwr6QtFWCJkWkKQRIwE39f1Ys4WXwFnN1FXBdj5NlhiC/8ddKpRMcwOzeCep6WPE
uoUaAc7+kGmdcLVKKXCXG/hwKqm529oKKXiLChJk6cjEuVIpmuEhGYYK50yyXUQe
BSwoTDBmyBx/SnRskp7ZqBpaJZgKnLElnEYre9z5YXyi/5DYta4Yp/IAyLxRAjMY
I6R4tz2uOa3ATk9t6zOxf8kCuGwuRp0fjFPbWR2pIlJ2eNlA972JsjBl1WnMWQXe
nfpj7sAghjLJHWL2GCQQ1fyupZx+FXrwY6S9xPnKOqBJM0qcEqAqGz5/uX8zqbUA
Fjq/HJDS3IHix1fLj2zGnX4kFbsEyBoZ2Zhu3cmv6FfPYBxZwARxJrA1UdElDNrU
PIs7unw0KltfXxAJBcV9xD75vG2d1ILaCNyEp3CiQk981nzlN5id9OC/Ie0xFzo9
xkFBeG7VWVBV+5MTXA7EMDYmALR7H7hhGrzZNWrV6E2YBufcA91L0BBBmVh+xlu9
wcGk0+mNZzi7ZgGlVAUS16SvjD4ZZAEUm6gy9SyeaHkz3vRUorOCBXoSM0ZKbGCg
XRMolZiOTA9ps6iclg4xGZIdbQd95DbIFL7xYNF0UB9Moaui0soChuUjRZasd0bi
Rg5Snoa40VB90HoUbtyFkiB2vJcwyd+L5khZhZiRgGsEn/TuE8W2givUH7tOdBz/
3V9YSjiDXj2uE3F3dLt6RjjYGTgeG1Ggsmf4GK9n17IR2sMBvhfJpO4ehngZtPNk
f70mUpVxHof+YgcyTD58eSeZTxTKvoIo8kATke8SdzWQrH7iLBYkXckiRAlkUe10
3qHt/A6Z9Fz4tDJH8oUeO39V66cw3G3jvNoWb5hA86c5trnzSE4am6CYJBx1GC6x
kuj2oQCE26BOUT209a1rSboBaTTeCL2017MjJfhkxW1owaImCprX0Cw9lbVjfh1E
MqPQfjrFI8NlL3R8lqLolWAaAEXzBqpeSaIquGBIhU9B1uaQLNrjG9XhbIy2aR1w
I/3B2XBq1I13527csxZCHXVU3aUti/Dhn4K6gAfdem9d93v3ETiFj1QT3uXm6ITS
+Wnw4ykq287InSR2ahOWjB2fBdScz9CsNdnvYjxkCH7B5ncz4i1sU1i1KeLI3RUN
jXrvmQTtd1MZbXxGIKfPXLWdZcuLqpwHxSoN/QCzsEgoqkQa6BDq3UktHJ1uOQ7M
LPaysUeVbPUcknpF9eZzqlLR56RnGUPPtvKGsi70JaBWHailyHIUfPZnf2G1ssYO
8t0G7EKezHUaxdqyt49R+Fl2qpOLYTJ+KPmwcPCV8TCg8XOSkZ/otYKdNczgHXKF
a+6E56tl0FXeXGlBLxJLDCMDNLqfKYs1V0hQLBSOWDZjJfkrC3Fn9uaHGK0ipkpT
JmBOiN+bNVQP9i97Mr7ynIKnNA2AZnSXx+5zJ9TxxcvcVfrCLOuxv5UnKj2xwedG
lETnX8Cz4LQfLEm6MbUPt1DZsECV01JCPVc7p97Q6NCWPDXGR76VP7P5xS5lpjYW
62XYWMcgicnb0AWYo+0EtLdb/Y5YpWhX3q5r73Bf0x1iVXjTUFCB4qN+WcrABg7z
HGTidGL85256DzY+EpRrdJ8sm+PaZ67YUVGUjtSLvvk5MQBj65rFtjD59VESgZPs
RSX7w99eDyM3lgsGGydRFzDxwRNFJA0yOjh1DnMa0aYbgo8fMc/RGZolfiIGAp6u
2/lm5cNmvz+XIv37bYCNd2Ku3WJ2JOAcO5LIsrgJXABzsAmEM73buJbmpmPPKpd1
kI8Z4gcaE2DQpZlBjoc1qMnKWRh3J21e37MI18WNB9xIb0z+6ZyfoaV3Oj/ic0G7
ZhvmLMWFk7eVwkG5gB6Tg9Sqe+FLo5f5oFud75nZO8FLf4lJI0IqoRBabhcUhbjB
MX2VWQCa/ZAXXw9FuJF41SpCzffTdgsQQbv8xwI3AbeaB5JmXO1guZdLbPwhM8bD
IJX+MPcnD5wPR5GwzS0W8niBf0LOYLMQ90a2XN81ALPfC2qxpRXsZe37VPrrA2dB
fmnF2ET/GWiTT4CeaWQslMmO3pyCXqIh/zJXg5alfDlSMjGhzlve1jlWYxoB9BOV
jqry74IrDQga76LvkuZpXIqe8OumU6yyWo0DptKaXXogZHc/vADGC/QVKeWWAODp
7X5Ch7ICMT4c+D6sAOlicnDzi2aKrD62LOD804HAvkUdYSxEYtH6Se4iVgs4Ed5h
4ByHNrhNKP3v7pv5UQoJ/EQJvWeE26RpKblU60d5brC8Cdh3uPtn4i18n6APTPJh
wRpq7jPKCK0ZKNHwLo9XoWihtuG7tWJz8lC0wSgz5qUww/cHi5CYl4ovYOgD5UBU
L6KOmVEVpEEpUbAytpo5pyFjC2Mb7KidQwS+N2d1mAKMpHvv1/vOElrVrFr2omvd
Pl6qiGNJAXRim6X7/4ej1ZaecHLkff0tjt1qcZPPzlXZhbcA6hyNfF4bMPW3jJKF
vj4wNXab/DoIukxdqpP/fkQt2CMgUh6mA/bDfjr8DBV1EG0/2wEZgWvpKd/fqtq3
vk4PZjWA3fk/4NdQhlHVLzivHBTowh4UAZrbh1sVIBSuYna5VUlMarb0dgGTen8o
CoCti+L51llNan55LYDFDucpdpF3ysoCoi8UBaYe7amiuMcVoS8CQfzlVNqrAd1W
0VcIzSOUUX/qJtPkTT16cIzMgX6nmLlM73F7K6LF11/8unPdwdpeAjTH1vIdCP9m
D9G/CpSdFBdA3bLgLEK4XpDe3HNWUosUoIlqtKToWoMjTeYalP97RkRIf/H+NJ6H
VTCENBD5t2qDjaKRZr86wZh1u+msdXPwaGYC4REnfpCIFtrHZSpGWWrh8RzdFPWm
eI5eI5qptWFVTDqSMau1xytcCpKLPipLKpHY6eotWk6YnDgo1l9Xfm1SmD+B1F+B
tJb/sA6ddXNZ87mahecmo7HW/HtRI7YSi9Dqgk10/Y+4e23o9oFHgc+vgshDIi9e
EndEc7GaxVO8xkxA1baUnwyPsmgOUAd4EBDiGs8RrrfteGhmqpw94cHndIlkgM4q
YkjX+MxFJkCqu9Gr3EXWYUPQ91AkonSEDlsl0QPSFWoQ3qUxtiu0bsTT8QZZj5sH
iQCMG4ZB5L6k9H7v8x03KDvhZZxFQhwYlyNw90RwfRXmljVQrrueXTtiL4QdHQ1J
zaSXWSJr2ICtt6EcPJSeAwXsFsCWdMfq/6lrmVPVwqW8ZdxvVD0IKyYuAjwOzfAT
yA+xD/g3Lb77hLA2shZhSR3oR86LBrdud+hR//gtqTtbay0ent3/q01CWYwQk/K3
Q3hdeqiXrE9+KYxl8p9NN+2UG5mDsHD3A08l7fgZtyBGVbBc2NV/oddiweBxTRUf
mQWD3ik2Ty7eoSKghPHQhGYirFprOqBQwhwbCPn+tGyZtrLjQ44cXVXn+qrMToBV
QIMw2t7mbut2kGh1SthSyCq5idrtYvmO7quq29hOX/AoSs0Egj+ao2qoh2d0msVQ
pdWYD59c9RrA2adyggD5zGKip/a7wMJNXv9NRG7XEv5ER/g0nbGG5hsbqJ0q/N9l
C1RHmGFgeVeD+CkgsL5gk1BBDzRrjv42sZOxkgg/N6goyMNYhj4rOOs/F9NX12Pz
SV096BrFLhm/n5Lc45Bj3jXFpWoqUVqnHJFBAucLnjg9j/bywZPiyQ47hdM3+6Ai
vdsbu9BTcblM7z4OFYTl6oU7330VzlNSG4bpd2TURAHfeOCZKBWBQ0+xIRyQbKWK
xgKMwJohQ8kVIFCdipTAyJ8fc7E5e00r4zi28CwRxRWrMps4VL/utNU4A+xbxzS2
f/WiMk8VxI3eiSOBtS6URJrIGWfxKtEOFBXFQfh9NSsX1YPckPMeWcViIoX86YWQ
BrHbL72UAfuwad0m3VlmNI4QAz1DXjVp96cx9p47LcwhgzS3IokOuI3FzySly8LL
HZ9SK3IIePaHR0Grs1owOCy6pO8wk6LHxKjOD0CssgtpF9RYo8jxqa+JXQQYJH4T
S9RPIpKjy/844WeEDXPWreLdMb7io6ZK4g0A7ocvqRUjeTXog23pg4yY01yQ+NsL
ilzDWUKNobpNzVxfABPerPdRkczrivZnPL9hVEiHiCMjFkcqun9oL2MozbN2UdEX
w8KTsJmKRzD+80IySaImi+ZT4SpqSSguYjWo0BRBOZ95G6Ge8cGKNrYKPmgnnbAb
+5uD+g1ztyNEIebfks87BSD7l+Lm9l/dDsxZD7cMWq6dF2I1l3c3fQmVdx6+SF0g
QKIFYdYlZer4WfABqNqLTnNp26rEc8ccHVZmZ3nD4iydVObr8deE5Oh3Q2nrctGv
PFQ/3N4iEN9SxbF49/xA06MK//ipqxu9F3tgtvGOfo72pmZxS23J5zfdY1Bl6nO6
lFvbgORihI9MyKVmo79rNOi2t3PoK/TfRtme0t20i4poi2LQGgnBbJUE4ANhdNoL
Gg/dKsKazCGF3BBmdbAUvZ7MKnJdtUrI7DRhynwYNl93Hw4sISiZYkRDYCVI3gZw
NkX6opN6ztygxjfNWZqKcL52KUdtqFMsRtFlaQb9OlapAg/IUdQ6GS/334L9vnp6
PZC+3gQpSAInnelDMSbs1aMtM2QPmTjenWEKGhIseIwxyXwVUveK2rg8y9V0wVQi
1k64Q3/XXNSZSEDnLMAebzATFkxhOpmOWSAqaRMN7N7An4RRWQyvoZLZDQRwqW06
ByWxzDswHJQM7ugU4VaxF3bgyPZ6utTrDwgYqkxSZrFo1S700UUM7BYC/zDJqGIm
z+ufrswk4Fcdv3gZxpN1UAAKVug3Rsrt0aZz4Y6rzpWSva8NAzRMRkjTd/Bz3eCg
jV9GJVdzDZTnzPWdu64OfkrdF4as1tRNNh5782xGb1uJ9hAiSixp9+WXFkI35ADG
N2qyfh6AiPMlToa5xsaC8Bo8V5nB1Ho1S3aZNyiucpW5sXXp6ovXlhHRLZVqJ1Ed
zLv0o0DgbX/aAqEJsUCHXbEmcZAK2kyyKDPeGLOZ5yq4B7JVXBB3rQQikEQMI/cs
qYe+jghKf3NscqrkRDRx4S2+GaSc1xn0pSMJABGGronIWG7DGxUEAGqF0dRq15d/
x7oN/PcaKab8Fv5m/wnRnG8OE3VCVLT7OT3pS6/beU6d4KvxSzZgM+UIBhRnGX+X
A1+fD1vyV5E9P4HXd7sguI9kQ5DVegQhgFGaQxtB4on96W9Fs7qq4GBmB/ZkqbBV
ymBfEWI7CHjqW5LMrJZuUrPPtkD38w4+KKf91g8S/CULZosTPTrIM9Xh63pA4oaN
97AfURgyo1Pfh7J1hCe2gKEi1VufWUaBbdwFmkeO3a87QL7LgDd/+TLgWaUE7iqr
Dn2PCKpmVtIGjowk08o4SSZ3xoJZsRQ3lbcWwqS8Np85Od1gG/ZIR0StwTsFiX0g
VdN3HNhocAEY6M5ziGGTQT1eIDnRCqWIauvUSKYWqvurdFUNoDQrSjWUywWK/7Qu
Kw/KVWFxzMuR941QfRbUZ97v4p44TYNaUnEclVVqqQeBMHRrM9+Y6YeVNgKbrxqP
5mc/lEjgShqe1GK64Dq7qKTA/wFm7EJILTwQVmpzGoAPWn1iU7ZgMtutGCeZLY0t
UJ7d7jS2a/umxg76wQuq1KvYDnm4qZnL8dsO1GGhpc3Ajvn8dMWBtK2W0e+izecl
v/l469QUE94TwtvEvPcdncImcWVhpQHZVb9lLeChsqnYBpRXq1847Opmu08b6HZB
BXBRgls5kg2dep/ABDe/L1yrvAOomaJTyaw0gX0EoP9X5OVuiWJGNFIjerBhu/wC
AYXEMNxnwvjpH3PnkNDflW3TOvIEjGqxnqtcBkbfuFiMs1wyFask+K3eONAAG+NP
KCJ7kSw+CvWMy5BEca236N+9rhWE/683+n8na3jlV1R7FH/8TUy8yhiQChXjdfUh
u1lh3zHcT6R49SgjekgwqG6BirGK2odN3j5F5uxahkvcXM/6DR00Wq2Gv2QLRzRD
VQ3wQh3XxusmtvcUkmaKyEYdyuhZr+RsfKncZLU4pz3clMwrbAOy+L3JMDa5/B8i
/Xy7UPW/zZUzD35eOnBHXbTxsTW5IL9b1qhUbrgLZfIBa+7tSLj5auETQZIq8+cz
GhwTQzRJHxU26Yb6ax4LG+TuNVleMlGJ+NuEXDLoFwr9qcI9cAHRuu0jFgzeSfJW
0DhpVHmPfmXZlHPIcyC7EC7SBlgiTQrrOBrSJLNC+bUGkDPp/KydrnWkUd+6HqWX
rbk32d1cn0YRlbdLgpWlaLaU4m0QS932rFGgxuKhTKQefcuQFGZfzqtlOmnobnCH
Pfbc+f6ufiP00MPShaxabditDuyATB8GhNxT1g2OSHiSPrR3WAN0YRENd6YiOC6+
0UJQE8GEgXVBitZlPcKTi+FttmzG2zF5KgHwd7TTf/qcRWMApWwK/zs8jfZp5f41
p2pVDZVVs8Bt0Ht975hwMuoQTDDLW4pXsFrHX8hf/N9uWhm5lqNR9c/Wvy2XJSVy
wqZ+/CKpKTMWP1iSksqSCicLdR5H0OvFt44bqao7h2OGHB9s4ol0+xaOHE22izLX
G2to6F5IR3adz4E+BJA1dv1RKqSmAP6EXGRoAByflBJGHSer0rpvNK8fmiKKzaHb
H9APaKNsCsntl70kKDS9cRSp0Fk6VE90kj+7Kel0QLvLIOxxmyRDLs/aO/pYU/sC
rIXBNbefC8K84/dWSJlft3xQYo0aq2V24VmXQYLpAhXqPhYuYqOodrUur6hm2LCK
AkNixBRiBCwnEgTSUhly7BcsWNdqwyUNa6XyhFVGdtnxoSUuWhFeqsl2h/QqKDAk
1CInn4fvQRSAtQY7s1o2/ZHq/pLqUu8UyrYa/0hAtYca5neR3lxOGBXJzIHVxjGK
8fSKz+pbf6h7Lb2OkTX6aV5UUFpUorGZ4fVBvGZJ1Y9jC+6ApMGtsVX9++AAKBaQ
tXtbC5TiH9H+1DZ5sIGQILx9wFyXmz2sSk2hGxpNEPsvc8kNffgZeCbXQ5Pyd021
cl25UGWSKP9fkiCtv2fAYQi+nXOoaqMI2qlVzyLXU0d0WI1ehNeGDkXxZKfVuo0R
oQUkanElSNUObSt1yTKQS5D/vNiuQDhmobhcVVKPQcwUTk3iMpki0+47RT+K+i3b
KQl9pzWkmPLWjOTek9sGEwPlOujXsUuYob9FczaeYfNz/0t3yrp45TxUJ0ggOIsS
WJWQokuuQTmhbbpZW4w+nXYZStTKT0OefBZckpBhPQ9mewkMmMCcun7pIMzMf+RZ
B2+btslZi3cDALho7233qBXv6E4LhBOe80ycmL9fRVTiKcotb6TE3membMoP3qLp
OWJE298+18TkEbVFBMp2gJ0QCFbSmvMrEzNO+rh6SckC4GJnxw4lfZ0Dk6iJX2R/
8kUF0Ly5WCIci0ZyyDN0qKhGVclkWkovV3SjNQAoOTWui007ujw6n3nOVjfQy8Co
zULDfQCgbAzlpLxEW070KCW7mifVSVy2heKJMoWbStT93YgDE6rZI97XHPifdIyi
tFvA3UXTE+M6Ihn5w0eW/E040sfwnpv3VGJ9ZGp5mqkHpK47/uVvqzbx81kZMAE0
f2XsYP1TitX7MeQ5ozLI7kDsI84LKoXGMYqR8zc2PCVP9vmXF0YWLyCvDjBJzJSN
fYG0mLfe70qgA/NPv2tWgLYRm832GZ0n88rlqWtyfbFAvNpUJoMRSa+agdY5fCTR
JhjaBKVF/Ug2O07ByB3SkabGJwcwFOFhXPg5UmzZduYf6DaM2OvJHkihUPmQmRxO
O8udMSQ7Awuc/CIsFl1+eNT2XtxQfQMB7gS4Iq1zocC4ONVLIV4QdMIozWNibGjd
k5JRKiFAF7uRa6XoVp50i3erBS9H0Y6r3tMw6rgF3Gdcgp2K66Kx+ruPKfiAMOc6
7jfkHHSawHHhEfWV4YzUXGaSAzknNFs0l6b6QwKu8ZEdA8mVln5sW8pD1JQ5t44u
LujPN/BlHjgJeR9UmkbFX+n5UnCEQ7Abw5JY61ZVit1ueoFi2U98pOWffX/urQEF
ggp19EEywcKUJ9ztwDZTj3mXHVq86g8z+xHLpblxSdjhJRr5RTnmBbNfEeSxowSA
Jw+SIBDLMwWL945769oawnIdsyh9gPtmK8fjCddoG0EbLPhq9dcZ5mC4Abvz3a6C
VCreOof6diANeIcUKPlJ/7PEIIh5jXtt3Urgm7m7X7FuxhVIAppDfsGxOan9yEqs
0SwGx9ccz7msQdbSNZNXPeuNMdhbC35Cehc1pcpPoebr7sDxgvqcmSDtCszs3HLh
2E2d3FjyN/OHZ6hBNY8wSpWC9b5YF4kSjj7b6PR0L57Yu9Ee1VzZg82q2Ek/WRQK
kg3bx/4TmE+/1UM/x3Dvi9NzZygUF2buEXMi/Rl3+z5AuXEtDNJgzsw1vftWnt0K
MwfXTpRihutm+NCHFPUxgwgkpru7sYe/x2lGAb4qPDqb5Ru0oJI/q9QjfoHvB22w
KWNSMsv9YlxAbt/MwTfFRtljjbMRgtHjbQ62KCKSJKhDrAujTXnPnkns8agwGnLh
g6cIuJ7g9ZwDg5CmOiTZNhSBYKUuqQl7z5AI/Sd9E9PfHe8cfU1xGv0IdGsyhXHE
nMp8fhQ3unRcpo2vXHQgu5oy6CnX/I4WibGNoZ56Kcf3hlWi/UCEfbMmzUWrMAlK
lcPqq6TYsQhhNwdlpkU1R84Nr4wqqJArw1NhtyM8CUJLjtukhUbce6VPd7srWHNs
xs+K5NMZ+kaq9Kpra6QnpdRwGjs2e/2d58xm15ayBt2Z/mbOHYSL95BoC2q1ati4
+aKrI+Q4NMi+BnMNkCGRPkjBzE5UjsYwVD8irAtMgVmTy1LQU6gMRJHjb5Jnesdx
Y6J/2NyfdSX7YSwRQpLr5GV75Q4I+0Dup0drArnOp+THedsF/sSSgnY0eyfWJXHT
FOcRuPKvd30u6d6Am+wADrtcIg2rURhJTMsmWYYj7Ov9gjmTsXcdw3LBSF08r4pU
NbHWSNgPKvjsaeeUf3fGVA5VIv6JBIihBtS5LCNX4ofhVsziLIDFxHQB/E8U3M3J
buNxOdyciw/OMooS/Lr1QWK+z96lQQZFHtmn+MiLexTv2QR0UKzO/1s5RGRIXdG1
WI2iZDzykX4scB1qsrcpN50u5RXvTuI1/TmTg8Vhv8XmV7qEWvpRG8hmV3iQ2MvT
8X64p8K3yPe31fVey641A2VpzMTUsKRje1Z2RWpcp16RbAGhBdHC2nofV3wvRFCJ
yVQNxqrpWL3WGLMQo6YBMLxJ0MUohsDHGOixDFFeCmJCm8hU1KPkBhXZLmX6T0hv
W//YOyycBWS95yXfBoQKb3DHp9p2y/QeRHkKuYU0v9km1POwjGLIpV/oMEAemw50
UsbV61zT3Oq3FKrVl+ogDmO/lvvDXacp9iBR8jbA1EonuL1NsfNlX4FmBUAaCYy5
mE2MXivuTCE/7DYTeVohml5uGJ+FaisEd/FO0s4LDhT/EJGOO4BryIS0Kpdr+uOe
36r3RF6kGbNwirzdaFhHhEbOi1rf6komiPpCQMpHDqJf5IW5lJDZ4rNLInPjTYLa
TbzJXNmxq4gDbWBeXgSdpTx7MDUFScmvcf4ric0y2ueXOkyfnHdRGxiYvGJxW62g
GFj5ygHbP/or2TNuR6JaguxvpfBbzxX/BS0t3dDGXBQGEmcL3AI+Qt9+SEGS2Raj
Aw3sjR8fDaW4kHRNkiZf/oWCZ41XAO786ZG8SGPiQPl+aYCS1gz12XjK8I/6FMW/
S8WzfrdvTWe39+RJGi+K5PDoW8xCjlJkECMuyc0NI0a4vgON11J6sLeuJxVNNhqL
YDQYvWM6KMV0Yz5uc7W5JYvpS6bYqZpVQbg0aHGZsqG4Jowc6sZ9oBIlJjZxDBO7
cYiK0w6MHHF17IfY3+V2EEvTIYFmJIAIIIMI5tDxqZkwH3GCfdKmC4ppVRhAYuOT
LqlCdJTIp8ch7k6gzPRh1u9bFCYV6+wQ6mdt7Kr3v+owpPi+F5KIvRKt6/NMAyZt
SgIXbvDuRhOghQVo70fZgzpyztgV61ICib3+lOWPhXmAcKuGutgyh14PLxKxUTp7
9tSKHR9fHlZcnhJFY0ytBT+1xJPtlu9uO5dInnXyIMd1OYfMTwuSAHMZTxZ7S9Hi
mCbdT/MziC2KXYxiZLMyJZOueUFeZ1HxI+7ArdNrJ7nwUz7dzl4+A0yRX6RRxR31
d4D9E9rIZvqrkAJcxqY9RlTlDo0Enf+GIckH5jpC5U81Hbz96l0bL51LQJy0Y1rs
T9J6UKGD7WZW+vZqcDuizK23hd7CvlaOnDtyeFNdu/NyDPi7RLxwvGvaJRJjn5Wa
MmYWHxdXjwS1AYsSzF5kd/8nA8Sd+lbCucyMCFgERTgxP9s6H195SdCq7WnjIG5C
CONYI/j0z0pOFGKyMgmDJzkVne1Omjv5/m672G8URkE2AmE6rEhpu1Ql3umvKmEE
C5CeYYwcDf73hQtO+xneAanotWLwVFogzxBzUHaa7iXrApMmfd+I+11QzQXE3IKA
FCpmwUVzcJ4YOPja6sG1jzrftY/UM1dZHteK09+j5p2V8NHxNcoYePJ70zSZ9lbd
RaeN+wt1EpVnfdRLjeqYvF3KhHn9xzw6g4rtwJB+DyEG6W+JWAQ+B2PSf+70jBt5
SsDwQiQYviEPa75Q33/3Gkl+KjCg2Cw2u4C2Is6XpMXtjyzLRX/zzZNRWNeHO/wg
1kbjkbkDP7QOfkuk/myzCABiWnlc8Ncsea55ejwJa8BpHAxE9L54UkknHUOeRaD1
9BXfjc8xNnOltHTJDeY6YCrubqsaECUCsOzIL/K8IfS5lmTa+vXg4AlkEQPKSL5w
NqzOnpFdgAyG8rhDohGb+Ta1BTMz44qUsuq7XhuNHRRAallgE0o2vB6W/w1MddYg
lo0hvnlQzJVWK/rCUhIkOjJFO4FXLcO5EvPTFpxXQ7DL87PMuXr9WROs8nmxMbj+
08CBbbZ+kC1qa2D0n2x3JZVh1DMPEf/Itdr2fB+H0fFVTM7GNQqu9pr76DxoJId4
GF+Z6CdZb9r7xVxA4CWH9ROp+cmw+RAE+MyfDIxBK+fx08dymCijVmFATmoj5XIG
h35G99ei+c2I4y0IZ1Mb+9QsSxKMCA7hGU9hzpjma9tHMsXZanUm8FKGx8dAKnGH
JIvcqLFO5fR3a0qcE2esUzg6LKwco0rrXpdjgO5SQZlsN4V36HjnL8WhD+wGmbuz
mzSMS+Pg4JGMQNgtb8zos1lwG6sxbHG59+TinX67Vyx/KETtbvdo8MkQERI7untI
nR92xOwbr8o+Sann/8/DbPqUksi66cZ0clWzExW1WDd2ksszNF8eOBh4EGMB8yLu
dNjMsZltGI+q8oyjbJxXcYgG85F2tvBz+vS7IZujb5vcAwmLtK2rWSMvjunEQv2X
+bfNF3cwRVCIPMb/HUS0n5CZC7DguH+WnvyHkt6IQNjztJ9x5YDzTxC+jvSoRDUa
a8yQK3cck5Rmi2DH4HtT8tAbOR2utFajaaX/V0d02nWlAsmFMo2GnuCrBsssJBob
MyN2KcFh18foazNAjcOsnaWT8MnN/OInJpwxMXEUsmV2ZJtrrS95uMClMl2lj0b3
LXRNe+xUMsfxB94L+yeixa7frLngLhf5fhbd0adsCg995IckXTrkQtmfmwvk3pT3
vhWxj6NPGfr0QWANmrBu1auZM2zr4nU6ZyiGAw3T9WIn3qvZapXxROQudSmxE1KJ
2u+tugFpFnJQCIbrMJLPCgtk9WeutO5F67bw8DGXtf9ziAaHLSSeknp9Fs3FLZA8
PYPg2/dNXBzDaPrHFwxZj7ulkb7/kAWuDgV/LrmPZtuCuOGHN4haCcYXhaP4x17k
DSeFtFNlz0uu05ykSA1KlGyfgIO7hbRJdRaoy/hgumtjZivgiXlXWNWMwPsNqyl4
uMT1jaYM3dqE2djpzd8J/Dd0Xd/Wq/p/qjBd7mj7ddFbC5hAd3xucdoJqw9IhSl+
urhk3zXPL46OILqe7/hEUP9CzhH/ZjG6KHUQsxbIz/byAyJzVgGhfkR2hVx+hrU+
fKBRfQe8U9CSmJufm71V9f6Bo665AFr6TZmHZWT+bu4rn2RPWXjckXLqFHp9URfx
X8vUFMgVcj6p5C2ZEVOmvOnOzOyZAZgI3GyPrEIeAEwOOfY1HFIn+JCpl2fAvkzW
uNc4CNtNDCsXs4k8gEzzfw6its1ErI6b5pKGQYhlrJKSsjiPvZNbgt/gVZqjG95p
HVEe4YIobXctCaROxnE7jF6CuJvFbk8LKbsV2bDj56xkUvRc2RKTGpEzbLOi8wDr
gMNNq4FE5pQ/nFRwljWDLOW3X1uJeiflXxu2kESXusuGAT4o3TaaoqyXO9aw1x5l
YbqRDqLf8NIDN7wsvHTgLUuKrhMqg2UH9vN0ZNfNqujWJ4f59kon2SMTUW4UIRlU
8EoR+xT5XMQ6j4KtMa0wS1KJsnhpqSsUQJbyeQqMgsqZ1GLF43w0zPnPHjIGy1h5
2yDtDicQAnv5X/mPsZophfpIJP9lqDVfdoDGNQhF3q9t4D/sC0ndcBuvFHRfDwxU
oQNzzobiM9zmaluMkxB6IqzUfxwxoJ3uhJEXKCwle1lAhe2GUTnSXtTqzvHqLDkv
78+LKCr9u7pHwLiVq9sYIeMvydtaUkqVWwi0CYmmjupwrO6+6iYPxzoKPEmox+IE
hQDpfh5nwAolnSthgx34/dJYH3Fjf7OoqHf93NN9teXHg5Dz8cq1gXdUHQUy01fs
4VHxOOPITu9QAeFcgQzAu3SF+Qe72tpeUeV3tBpu2Z5ZnMmtNbGchKQby5eQadl6
2pd17bhQaziOdL0678v7LTKTiAPK1E1VS2qEg/gsAnLR5WfEgx5jeqmTh3ksjoAR
4awd/ytF9oXOgYzFUSi8h5G82ablWuQm/Ff9gpfqgWJcpSE2v1WrFr5eGIt3DQGd
aHEpFN8wF/XHjGUTZjH9/ueVbnX/1pl6uTgl08zPvW52gttcA8/b8tlEZHKeaIRt
k72ONayoU+JXVZyCTkGuFp0QudOC3LYiI9ci9O5Pf4vwA0DlAcZlf6h5zlD1waLg
kamayfmdkenGtYDErvpEGjKlLMqh/f6RkrwCCPrBQV/6vsjbl1UCorb4PafaC37l
QcFym5Aa9A4Qkmtztghw4ORxB1AXkJm6MJY5wJI8zHP3xzcU4AhVv8z8hC5H08uO
QyThhHIq/j58Fg+JhLRX8mnCsOulDQe6kxOFZkfPvhPL8Sh78D9W2d8DAEuLReeV
1ktY6MQChCxwZYh3iQyZ9p7g7yOxoeHF5kjUdPKEFyB3UhlCipFqvOT1dwdxZm8M
GsDEkFjbsmhA/6g6Vhf3LuyRVohNYEQnw/IqwAMRmMT2FqPJ99Un78TTjX/YuZYr
JK5P+SqkXZo5hj3s2Gxz/L+nCuVkKkDxjWJTytopLI+5sWJ5oe3AXg4TAQ0D7Kts
NE4S30QPY/KZhplUQ5DucK4/K/hgxvw78gxLz/XNW6FCqai4w8i+xiD4pX5Z1DQK
5qeLalTwo4cfCVJP8XE6QU3Ps1K91qoQ0sl4XrP8Zos9Sj8pkFVHkoD6CRCyc8qa
7LRUo/tYjLTHPIE3D5F7o/JQ06Rmb4hanhgl6EZF1dOu+srJo80QTRBG5H3YUftN
Mv63/MvWkhPKW8lHwb3VL5Xn8JZVQJ90jpY4hYeLo/obJLNGYMb1oZ9MbiOS7yHY
Pr9L/VjvWyPhpDa7NxCOmIWLvovUvpsXJANt/HNSF5Gr6ZasxC/912oj8mzEzO3h
JddKY8n1FR3H0Pke+sh19fgDBQ6B6LlQEP/6SQp5NpyEm0C7bulKXdujY7EqUYdA
qbXQiKuVP2GPIbX9IJhN4vIwBLVJKRBphrfVgmakw3w1XJxvxniuCFTwU9P3D6QP
l8FkgBr+uG+Qa/DaafzLaFbhCYxov4suhFgp8kjZOexK66QBvDcByAo/2EY4Swp0
lPX//uO2BiTQAEMGd/9BDQEnHX6+c3fSnfHngLufRzVIKcjR3vzvPvTQHN/N9I5V
1ZlkHvOnzXE2lynDdRGUD8smCiyNnMxeVYqmHE9A+bhrpgz+SiYlX3hwkRJh87pW
uhHrLySSiheGpM09ZtYSvitoOBvHMLdflj7abqmJO08H7z85byDdtJLHfTVlHJmc
wXcj76C56/Wc6ZAshOCsgZCjthBi2MGUS5/l+WyKXKjPVUnkCTtGioA9AqmGIaV9
ZM63qE85vacvWM+QNqVc8DMT1oViYp908eF4XUtpqsn27pLNkmdzK72CcBELPba/
B2TxyraIo1KOQqcMiDHfWHQW+ZuiSO1M/xbodEbr6odbb+2BFwcOfoWECL6tLVM4
DcOzQa3ABkD2TkyAbE9KxnPAHnp0Iakqkgc478To6mINFWyOwbdjtCDRarB932VN
GD0O40xi4k9CTHRa6lkEESxkq4LfVRuJUoGkA4roRiIBb2D3e0J5zI9Bx69vyCBO
h3WgL07LYoIhqHbderrnBFMckCqYuLlU+EUBXog10YWxuvJucCeszkmyyZX1KSlg
yTX40kStY1SmGKQvKyFZOSh8WLH9NVuiPMpIEV3A+FB96uhBZssFrAYDwQePDWnh
xoI0yNt7TXRhz2kUEgsMv7KCtSc8wRcgnW1hwIfPL8n2iuVZIyK02zWOLviRkPlP
t22Mi6mUHRpKYruKGGqixnvwC/gqfZtb/YVlaYJZxkNyKS3AGqBgDrofhvaEzIVb
tGPI5d8avhOl42sS6525N/KK3M5R0lODstPeYJCc+essgwBykITShEP/tyzFlnnP
RnH1j+AhZ36t9+6Bvm9q6qQCXabV3/uNxAaAp/t72n+uzXtMsMRymK3MocCIPtYk
1xSPv/h0qXSN87PgC9i0bplLP3/A8tDM1PgRMo4hs1Nf7dak39Mcq1jSxfZd82Pc
Mh4X34LtsjbR8zLfrHsfeB75dGJwj+Wu54Mof58lN8N/j/dn7DLj30NmS6CdnQKc
K3IZumwhNyp0Ib4J806N2xLr/YAWY/lfB+e5+E2BWqpIcrk0qq6bGcHJv7lyjBDE
DREZN6ko3bEeerVcWzYdXfXYYDp2mQSxKTIxgZ9Uv7BUehYUpIO219ev849m6ifb
pabvoDKB6gfcyGXpmcQULRpTAaw6gRnk2v2IuLKPAceDeJKSznGaORpB3nbp0vhN
A4dQBb6yJikibSdm1eUIU4zivEm/mERDOD5ghE6shhur8X27MAGrAn0rqesRL4lB
slIxduWX7wPe/B0RMmCcHCkZTdOkoGepY4aHAiKSSJGS5kgo5buIf8wWGZmABj/D
2iT6hdLeBAeC5zCRmNpDnC1IWLApnGjC0C92wqpc68p8znCipvW1qG+0CNCv0cNb
Qp04fbbLd4K80ZpaKFtPm7eTy/poiAVmfDwl/JFZi72ws6dhux08mOobHpU9aeZW
uzhxHyelTV66RHu3gyDfo+AubHOLDLwUf2zLcxeLq1eYwdOAJn4m57a9l4PcJaWN
jLiTWzA9j3K9dJy3xaJMMXWcXd0d36VsSUZs4UrMJCtF2c1V/n5sVTDT4gzRh86S
5Rwp7QHRudNmiN0JlENuay9F1Gyggp24gxn6bBqhqJiEA296GgkCF9vnTWZtYBYp
KXRUFNyHb6l+agBRU60ye+Z7hbvb1bJ0aRIQ5QAJ7PrO3+VhXUtIu3XL+OqHNLv9
JA/jVo0mZg3Qj181ZFOF+JueppxM89BrUSx6+wE8OoEOM8Nxz8BuUgfUStRTTaVu
ANSWm1yDR7A43/u0GbCmN1wChRNkyyIJzMrX47OdeOYZfrvWv3J9qKwPremgUv9H
eobWziLt+q8hWLZySp7n4ZHgol3R1uS95AO7NXqdSiamEsy7YgmmrYtluFDKDgnc
WdbC8sYbELGfsMb2bVdJfJ1ZjbnTvFABAzq2GOhlc5FgQjMjgTRzh2dZoPYUNkbF
9R07P8CUatSnJkSN+IN9J/svZIelD1hbM65wITaGqPvn6anDXZ05joGNtOtQtMFH
Sl/A0q/413HIR6gdKRo291GvRL53+9My0yzcocSQVceNtq4Bw6xZJ6HH505cFFNB
IbgYkhZq1Ts5lFxBhTAMZLRyW3nY0F9x0Dfrzp1fNy4zV6iRd3eqpa9PAmIrFq6a
OWBX/rOiDyfPqXGnenCY7HU5u2AKrS3CgAseNf+wd2c3gbfO4XtNoKE1l9d7iKV9
ylJdDlJ4r5Jl8qW/jRFacWGByQA5ToyAgLz3QjZU4I/2RE+s4zjJcS/gK/yK3KQO
2A0PkEJL5KXHdQisEFi5reeRhnes20nP/35tA1snOJgNaMvrkv/VhDf7dAAYDEzs
hf91fQXPTsp+/kMQDlsZlBD9HwcqJALgHcodd9OjTPPmT/WJnLSbQhlZk1G81dks
13ShVC0rIMlUxXVi0mqkmbqT/zNPaRzDF6yhPBV80/A8XJXJyEhf5gQPW81Oh/Rv
cUxzeTTuVd4SnxezWdP7bIRgOC/dDPq52NB2LUYp5Yxub7WR97dfX/2rPbq/wljS
IRXlTwt8qiaaxXff6hldaDeDaomWyWPuGRa/t/DCRdxSccVrIN+snjFHfjOMmov6
kPbyDSWEm6UOAiS60aaGHB4PlAtD5wMmooFOIMUNuGYfOnneRsLz8HffEVn3cLS6
I8pTWJx11CDpwYpbtrBKgi88BTCfh+Jtrgwep/jIX3PUL0oYmWhOIpwDKZ/MXo/P
yiffgPc1N2AWy8PcEvpdxsS3Uetf8SiXqSC9ndq1ZtvkGrvxg5k0wl0ZH7c987X/
Lg+wdGx2VwK7c1exZfX/1vLj6YnJxCt3QzaKuvEeFlO3S5m3gDRC6oodEfVpzuhc
Z9iqRRHhdnJShUCA4nLy2w+7e3uIED6bigXxrh1pabQSQqaefPYeDP3Bkkel7Rhp
zpl12CmmKhX1F4cGnVX+AsvGCMf5hqVFzbUBb7ic9T0K2mrrDdF9fvI6cCSOfFak
FghC+4Q9S5yRa8hq185DHCVHjM4Zs+GD6E7h6m6pQWHG2A1klxWtG/uHQA7GXt+Q
SuF3EXM2m5DpzF0/YEMi9uiZp1rWyJNs22hfONzHbrMOrDINzB2RPUGpjHa2SIFx
vqAHdJtn6KMwVk1C5iURvFeUylUsZeSG8jpM9DMhlAh5AOjLIGK8wbMFrHvPU+Rp
I4QRFp7zIqDbdx+zhALvPxbMWIw5FBSmAdcpPtiUWnLsaPwM9IyUx3nXxdtDZ21X
M3vXwFOXeIkG9uOrJdFIon4aK21kqb+ukDaPjU9BIGCtAL6vbQpZU49mmmrYhPbm
H8c2Af0w+jGKM2esazY3u/OPBRRlW2n+6R7U1rK7AlFGHGTN7psK6niTnEM5qfiR
/vLMN2LzJeZA1bAf6qSw+bQhYqtv7efNghkm4owM3+HTo6rog4rnDwF+2oAj6VA8
lZ+Ys5Mmlw6Uu/qc3J+I3MWHHLvhPeCKHLhn1rQjkaIWdMSh+Gjqtxzk5wvkTTFE
munq+0Yt38DgPFka4pkTohs0b8b4AHCoNWDRl2vWirksiJxTh4KDZFXlCXTCRS4b
QmlnMala9Ln/YaBr3L5cCRM4eus6bX//ilX2J6lX4E/UQNOZp8fQ4L0XUh5sIHUo
aVtrAJJK+FwWgJ5XE363/v+IBF5vymcvcXuxVSnNWqHa2TjItbP8rMlBKVDntfiw
/eGdiXpzdFWvPhffYPyttF2KZUYE1tx/Tciu6Sj3B00DxpOaqvO6YiUStvmMkiGj
FD2cS9rFKKO4K/1sCrKwZUY0Bn37hYs3EPcYJGxsauh1UuAPngnytXBUwh6wfwHd
BPeFaLKcPMZq/MJSIaEJ3jnWIVRuGO38ezHlMXKYIX4YiTIl/Q/1hf+MIAWGN2GI
3cmX1Awyv+T4RtKeccNOnhUsafUdMq0PYWbAwJXIbjASMkvQWKn8uzbtem90mgNt
vC5Gnk+S9/kQRB2JSaEIK4Ulkr0nMVKCEpF+g8e/s4hsSxm8Hn296Yi/JvRVh/M6
j1njwl0LwpCpHVv+/QhfFcLJXM+AnQfl8917IhV1A8CecYOgu9qWlEPcNXE3HcQu
EEqdPS98bgGV8zyaNVES6hHtszw701dQRG2sKozgG6w4iGgB53aU7bcwOGcSXq4B
tOQ8rLmBBUUU/gEWYPsewMGF46Dru9Ao0mJhkyYf7W765Xs82AwIYArQEOzS5flp
rSwomEFECQjN+abwSJFHDf+SYCP3uk7Izaro6Sl7PGm6LP7wLagRNxJ2+OCgdr4d
0jErnZhJncMWAYe0573+xKjmcw+3wHJnKTsO/Rbz0KSQDiqV8knKHlI8Wl2sLIoa
hq8EgPVy1rIkJ2g1UsGhvRc0w7HZfDXyQJaXfi4Itl8LR83KDdYYpgFS/lmEyfIb
EhzialcRRyyB6E/Nrpho3IiAc9Qg1fYULFtIW3WoBRujIocZnRT19Iy17OW/8lRw
0o0UfNEEqpt2n8GNp2h4hmXFDhSvQfNERykT3KTvdpLud8myW21YLHIV3na1ooMc
pjFxoabxxiQ4LmQ2fRQDwz8VkqV9HGR2CfBSb/8FLkNaMzm3uH1fXpgnedLiSqIT
JH8U/FCchl6rbakf08l8qCIQFOcP/kwnLgnrQk0+3TeRJne3A4qMtBDY9kanOt3c
tgJUySmhx9bLSa4yGwemHj2q6avgR0E+GdNj4LvPD6xN3ESNQ21qm7ohY5vDwEk1
6oA2ejPzibSXFpKnKqQ6sV4UT7UZJlKzJ5R8UE8t6b7akOSjTaD9G8de8SE7TCZ9
MP8AfJiMfwcwcqBbSyIK2EwrvIiCN8/2FZWn7UJlH6mWtuMsFVmU9HnnMMDMqpuN
bEa0Jx83mByxqdBEzU8hiJmeC3f0XLc9Vfs+9ctgqJX/8eqZ7jR9fh3zfzalfBZh
N+MKryVsgm6jAV2Vm28ijgb5fw+BKJhkEqq+aabfLU1x7WMF13Mb1WOwnnoZwnrF
RZHNo1RShO6s0CcgkTfAQ5y8FIqKtcdQaL9fduQBQA14QEe7zKbrUlzL8EhOnabn
UtmhTzRKrxgoF7ThCrsBAuUeVLUn3+ZknDroZER90DCiIbUAkLYk/9gB1PZ9dXtE
OJ37KbgNs4Org7Z0eNRyBrSmTA3/PlwXVRn6z7qSrU3bTgdiOHdx3SZNa67NT9BU
kcmlLWdF8MjPN65wuchqmQXT9MEtqhMQjUP6kEvmW7esnFoNK4YJ7B5f27hnUu/h
Uiw0QBzeq6wiDhiH01/uBOCr7oIBd5tT2L6g4lamonY27YcqZ1PxQfgTi+IWQzjd
wsIlCzyKMYCRIWOps4FCV1j0ur6N+OIY3nPeGH8vbqYFW548YQ7XCHwMUhpG1ia6
xq+3rSJ0h4uzdjhBxCtVUr5AckdnZsN7uJoHKlo7lVw2D1f0YwFxyP8sWii2/fZO
TEmVTCDCU/0KsHFAzJ5S1s3p08bypr6AWrQDcfz4IWweXwzF1ILWbFZsvNcxKal3
u29uL9pPA/doOjttjrx8UVk0tNw8aTndSvERmBJUDJrZ/X+rKNRFhwGOujHKbEjQ
OnZejsI5AKhiz8Q19Gd6OlHRGkmi+9ztlozQBImNuXFfJwZSuhkOTdg7NEB6P7ZS
OyNTf9xZhVWBF2TiFB542rCkSSFkLv22IfDyIrAeUf2JxnGl/VbByaSxXGZHnES/
OqYwyIaBA7zrPnkILqmoKWVTNjwYl2qgozy+XssUs4LZKd3hl6hfWcsA5OcBCbzc
zi5LIl8xuwmzKPiWio6nMtKzhvAFLahSigOGM4eqR375PTNfLWlXoWh12WudBRrO
e3DrjdvQgo6eWikT0w3MAnbYeZrYw/YhtaXizwUjx2ctBXqhT7QyOVaPePi44KVx
Ym0RTp6MIkIjcUlm64svCzjaGNAsVN1RjVMLStTRL0r60YpGPY8eURp2wYLHKnR5
a2m+cdEB9K1TRMdVs4EL3VJ5JECBe7wTq38PL5mYNrWKGMWoVVujJCmWH8ddReGV
9hbkV4nkWTG5AhsasNFLUNFgBA6gHiB97JJgIanj0iuIDz3a7MbtBON0HSjzsleP
ZaPXrJREZVp14hvCEf5YtbGINPgP1GHZYKFfYmMCatyLOvLrPPD8SNFEpnvSiCw/
77t8yrEWCMTF884G9mTPfZQP5GW6N2WDgcOp/ZLdFzybxKKocxRhNWZp/NnKQhcc
9g09LwIzPR/Jy93axIpbidaYiYGsCpcqKM+wtZvW9V6Ac1REdwu67GgNMNr38qr5
i6PeZnnB6ZTC+hQY5CfwCkViTOV5bJ8hTrnRPMXeHXtsRkoDmpA91VxTFqofpl/A
TX2BIqodwzFggxr2lqS5qiGUOXR5Smnt+kSkKjnCWilWM9ECRw482W7jf/o1UTBS
MSbu+d1t6IAgUdoJNEd1FZtyRNs2Um1idC0/d9K+DMUHO1AV3tiyzF1UBtKGpWZK
ovvSxVY2b8dXZTeJWhXryZkdsOmEE+jMBDzCAqaAj/9IMQ5KopuPXdJgeWU5EYgL
a8T04U6mJePA/k+ByNoa+dB2CoYTizZZAWIVksE3prgvNICzu2ECKpXcmIvEqpMQ
rAJRM8UzRORZUTWqo/jv1E82clD9kEg/GMazIxvTAsKnohO4vfz1gwQzqUujda4F
pbTQzBV6EqgnTSchIAC1Nii9ynIHUCFhu9ipcz9r8NcBb/SI44pE7cGCW03YEIS3
bOEoiew57LViD1ibnYyml0L/fS+44G4nRMaLENM8ncUc9wiosRKxcS8sq5nYPAzY
NiOfPOKPpZe4UO1622N6xf36ZgRhcNddsBgv1lUYTIiXYUYMkR3VMCisWz7pSlPz
y2e40hqJ+wN+c5Tpwli33YROH0s69hdZsUr+ZugcK/00+M5Kd5uXH3MyFBvzmftg
wCm4woToQ73SIOKfnKIs0Cu63Esj2yoItXukkSSptkgCJCAhW5O0XRLrfd/CW2v5
dkJQgB9aNPwtszD8EJm3MQqDEu2UvqlcwgOLFFZqw46SWx7Ma+25VchWGb/slKlJ
z6ZHSesehUqn2M+K8sxCDb69BKArenHKth57xkL4dCHz77fwaJlbmA/AiT48whRJ
jQ4q+gmge63eHIlfNEu4gfQdaNjiSDe90xmp2bEbMLUAVaNvFaj9fb9/dWL/tZ8j
jnUZCGR5PFkjzM6Gk6toKvsIvYCDxhMD4rjVo/ZfgNMzzMsYMEULbYkBpZ+6mp0U
iGZzcHnnSlpyUD8N9uIQCtidH5OuWkcgsmal18cNmnd96rpz8qqZJb+3ImOk7McO
lHlRxaXjFxjVUKGen3NTz3G0FbBHVqRaHC/P21M1avbhM+2mIkRpQfY6bqmYlriE
4ooySUJLuZCM1XV/npxo9sjU9hIx1Nsskbuop88RXWtlQcZJL7b1/CpukMkAhUsI
M98OSHGU9w4bg8++wtqk+cnIAYd9b0JIMqLq3UtqBnvUwRLAwaUOAGsYqD+alUN2
gTqBqm6t0Ue2y0BUxfIrMZ7AxO4inUuiqBQUVUFFKnH0us/H2YzhjIGnLPiYyyO5
jeghgkdhZCt36B7/5zfmrov9eTbzE+A/Ua6h6IZfjdMTloD32taghHE0Liws/TYZ
Rvk8ZuMW/98Ey5cTLcJ6/cq8+1IVU2Mh9Wy3bGWTk6u/tfJ34FC+XSGDsoCf7gPF
R2blc3I1jYAw/TMJZnPvUImCS0zpA6YNs3uSsBVnOaXn1tKTX335eXLVhtuJCFjM
Vqgdz6TEsyWGd1RTVn5NnLHEIuTqnh/KMTWv1FoU0/2sSl1EOoCwKTlZ4DYuc3m9
bnuU2u5M9+L1MqIwwoqLt5KC/HSlnYNbZmnzRZCx/cJ8wP5Zt7mUo6gPieT/J12u
/8C17UDaEegIj55nR53sSDmYB7qCaEr1WwhBGO6CmoJWUTWqn4v1Hx1dwiMc9utr
TkLfi2TQGaFIgO4r3UpBzgl8jKoo5p65EmrOQeNYix/78aSl06/cMNDqQMKlqQR2
VMNuNjT/VYtRmfXpnV7L/mpwWE1aA9fgPas1l1p4Neta47N5uiz0xVTr5e9p31Vh
Xob0LPuyDbVmOaFTkKsKazgWO+hryejT8KGnlD0tSjOq38afpP8+Rh3dyVD8a/9D
4ihd/U8wa7DjMuW7SuK1GDNbtmjxW1NhVmeIXT7dbhazPSVoW0ZZ/UNz2apmcuQE
GXUph8p3CXGlkNAtYKLhLemSSmBk5CJAOIcP5ophY+0VXxYAXwPKx1AU2twlLbre
3H2croxE9tMIzd7drNfw5bma+j3i1jrFKfXUuBrX3zWhV1Wnr/OdEoWZDi2GiFe8
8XB9uliRrIZvn2XHXiMQPYW9vuEHtvgrXtb9cIog26n43Nt875qY/MTj2MLvQsGH
OWIyfpPyIitHfXg+8epLLcwe3WAsWPdpMSa11Uu8d5vJyzXjVBgzgkzqt/xw4s/A
V95P5UhxAN5+RZ5EqhgSFY86jAEtBLwcz5JItaTG/P43LLo2LNf9Qy3FfNV1khiB
IQTZ6RBon0hY5Bj3Q/b6wdHT/glIsA8e+mM/MrKzyRNX2EOB4+ou1qDGAEMe9G/E
Fn/XqFiabBNIX8vZogUYxrn6W4G+9lLZXFFmCNw2hgG69ixELjrH3hnqKdL2BBkj
IPtbCTfbZtQMOnXCRS0wcTdOpKSs69AsWCAIVbzq73MGr6uCPJ9YmdP9MYuVy+WV
6UshAfleMng5zhHX8h17l06FtbVNlkPvC0Uy44e0FPWjHaMZy8UOa+0nk7O9IYNY
oCDwX3Hd3P4UbeAepE6N58/x3neCeR/PIMYFYntdBB/Wjc2vmSWo/oK7fMcW10Kn
oGuCqyiCOkLYdRbRFgdyeoWRacMZCHG3UOiEg2ZXhZp0T3POBOygVt802ZXpUCho
a7Qb+e/d41yU4RRvpqm0u7IKAmUe37L1+vnQBJYNWpTwHOLoKie+Im57qPDYNCXN
lHnAGUu5D3s/Mhrtj1VWI2HrHr7qp+tgM7cJC9VDjA+50wKRXwK67STlyIbYfGz4
q+gr25VIoSGw9qoCDg2pGpaoACfEXI9oV+u7vkv+0KpHm/ysonWKfUfXSUe72iQ4
PDhKgGAaA24xrQJvt0tqg9gDJ4Aby+RxIO5g0NHLySZJRxmcAwiZXTJQ0yShcjJR
G2llu+gF1uAGU6VkyRDI/qocMZ5hfclc2Y9pI7SmWl0KNddbIWt4jByeH2CxC73b
ryw1btPS6NukP85C/fOddHyhSTEWGlqgyMuvUo5ckNforeCM6TMxUAaNS7HjkvhG
yLUO7MOgjkC8G60zWk0AkA7gRJz3u9FGvx7/BzC/BlZwIS0crpbB9A+zZb5CKJEZ
cJ0kptOZTdxV5DOg9h3rIyI3jfDHmfqybX5WRjqC5KSFrnTdmVpt3MTYN2Hi1Md8
X2GgZju8KEK1C5bAvTMx3+AZn467oGc6iewVTsV70sJIXHLOjWOAfvcEaOYR+w0V
VAmZ5dr/0buZa3iD22Ehpf0gJFm4RLeX+aJ8OxIx2g2FebZX9dTL0PVG9cTzIKsY
bopXkI8agnboUWZn+TdLrQHgL6OWOKgqPGcFkkO9Oxg4j1SkigABwr6A1NaXZrJN
0j3ZTOsDFUVzXFcWhOK9tF3VnGbDmoWru7rQCA/r02nYQCEd1G56KI4J9p7581QH
/oAVdZCFPdHmqfxmOxbre1USe/3hmkmx4VRNli/jY6A9zULvfg8FQSwcOoTdk4/5
0jbhIfbAZaWFFQpLXnlFtPXq9d7FqtDPOGn8b8zWcQDXCu+YKXb0SkXQpVhP7WGt
NUzoEyU1r0OBiiKQsWCVq77DsTub9WN+rFbAYg+rCmPT0YnwvgVijiNHXO59OsUr
FzINXILPom7PYB80NbWwloxl844JNvl2xdd2hfEmyZhGhnZbt/pO6ubhR4FVB6Fs
E2rBj/gIDqZuSmT2wf69ogLNzfyl8sMM/1xaeWwuAznQjJGjy1ht2RdU1kHJuXfM
TVIk8zu5w42JTnny2kvdykxB33kysjPhU56hvdYBUjqEv+zNL6RWTKTg7LkQPDNr
SEzz/ogUIoZh0dG5KxKbGrM+2sQkyQsHbI1vmTn3PNQ/pe5hOaEfcPTPLf+qw62s
z4EVugnUq7Z/LHszrZjIsDCPAcF1xUgz3To4cp9QInHbrGBjGpfjew6bQVvzIqoG
UlBS7lwrh+V9Kx0UuqWSEmkZJZ9TgUldSSMUmX6/sbfQgXfUYxuv8SlUVd/+da6M
8G8ey77kM/Le3NO41rXTa3UjqKrA313rq+9bgqF+vjUwiAm1WPwPUOicXmGhed1e
fe6UF2OY+pvLPAlftInvehUP71HEVoPd2iB7Ces1lKgFepFhqTRHCzLHrpv13kjZ
5+E7MO+6nMQl6k7eJWw9L/mLX1/rOomU4/viqtxjJcBz6bZc3Tk/mJo4VoCLvfTd
pxPSM7jMhmf++kcAXzxUXrgjB3qUf4l9jiM3as9y2r+iacgzPZ8ZGgxONGaYgjN7
cpR8B5vPmhP+bg00SPyioqLIMZx8o8VMueFpdttDJB0eHM4mF4EntU4IMQBrRSdl
sreZNfg9OaQtAjqw0Dw9ejRHHG7QiZDAnTUSJo415BLkWm471XML7FYyaWz6Sn7I
ogqqzCxktZM4ClcCppxSCGujIR7LdpoOWBrTe11lAdioSIuEmeGCI1kV1NbPNFyI
i4JqBhN8FyLk6BzzUMZCfKlciARFjvC5BOYAjd6kdpaxEkFk06d2C4rN4KNnl6cV
irHk4kN8w625+gVkAjTSkSpWk9/fd7UrHubmIH7EuT3ln65VoTA0AJ/odsMq87gD
82Ch0Id8TbU2oq90cq7/7nL9XmBb5qWxtuPFiYgU7MTDTiur7ZvbvEevcTfMWwgK
2m41OzeNYKUKJNQsm8oxA8JIBO6rS8CbrFB/1GfbJTLuxl5iDTYrAdn1byjxsU+1
WvGwVT7NPaA6NKxFEi7iqqpXxsNlL0xKatOJaEO8+TrCh7pLpU3pLSzCOQuWWLjD
+VqKmoi0I+rbxv+EJDFi+0apn/oTAgIh6FyeVuPp+91YumbIS1oseEJaqfZpOVOl
of+9HObA1Td/pMLdToj3lxuF8zFQcBYW5fqjpiCBEH0QUpoU9tiRbH9in6e6SNBt
bkRwDpnSj3PvDnKEIRtMHmG8JeMdvE0sJl7ZTsePo/j4BVfTcAnQc7LEIlkOWbCx
tfr1iT5gSVTedPWllekUQoHkK36D0UBwEThYhQ7BqQlfTZWVJCGHEHO7Pg3QZ8oX
raN/MiU4YJkvMz3gCz4G2eoh6DAf0dlwmCEgequ0bcotFtgJ4yIwRBkXHvHlk6Tn
neic2Dk2I/v1Zeo6j3+H0XD52kwfgn6l/8c2R6ThmUyBtFF73USMl6qOIshUaDwd
7UrLPrv8TGzlPFo0W25hTLnwjedZbpB8z95Md7NRXTpFnzdQEs6rEL7baRikCgL+
QFIuf6b0JpImP5QzXsOCW82l157SOyjHOPvdH6dv6Lrd++a7owIVS6FE3QOAwGSz
s5udrHmQYVGBO90NwgTbBe/eqXFmAlh6zrt7AM5Tkfz7GeQVesJ7EibJLxqJXA+Z
n1Ic4G3V5g/9J4MQGgr9WIstZ73OuCLRW8uWgE3Ycu+R2foLQYpwHxhcHu+1OBum
kHuE6LU357rz+faiJczti8p59Sqf435EJKLIR3hD3LyMyUuEdr5c4a5utlaQltyS
e3SRKSXxf8xUM0VV7c2GI7vCdQoYiGWPwWY5XHrHVrJ2khKPZFUIolAmEDrVk6gs
z3B7TY4BnMUTU0yNpOAVNb+sd+Vz030OedidpbokfhU+7Sg7s/Chfs7iaUJuBx3n
h6+c98E/Co3LzUTiDK4BMiWw/neeBFNJlPK89DbaaIomQfW2qhSHi+86tI3DszpT
ATts9RvWK4a2G0CNdGuRgoLeuW5RFxGuB325pvUqWFiCREPjPUGnjfM4XS+vJmDF
JUUcav2x0wxxKCIWfLlSsRiYq01wbyKzN/2KhsQXhZstyXW1GXfi5kYrUnOVZKr4
wI74xItuYysTUY2M9TuLbvZtQTWI4sKQ0z4maDS81nQ+x6rr3DqBxt3m4oRto9XT
nAJ1Ciax+Si7VGVq0z5QNNfoMeKiU8bPhjq87GFRfor6IJkN2ebEe0JmWzQWebde
X7cm9Ggly+YRhN0jACWUhT83N/Sok7xGExTCyuyjKnm69HChSvzU62bbIMNH8SYP
umoQ3dSHjQJBAgKnHtiievDrhlraH1EOZgNmNHM/dONLYRLIKJC8OilOeH4+t21Q
m87Rn9OH6+KGFFnT+3sB4siPW6AKFDHYMNnC6NDZMR1LKTuIZc3duFx/4LIX5gJb
lIpxil84t+NCsxPFzzReWuMUjVCH8oWeKU69rcrwoRC5EInL54X/hf83TYYPI0u9
0z2dUX5OmicM/Owm4pzujLmxEjQmJ2ayWpI03dFxvxQbH2s980BdCneaYH+VXqkQ
Ac3R1xkf1Mcf373si/sHOiXix5nMSViJy9Xz33aUfVCRuVqV9+pXAthH15wagu4l
Z6KmkntB/ldlmy0Knz4T2+cEyJG6yzl9iN1DMErB6rvkBNsdY12X5g/T3fmCCM/1
tRSShzjgEBmNRkeA6BIYhOzme5WgCIgL6JjRmaBg0cVbnGuXFqrqmdtMtMFOboiJ
0OLwXYzASZpfPGqTs/0xWBuFirguA3k+VUZpjJalRLdcqo7Swt/ISA/XtY5DZVTv
D3pk54xtCCFucuNjyF+S8ijLhsMuBid11T9cOua1aa87TUzmzH3DdBIUJavFdy6D
w5Mtx1z28yMb4HapeJLv/DBxthfFKTJo1GVwhXNSGSbzzVdKNOHfoqZk4DbAJBHz
10n5mXQiZ89/tts3y6h6gIVO7b2PtSmmnjl3j1WR6ufHLr1J3F75N+GZcRccVko1
zL+JvbyRQHrewQCeSMk/7xw7T3nibwRKgJw63WRbCCgNK5JBlkc5nVaPHztk2SP+
B+WVSEG1pKDCYyOB/xStcpXFvNnz/xpVaTS5NkpU7qkxyXURqz+YgsdZjbfF/Rz3
ZUx3CVcnUjfIn7LC56tPrKIJDVddjL6OPzvQcoiu+cMJD7S13tG2/ul6AJQkTc9b
AJ/TUkIQ+yqibF+hl5vCSJXsEV2xgALuv1BJPA699LZF+XNW13fo0XC7JGRtZvRE
QtTvLqNl9zH3YqDU068ibGm+4GS4r75PBeivYTLYybv3DfFofZxyF5RjkWjRb1s4
pmFzs4kVcl1nYJOlO5ppZHmn1+AUHLcqmpL32fLdsG4kwdixvW4uRYNnnkrIN8aF
TfRzWyUihiCWSKnGf8WIdw9dKGkzka9zIPYHNKsRljqDtOqewEndc2Gl4V0GWm77
3OQ1dcRDRNvgaY6vjs4O6rXiGfZs3KgzHIHKxsbUf7IQ+zlFv44eQbH/forCkXeZ
sfz/dmx9G6kIFagAZ/xk0AbHHJ5VE5mcxCxLoiNN1ZBQy9jy4gemQB71D6tJ0oqw
DaYmhgzm3Lj08URq18xfDiR0c1PngWqpJlR19vhQHjd1kbpB8gPyzpEOaguYf/Cr
os7uG++4vTkY/gghvAYmMq3SKkd4yHJKZoL+TlTNPOErkJHaq36ZJ3RVje7CPR/8
9+pYGa5dK1BsH5TClex63VqWc8UZestaQmDIPyPFX+z49uadFo5kpOYDZ6KP0PUm
qwrfQuaC8tV6S053hqhATgXzI5f3Ctly1HL3HR6aw0NLZEcT/iGAX41kDFh1UXsA
5SLt113puZ1DP+BNk0ZVOKw/LYvqDhSn/Bs9K6bWsyauB9ElNM5kD6PtPu/0l/fK
IHfUDSmUX4FAbd0L8wm8oi+Lm9xLZ+zgaTVeWblC9fSABR3hDTQC4cz7JqxwDsqs
IlUUneGniN/nrDhcIv7//9N/Ta99FVndowhsWrum1M/GDe9uRhiEdYrmuvFdIulh
vaw40HV2Zyz99KVIhQjNArPZk3xzEdrK+6Gkq6Jec0wNSeKQXroAEKPHMlmHhuUy
1u2cfeteAWEK4C0chjn50lC6R6SIbt1KuC+vZ7wKyyR/dm9YCoMHyCqdBDkYGOVE
gkP+y7jbfKQv8vImgAJHUPpFWqKhTVcxVqm8BeZlaAHTvyroGZONsTiuES0nO5TD
j39I3YsJTsLs/SgZ+3B/Zdsp69kafg6ndajxhrG8INz0CvGLWEaqNzUZ7SgKfKHV
8H/LTnHxWSW+R61zpVgdl5z5/v9TqR9KBYxUwALODXYEYPN215MySqwvfu/OZ5y8
EPEgWrD0V2keXP1tTSUWLd9hKrGdyB+fdnT0veZAldcJGbY59uxZHsYeEY9+AwmX
vPGQAc2KXXaPKNvx9kUnOdAVNFgtMjncJNWfoZh5mxqU+cDJSHWkOmEG4LcQefud
D+nB3A/5t/V2dSyruEobPWoS19G3xIFW2q6BCscR1XeRTnRrvF2RWV5fq7slzRio
kHkzgngoVqF6hPiCaPpfUVuehbcypjGxWQBI2GmMhYbkHcMkTRK52WgDEA0Vpa/2
6Zwsxoh0g0zfZRD1+V6F+TtNRReaSRdGTHe6PVBxOoAohCLxLCtxX1YpE8uTeb9O
kp6+RQ6Q+O0K372orFFGDlsYqp8eQEiZStftWxrK3nFpicjkEBI/D4EF8QwKijR1
PdPB0wry3Rd9ClbNTfwBAAQlLEQ3NXtHiCg7mdj9gFX+uSbS3adqXBfIXm5uk88/
+rJZt/Tg61OF3aGVbisFUEQbloWubW1W2hqEKxaAN82wG1P2IVmD6P5h7XFkdPev
TG5+yyeR6AcZWCsJIeC9S3Nyx1oGymmNL6afUUukaiVqeG9civ3ReZWls2P19U1V
teCg+3djQnpHyc9VroP2+HvyFKED1lv4a/zSluMoz15SlXs2d5hDz69T1GZSzuzJ
WxHl0ObENBSyOGkvIEwaUQpePjSE66y/SgaVyQSgGaQLa4kt1eiobYywNG2qjWoa
67L4EPnJKL5usrU3MJvdihR/FjqHSTapwYEEf2vuu8PqppvrVF50yGFWFGsBSDIq
6QONTujpo0Ooo2PPO2D5Pfe5zCo4cUmA+LzbpPr9I1dREywjUpHe2sEEWJCVM75Z
d+tKKB9Sjg8NRfDt1msfL3Tt6TXNamTiQOY3bK2bsIvW8stNvgGRSVAy3TCcmiH4
7iX43GMw0cDdP4yE3Bwe3AF6JvQJiTi63cyPGYiXF0AiPO68hSOIHzL8oDLJ0Egd
JxEvLs3xMSAO7S8wchPZhm0nlUiyDo7LHoDYUit2pPGZmX/jf0WBj7hoUYMBoyHZ
2MJuJSdPn11GewLC7h30aD0w/equeiI8oiUmXPGUVpU5KWuXBQHIgBPAzgjeQ/kE
1UkxMMr0eifL0O2Iia/3uxz3ZRTU/yGgnhDmABpmcWKyphs/rm3vjsdBPVMPTe24
sqQq45OwgNFdtysHdee00oOB4TOHIqsU5JAPp/LSZXULZ6d0vaQGunvWzBop89Ij
2ds0H6rM/9coE8SevLOR0RVMOCNm4zck27Lp360NKxKk+Bx5RAnyNq55rr6vQ+/3
4IZMacIPVwI2wDQJWTm/T2IeKFNdXpcWCJfnAd9fbcaemV7GHu6cU7u+WNLHp8XQ
VJgo5w9KS57k3VEr20DOYNA6o2kYltdMLlQ95wLy3chG49O6wAu08fGjllLsy9ja
jGPAWc6WrOs9fKuwu7iFH/Niu+Xn3tgBq1xJlmhwz2fJuTPUSmjjitZxgn8zUMxq
XMOQIZbq66sVdadBo/Z8l8maosPU4h6z8mDeif8Dqa1iQv69ZY+2bSGXR8jSULwa
OtKeiexCjsv+GoTPHRFrd7B/3b03UmGo2ehoXpiu/ZZgcgI2uS6VK04qQvbMcAFi
v15mGqE9z0iKKSZTkRMSDHZ24Dm2X216KCV5Ia6eHYKSib2TCbUSGy9yObURoRp1
Iqy4UlnlG1AUxYmoFi96ZJOzmcpER1Hd2if/tnrr+ZxTRhtVqaJtVPyNFwbUERuI
weyXcQqMsyPGVWteYovXuJrfrMnSVWXYnM9z2mXZSR8A1Clc9fXpf6Ts5hxdr/rG
uCi30Q/s1gbL13O4Xf4V2qlUAK3EnGCp/4VqnOxd6gnNHgPwjYk0LQ21PdlPW3Bb
M6jHjspXotfQFHyqu2I8knOVGnT49rtJPXXp9i3W5il+nMVGlclMwnpiUR0p72I5
zSwMBEN6T85/VXVzMHSICih1AhDvIaM1y5QS5NfpPGu63DrmhUckI8JmoowzKbwc
ETAx525EExfIA2MdHe0Z4CeVvgzm7dHFNdKEkMjSBAsNX+R2fiycgj02y6qthqVG
chv3o3R8iJuOM1vo92YI7RVK/I+PFZHGf6c2Mcsnii8aL7Tq0chkX8RWkMklszvW
WWda7ze2FQ+44Xk31i4M+JkEDIsLyMIkUpFUy6RTmODPSl6MtCrZAr9xQ5b/yJg5
p7ithJwh8eFM4y1stCKhx04ueuQBuHu7TQUf+vFG9siq0pf9XvavSEOwxRdFGQeY
jr3f1vLe2sxUvnxVRxarBnr32TpO+6kQBycEBGBUjoH7IKxK8lXdatc1XRXBTbR5
CpxY/tzU+Ydq4ssP2EVBSe1ckSVQVZhiLT4Y4IWsyq++Cfb23NfQm+oRmzCI9vUh
D0Rht00qo7hBFgmBUH6LBSb9Le09k3qe1wpz6kKkuE9JgwrKF3FrVpszCNNqgHNT
2DMNElJmR0qQES3SQiMnGZpK82Kzp/eRUldxFxcA1qKCDqbPiwfoamZHG/s7KEuS
HcfljTmPH9NVWbm3zvZpA2dHb2Rj91WTbswNGClm03LoXrRb8IqC5USiAydiY4Eq
IIM74S9EXCG7zeKpn9myAbvvBG5n6Sw9/r+rGrxfzGOL+ljgfTupWA3BjlGp693X
0catMQqvi5BdfH+wKjV9S6UdR2dtFPl2HxTqCYaIK7rzSKEdBMrlGZ0wldiAe4/O
U9qHd7HhLth206rXSxW9Niw9dMEKlOqByHGV4wf4bXOGvmqelvjnlmgYDZWAfopp
bg7zdMeB/esAZZVZIoFAYpISPLT0JPqeQ6bdCy+47R9mWKzA1TSgAswRxTxSB9Tp
dK4GbtFOBSpxYnG9dQ2TM8YuoKZisXv+/TcLOSxoTuAKR+T3MrUe4lYNt3bUjwAe
+2KEabKgl32gd/B/XNrXMvfJpC3fESdtfIWgMzoCI4ultc/04jwrAK5yZ1bcK+1b
hpGVzrjLIzg8guLL1rn31PqPyYO01PCYOodUbiT5nH8tnxJsd99u298dempmkNg9
k2Wk/7/xR/9LbgsxzQLSUc+BBxP7G5ZpqbsCLGhAjcl2kul3AGTJZSrYtyUEIMiu
tIY/DuFMsDs8Ev1zzbnMt0O+a2oT485RHjzTM9t0K+QCjgXQD6wq3Flxznhlgq3i
5qc2KEBPvS0sWfR9G6SGEu17ibBp9RdKqUGQQXepCy2TYzzIpJQFKGbOn8mbeThL
an0HsOotJIdK+jcKXA/CkfGk4qtQOdrePuO/mmFRplGBRRWqkEcEM6KErlqOJN78
X7MLrv9tJH8113HH81M+cCjUdjq+0zlA7sW3g9/Oy8KJe9nPOfT9U5NcFoHt127w
8aFQOI1gofCCdrdXg1I1WwKo+iyEVdYLNldaenF37A1/fJqYgu8KnfNy06f5IJtY
MkoTqSJuRmiqByaDDh+jPraKiigMVmZ6Xw84vrR0YplzHoZvv6q6AB56ODKdAs3S
qkmhnTP4+nLl7yvCSHEbJgv2jhV3OoSppUWyc0WcOYl0QmXJZgmIqluVK+A3ykTh
HXDMmczF06TVm+e3g4WTPjJikkRwJydU4xRawUpmJTKq0sQwK7WazGlRWTdaaG8d
a5ZqNA3fgIl0eLrW2Cp85cPsU2sMZuAMllwsKfYDg2NEkK2WNT/QA/IWoNnYyr/7
DqLkalo77I3AsiT6vzb5R4abMGN3kzTYiFbp1bJMphZAZmO8i6g5kBy3MkO0i0q9
tsJIzS38IMRU6QX2/oU0JrvK579D89nPAxk6uJ7cTbYN1xErwSSTw//2R+flZZng
RBrdkkA4Wga5CyH1McNa7mtJWpb8CwraEh49mxS2Rdvr0h9aoHpvXl8cODpN1hfG
c7fNDT0tDnXsWEPqPAbKrzXGK5T2V4AEo0qgyTPkASmdGrYOc+8ykjx/wV1qeF3s
jgJ4Tji8NqLj4gXaXhmD4qTM60EJ2NBBoFq+Km32J+2EH6BRoC4uFn5NxJqU/Ozy
I0mpRKr7Mz2wdmA27nYVlZUyH4NeMhBUiBCKNkSwdMidEFMtI9Rc87pNF4xtJPzj
Y6TT50wi6Drsitn5HT2BDHOoHPT4E2okME1EshVPPbMru9dnLeNQ7ijZoWczlUPD
BR7rn2oMY+ovcJ4RcKYFrjamJdHyC8/CllNXlhYATqFIyoAaWSePGMh9ra7LBqvD
HILYHs+nHGOYc1MW177WQHzT+K/9QH2QcXxsquq1WuuM8zDnonocuzSUwJl8A6DL
UAFhwXwoxqAa+4tlxd6TbmtMN8ty0vFkSYaniNDM/B1FKTE07iPge2pgNWXz5A2c
uEpwmo1GUBis8ENWq6rMCLMuPQ+2HEo9dWjnaJFXa8g9jBkeMTONDtxT4n0Zo6Jw
/q2Rqhx964bJQtQE7dINCiJS+rBJ3tw5b90rYu/nju9vBFGTYsuN0YaQJYO5UDyO
8WTVeBBn45k0qMXkOte3mn71/LVaAN1E5xOWHqBaGIC3+ycORtJrVEuZOt2qbFaN
oFXeFhzxVfQ79YL4lZSgGq0k8AVm5vH8vn1VspOO85a/KpzCsh+Juhf9CGkeoOZP
zDIgOHL9ziYds1fwsN/o8TczFjbHE9ITzvWNI0KZZTOHFFj0a/CDCn1WsYaBRrRH
IrScO2OeOpqyErrQXdU2ELWv18UQn3eLkH0cZUXmBJntrdJd0XFgg9kfclmUyspX
l8aYo05A3FxvojTyvx5/DwSzyPLHDu5mdZ3oE7gTOYFKS9FerDSMn1lSgBVk3O+r
9pOdGl2o3eEKuX1J/GEcixV88K4G7+Ua+BPcbLcpdVAioERBKpfVBjc44kIFIAzG
+QU5bT0Ae1pj/jLpbuQWhhDRb3/MDrnD1jVd06IQhw/9KZ7Hcd/Eec/EKWMBm+vC
HkFftXAaqNAnEyWAxsaAPkviOSxvKJJsG1s1a3NFylEi9U3jrgfm+SKldZB0Vp7Q
4UdOCrK2IAna1T/3enosogP+YO0KnPl0LCotQ5mUZ9gWZ9waB1S+bHgd7OQDm29R
SQgx8AkXV1YHYMltamtTEpbGmxmKgUcR9HqAN3xMys0Q5B3Bly5lsFzat9PjO2A/
6G+/Ums6iCEnq2H7XzDzJdX520TbsO5rQe3MzQbKuDiVDU80G2pNPZyJWaEWr+bX
hRgJUSI/TQbaChdBuQYZWSRx7pom804z0RZ1Ei0i73AQYPe9KO8pVnGgbWnx7Hdz
t7CCwF4ZoCDgIelsNUDdLTWiFoHwDFKoRCb35FAegXl18QuTOGC7OG5xlHJYGs8r
SR65VxLPwFx1Gm7qxWifdI7VBY//GhOOcg6ipqZyw5TqSfC7lAXZmuUWjOOMsB0M
7SHjird15W+irD4fji58nw9SRlH71kudNBRhQOcz+frJP6yLAXoufVor6dvIf28W
+ZOKOumTyqsimFBmlW5hpBrnsxRXwBglmwxU93Okoh+aWYClHloWis/HEzKpXZ2c
wM3EYFB2lvzEDBU5A5X9ZXJrKezxk6p6WLKLW2oCmYhu8vGNSSy8VTrUlRngFpBJ
FMvDRTxLtRkI/lIT9e+4T80LqqIzXUiG/2l1nsJC9xQVn4ftF6dsKgcinDpVj0qs
Aqvmvd3bP30fcWw5nBfjmI52DXLDKzdYG10Ms51BNQ7AvULT0J7jixQdBRBJsBob
B7vQI/lzuPf7xKpDtr4841cSb2/CNbdvHpSdHN4EHhKXmGQ9UG+o6SZAwTvP4BGF
Nmp0P2fjtP2BiMAZDxeW1b7UG76FcPezxJJx6BWAb+U4zpZtEdQYV3JBfmKM6G+Z
Bax+yQRet42374oiwqNyvSfIWLq3k1OQ/9JJwBQ0iotL5dDRu7OOiouLbQwz8c5q
MaszdyJdNmWlJkgEABoyORJ7xuCqynPFeSlWSZk+hR6E7o2yfI+2N5759P705JBG
o5Lgx7vp8NIrEBHZ7s0DIrSMA/prXoMzb45wpEYHVMShy95BWoQITzZmUvzBjLkD
/h/4iFstUrFWgf45Vdt8zaNrKJJxyP1UrnlHkiVbq4OPXRrGzCGkDvPnWVhq489O
TNbxtpqnVORRBW8KuD4FNZNAb3CmYNIu9XNOsFx7CFvhk+H9HfNg+74KCS1/BuYV
hC1l4i5BllUyQolw0c/2FZeLcpTCporKUhdfQVGhFI48ui32VSji+xeZNi1P+i+J
+UmPtSFkkKkiMMu2Zyl1Ms/gQ9ja46xtYmwN62KtR7P/0OZdgF456WYKY9Vp0H6D
yrKY4HA26loZqkzxF8u5lbjsxA0QZiU1ZrgQWu8C1Xkgu3SvFt2lhjYOziM4rfDK
sPekix5oJnACjco2dDMSf9chMvPPsXZC5W4xqMs74zDKRKGZHQkNuyZQbEf+g9uO
TyYI/nXCzbLKtNQ6993HvoSHZrFpNPSSEdK3kiQRmfldS3qM46JowM+ikjtkT2yO
g7lErUqPuqj7IJh8+07843hlGz7ur4xlHy+PAMHrldRR80Il34tq/RG+YjbDFWoW
m2Tw1OjGWRJLwtzBSHBAAlt5KdLjse1iXjKWCe+/zAQJuyaOwRyRFCIdYW5HS1J6
oGIsdOnaBwNsHVY8wM/x2atu5n35BIlXumD2BN80OL50y8B3Vq8BTFKRwRfSyLjp
CDswHO+gulzq4YKPvjZxUdL1r9b7cKC70J3NPPG2Z9RQFulsNrFxhmAa4Pwp7TSP
jkOA2SsG6gITckrIvHXlFUle1eEOUE4w+Yvqej5sRwdtgF1QpwePoauMPcZp9mq8
JVhfxtldYrh1tqh6fossOIEfKffy170lFcsxLydozeCLBO+FAWR+I7IVw+asLSGD
k0GIxyA1B3Jr7Xur6nxi5D+T1Rkm17vOVhE3L4O86InP6DmN7UtMm68UJ3HAd102
DBv+84WqNJ9i3NwtMjF6NRgYPN3pr0/D+kFO6XKZvDUr4Nc7MCeGVEiiw4qmARUI
GaSs9NYjAE5epJ8nsGhEe6mhYcu6qRC68kcwgz7GlmgqYuYjnh37VkhQuIvoJit3
zWVWMOYjDKE01dppuO6MmiLr5dfGJgUhSH0mbHZtxIGQLV82iIzjqjQ+GdCYrmwf
PoheCVZ32Do3kbWzuGbF3N3wUCXTi5qUAF4QDXYe2FUmUcoc3f96tCNTYg8W6pHn
6jZRw3aCk+3UaYjl3+OjDbq2mrDeB/1Fcc/TWOIfoljU1WVXPXnJB+Y9DGRUKJFs
haIBMV4SSEJnztXGo99pmV4fCeCysGVn8ilreGtjMyQ4OH5nOLH1uHERGUD9tckX
LGYUJzAsZOTfU9RRztQSwZzv2gcGyqPBKcJx1B5nqc0R8mwG2zzK7WV7rSHaihO8
qlZFNlPzIkpu2nKaPKeshS6gczL6YUTZu4y4u1+J7hMG50DKrBfGz+tY8+pD3Zl6
S13qVCtyFYDRtW4WhRv1i4UuuetSKz8q1Y5V/sW1qAWPUKayO4g38rfNgLmfKNWZ
CMNPLqAkybK4+Ta6T6CMJwopvsWv8CrXGE9nNIs5AckahG8igqsjjr0Y+daONLQk
d4S28SJnH9YNHmTOs7hx9xLc71nfsngzV7/Em8MDpvwF/cpB1RyoUZ02pUnliMdm
IzsgQYTgJt7kt5psgSqgFaPnOe7cGFJ0dBSGtPGpW3PumWpHvmBaEITgMjPs6COQ
RwZQU1SZ85x/ebAG1TFRKt/hIRGJoP/KysV0DngRRJboO8TmQ2uZI9BzUcY7aQhW
iHPJDu7t8Ku8uX/KnKCnSE8ibNHNBZEtb1j6xHZciHkH9/Pa1/a+Ar8DNF6G3VXu
HVKEPpnmwmNyIMEF62UK1k9ZbvzI2Doz4QGYpwfwWZUhzyx9Ej7NDdcUpZYmoR0H
J+HssCesFKjzZssmFUH6oYcswFQ4HXKKRDHRRTiYF2ynnl3tXsAW01J5iZkPxtu7
kVBhlCj8OaHrca86JbGH2+NvYhtcogfuifbCWLJqClNLPPym63PYztG4vKR67Gui
plCorzth1KTJTkwc2Xnp3IBLp1gyWI+ysGOgpa6d9CkIqbaJ0tlPTKJHQbOxaI4Y
GVbYpQohieBy6MNE4psXYCcdOaGb8/sdNmwLcU44RfgBJLp9puMeCesK77Jj6T7t
rDlP2x1IxdQVGTHANMOdtCtZiRgBKDvVLDSdhxirpoe8zzIzCR75A2qL2Nvc46rA
sr6CRn/r7orCgTyMXM/mozzbDLie9s0ew+u8CNDa0/vqG7gVaYn3d2jGkqCqJ9cS
OnH+cFzcP5Wsg3qdRHcNRcV8yJwWURHlTIijunm05b0MR+bOqu4Js8DDQOlN2Tsj
W+1esrxxLnBBFmxIReziF5pYz3LNDyQyftkqED896uhBBzrIQKOAg03Vn3X4zyM0
TRStitYwbNkNUxxIvhQ+M7zk9O+Tz8w9pH4t1xzlR1yeckLLHYE/vSuEtSdXiOVs
Z7KT5FE3fc9gZor7yDpxt89g2RSRxSH+IVM6w7g/YPv4PVLBonncA8UBlLziRyVr
cW5nlZyfMxbRUezP3JEvAYrdK0i+EplbvZeQ7+apyXRFZLheSzm7I8TCp7S19tsN
sNkLmWN5BYP8MEcNW/a+8b29lmbxOfSrxQkpx92137HAx3fgbbon3yhYCSJh6Lwa
6a9/Xnz3O3Bna9q3+UOH3JBC5clRCVxxxnUhL3v0uxynrp1Z38nzQW6fJguxMwvH
pDFv2S4L/uueaB0HpqJnlc/VtimprBtriD06LdlrrH0zSqdTCGYJWbfx4U7ehXcz
1BrbHilPCFNxJ2GOXIbd6nQtKDtYL136zV19zMHEiyJ4hEcB3AN4pVSEDInO2Y+r
RcFIjey4lj8mtfb3CE577xBzQcHT2BwZFkyBVdGWbuMMYwqniV/cdeDo9ZQfjjUg
jcWss/Ie66reSW+MLHhL1rlX1UqTSlXMbnu6Jcww81SGvF17/SjPuUxQpE3ZksIX
1FxKK4NamCnPvcibt/v2fA9P3RnzVaPb4P4IoLx4wOOzt8YLbgzR8sm9TLYDkwrK
kxLLIob945k3xoyMQn/k8fnOKPt0me3Z/j7x+RCgXVYAdRzS8HDTRI6IDZbWxYvm
xOsqoSakv38FdYkx0a409Fc85nbVJPbQwSedKMb31EeRocotBf8+uO4z2vokYDs7
fNyoi/C0CrCnyZmyT8lFRsL4jKLjTmEWcmfOgtHWUjtigu6FlHOity38yIexDDdZ
n18zsnkv+Gl8Nj2UOIxYn0hsix9mUDiBtIy0jyXe/1PwuYE/vTBNxtLYaJslYfP6
bFO1+nTocvVEkqqK7wxRHjZZNJVIqVVX0kP7+eEDYXFx2mMjwk+45yUQMd280IP6
KQyMTFDVCn6SxTD0OkU5gtQd580Qb2fLphD46HQ0XS74y5j2Oe9UgCE65JEdmEMr
Py+jA3ruidJxMGPRSFMre8AXbeLLBIWfCG7aqOMj+WUHcAurUZWhLSMLXN/pyOuj
PfHaZ76XOmPmSKD/AAbCJkYFvgOHzXlL8bFEax0G/ggZ2aGE8Oz3FqJQ1yk2Y79T
oZXI+CC5GTtjpxXKRAMha8T9LQZ9efFUr1dXH6ZpOUoB3FLRhG6sh5DWrYJcx1MS
5rv2NdrCKKP+yWEV5nG3W9Xd9p9MI2GNWohpjinQF+x2LQ0cD6RL77FkkuPEyi93
2K+7nqY6A7GdjFBKfHiJFwSKxPju1Vh3Xf9F2VY9Is5axaOd2U/Q+OEg6f86PHHU
nLl02La71yUlbEGdaSYS7mEJJ3S7vJUAvH6hlQ1KfG54eNCQKnwJvQnRTT0cZK55
+UK8wbvtnCJTRmFLi6LBOCvaM3mydDL9awJANjNYhcaDUHkLgdpHYXZlEA6Yllxf
QYDNuXgIN8r3Cxo9t9ZEb7sdcxOBpwp5x7TzOLmkeDskGWfSCL0E6ksB7XBqss7P
p/2qf1uL2bzpPbkqj4cJ+GWpugYFM0BdrYyRbUplxx3Kq4USHWpoBobEvGHvCano
kGt8Auo4sWJ9tkD4FmcUFpdYsqA3pKY0eaq+moxBjo9raCVKrgO3A9twWCtDDf3B
Mii9APq35x6FdNswVsNzOInNYAgw3vkg/cSt5aVkVvHLjbcip3Ep/RJBTScDzkKY
S5GUWndUrwtkAx7nA8VfxPIAfGxoHhba5IRbCPcpq5pzjIRA68rQiLq1LuNpT4dK
qppEfgy+dZkvWl1z6RgsDRtyO8oKatS1GcXQMghvrHJNUmv1U4hEHTexXyryHEza
LtiqdtUknlAaNoLIQ/SodCM9CDlNXmuk+oXFahBniKWL/6VgHsmWAUG0bo2HPyes
rW3PCIne+QdSGuNV8rq2eUIrrxbhGsIKqSyctQV7CcC0CwnSRBhB3eozJE3eEOYW
RgHDUL5s8Si8IaWtvVBzcxlX30C60n83dwtFP1yHuQBWxHPfFNXu6p64msPJQqLp
SKrVeY1aIUV1PBNE29taYSaGxEZCDY629Q0b9dV80zHAjOAq1s8IuDqKwIizXeMD
e+tJBlHhiXCQBGI8w0159a8mAY/osJIT7hyPVXDiYwwglmSNB45QKnKoUSOO3RHC
9AnZmaRf5bN0vQ2LNrbGoBn5xe0N0HEHh9KgTgdfFMAwrfDGSdoYpOPWgqg/yeBe
zWeEE7jHhSyIbBD4qQz7MdG59hJJQDHCfoTr8QT8jIa36zDhCGXZbhoC1psH2Cj+
Vl6BJc45pQ4oyZF9ebDj5wClxBiAWEqF/Klq2blBysgH18is1N7Qab2qpmZfoVYm
Ce+oWleOO077y2cBXEi/PUcI5z1rjyabpAnn3+5eqmKc44z9W3nR5AGPJFkZx9bZ
TfjL51teNT2vNfKs1GEyT4baLvRZUfhOEgIiFZFowNO3BjVTE6nHk3/9F0QvvekC
ZufNCLsVuqfiLdDSJJ//0FXUQQpOLXeO9IDpuCO2ZDDKps0XrSk8r92ZhtADGbzq
42vV0OHzybB/SFveJewC7fn8a98x+p7m8mm4ZqXCEYondiE0/Ww9CzrU/KLS63Ka
JH9U0FO+lerAra0x/8dNtdqr90XxsPXE5NKA10UD0Ipipj90hA05hx1t/01fbH/7
PeA5WZ+srQXMQHkFT+SIJfI6DVdg0k+8vnnYvQv5VCVEK8XFuACXoHicS4YCsRHM
McMyGTd3XPXILyE7Sn9USMIvRZkMewnoXEby7/0DodrQbLCsTDemEZc1TX2GvHWi
PdV7GTK85KgDZaLbe723KK4DDfiYz/QPPFwPfoXlcouRzGMBEPYH857ZRsbjM7CT
NeAD5qxyctWLNAjNfRJS7kkFyOlbuUWalG7c/7+ip5YgxalfwNWsFLIbyQ2i49D4
Q8kHvjmp7qmkJTkfaIXQmOrE0wdZV0FjXFEJmCdGbA4VctLmM97hhsL1FzncDWC2
pnO3ux2Roe0a/k+sF62J6MouOgSBJtA9NAU4fGKQC2tQmZPAOpMQUhhy7gZSS9Bh
thUCrXgUXaeUGtoZDT4oWG3AD4bYSIVIk41FOACWDA0r0eqo0dD41TeM3DZvzRwh
TYDPGjLrgMbQLyQJf9znf+Esfh5i0Rhbvnmn/fLo+R8J5sea7JWuuta5+sZKZBSn
4ETcrW1sjD/mxF2tGq2ULO+amnG6Cr+OGQnTqTsqpZNXTusoTp66MS/sH+BubqZN
dL/B4fVcZP0kG5B6mZ0P4/veiWcwWn+5I5TJvWhot2dBZeWbdjOg+Ltf7X9ro8H6
VCcFzo2i/RxtBaI2zu8K1+lUinxiElld8/3+28M4k2ZrwMOAGt/P70bxgeWT5tPP
aIPfTrwWao1LeWTTSTbM62oabLDyqC6GqXArHASfZuN1T9Lnq9AmS7ZLBW79zi6G
6PLq8xBuc2MbMNCXCjnBjPJCR/N0R8pCY9N6GaqYGUGZT6pKykb/wpUlzrSEioBS
3jg8ZJVhw4m4x4oTSkAUIUk5n8Y5DFI3geYwWb/bTZau3ySoZmig6wc0Fr17Vn4/
+i5nPdUV7sNbipxM8g8npVAZhF7Ni+QYLhtqpuAJcmkrdp8TWajbnKqvgf0Xd6Ud
SQ5p/+vKs0b6M4B7EWBxFXUsGGTcpqXADD0QN0su5GKmpCnxq2OqtfvU0zTOkgSA
yhUBtoy5Y0pYGhtseOvv8NPv9mCL7MtVetB7rrvqpsKARhfwFPU4Gp6k0l3sa+SD
BU9UuwJDYi8AKtRh+2uJ0thUEQA8qkEfOcuLQWIwNeps2c7BB+AadWzPphrKAmB9
JU++ci9b9eDBEg4Gp0crr1sERA9Rg2rrw9YuMqf3EtLtcl/Mih7PRrqhj9s4k+2S
ZhHplzRIPVSW8h7WIrtl+gja6ymEVD2HWLf6d+VUsnzs2RxIZEuQlkfzhbA09/aQ
mfIvTGazn2NkORMJn8Wd3lF5459gg7BRRB+AtDZqOvAGd0KT3+cX3DVQxikVG93k
AcUPFDHMpOXh2MYA/ZSOKQXjtfd4W3Ag6BfMUi47dZQKNpiurIvJ2fW6SxEthHR2
LUe78uosMajVYRUsCXxB8dfhsdwYG3EtUF+tPyQleCDKY4JVZCI046o9ecoapws2
pRfqi91LPoErD1SVNymL2F1rUVrCL58Vg2kedEiSvCSlOLHougZSlF3B7nw5kbcV
dBJWXYxqgTYZnuQRBmcmLAbrVPrzEoFlqWL5KAGEu6PpZ1ynA0Xps614Y4zSVYmJ
huceRBHVZy5w+SadR8n93NL5QRFu7zqpHPtc6xNP5OazhomopBrO0oolvt+VTeNo
jVSur0Ycy2FmS8fNTPzKFZ+QGww7V2AYkRP5r9avH2aVs6r6m5G9JQrQIeTrGfLf
UeHcRHwOvtEJusx5nXY0G4mLSjIHSDBV4qe7QrDdSFaAprtTzDK9685pBGOlRra8
g+QT3DTYhKzask8eXkwufcpx/cg2CadnqClbG17RBWwxAAoAnSFaoLh1vd+HR5Sc
mUwKwSdNAMuW+HOXeO9HfIZo2UGPBMtv6ngYsD9sdoTKzT8S/OF3lctLMQ7VXFoL
gup4S7XyPgDQi8r9yIYsu75c2gj1/eLTqaNzJbzJKm81dtImYIWDYtDim5/na3Bh
KpLTOV353hRtT0ZZIUkQodhtjc46H10bFfF1XW5bmmKmptMztoQzA6Hu08mxnUfH
QxO+DiGJdp5oxvVePuIqwgVZbQpt8PXO4m8JrEpuH0uoxaNvitD0cWmmJ/AH7Wja
yE4eKMfN6nwKY64E+flVi4TxXBfphzr6cJHglg2hTnhm/B6w0JhSEm5UVspkEsqU
VmCnEdpSnayfPXH1wE/jiRQIT7YtZD19VHKGb2vjV3JhhYBjWYfg0X+CxLnrftv4
yNAANVOi8oudGCSfDEuqMOFxkLwx8I5mF5OMu/MCxJqFQx7hwkzhqsoMt7R1eM7s
IfQz+cZk+yPVdS1ECvw1sX20MEE2A6PYZBR8rm/IBHvEex2riIAgdiLVdAewm3nJ
bidDMZbn13oxHvunslen59BcxF6ojwU5i30w82XmaVLZCzz9CP1Ccwqj0Qm45aof
RvyzfLcn6NJmTeVN+zbyHsjTDYHEl3JQkealc1vd4yC5AgwChgb/P3YbnpqQjXfR
5bvnUqYYDHmeGxTze517ZakgYpzx1bM8QtuKycnSneBuID5n4FmFZfOT+ZHnuuZd
kWhdHFE5g/+ppPZD1eRdhuFlHLVLaOOnazbe5+5iXHbLskgU1IaJCy/J7Sbg3Ar8
6347cxKAP4Yo8OWC69fD1aApKdNRJA5VuNOmVLu7fefYO/MVthB5Zr+XjrS7Q776
04yYwTl+IkrieK2+In1eyzS8ADM5FroPwUXl8FlnjhUXj0cGXHYYWQfhqcJgyLyL
REPn5oU7TFFVRyvjQsLqynEtHelOTxN2IiuwyXvtVBLtujnSyGt5Hj2cdmdzJeCU
lPlxuyvKHX9jVEQCpJRcATXgdcEGpeODMaKhDZQz0TATHAk17IXq2enXGYetbL6g
y71ytbZnxdS6o+eHOhEXK5PR7K/PX49UjQgcEa3SX5jhx74aQIrrpJk8+bD8XjWI
5bwsiKO605MO1OsGkeQERWuZnBmgE80YuucpFKwJRh153tcE5ruGaT7RMJ/FRJWq
dtrpTQ/lxSIk83SEZXC1i2PeOkkUi4cImt6mOzUnTbfr6wA7THA+/Xoy7baQMWrk
zd47ysyuC9aDILcuAdybVfHofZqxPa+arAb9rtpXMklD3glUPeZb6DXyIWUkQcN1
1EBAP3a8JqPv3C9dhTCnQ9PGw4pGXbfIbd66TwD3k/83mKF7T6s7F+fhqMEIo+BF
fe83ZMFTxXNUWve6Jg2DyUlHXdbVq1LU0ix4n//wBDTMfN1KGrln+gQuSWWneb4e
aRY8d0ZaI2RFJD6gdNiCRg8TY+/sqn+RBKSyS6RewTgx/wYDUC2TdagBNSIVamhy
p8fls/EtZ8zffYlDVw86+wFHNuv66fDq4hGk7kDtFX5D6dwPwdS9ZcxXY3c4bLE5
sZvc2dn32pqpzjt5jslG4KM7iHcY/ndJ+nKL6g85O2dYrcFqpw/0s4ivJ0QXb5dz
5+cZHOLPbdWPS1JwvpNm6ix2SFKP3xufTH+dGStgcrAAljuWNyj22nBVObsVqagX
t/686dx1YYLtFez2rNIM7IQLlQ+Clgcc420lyklRXkRtzTRr0e8AmmLhpIKauzjF
sFWdSBgtsCXDWh27dBBNZDz3pgHN4xjpbxiFbBFS7mk=
`pragma protect end_protected
