// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mONRp8qSZrFRh0RaaXv3DBR0xSZzLBdZfmCXpxrqTXriQZuHpa9WO4iHUpgC3kqO
PttiBS8HYEbRQOlrAXMB/XTPniEqH5SQj2bEFHg25Jz8YU90bUMZjoDq/oPEbM1y
IQzDflFinkqEMhlS+FzVlFPVAgK6bYt6ID9xbTvfizo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 86224)
44xviQa4AxrQrHLD463vqdJYVRqa18IR/WglGR5y1yA9R0FPK7LGa5vJuckGjJDB
a7Q1UErmTbAL66B6loFMc/wzht5ok4RVYUPXys+0Y5OriInAbS0Jm7TXATTdj9EB
6YFvD72vlIprAuaTFQORl3ViHszQ261dKQ8H0WHWIYjGKjb9wO3EgXpHCsYPZKQP
V70poXZ8Qdzy3+c4W12aQ/YkIeGEE8JU+gxjOZ3E5ewLo0yowfEZhssu4QJJUo5U
nA62YYQscrCBLrdQ3Mod4lgrzQAZLOBKICSJi6NSh9SVVnFZklKF75AjVbqVUGSh
fulrxJpH2bma/s0+Ntr8mQz0f9f6lwIe2Kn3ac/D0Kwwry8FhON5dOeaklKRNtbD
nNhq12i769B+jzkxNCK1W068a9tgaoAkYwHhvIxtfdO38jpCpvRl6LzN9nwJZ994
KgvxonBc8Vn5ydjbNiYpCI9s5l90GozJYOFC8WFTCd8ltHih2ST0C90z+I5jo5O5
e5Wo/TeqcYhHiq03v+UWFlwpNNFwJm/azI8XkXxGBV/DDniEW2l+UK6Bfl3Ir44X
1ifC6oAnpV86sjU+e631wRGk+8X+hgyq/yId+x9+guQHjPcYWvO4CZo1TTAMhfd/
yx9gfKU8pCtpBss1pP8jWpfKMKhHarqSRTA3fluuNC3QWZOi4ORhNO4enTglNKjR
lSo1wZahSCX/27DvgXVTSMWg18fDksdhDl/uHeBFwoaeP3FGnnTtHK+IAcNlEEhh
HjA1Ue4sUe46IFx/gRVu9/gk0Nt3aOINtCqu1i8ZMDWMpElwe6YQEgK2sObNvJ0U
RjFMeahU0ZI1GQEe8//N4nH2vGCwY/EW1y8y3L18J695Z2mIDbAb1NLMF9RadA59
hFmlmEYNX60zfDdqDL4edzq1MYMNkdmIMyLVRKZFa/z5Hw3p/0y1mWfoPegsK32K
oTSZJYzYJuPaTtd8mYWyVhXcuSwxyTZeRA32B5k7ExXNVKoi5X8SmCz5/gdpnUWY
Uk7aKaMk/y/NRJ8HenRBPSSxjdv+U8jh9hMVuJ6oMjGpISLsDlgwKB2xwz+oK+AG
EmfJeLZrOSCtXyr38pRpr1Exsi86wpu27HBg/XXhCHf/Gtc+as3tJbtTM2/f1J4R
uRtrbz+ar6/Q+jbinBq6o20J9EjkFsAAWhH6GLD2nxEF47+6jDR9B8xaCRyWm3NB
OmzRiajoYqel1xR/d4UBY1m9fdHqXOgrbNwNsqIo0sj6crbUD2wkd4Tzl26LcTZ1
6YDGeOgd5idvMVw5n+D7r9zKE+MEF5oj0g7SAIUThl7pjd0i+ID0D/YJKmblH//P
+DkIDQBo0yJ1AcZwvZ306tDcqi4BcTjv/xVbJGTcFc7OtiKZTVQiHbkZsK8jnr2I
ArLn5XzNUNMZ89iwIEW031ungt0mK2BeEAYESHqnhTFl2n1ys+cwgHSuGM7dV0DT
rt6yn3e2ubdrahlIJaSE/64xOc4va4FxsNONTKp78NlxZnISSzOAKIYathUxBu3a
0qfZzTTLYYlpsrlPpj+I7UKgut6dgQntu1JEasOG7+fSCt9ivDTnPh8NgYnQPfVu
52j0+qfz2IRnspw+CADZYsnZm5t1oRzhjyoCjkhelbjKqpY6M0Vnxl2PUx/7w+CM
dePTbzoV/KbrXEPKzV9QzPkgQDH8eocqw3chSUac7RxYErWyUKe7e3cJSXPG1+dz
MohVkvtHIgbcQBplFQkLkh1eVdDQuCMfzyv95nNhTv+6RGrJSk+7E3lzcEP9Hrfr
eZElSmPD7H8mq7khtlurnROMZDCaU0a54UyrZz5SPV5XIfAT9/FlDHtN8O32fuSr
n3/ViIlqdwD+onY4BvCI6bnoxDclaPJsoOmI8p6Hx74Iv1vsU8uPv/xBWWudhrJC
4e47B8m8jG/EaoyNhNi0ghk4wUP7AeLYQf8cnVcynMwPy3awe3OFjIqm9/6Jreuq
WvcUrYTvzOD2GLxbCPOEURZ5cQG1oDdbsccJzuNa69xI2hJpw/b9UhC1WfAjemOf
kKCw3ZjyjFLLq308tu3jWBHkmwWYG1cUWycpKMWkxEdWmPJ73nfpidNXC8QCGnOJ
3Z6auX67RXN7RidbetrmghaZTopdzQF+GXy+3n0WkdQ0WtSYiRvX90LXaKXfkmbL
w7Yo1ZEIgeor9DJXHWn2hZdTSFJAKHJ1rQei5HJk3NOY0Qxd0Ylbhxvxl+qp/GSR
6DL8RAMUGlzi1K3r8cYzxijwsVZoLZvciIRioDGvAgT19I+e+PGZzpEAJ508siqQ
PboNGxK4B6JWTqMmgAGfHGmJbZh2gfurP0jSZSyMhDszvhO/2D72MuqHCsRut7bH
Wv8bq6Ax9CRWM13lobjkd1aTpA6MWlhZfZWij55gt02JUFec9PEokfUOGB+LrK9f
hw/JrlSA4I8GNm2tAIvzmnueuj1+bpiBd/hk/RU8EUAl1IXRLV6ePJyjRU1+2ue4
D4SD83amQbZtbNvOfHFqN0PYCoXkmiz8Nc+V6vGgh08t4t31jCbKEhiupQ5YrTOg
LS55habTiQLmqwvxG362LPHuS9m/KV3JMwWc1Nxd3luD0f262EvqYDBM0UO1h4zp
dyJXwUzzGGhR1a7nN7/E9qwwCiplxJMgerWpyuZhzTbLsOmO8TVmhUVr3oqnZmuI
rCYETwdRC0IoNZZVdVQ/s6+VDaIaAKRA5P5tS4LxWHEMaVUxscjyxGpMA3dYvA1v
xOF3xWaeq8JgOI2jeN6Twqf/EkG7GdsdDT6/dcAHOM3DRZXbnNdfd7AS5RR96yO8
9z5a6xqw6fK+6pwriPWMa3GBFAFWUU1NU//+kEgQ/bqbxzxZz2v4hoyhVmNp8Cwq
m9YX3x3/1+agpRj4eFcaRCd6IoPW9g3VehAHBW7GHVFgXHptOpwfdh19kMlOr0tx
lfZC+K+TnT2ISpRMdPgxLaJgpZhXeGIe62YAQ7KqyqXERioRdQEY2NE/FKjDFwJV
FNTlqFj0EBQ21jpeX584HKPuCrZIZ1PMMH3CTG8yo/ZZQBOiNL+q5JNWkuZn8WpG
mdO2ALTSuhDdkKjcVbKzNXT3gfCfDOyl+Ow7nAGEJRAi8+mPCdMauARfur/JtAt1
InJaI6OBN0O3BiHmxqLG/aZ+sbOTg8qEfkxzuvMkzeinyCwnqdS89IfmyHvr9j4c
NgVU+F0tXgHNnp2LnvdSr/SAVwTf6gS/yEklVp5YwygOCkc8hbcQrZPn1q6gM+7c
HtDHB1QWfeSFU+pHScmLyy6FKJC3qT/3YvS2Ayw60ItWtCjlpWxOlTUka+cEk/1m
/2DQGxdn4EV2v+m9Z0RzzGfcr4fEXUJNoAjkL6q6uOU7bYHJ7LaFDGUuz6bbRTUx
HebWi5DtvNmwWBAuzOQSigSDqMykaV2z4NYtdXslBHfXcohAUKGRKR/ffCcpH2qZ
AU5+xBmmBlbe6qJfND6e2FHGcT+iljsY1JxJ+qrjnqZzQZDAL0rnS65RM+qtOuDm
I2YwephRFDIz6X6pVHa2OORbp8MTyH/1CWKs2F1fnY750dxVxEvHfrj6MHJBXYQq
hUbZT+XMf+UNr/tZi3NbQnYqny7cNIc7Tk1YLwSG56MGWdQC3ZLMuNsyjSMvo02L
ZMo2vmFEooenknkV2mj/RsO9XEPNdbaZxRJQM9d4F9wyFiL0DWU+sle1907G1ZFu
px0q7xuJSdT/RAold7OB9ss87tOjNxN/2sepyJVPHcWx9nJ16fF+4QLf9o/cSEKq
YKIAYIk7SnwJ19++yEhmczPLVM6NJizf8ckSf63ce9Y47SME13Amdx3gXPtVSP9l
aLRwsIQl/4nSgJbAzWrrrU83FDLJ9QnnLKOaLrpQicu04bLqbOdIpr9lFPiNQRSy
lwpnfaacxOoWf0A3m/O7kuNeLM1qjj6zpMHC8bNERtBhdSREi0QxCre13GdtzkuK
JBTcqoCaw+kzoEkJ0Cedkcrt0XhzsgB3I4jhxA/KBpECieR62NDGICuGOmT2M2F/
M0wx0HlYT/g6Zd9lDCStVIW0JaI0nLDHAhiNJPeLC2KaxAbgUPZjHsZIt32sTfa2
xhTjEhv5B1HSfR+uUag5FrRX+R14Yn8BASVeDnuvxMVk7PRKMFc6/h3aEKLen8Ez
k4Ym8FMkVoffLPN2j3a5cBVsKtlWtd7iiETrmHnuceEiXypSzIkldZdqR7qO/e2F
A8PwvAtA/XXJgOjUyXUzkjurAfRWPweM6AxPgwrL/frKlDqRozRXqykCjSgP/Cw2
sE6huLt9OG3WuYC714EVjTCEroIjObBDJg4GyhU6kuj2aii4wekUhvsW2am2NW9/
Qar37Qv+NeWftGxAIOK7FCYf3lIixXuX7C1zuwvB4sCn8/dqKIGsZdFVq0W8YZxA
FawudI81vbO76T87iuj50/xjGQo0qtOcYwlqRvxOm8NtuDY5I5GnGSinByFyWGfG
PLcpIuToHRaab4oJ6skcpwNelHGORHHnglhkGq+7aSr7Qfuf9vjx9xGtlsdTIDVC
lGnK8BgzmUsKY02uthMfPh9K5b0dbUVxvsqmRwTnLERtonbVTmp1tT25QpquDw/S
aJF99ITktq8y6gkWbX3sSlAesi5nF0uFysGtny2a7+8ILztaUodHur/YpQjHcuBY
/pypduwhG46Y6bsS3d3TMI52HOBX/R6VIAfljesrWfBCG7ad/5CPOEC+LsQofjkc
KcyRueSP3ulARb/3watytBhcxuaDUoAn+DTelUbVVjlchnfe3kvtGotv1zEYV4BM
+K0kvntito1HGaEMkaN8bdh1Muo0gWvFSrzbSLTyObY+n3JL5e0W0wViG84WExlh
oC69b0Q3UoMFKiASS3cw/KikBqrw3VEzmt1NXnsoGCi5WrnjjPHe9MR7ASq51ILC
3jXt4gYrLCo8OAb4v2J6YYz60VWw0X1AGIwFlZRwbTj721DDt+MJHDg5kokgNL4c
X67D+5XnMuR9tZTNo+OZR+4R4yVmjOdmsI4xT/vKONuZVPCd2mpPvF/31MGbY647
Y1yktQkG+wbGr2unq/V1g08ubaYLoi1k92V2zcHLAMsiVDkAOOEQFJ7v9sy+3KBE
ykBn47mD8gWKe5gKnMLDJFB/i77NohidnQn53z6BAzvtc3dQ9/FV1yWTXVjQKE0d
28ywbEqxMN+iuVd4IGqrTTyeuV0BUZd1S+xkBjH9IJlcL1PXYvJUUR6AyHO9YzBr
+2uj1HMsE5VQnUC6Xa7LyhWd0if0L5r2GPwuCQzfrb68xXZ38Gr8YF3MUcHbOIlY
eVF8wy6B1G/JAkOcyg/vgxUOXQVhasG7rwPUNywlHzF+OEg0tl4yRuY5mrXkrOZ/
prwwadwopd/uTKKaqgWhDgb7W61+DKjwKyXAxh77C3AzOJc6ZH5zZDKcUmnx1iaC
Dp3Nu+Jvkmhyi+CMtwJ3dbf2pkGglIbziCbtVcPiJx5hT4mX/o5+83GofoDDV58Y
R2Jmk2o+2HeCfZdtYVFhyIS3a11wo8gqQ9lJGvto6f49KvGpzQ5vaKM0eZ2RpmWx
3sPVmIgtkb5EZGKZc7ovOQ3H8w4uUtbxbZqWXTWmNd4iVB0M4IXSJbyUKHDHqh+0
NRkWiskwH0fjAGwnh6ZQ36q+yorDx+o/nYZM6G5oATU3IpZPD5DWjfngMtI3et35
uiyqlmfrwsRBn6sjk3snepvon+Cu16/2qNodefu4bGRLnpYWv9kF7o/sOr6XTN1W
bsBhoGXGGD/rpAkt9FAu8BPM5odfYqGfL1Is3YxzF2CwLnTAda3X3cwyYj3HBsz9
y1JfKFwXwoJ5YG/BSk4uhEOxvyf+5oqKSgA4qcw6e8axSaUQAgwe8LIppTBysmXA
CX56VOsLjHvLPNbQoqEL7YBRepcSR0sDGH8jSUE12M+2ITjh/OcoKizmfVX7Szpo
C4kFdiDwlmAz+qyAzZsgwCmC8zYJbKMGs9H/zSlSVb7Bt60kAMKYIARqo2iL/2ld
mstwSWiPIvJLA2APaRINYzFdgNwUBVtImr63wqHuuqonCAMlkz3G7jcmZo8UnXe5
VnMNaFPBerMxIupJNbNRGnZZl0Ml7JKKQOV3L3bAx/sW2mHm0yvzwFX01u40bqCf
r4r2NA6gNOy5CEzfbQdCjmAYHVMqweEtcUpmgbRAe3UOcwHjBZt2JfqJQKslFy6x
6LKLisvlJh1OInU17DYKA6FYWxW30HL3GrubP5b7HzORQUDVmXtN/DG1diANZ12t
IIF5L+dkB8P3nPDWMEKv6oLObaRGD4WAmVglP532gt4hl6ua9m/ppr4tf/PUBXu/
DU3puzcDcE+yZCoI5ghVcNQIHBz0QdsGlgBz0b9krmetT2eLnVP2m7btpwDbzFlU
F/mZbZmED6mbbhv5QOiFAcMjbx5Oc0AqAIAP8L4I31GgR2NUlwNgqXAy2PP3h5fx
YvONauAdwtdzWyl7HGozVSJPzt9LAJjiYuws6PskCdwRTHxSE1zI6rFaNlkfWzot
G0TdfQ2hgKvcjtV2nlgDeNJqDt5g/PF1tMGdlNc+UPrDkyEhQdc4W9udmV+TRtKE
9IGEb8OfFgCR8TU0CB1INVG0EIwvl3qpjvrYUdT0COl4FWFeDE6JSXsOfPojfIup
3VfvCZJic6t3m1kd6p8g3eUfyApVRNLbPvZmjg29TkadVhC5SyWNbjPW1ajE2fhb
hj5GmEbThISQMyZpK6s2GX7LWe5vKf6EAAu5g7fBGYrjes2j52FymVAWps8RjuQe
YzOjkftJddW1BvFSZdjJyqxV6FFsqcwIe5qz5gBsQLrbP/3B5cfHYU7KjtFTXede
vyscbZxvZgneRKsv6KOT1z2zrRwoiis0s3wt99E6/HIgMe4BglqHGd03XPYNaxTu
bX6tXTrU79eJKPkyd/ZJANE4OrWUUZ3Wpy3fC65cvNbsgsmm4Dkqqjxn6GjJKM3j
kKn5MpVhY83odF4K/R1jnVbv0nJYr6xQ1jzSw1B/Bp88vHWj4imrqcXuAm1WHwkN
y5nhAMq9fh1OYNT3IW60PMXO7YpzfIM13Z/pgQspV7FsFN3YhFMpn05TpuDvEcso
OdFOeH3lV7YNHzBYZhiijO1x2mcxfhuLh7nvWXsA4H443lQ1CvVtkW/NO0A5hXlE
leZN7MLW9UzX6cMLOHw6FRgIedTKqEYzq7FE8aS6FEyw33uK7t/DlAVLz7qBTBGY
V/XOFfEcO78BHT236KYlypkmS4APr1TcG3GxSq+ofWKdbxuHZUI2dqNEJr2Uhrf4
6eNSICPZrdOXdj9xBI1yLVdedxVQy+n9D3dTa25caFxKiMq6xQ+3k35jCJetUTOD
OepfzGGe5rW3PNJzeD457nxiPNEnh0kLpVkT9Yc7sZw2JV1rIaLR0pkbgYaBd0DJ
/YNLlh9mWAdE9RawWRJzC5VagMtfmU6AHOzeIbZf2PQlPxjE0VVpaI6waay5KEcs
G9x7LhiyC20MyhEzbuFe9EPSOtTGu1kKe87Sq8PEL3YBb+RgBBq1b+fZYjr2/LL8
hBfVTNB/OD4vMYEKoN1mUowY8h7+fjNjpZwu3SNqLbxoel9qsUTnhVhnazCgqxhK
gsCPi+q2r9FWUC1tw+Gk8O0LqW/X1XEn9MXdzJbqzhMF9MMIQMSXKq6lXiK7+pBI
refv7C2j67SR368eXW/nBvAnDcwabCS9srEmZS+yFT90cqPtfkH+TRgH2ZCGdJ+o
t0Iq4GmaFxnU0GiDzDU5PURGKoLurs/ZAanvzClFwBSdoRliR+VXoBDfmdnpeATN
Q8VgM6O+4BFOw0uWKZsZGAvXjjkldCky9LxIWCY2jdTXN7SdkJwFn2DWFNfTElUc
/5aW7V/I+E7cuYZKN03I7tbzKDfyXRXfgtADvHpoYz+TvuuuvrVRARasw2985a6u
2fWnEuWo1jZnzgi3sfpHN9dXY7BS2h9HEnKa3WbBqzZiDiREWF5+HAhQ7vYjN050
ru5UYTxIRrhjqYLv82LJyeaZR7Jz96yd4/W4ZUUP8oKlCYzMliDQM8UHwjvRaCrH
F8r7KhJA+zbJN1Ox+mOHCSJbPDgFv8WG/VoOEVHfyUiqVD3tDNKE9MJ/BaYKXUE0
b+EZUKFcOg0zZy/313XrVXZmr7YyN3MTIWvvT+d4VVjc4R4PqDy+6jjLN/uCT1tn
NHTYES7oejVZH+5dXWF8woA9/LL9PYnT1f4+pIA79XbXR746XpN6J2HUkJOyPFob
QQJZFNZ/CqGRwTCAntacQFpcNSPvTCva/nM2oaMnbnXp2MhO200ez9Oly3G8tc4P
Iu9wJbprrMdVcQwlYLxNYD7tnaj3lFEOjiisppVEciIcqZEgK0zHWsR6kUMhbFaL
EVqgllQO4E9Ldo+3vPuZqaMFTfdbJtXC9cn7Sbbuz0ZmFAUSlyWjq7tkiHvCFDfJ
9BPHtf/aPTjdgqIPlDtNyHu65OpCb/ZB53cNgc7RgcQ+hq0T51yzTyMx2/sbdfw8
qsLMsFQr9A3NIR0NY+WfbxcyDbaH7y3OK4wMeZomGeNxGeVNcFrqJ6GrmDXruddA
K+bARFGyrQDTPjxr77sU+DLricZUcv/8B3xxlef7uvuo1x3jvDB/MpWxJISPOgbM
onKzZNNaRsZSSBYhQb+Gku6YsR4xU69NXDJOehZsho2RehAmLT67ZZUQUwn6KmMf
NihBHIMOdcIDg7bXg5pe1lrYsJscSMFgagHqR6nTJAgc5wxxCjKzKXrcMQWeOEE5
mm8wkJMmNg3XGFnedXFyDYw08C3HLqJwhR6HrkjIdP8g0zw+hNWwMoMzIrFuXHWM
9w4JU0toIRSM0fW5K40DoevLf6Iba41DaaEGjCQsn5IAIGzJiiaGQK3qF0/mojxg
Ux9CzPb5dWW6D0VgSuQT7NbtEzzqkgbtqjUcvyZwGfK6p6xbFWNJJtI5DnDNA/oW
HPXJCOmPPXdz5mTE/Ggt7dX5OeVnnU1b4DvVzLB3tWz8mppu6IFVhAN0Ix/Zc3ym
fZL1xKhDr1nfyD22stSr2iR1D67cABlAnShaNfo/lg9DLM39rtd/ehmtq9i2cW6X
q7GjcDA5i1qr67g6u/mbcRpSZbtMDd17VxHMIj8Dt8oBDMQlbvdQTg2T3V4mZgFL
gqIL7bq5g9tgzqjcQsrrIvLo4ZT1sgGBoZjyLfvauWz0dN8RgLyhb8H5w5iTyvgM
Fpup8g+xfogswaPyJQstqQ3p/YMACFhsbfid7XynnseETpRrkBVUCYuWJs1TeM/g
6DeZC1KpKb/509EdYNjeKCDWEpxarELuveGFOprRgB5u1dnLf4wqq7VjDd1jhlL4
R1fa2vlTalAqeR59lj4oAPKPC4BFeuw8ATF7REW1KNp8BvP7aONc/kJ83mMo7EGV
5XmRa89HDEW+1Id2q9zvbyQXoKgo5u9MOQU2j2TLfFOA1IIFCguijqEI7C3ERk8w
N0XOkNWkOPVbSXLj3d06lQ37vQNzp17ZyyAsT49ZZp+Sl5DBAup1Iyp0p7UCz+FJ
PyUpPJYZcKp2rnYxosLaWI8dfDp8tjRpTqe4+QEoVXlm0S7VJFBsh6fzcw9p1nGu
30WsBWFIWcmo3xaLgvkYZ6vIKVHB4vxcY6ri2xFUBWhIREhQKbptSVNKj7ORYkue
8x+mQE4/bJCV4tbCPaY/j8NWqAykrpCMJprHCKk6QyzRIqdMcdXqsbzPkVQzGe+p
b5VNyIfAnF6lDg8RYhcJeNae8UPI4hs471rpC531LQclzUwrt5SOeQiCgqGQKPir
qNaRc3WMp4wfX1aL74Xfr6iAgYNW17BPhNIcI2oL2mhBnfaX2u0tIFy0wMhbM4cR
9Op06pX16QGLuRRA4R9bJU0meWzQRnjmKYBh51fTTRTmB5a1FjOzRKiGUHu3vnHh
qlLLyJBuYcSXWuXI1ZspzTnLblPeHpby2cL5wqPKxNjKYZYzbKrQ9QdS5/ifv54g
M+SaqT3HYrul20VNxJM/r2PqomDKr9IUS8+FYnHEUe8Bb+hdDgzUJSTSefbmcGl0
46mqdaanV5USzfx+bzkRyT47grq7ERFBGZ0DdJFeTjdmZqXccxpdSARB0ZzLBF0i
gI1agq1bjg2Z+/KgAu54qMRBI4vguJWw8tJ4+Yft8slhCSXB6nxa9q02G6+YKzWr
FSMUrNia8zlmn31AaaLLFMw1KVugokOjOD+TI+L++8iC7UQK5ys3bOZlOEW0NuBY
81vlC+NHEiin9I7d8b27ABJ/aKZE7Fbi66ikVL8TkCAUH676vc9twwmgpNR7FKLW
kGeJ3h3KD7YLdMkED5U51EoYXu9X8HYuftOTqULyLIY3Zav38ucs0Cb01FTQ5KjZ
aU4ryLQfJ/GaTz9spy7PwXpO76/IQDtUwRrwftTXopDDeMZKxRoCnhJFjAgqb2xa
CJW9ckzz9YFOk46OwWy5FVpcg25CeeuyaeyRabZOR+585fRdpemRIXUJm9yrRYlT
njxTipV6A0z5DYng61qqC22QzEdpqYgOFBE0ZSfKrEozELnNSzByw6gqXEXEffIi
N+GKinxKIR8cu9Aehis9/xperu3updOWvtl3ZzbmLDFMRAKr6YJNL7RrPEqMvcE5
KfoBA8PBv7vxmERy1FufZ4pnoB8btTGYfHQ8FYgtOFZ7ELNbmZ3T3DWDfv/FqEPr
/VjmMe+iyhKSiq67XQezJJFfcLHP3+JmK/Cr286Vz90gOWJmrQmsuYcQKtc++dkj
s3dLS44QpJEIh1hZ/GlDRR68K0QjrOPW1sw4fbNpVVHQ9L7SB20qyG26MmxhTn4c
nG2bKcCFSrbwZeHuexm5lH3YfnGLTxGNFnScOfaEbJu+vzE9doC/7CubpZ3w7O7b
0hUmhk7ZjewYggL4LFO7vOgjpM2jUU9M0AnNwkIIAgI6kWeU30bOG4ifcPxGg2XV
cq5Nhr7b8uKUV5cGb6vypTzbk8FuWZFRST0Lsln44NaIXgfOJ0Wly2Hos2jNY+ib
t2rl/YdgoVkaLcMdh8krKAEinFBVPWCeTx7D3HFcIvApBk+SAnZgv5HS3Y8aPQe4
OxyiQZF9bdCszmboBkt6ndZOUx9pLnzQpaeMWupd8T3xMljdOQHuRHq94Y84j5ok
gz03m2rg9NGq2OQdJrhyiJ2XYdMYIkKfhSHqlg+TNyzJoGQqdvVbiVT0tj2GG1R6
Qvmt7J3vTWANozIJiPAHogDWpg/jgmu3hD8p5aOPmjxPOCsL7uGru5TqYh4HXhC7
QILalen1HXrWOwNTnf1C8zI1BCci1A2a+IINTeSbuAH7OHv6lgrfXVRCqu22K7ZG
IusubMq49681e93xecSirtw7vmn+LWzxqD0AUTJZ5AuHU38LLNSa4g5kW1S83N1g
o/wqgh7/dWiTYH1pY9kZLk8iKubO7yxmCPpwJFq0jT8gDD5Hz7I5FvdrahVZOat9
AGb7HTQdqc3DDy3+5ffYaoiN3AT5uTmFEvlWa6yuk8t84WCuqLxznYBwZqEC8gYD
Iwx4ILKhggfDEox+w3BciIE+p1GTL3evDrqsdwf/l2a9jdYyFIz8mhaaPhkb0W6X
6rqI64FQ+4UuRgELoDF+uie5UBzaUG5NfRkWAFsNm+bKAOC4/gVRJfUQ3qJpG91n
AC1tuj0pojsPfz60d54BxVCVVaA7HlXsaQ9SWtVPxsfNeLahIMtP/5B5z/vaKWpS
p4dz5f5WsOy3kzFYw+vQii3cZ8GXgUYsiPa82R4L2cqmLwqBZ70QkishMdKcOyLM
x9eOlGT+Hjt8+YEz1UcJJVKz3T185XlAjaL9NT8InEHUEdIgmrPwRVddIzPh8aXt
pGrg85eESnQ8w5aZZyQB9reAoAXvJFNYi67npRJX8ziFuukj1aoaVVVyMKaAtX8Y
TvmfWyzECiK9xVu/wuh9VmW2UMWtTNFMNfkyHMkI97QEXYVUsYXlcm6zQAzgDjOD
fFzSClxe7BTdThWsLJPXf0NZe6/KUxHUyIXx72/grbhKP0wIfNrb5dh2yYvwQ1NC
h4QDrdWCh4XPI13men4JTZSVCydbHTrlEzGaKCvs/S55mMqqvlpg/evXiByu7ald
7HdvV95hIk5nAqdkSVx4jMabsHvUHRJngIrUqceerPORHamdDqnvrUqzbcApZ4gZ
+QQQElNTwr2UU46Jv6/FlTjEMRFjnUciDsqUfDnY1Wy63fuBiUhhTqh6mXjOAeiS
0qK6TeUmoS2c0PTlwvlfxd6bXtnzvgXat3D0pmKl9mkiBLbxPukkl3rq1MENtTNj
1BE0aetCMLemY3f/BykX+k/jr3WxWnRKkwiPdwiE+v/EJkQ1TgDkjM7sJ1Lhw5sT
i80zrIPrNARGD90Ol1vUNRSU6lVlMrNqE7feVrYTQ4Mg/mUyZQKlZn0Tq4nbMzXe
oRk177VWmNrl5psLSM2EyJD8LRhKh2WPToFt1aDZ2xw2N+3N2ANipAEsroi6zRqm
Ieoh0/iJdBPew/I2bWK6h/mHdJneyJf0VmpcgO1B96GOQ0y96z4it3cmzyLkk+YC
m3HIeb5pVXyV2fr+w1Ee5Z9ad7I3LQzgy72bYRIBBct4M6oJ1nigEx2FGBSuJlym
NmyyyIdsJ/rse9DEA4evFPyH6cSzmbSStJpnw74US0h1rvQMeeZ7dyfS5PMAiwcY
mrkLpuiDtMi1kbdd+oRsuv4wKYD4jIDFVZEiZMjKMqK3dHg2Le1bwpHfJd7Y1CAa
JxJdvlW0GRpB/InZ5ebfpZGtWOp38/+/RHDBY8cctezL3ipiCnynSjV2tP0+sBFU
yxs+n7lG1xJDF6GKMt0DknwPiccRmKZDkL+dyUz+WQMNTg1OnpjaXczyy/15PSmr
9JOJZIjFGN2TaqWOMCQ62yH51zbShaVX9JRIu4Ene6EtfQhkyhn0tQ9pf7sy8g8d
TFFG1tUokcRluHoW5ZgouA2TcSZKyw0wQwDAm6Hk8K6hUgaYuy6KxXM0CPEk6Xah
D/uwYDugCKynquYZg6g8p4UtxHMMXCJAyC2Sd3mLd5X0PcjlqYEy+AOI+mrRq2U4
2PPbe1Pa+qCQ+ws8Uo8mMb783dAOHIyp1g5V9xsqPBN520sUy/97xAdDlmW5pEt2
7JME4IwXreekl0x8RU162AdXWn6cRmLUtI/Ik5kbxVinPRondkWtAFqEtUA6am9A
+qcMeiirAmm+VX1Fg3FxG40JmpVx6lBenCIyhsJIGG3YHiN19aB2lbM0IDJUmV27
V8HGCYO4bLR3Pu+PuZgGSTGdVaOuDJ1TKMbBerbMIYQ+fjjvkeI1zpbVf/RIwUp/
crA+j/VAkYFt5CJv65NHEkUGR/M4U9L652ws2O8LRKAuEjKz16egQ1dUhswr2MAN
sItIRUh+oR+fpA2XsyRc0yvU4n6+SZNlP4Yxk9i5k5XUova8eWdODDbzfZVgvPFR
UZtn/g36sVPlxlxmhf8GeKeaEJ+jyS0l6ZQ8lyCdZzEli0cLMauRgQtZFtlGRgUc
7RwG8Wwks31/0h8GWXT+j19UZEfJosLc9z1/i0CWzY9WIGQFmPqeaKcOi7x69itU
A08MVLC6uxHoplfHjyjvoxctJR1wLSCgD2kG+G7nq7ovFgiipKw/GmCJD9tlQ799
bx8OUL9qyOyRWzuhy0KyKONuPJ6XK6YYgqo+usGsUQm0DQP+1GN5md5ma09pcfEE
ca+/g8bWf1ktqItdePNBisxu1DwtQ/xVUwIBI/7xCI6UwbFAlD5/W6WWXQdm3Ork
wn89mPIpIrtcO4xT+0pAv1BnCC05Qg2yG/8v0boE+7Ap+BKdqQs4/qnn2mmjdIfH
uX7VwZuPakFEmZMajlvYKOv5LrBNH0a6QPYOOsHg+IgKElQC+MPxoD8V+Z7FI303
OymbasISNX7Vj9sa0isUUBtEflc/rnUV2qeQEt78c0BnwfObCWuMxts5VREx6wT3
JGQdvVnNgt+kABjy2WHLxeRtm66t0puWVhTFEDKqdjcAInp+ppoIgW1D0UxkjQ/o
8M/XwNbeK9o3Q9e7Muh/uSuUwTjNTuj9MCkvbO6/YN6dAloOV+zkawlJHbv8aMo3
FT+R6n25WisBcWM4dN6yplYmVOqONI7bya6dUMZqlxp/vxfkfhRMCYyLloWEfhdK
kXSQ8HUCOruo/zH1jnOpCMlzVphVMELSay0KD0UXUtoGVEwdWBxs/8MWJ7bwYDh+
bj4a9iph/m9Rx1jJJLvk89mWKsyHKBl7TJwPu3Vzo8vpwAYD2LzM++hiJemsoyC8
evxi5xLioyPvguoQcF8eWCXVlj5cAcL4DdJKc9CHUl7NNLXJ6q1MEKfxrOcyURDu
dZqgDV9+wbcPrKkPNfnTKAzCsPjlz5uqC5dwAQShKv4HterjX+2SAlK1qJ04YLxu
/KuKuCu+J/l7vTf/zWAgMJR1cfuSSowmazMgnP46c0yZsbkvl+6QBBYg18xd9ZvK
1SdA0k7dTSWaYdJiEWwaf1OuJMJdsC08dbEUkb7wjgH4ql5KEmfvYhlSAW/7khjx
w5CWqAhIegjfIdmyQqL+4tfnv9e3pnzH3N0Jg5whXzisuIEQN2HDxJ20ZaLeC3cs
ePnvn5F1cNyKqUv5Nx86r7EqfrgSnWa7q9ZzRNpCj7/SlsBDg+IqWnz2DLDYp03x
5nZ9wMkjdcxznHb3pV1hxYemqdoHmWNrbFaxrBiqAx4/riB5wsq+/ow98GSExWmr
hZo9QiYWSvRiSa5FJ2YSYFPbiqOIIfVJi4shYdCSzaMfD2uuDDrDXVQSUVmJM2Eb
jYMbRgKogEvP/e/+YetxB+gu9lgWPD7NLWKaGflyxUahfeU9ibnWk7vCxC5R9oie
fNDb/fWMMIbOP5XkUNzuCeMp6bVeGp92zSXk20Dy+tPJ/Vb9bY7BpFREXMNSq2jo
QNeTC1woB4zuR2NLn+iSNo8UQX6zhNzpswIpYgm0DBxfPqHplec4/o3pYaCwpeW0
cnjCQsCit5EgeBndhTywuPfBHduzB7p+vPV8XKYVeX+uNGSmI3/07GS/tGn9jqyJ
RBFh+9n8LHuVI/Emf2CvcyYm9ZE0WACHLDn1MTg1RJAZLPwHiQ57NydecHt/g81P
hbMx5D0rKY/ME+JnXH5pV+Bem6EqICcQ8NWCsrON/wHwWVrwPo3bYjE+cFcLPVcy
cNo2a4n9euqPJ1IDia4TI7UOiNvmPvwlHBA8JMTvW8Z4uKzBQUxUK2Du1Equbdox
0KDJ891AUHLQjHV/EFGPqmbBaV1qMjUr+a8QeA7s00m41p3dCQu6dbgxRv8BSEwk
U32ONVQFQxQHk1FDRNb1ek6XK3pnrL1+neWi4ufN4I3qiIGiBnO0ZzjLpcmqzrjc
HqQgb4AJcT/9Riut5IdF0oSOL80/Pv4to9Oa8ONXMkUD4S8XQqPZVBYHuWjW7nfR
WN1kU9W5X0trApMTSjXn0y3JMuUcKlOnXur9mbJSUJLl5N0M//65TLFYOM9RQJ0E
iTuZOws2whx165NcL0U6QtQGczto0ZUlWmzbCusq5xkzPFOtNkLwBUujGBT0ix2T
NtXyzZ0Th0FjhJz6YCiYV7VFXdXUp699hluha2u3x63zjdyjKxfwLz4BRPwLRo2g
1GHa/TZ6cqaHfODWHladecFf/JKJDrTcKX6V3Q3suc0pLm7+34843sNhDmGhz7xL
z9SdLUFr2yxfSkH/vOeHNZzxZopBfjBaUVIFT37+8vDAz4ZAv+A849y+5d10shP3
qr1IST9XuwaGBj1E4nkZOb0GG5wzDyii/+UKxn3mpVpYeo/DkUnZ3exzrf3UX25/
scrVhw9e/wp907KjZOFFzXUADl4NW1S5roREODynyUO5jRnAl/DzusNbolq1vbhR
2mSP2nV6nh9jFcuyz8pxbqfQa3QOm/W1aFD0rO2ZdSu9IVVvtP3tUj8SPqDUbrWE
XRksPWlUjHTrfwM3aiYYVxH6l9t0GsN3fPBDAmX85l8tXK2IG9JB2LSqbMfmg2eb
rPJYsBjF7XfC4r01qWA/bFN41DfXDMhEEong2bRiyoDEWhmM93bqHhYoKvm77w79
CQLeE31eqgow9LLSWuwHaOCKm7hQyDLk0CoaTqEf4V/wPvYcoWz/94fS1CFYCvUY
ipS4GiTtvEVtpjRQr6lG/6yxUVbzxuO5KOxw6jod8nwFAf1qkegb8l2JtC7iGCu5
pbybZ/SXsXVsfJk5MS/HadvZxada1l7wZSB5b+PjAszK/3GOekqAQ3Fg9rHfaT5e
oGyFSdqyyG7ORvZFFXvfGIylaIcH+XtyEwgZQF5B02r9NHygWUDk9/2R8PONb65y
vWn6G5054jPzV+A3VF8K6D0vjFD8tzl8Sq/FFzKNmDMfl/UeuqcJfOQUSxeV42I7
fPIVNCtdZL9v+SD3F+FcwoRrtTcD8rHCIxU+T8FA2NDjXdxrdTc9GedVwqIDpk2c
8lnr2WqIdmTv2CqpXFYi29jDvlAVJJjyLm5pEUrZhF8FFOq6HTpLUZc13P84MZaq
myjvE5XXx8Z1tDjxJN/f4BE/aW09AgLYlcjg5apOrQKCJKFrPpd4WEYgcEBHjcMv
wal9ywp3kmX16V1BH9+dPowxbVV3+CjZJOz9pczqaZeEu4hHFyPhTI7sbVFdrA/F
C3Jky/F+5VHnntvs1iXkhttlUbQnyqcbZzXbU737KnkCCk2NwZVxhuUpsKSEb2c7
1dvwk5DUPQhXH3UFdRS1wDoTb/OeT0R/vdjYpU7Vv4jcd+Ky/BxfnfpLeEaktmC9
kQWJRs65W6aiAi4dA5W3SJ3FTfjWkqHozuXHkF2u61TKvppiuAmP86xt1g90PiUu
LaXOjPwwjiQexdlVLIHLKA3l30j5eC91TVWmFEwBafLqO9zZh1/wX0WLruwIWDpn
6Ysyvv593xVQ89JwdUZJsR1eFJfg/Ujrde0eBSOL+S43DDu4G7vLgQ1niAAjVOLN
2OgmOnrrylvR769BaVQ8TAk+XGElbq0uFMYNko+kXlWNlpo5RVEj8m0dvGd6u7aR
jLjVSuH4MM7Tp8pXpj5/9lx0jC/hsgRm/vlwvy3VMG1ftSKNsELAm3Q1zoaqdP5P
pzVtGBTioX972CUs0fLJXk/BCe5hBwMPWBM2thQmXS4gBCh6rRZm/xy5kB2hGRkH
eH0NHbtw12PXSvqTchzeCjm84S8bS985CPLcLTvAODx1y2K+GWwcqgnXapWu+di2
GleKcV7nTyViETmbfzGtDPVBGm+YyLgULi/Y9RB0sA1Jj6qT10uZFRz7RFYAK+JJ
LI5TNl6kZXM0SYTUxrkGUCCzfov3JqiIO7JO+f+2FIsWlFAyWOnMoGsSDQue/oI6
vJOgsqKr/LGflxUfUZVYELEDNXeu9Gx8D0PEWc+UsYuVmrA0KxC0mQFGjl23na3m
P+PotSj5FA0SBjOn5WEmrKZzHtkK91fxqD8aZ1OGKTLT6aHLmqjIKZDjgCMZx6PZ
jnAblS1TzqR3qCLKSx2q5P/mpN1mjIA8T8doaeJIHfTl2mFGcDW0y7OC76AhhQEp
zj3EWomX0CLU8axMbOpInPRWOU5j97kMlR8ias+M2erFpbowb5JW8bnH1GzDhuh4
EogwURza2rOmvd7XXTcSVpFJwU+BBjJP8MLnmWeIcRHBF2agTjMWc7swYPQWELuy
1nhYOKpmTCgzfOP85TLkFB6IFNZpdHk8QK0cTk2NwebMCMCOuWsDABFfnlAVweHt
9Or1ry4O49HTCtp/vZrZSPoS/r2WLdZ1pioEFKQ5eRJGWDHcvGYf0wGRjww3hLc+
ssA77DxENp20IRwDuU8uqhy2dlFW3TPcIYLAJFNoq0Mi/Ct+sEg+KCV3wxXDN5r7
Zn1ZpnjNXraqcXIxEhsYaTNB0Slv2/cjti3z5MnkWx4ZmQgV4H2TPoDaeq8HiYKv
R7Wxz2SYaKF8CreukRLA/GKb4rbvnanPqeq/sZzS5H1jb+PGwZfmLZeBQ8gNpPay
+6HjFsQ3djmsdQVytum1gPMasts22mU1daQ63wCCmReHRWmK7Vnlp6RS5ruc1waS
sylPeJsJbaP90ustSW68gBEQgdCNyaerd7x5PyHBGcF/IjcpRlj87RBtA+YtXhv1
Svr0q/ppBknFAXNZI8uMd+i0yY+PKmIL/RLy9jaZVfHFVE+7CEpEDxJBJEUcNYdB
eDys7cv1QSS1QhvtxrX4xNW/USF7RkcbD/0NBG+ThuCL8twEM7NB086+ct/k9GkB
itlNAkmpadHyOQqJ1ZS4sXID6XTUB4NXlTst8HgQn4aS+nzU28lnNBDVBPO7EL0R
OzEaIjTwi+RBW3MG8efRshmPFEF4n9dsgYDMUhjcoD9jr7PZrXxyP/Eg6WJkTnpt
S0ja6tCQ0LGLEUgjee5mC4TNR9HrjgwQvGcXrWSSaodWJKpgs3Wy3ju8+EwC6QG9
sU1E0CL2HtwlVF2u+tkC5i7fgxT36AO83KzFZAXTWuv1CF15QuBB+2pqo8F3g3MU
gpgFa9rEp6R+4Abi+I2h9I666oTk74BCz3/rLldOTiFRMCJMAdDyG9nNIp15NXf0
DDMLpKUwKGOi+6PTa0LNNa5LoqzC551+2OJigTBzDTe4YIzyjjPCHDw6ns9E9fPt
/6KypUP1tV3dfDCu7yz6J1xeC1x+lEafI6+jpLAKJkEZEqdDzUXB/o/gEWwMZWIx
BnKklfJm3xKq8RcZzp0cZrD90LcqCjPzMUJx05dze35oGmbLH2k+BPoE+soiqte+
8QfLl1IQl8HAznIjKJnglE/w7EvTEFA6gedNT740xbBTO32D5sw+NHAZhN3A8nwm
nJE64FoPiAX5SPwkosKf2PYUfFZWGk4dKj5NokGXtDhn9c2h1yW5cVIjIKRotFCQ
8zmrKw3WtTyzjBwGP1oTctSPsNmwrgK6qawGJwH2qJqIuLSz/UdrJQSK0NYkaced
idbs2oEUAKrm6IbcK3ajem/5O2oyEdX174xrB8e2af+IMwlRPf1Nad44tD/VeAmA
dpXIr+5wO9EdkpLDuRUbbI5xrMLlvukKg4bFabsuh8w2gzLpHoxJ++E+5vJGG5tQ
OovBR5q4Qk4JFwDkbWHi9uEaTztbMQ6LnRZyKeFU3Z8xFDDFvse9FplInGy3LkO7
NlzUwu+VJDd4FXVvCp98WbBc+25hPHVSLXWQOJ9JoyGo++r9dkLrSGTFq+Lq/u79
fLzg6rrbQUELVmiShuytXtYbLQYeHwuolXCcOL7zlzlaZx9dfPPtBO99kALE2dYH
eDuB52dlkXLRKFMECF35ClNYICM0FP6K62dy1G8kdd3xiirKQp3LQ/2l2C501zOp
R2pffFOwWl6bQlMJ7sp1p8dTefh8TEP6HXj0S9p4sqnjDzW76ypFTodS3b5sRfsx
4eo98l90EwVnOGz5+MkR1RwehT/Ube5oxfJedAWVPzc9DtEV6uwxX20hb5UIGtUn
wR2ypN2dw8A2qI2cdb/Azr42WKw7AYAx814zngpncQT6gKfk8wycmQWIR/Z/D/LD
lMHgbuunBKmVCcggXFyvoTrnt1JGfz0ck9sOn0f41//g5GKFIcGABgliywHxsSNW
P8C0w6Q69UCTCgEhIwx+iWnyM95lbbMNKJi1mBwEihaBp5KHw4ip59e0J6niQxhp
cQ5t6WGgfOQdwkbw+3FYF31Qpzm75MX7AuSv+UMPNAxiJkNAnU+PNV5X0SKHdK98
+oQwSCaVeRLF05zc4YlmlncRreMRYdZp8mY2Yvg3Ih96/pMtFgZvLXj8+5hPCudl
u6FJ8hAMa5vOaBBt9SmF+TplNsm5Z5zi9o3/M0sgqdhHmr3NH5rz7yWNEMcMu2fw
1hy6LuVEiic0FInU7+8VnF3gs+E1vFdXAO11qBD+1f86gKSC1mx/W7RTJ+qreQke
r4znU79JMb/Hk66YM9CYz0yo+EdQxSVSj3g+hNUgwiLju5n+1QmxEWxDGEPom6kt
f2zyEIpulk98TNWjMbK5Ywpt2VMNSTXRSyA2QorJ5vBtKrSKcUB4VariUdI8ytCc
FAI/NQl/QvSgbTmh1iQ8rgiNOOknb2BjDGkt37acqf6HVrD/vn0PbSLcbcydG/At
QrPbBaCCqfR33T95Hy3+Ra8d6nqKbAgqInGqTH4inqy5hSn/DBi5r/iHpDapKyPu
PsbEySrJ9MzjsH6IOvBQ4W0UTyszfx6yBuAZDv2A+VKmIJ9r7FqwIbzktKVn4zRz
k3JTDR6+jk3kRveJ+D5kVAm1d9Oik7ccSxdwMnBMFj8SmCQdv9rUOM9NyzZ14PqA
CSpt5m8EaKrSkc42Yw956r0G1tK7JO9Uw3raqNePLwGsIeQpadmHUMo6rjPQhIW4
DJuNRKQWiqpCvEgS1cub+N8QMjqhaVo4zTmInNrT9tKrKzUbIdYtbIa2Bm4jIOb0
RenACGn13TgCRVCoOd4mBhMTO2PbLfvetJ2hQbvsg1nfA9yG93S564vpq9OVSsxo
WvxAEosOPdRkaaViU8Vdcwttd1lqqboUV6wj7clw1LvuYDJmtXAHXUlXz5yObVyA
ioWm8rWmImo5NuUdrzsUYaZsTVSwj59T8ujNETXHnOk3O9631VlC1jnG1eKR2Nhn
Qs3I2dKAwRQ4jYfGtkwCrARppB1IyjeOxgKZRx6Qkpt8cA/6mVZ2l5fAUpelYygD
n01s6kQI6bO3h5kl9mn7IKcROmgrn2QKAbd/Xy4JjwOLWZiGvZ0hDrj6Q0h42muW
+WQpg9pyF0A2FlHqkAiQl4jQLY0pP9eWoiZUWyNg0g2TMIOBeGu/fbLym3zmjDjm
+OWO0E/k96GNfckPyn6sv7dXZEo5f00eHK23HaJmq812vBSUVGsNxE04CogcXeqo
GniOTO4GDWmVnUeQ9smPsslBVZfQavrlHufk+Gb2dztVSKxrtRuTwfKzCB0bYkj1
rc6ufynyTlhxaec0SxGyUOUa3DPbktpurpgctgP5BJ20qHI/0fT0VFQjGBKqTD5o
r8LIUEGJ/UKl2Nh9ibHS2dbDUg1XMzk+j2PsjYSWTGggH/kY89Z2yiJQxJLxqfQh
TJit3XHFO8v3pBLDeA0dW8t5Ow9KAmR2HhRmEK+8bsvMelT96LVe/vunaufU59iX
MNf9tT5OAowJItsq3V2fzqYhLj0avZ95MQNLyyedDJ9jhAaSnUjauikmoRlwVK3K
aj08zme1aoDBI8f9qLPzTrBlJQL+D+h1/HejLQXDtKYzATam5ZYlHRpcGyRaAN5S
Q+NjVeSeHmiycAu6PTfGCDLJdMCCYcQJ1z5hVlw9Ofusnwe4OZkNNhRD9GNo7s/P
mlN+Bm/J7oadymlHZLk/sSRk3Tj29swUf2IN9XQuFiWcxPVWIEubcnEalqG7D8YP
A08MfNJUaQAfSrbwK1Ff+9/Bon8Lj+76lQExdUeLV63CdheAjaAAviwNqkp28Sh2
KHJkv+/6N454XVb9VfSA8WMV07VGGaAoDI8QxiMVNGpq7azV+MAjrBRz4I+tjO+E
nhqY4+OYFchHMK3zEDrznKmeHAdya/GWwg5+78PKtPA64DUfaiackIcIk6XUxWnt
/R1Z2yueIvq0wFDIHWuM2stlTHjlNfnejLuGw4FFZ3vt6gxjCgh36RfenMdtmafZ
mIhVdCSfoufbgiWOpbTkYpgOr4/dBgL7bfJcMgvHmGF7tzleFRpmK25D8CMRKiqY
4jEbZJseEFXqwZXeRZEPl3qmnFUU+9fMxyIi73h7xUV+EQHmRHmBEHXhxRByvguA
usFDNa25u3WF99KrhcAhdfuSqFl2MLeG0vTb6J2WvP+qwf4G8tU9PuHiogpvIWof
EbSs4F7lM3uIlFfOQDroXvv/VlFLRRzJmHODwtdjvhcaFUZIwu4moIbw0U39k427
CDYBHIZqjxlCiRL0BR+xAbWFgzEuoINX/2sibeiGRS7ZZ2fJEiEZznXVyG5yl3AU
HgPWzuz6lvaJuASDfpOzhDwisklqpZ2pfd+yeB7DnYMWSTG/0mDiYxu4iAJK2vhk
ZwmXcKmJRz+7pXYhw0srp9GmmCZxelKbPZXNW0q/a1gxHDWI4u+FbuF5HSbDthjU
XtPpg/X+5fMn/i8+jLgs3MCAWH5Xz0tLxYjgkSqoYdXZ8s7q7XndWjmRYdmaK4Cr
uKxbja8R1jo4XDMKnAf9FBkaUS+GfyXFzIj7b/2zvnHW/c1ThwLBRaUMMeHS+pTA
4O0ZOCI/n+lRw5x/A8/L5v6dOrjXHx1ep4z0hnj96e+s7kpg2+d0YBkDoXNTcrkv
i2/url8eGLo7jes8Sjd9shPPLH7ozYxS42ul0HNcBsdO5sqbDvrWrxGuiJ+J3HeX
EmwwN7lRCltuvDiEQbaVXkrdlV5/A39DH+mR+JxGjHNb1C1B98uXWKGx5D+acU3z
HhNEDvtcT3XLV6r7Y2O4CuhWmom/mdFMVfriMksDAejAZRnUK/i6FN9xuqRfxuXa
A+J/mBya8lhoscNe+jBVCwlMGMqi1Ncu54Ow7pv0UJzlOCk0M4Vbccbety5kYxSf
l24arv9/OiW6ZTOGhvFXg7yWocBdZCAkP6kBQaE1ARg0lH3qUKvaxmid3jb/6Lj0
7pcWi72XaVNuVT//dI0rcwxeE9xmmXdpvXM4bybXMNWvjYz5MbJJl7iCp6lqIlco
eEtBw3hNpz7N3x7EPAnZdPdfiaT7Bod+8GrDr3bbrf7qJshBYWFPxw2nQsNkBrqV
5KCk9yUojNQVGSFiiqj4WaVLYQmnCrdlHVUzqbDujbjE0uOqQOupYJHpaHTvFD82
TjCis+Uv4nqOFN8iY8p4rb3ODQIdo9BKGgrmtd3HFEtC2X3w6QYgTEh+1uSQjcYC
HMGc4+icAOzmDCOc0YoJtJ+RcufGpCSLYOftXWa3SEwaybuD4hZcKHHLWUD8ChEW
VraXmIhxtAaQ32/KWP2F/8ytERFYMbB/Sz+Ftoqet7sPbvgMa9x9ne1BSMHD7zCY
YEhBDCHdg25M58MRvWGKF8A/lsAVqTI0nisRTSSArVwe4RlSKsFLwb/IM1ka8rf0
qq6AwlgCanqMRnM3Bx7aGBHx7JLB8xlle5iRt557LOPWvESMjPXgJF/7mVMKZJU+
+c/18lGaZ9PsqOgbtOoUqxyemOkcDzRF33OVPAxvaYzjC9h5osf6qAHmoh99IfCD
r0x5lnqiPmH6Jpo7TnQQbdits75t5A9jZ0kCoyQ7CrjgtxbDzqiuTkIbfgWRREg6
mZCGhckQxqbqWxuhGn9nxlvSkPS8rN3ynrlMp+w9GyC79y7pBn6NJTqjS5kdniEG
yrpR2/JnYWMGDd1NGUeT91xn9zmAknEGj1UDXfchL5iXKUfmdQNHBXAxaHMlNogV
MZdL5s9kXf2CKcctY2kRLHTjqdqUGNGK38RkpGkLXPBRQbM+m9v0R9BIFCxl39X8
Ha+r06aabhelFf3E5OGrmIMwBEWWIXIDxiFrPkK9+zdrOpdJNotGjwffXcpkwctd
5phGHThtAUNX8B4HECKYrid/pyFuqzjtXWvwRaFF2O222q5AJ6lryFfYITvUhu/X
OqmOv0XQacBOiJPt6zfeBs7+qEMiYWZb88baQttT0xMwRLf1fz2ELI75n++BOcqs
rznEpellWbRw+Ilv5EsX02R85eHLL/i5H4sJzRiXBMJBtUDnF+cFVIk/mreOfZkF
5Uz5G5WBxbdE9fnAmni7E9bTZ8uicVy66kub9imaI+5qP3WHJnBY6UgKvQiqI7Zt
E6wDHjwhjAjNbL9aDjHaBa7lILJQBREMBHKE499oTyxHHxn/D/mdNdqI7si4Su3+
E6VO6ojTXM/HJY9jTYuRW+63bYlKB46+cd15rac2H/jSvxP+/LEoFxBGeLx+fLxA
exaJb1CDZ5A4Ddx3NoZmnwUaJ8iu55HNnI+IGFmB+6+E9EP2OsM/GyC92q0wgcYC
Bq2kkbrLh0pPb5Jb9SRfzGwMit1X1BYmlzHt8yk7o2mYF4BWoPFGS5ediOguBWIE
1slZ22qFsRWhSwVmq6nRATsha7wEfw1xwNevWbfPRetkydmGkQtgubFKAYm8Nkwg
GN3xpsy/Uo9CU58qMXuZaeGqaYt01QtYs7wv1GZhLdrYXxhQtcuplKshqHoiq6X5
RGHLWUg+sJR3IwkRSyKpvYKwJ4muorF4M+VS+yW02gE77Sne0NxZP92DaUZofHAq
+KU0mGyRu4nWkon+G3St+dzH9wALiLHz7A74zxM0LqF7TNxHozVSnTz5VV4VXgiJ
QlyDK12pRtXITmDm5aUl7dYiqNYjGABLWx4Xk5ciFxEgR4je3o+w4xqoVHqPZ5Gt
rWuOXnbl52IwJPqmYzcjN50Zqeat6woa4Q5XdSOLenVnzchS07L9gfQF4uP0yxAq
S7dfVRCxxUOiTDrsnW8fOKiZ57Wlv4EZYGbl3WZjTYFufYbox1hWl11ixhYxd42+
CnGQfCLg7zJ5LJxHg0wvRwPwj7zlTYVNgPgugzpAIb9Wan41PcAiUG2YdplBN/mv
FWjQtzgj7Ea8w7qIMkK8OKpnQirgVscAxi97nfwwiM4oO5g/ju/H311CK3RvOHMh
DhQBh3uo7WbE3BFS1OGJk62YpbFI4eCikuv3cdAe99LMlxzmm1oiLKAvGX+r2F35
uwX5q/D+/17XBrvgBfHbtl45uLwgCMPq8hWg3JvPcrugKQeVRrF2Ak7ozOwWnMjE
OCMqARtYcPDD1ygv8sjst+ig0LkKx8js7DieYNLik4P9fX13IR+lnt+9saLOJYaW
COJafNwq9Z4elds6P1qGUJIE/T5IcS5odK4Z4GW1BihHqZ6kgXf+0P6AnxRQW5bL
10ZLRMCRY/ZmrcIqcSZUF+CWuPVtAnna6jWP4uRy/2ZS193dfCx68yVBpnFgOfTK
qYUh/Gtk7dKJUf+DXLCH8POqcEPTgjQ/C/hd8wcL/hTAuVZRPpNE4Ilbk1kNB/VM
mgSiql6luBHbAEmX3oRse+1gdHmIfsXr9EZzM9EWnFwLlqWAoP/4gZFdpRDDGhRl
NP3VCrp+AcaZcIIt5op4r4mTHyvraY5k5JcQ6YPp9umNNOWKUtGg2O4HyV+orc6y
xXNtJwO9NPDfFIAOkP6wuHT+CZ3sFhYrjGMV8OK+HqVLahs/IiYpMMc9wKsp1wvE
DcaaygLEJvSm0Gth8fS9SpmD9bV8Kn2F507a/5R7aISRNxN7Cuv+gcyl97+IiZB/
pEpVwwoPpTO8d4xdSYnYE4ENTwN7/lKs61BYMaWyrA9CAGdDoL7BkNMAXAiA9ydv
iKIOWa397XmpGJaBDaZOVDNIiMUcLUFMIlwr4iJWz34KkubKdK87PT/ceuL4N1t5
UwUyaeu/ZYSZ55TaaKFc65oSGGOYHfWSvKTUmRcSjRcuUh6ibrUHpxmcRMwd8ueQ
j0qKuuNj3BtcGBPqBqlG5FIzRugmLZNXokGuCEE3c3W+dy4ihiG3horcFqukz4eB
vWF8haa4y+p9lbswla/qluwHzOYmOVueZwuiKCS3JUpJaPmjvvxcSpKiFhs4o6gK
uqB6wumvjgxi9ARmw96TqxZqzoLd4xDk/AN+YVxfBIUEYzYaIJ3+8wHm93etrBxH
zq26nsoLtHFdAQBZ0rQDW5zhV5hUhq198WAvgy83ksZSjg+Mad88MBqafgxvBC3I
XykTkDLg2pHGi88CJWsZL0CYwEKGyzF0kcLpoHwzmT5F80tvPliv957MUZ0Mdfbu
Lzu5Tx7Ij8XDR03tuRYbZSnTkG9oPAAFqsUK7in3CyomqgAEXuIWTg4NtN81a5Yr
7Zw3kkvhL563ckEUersZ2oZ3W3cFjzfqhMyPMGXyAvEMtvx2cBeIJndzKcD9fQ1Z
pVMtNVxl39J3hXvwEPJuIrnhsmgaOxLEiHuI6dVu2Zs9D/R7HBp0jatPmBokGDWD
Fs8K2btQ3YmeRj1cIWk01GPI48TqNSMdgi0ZtP4Dix8CEJ7u89wK+Od6NhVE5hZo
iy/3wNtEwYzYpRRoTpuHflgknO87nt1S8y5A/EcLLFSEoGihuh8GTDqtE6LTKEiV
M6oPSb26TiY3WW7ciU02mJV0D9xRFnbOTLqCLU2bE/yXamNzRD2SKzgeH/G0YSKJ
VWteJoJ846Ulxt51tmQG7AsUyT8Mu/uJAx2niKcvYGpBuyf1UbzLjza1zxK+2Yo+
SAAyUkXpZ0Br5ed12ZhZQkWMDZnzXujVqpxma5gTfaVfPpDbhy/0Z2JVUt+g29+I
NtA6BMF3PAmqkcKCJX5TeCrDrtrk+djJLso3MrBCVDoB4gK2oGwQ8CyjFsWnGDfk
Wx/pBd+LKdjcjHs6yIzWA1BeHQ4IWSAtYZd6jZhWidV282808M9qNhw++6DIwwRs
XgS7TtIKgkK7TwpBGfwRaeO5KwHXEmso6PDxkQqvaA42b/ylToHPyJjNUTePom9D
DVt60Cmc5UAaV3PO99WvwnTKe04qXovAz3NF4RJ+Fo7c6rWBP02lKghOCwFBwN4u
d2LEPLJfFAFCW4sPHrPkj/85oZYo5wgkxYjAYidGxQ5JrI0twlniuECRrxULvbqO
NDTYYUG+OYNc31e9zX+ENMM+cjflenfLv/y88D+SRNvKunXw2PudbYortRttyOHF
BRP3PyDm2IJLC3eragSmkmy/ZkdjX6KnSEzICHVWSWqTC+ESdpqBIC5qAxFer3XR
efyqPUqUBOdm2cJG0LXESZLdSOTl9pYuLxSJ2+QtfcqGqw5pANaWBW1oHL7Rful5
s9qBi+aO1dGqIC5xlrKMlGORwZHEMLq7Vrz9F0krfduRyvb4NGzu9GVnzIYQhz5A
VIpvB+T7cNk5D/kv3avV2TUk8HlGo6GXzYCGnH3bKGccicmksKvKCY1kjEG1p38s
Mcy2cwxvUeCIX7/nzgEooFLzBpP6ArAbgkk3mWAF/CCL7FLwJsTaeUC9KffcYESy
iMmotY6NG8Tpuro/YdUrXAW2P07wLNdC/XxKW7Cx6o2M3QRCse7bVsF27cacR1Or
w75G9HNRSuswuVZ2ZSWnUkiCfI1Fez7YUwB8flwVaquQki49kLrT1qgYlE+Yb89X
HR6MfiiVTZ8PPAKsNFyLv/lB57XmA9KUi8GmKnPiu9TmJbH1shlCHmekMZ3usxoi
yJcZvP71wD1Oav12Uz5rW5t15iIhXlOSa1t7a2NlJmCd7lNMm8RJQJbAg9FLQPy3
lcwdrNDnZU1TjVIqtojd/8N32USH1nO7z/EwBDOnUOn+EBL/Y116ggmzszmTzkkS
oCTAkwYwgO9vl3j6AKvs/xLoVwE/jSSiSCxxFeYgQYs7LKb98zaGWtnVKr3Ou4YX
mG59KE9zRn272pXdpdpMHMuciKcr8NKAET0kOzojuxyvu2rmMEfY27tB1d36HSqH
A1fFjWqz6pGvGoHVXNHBehu5QqoGPHiLPEfI00Z5uq2Pi6UrPjRJUbcaw08tmm47
zDvvD9GBqU+BZLgTL8fspeU0KmVdK2LjAPnpvmMTsDDOEMX+gdcQPeFl3a69OwRj
aW20UTs5ctxHNtGMOwK24zAgB6gN7R8cOAtCcIAiex+hriaAun3ZwGae609kgzfB
Ti8ycoo22R/2dYfGh8hFUZ2rGC+tVmw7Ylk8yXqmA65TOqGInVLnhEBFK+kEmUHR
e5hWpaHU7ReZA+RNGJq1/qeGzX4XZf+a93jc4FpcvJfP3RC/dkgm9O0F37QMQ28G
OsXb99a5xY5Z1dAYSwxPaFW9l5+z+5UzJgxsIQ/tp5BHJlOisVAD6w4LbkHNcfHU
T+j1WxSV0IdlWYnfoYjOY7pI4A0btte1lZkCOtRvpXT5lZRlhe6oZaYNUX+afTaM
JjAN+w0ExV40+suVIHJSdIgCl6fnoeJwMSmJlJwbetRFjrT5j8sgGWhO2fw7l3yW
NVA+LuDG/Nw9Uknw4bch78mnj3MXITJGxdVv4sFBT4mEjp4kZ0gMJjQg8cPnDfhK
OYFvnGV3qmTyVRciaWSjWsggmdPC2rYyWnwAg/QdH+68IUCpfljJgCZTPsYm1Zvm
H74ytR8QmR5rN44RiEEz9h6aHxBOVnlmqmO6s4oXBtNO/Df0W1l5Mu3vbGz8bV2k
4yf5/TEzBbf+skG4c0pbq95R06RACOPcge8PkYXWiJERsTrAQsb95zUMcefMP0DZ
7i7QkDaY6Nh59mBh3SIJc18L0+8IIv9U9ctZAcfqPlnbZwqrciQVyujM1uqSzmpO
xhYN19a8prytMUrfdSGtjd8ANV78XC8lw+7IQaLCsKtDk2L7lD4PXWYQQt4mzclA
MczYWDZnZ8d4w4jzp/z1cZjY+qCLt+fso8P9DBFasERt49EsapUz6MIYdBWOEFZN
jIYh6D/9UA+3yYoCdSuD7kVKl8R4D9h54w79toCGwY5jUoqWQlqlvQJK1AIZK+sR
lH4uCdemePXk7q6+f96lG6kl/kD4Ol8/jZ8N6aWzoAgKFMAXfAnle7wNiZHabKxm
DhNHqWG5R868pJLw8+EMGE5Wx4qPruFm2creU+Ayz4vSfZtuaKJ5bC/siNZRDFCc
hctgTpGV0vW4UmXo883qzeJ5f9DQWC8gEHXf0jCwLlI9e+kVbaK4JTf5JQJsSZWU
ZodfPssxgGAci5y9YvzsoC2H10ZBNyftxivouRHbkiaNH95AQDQ51H6n7hPuLQVR
q9F11hsADgvggxW2rNkCGSmZPA2uBP2PJ7lPpL47xPyJ8soQ++xUrRT10aCzVWVC
vNDETUsV16tkkasO/ueX9OF4S6W3MUexZ7oP6hgKO3NekIbPbfCW0wkLnlPHHo7v
H+yLrJRsQ3X3Tv2CfSQKTQEM8JhiDowihj7UO9Eu7E4gc1exuL5rF08/NULzlJJJ
znM7e8eNEp3r1vFUDNUunSsPSqOkRT2YwyfKtxSoM3ATHtbjRUnNzEJxwi/PxZ96
/dO3hrvNhRXxB9D/59R5GUJZUZF/rdVkKebHhrjLgTIuDzMQRsaDU5ea1UKMXE+w
C+skn+W8EaUmxG0NLAB6Z0VWfG53Kd2k3QIeMbCwg8/61PoVDqpCSF2xQWcPby12
mrhae6aRWZbHhyBN1mjLX959WmGGmUVH5cUx0DejynXPtTfmJ+UAqe6jLqUfgFY/
iuwyjd9I91+Cjwl0zf7KgnHtxPJ7hJhtlJ2dAksxmqQEHKYYIH2FcY/LZeldM8Oq
dJBpaY3GM4l1ypovVGjKgrblZNZ8Zq3kGwl5N6RZM1ho3Tt55kRkbsP1iNoVnUge
LYeC0guTz6v8/d9Y2WDYaNjC1Mv36PBttMFoJrjZpANd3l2bgEDLaiVfvahqqljL
SWFuixkrPy8gJlNKUPmbY3mSxaOKLyRKCQ3n1ocgEoAhQEhhKkTgl4FNRmecvjAd
a5uPKu7TFmqXE1G7cNCsvXBo2C+wi+Qy6eu6B+9jW+bvkL+kNBI9ooP6T+Gis+iF
qsSkBnrhWDOYb2Pl5khFJtMuTam+gP5jtnTl9yW6gaLChZr0aZExC+lnKDvg/s+g
mlpdtIz5C6wh2JGRDM9EZuYBlZbs2HYgt3X4CrPQj00LL/mPlB2AKnkJjH8uKeIX
nEPF4x1sGLwJaqqHliIz59OxNhjrLD8HkGe4H+aBa37Cw7NvEWi2iUh/QDZ8/LXK
QBk19Y3DlFsAwEYwgXYAE4PtT4WVmKXyKRAxtc3wgbMA0jvXLkJiPb48JiIc5Uag
v1Kw1pHbVrkG+3S8fAUtEFjidI2TOnN71V0c2bpHW8lVj0O7m/amCzTsBBUjglAk
8Tkq717coP2vJleWtUTqss+pIqqzeysBjp83GBCU2HaHCf5Q9MdXI5yhD13fjkR/
bnjg0SZL/kA1MfYlL8iY94PPi05OXpyNZ9qCbt7j4KqlFAzZgRPfX/REdmgMCdZL
y5hsYde3/3xEONfBgvbBv4ohO+ZEBlygYB5flNW3qN2JGw5g0ZCMoMKZSxuJ4CRK
OYaJosLBzOvR2I24Bf4ydY20LRYCls1006irqPaW05Gg54Wr9joplE43najfSouM
EGj0CposncF2PnW9mJaBdyrwQEZazefr0CPm0+cXHkp25YbwCxIQHaxz7ZVnG1xO
4j+hEVaxT6Cl4Fuimvv0+JxDUbBxs1xvtdkbVIS7aEPNsZQOF2sMW+Ol9DQid1gN
W+OaWnX9zeFHQtsC8j9Ee9EQVKny9P3PRVeRv6KeIx/FTI7nLTW4fYKF4DtJ8eVA
x2GmcRJs0uyMbbFLmJcNXczfG5PH+wsigIATcsXtNKOp6zlvKBoOrC1q5sapDjmL
EY3ejH2cN58MrlS0Zg8ChRiTHkwFeugIz9l6icPXdhguf2OIz1g1UtvtA1j6lvBS
p2tEwRXrXaj3MucaYlT1bxtVN3e5oC3Qb6rd6yJOSEhZfNeNCA/P9o2KXUu2Kapf
hJvI3Mp0LYshv4yqMqq8sJpBbYYCCaZsCjXX/Nm0P7/deeSQBmUd8zuW4h7NvEJv
Nxeun9Gm6LnwagjPPuikxm255HcSkwm6QrnA6blevHp3+3+2h/9qVfwiOFcCEjbp
g17G7uU6eLQ7g+GwxCELauq3xfceCVMQzW0j+n/zDs4sz8un1/0zaAtAEXE9OF4N
6//A/2nQG22iFrz88EhC0eksIICOYSQVPp4IgBKUNFhtequzqxGPXQF9Z3lvqEaA
nuWN/CkhRMpPnolYxTDufu4TzHhDkOfYt+0ZhAR18e8+G60AY3VjXbgzB3+F2ktO
lsl29Wp4LaxIVjt09Hn2SLJyboFlfvIfr9LaQr726jq/Grw43E7JirsehGTx4XdM
6UthbuvXvl2dOY1aBAZ2zJeAUJAisKZwZinCuvtZ8CeZVk8d8xPTWfpzTcHXC/ov
VCDZDMgxTtNIw9kMjSBqYDr5PA40V48rc2CSOwpPs7WkTJRobxmQkW+p84GotG08
0TMxpRem89QX945jxlt3NgMr4Yk9Xyqy5meHScfWM8K3pA1ph8VmEWHobAjLFq8i
p1DFEvB0LRJQlppMOJfGf1lMPUbh579Pm2IH2lukvdA2AImzuX/TN5Bm1h05oL3r
iKOGnDCVq50Jd/OptUdIocUUeiMEIDSr+g5vs5CaPUOh9gl8Qn3ONSWWVIfmZ8Pr
vtN8qZNAGeKsZvpWKyG+2A5s6Qef6Xrrg1OYBk304pA2B2P1tjBf9bsVXKvntZb7
565MrhdidjpJpMihbrurdMzk1t5C1guO//EWDOxVq6Fv3a53U0gIW8vJ+iW7cmcl
Vb7BGu7jfRNwpnYJgEJxLPufanEsKt/iPkurstPeJRZmgiuhBjDzAixbWSRPs9hv
chJ/yOLJQSQmj/EMahmx8gDSZpfktz2jYP9hPrEIfLBaN8OylcP8MtWVRg0XJwv5
OBYjFKV/4nkrnmZDHRWwkN/+WwaE3RhYkth70o24MzyhO7HnuNWayerFJ1A1rjYm
aZymep/zTC3laVutmI1fKYZOAMDGakcByoUMT9RKt5MVMnLMNppKRDTMkccMlx4N
gnBMUgdi5QHSuk4ISXz66LM185bCRX/AICwFLtHqymvfg5s3chNezbudesnbWiNd
WyehdM1HF+AVNnovlKelcFF/ClDM6KFuC00HsMvnPOuoo0FPxjvGugJhDufoLmD/
A9pKSs37OGPsmbZreP1US6EBfoqCiKY/hGsI8y6piLBmDRJkW5MMkBpFTuObJFHL
8dnDpP0ShQ24JC5rmn12ROlZ1rQsQfpHmbHSV5tOlJv09pcUMPCbV3WTHvjo+jeB
WyrGSNG+oCrelTN6ee1Yp+4UPelf70+33V2pPphSUq2UIf0zKCKoGqkBNiWRZ31x
qTff6xF9SKGu3+L13ESDWNoAzfVvLeE0W1NasXz3m/5FxLR4YZRYg2gEGhph5sP1
YARPCEy2uyivmPozPLHMxRS0uRnOKgJ/NCQuNJrX8tz3qvs5pd52NLmW1hjwLn0L
UXzTREnL2A9d/nNXUPio2trAw/j6T8CikpAcyUiJE/JaRePDQOhNwiubYdRavdHO
7pYOffbR/Pv2XTmiW1rbIxztn+POuC2VOFKoerd7UytRU5f13g9Z+hdjia7Mlv4p
NN+EQ/j/5jSTZ/rZQgMsezk98ZpU103x+FeFax96Zw7MIRIY1ZRXFj/1KRoYvvIr
uelh7iWBuCKaOmHA2GP3NKdyiw1bon+EeYeoJMbjSJyxhkAaPkQjbGgzxBQm/Lr+
oIcy26Ruc2+fcxTLza6qzFjd4V4TDTs4fvil5PG3XjWghQzMNsgUCw2nGPPBlHFd
ouiHKMtmI46BFdiH1+cxEor1fKYHu/FWN+E3rMWmK9QwZcdWOAQ+7ivGsczNW119
8KmiX+SJPGIewhL5vu5895ZuV7ppKi02oBvAf/PmhGxbL7EdPdvPybKJp/dhiXpM
tuhMHIRbAd+LXUVc5ytBDCyivvQa1civLKuYdYQu+uLmT6BWVSEG6T8yI3PhKRIN
CHS29PS6t4N1pm71NgKXxBNNjZcCb+oi1e+/PWsISqSvpXweEGcUWhy4FOeVUJYo
Lj9UuP6s+oVLfXA5ZyliK+IfvQCDkOae7DTSGs4zJPVNVuIgijKsAAWgdrTxKs8v
Wx6OaS6PFffAjqMYZDxjl8o+hNiBgPuLSzqaaVz9nyN4n0/L/dew248wux0FftoJ
qc3N75pBhRs79VGs8gF7LzHfL4DOiHAMALy74JYf44TZdPm3gcPrWySaVBmshsuY
45oSR0mVnjoVgOhV0snC7U/6Q9iTpuYXLCWLoFSowhSeFNhGaHHngeXb5lNAhkgO
TD4Jkrv2OAecFRRH4ILGGjIiI41GJS9Hl2LdTbC576nZ9vtOM7JN783Le/mKzqCV
/bAixhWIQMca+dOnLPaD77aYxYgdg7+mBVtNs/uKTneqeDq495rVny2deXwJjf3t
QCFeSyxJ1odcxJfg1Z0a8B0jQxJm5bu6l1+uH5ifYoDL0INiOOr4+EeuP79U+zse
cDErcJTNJGtiq2AMnr00Y3mh++Km1lgzTk7eF4PxeUpNdulM4W4Ljwj/YXKeHn4u
jsQORlciTQeGgieoHzOurglP91yHuNjVP9O1EfFlc7u8xflg2dZUA5EugxPyp6vL
SC91da2TPCbwcgkm8Ay5jYankY865CjARNOeDS/lnyryYMCp8XFC1rwnz2+iAz/W
T4gyigF2rk0GHOqD7AyRAiMWoPkUhyh45UH3nkD36fD8FFKrBy1zcHO3eBC3spWt
cLjcczx845ub45HEEB9n5S+CRhcss2U/O8v4Z0fFr1YLuEsPWaQKDOioQKyykrJz
JSJxKIZ8i3NPNjO2lk7nYgKqICEKSAk0LAAr1yZxm3Bzg8U0tvdhIYDdYtv9RRGL
zLKOlp6AMT6SaJfcT+EmZnUGFkUVxoNN+z+/AXJK+Tl/HEifPUXUCC0hczXMb81W
O4h/SLNedUIrHsobaXEhJpkX8BNjtTzoOqXt6F/15OjAMetz9b0I76JNzWuUo0kX
PytmNfJQcmueBFDuj7HC1FVNvcRbf1x3pLE049GxsOU9CPlfoHeijgezpPmQtqaU
p1adEpBPdp4teNn8VXW2iyKMmx/61WYtXsgcgiB02ipeMfsPjA00b7lIfSG6MRRQ
6VNkbV2nU7PJ/mfzUGl9ms7GT4oF+DnyHXsVJMapvvrzyQkQ5JG65EJOUE+vjTO2
AJkf6AOMX7Wh0c6RLQwD39FXUPo3kI126NCVfOYvyFbP5YYT1TZtUmWnNf2lbADN
VtM/ZKqgV+L6Ajes58KJaIg09PKnbHKAsYGxUjfjB6a85yqdQBHi9QYZyH44WEn/
bDyDpEJHOiw7vZyUaAyvUB3m072vgTUeNQEtYQTpQYYHyxSNxHHRXkBCkYqN64bv
jteqV8KndBMVm2T5riR2ZXMN7GP23Q9cbXgWVxGq0Pb00mgKMHor80wzekH1Dxxz
4yA4hMmjCQUjR9dj711yirzCE2p94Au/A48VFUgXzyJJCDW7RnTp5qFBYZLKqVVp
6LNcpLLdRCc7s6BadpLCh7I24FNO7Off6XR2PHHrPw2oythoFJN8JCQKKMRn1A+K
6nYV7HzrthS+724RrryJyS0qClv7bH4z0rI7kf0iCuqz0wD/IusKjfM89AtYzV3z
o5tOLObaY1DfwQYkcIxSxqaymq19naunP61m8FzzgMAI1TIABChCaG1kuW7yYUix
085Zd25yE1JywL43Gsf/yB2WHbSGbNM7Lz7wxmf8gr4Rh6RcubyWTm250oG5CPhu
62u8o2ubjDB7ay6DXPhlVjCMeb7/IxKDWX+KsigmJh6AQj0W5Qty6Ru+cMGnhCmj
XzkvKoMFgFtwiG0hcX2efk5QILe0fMiiCOoDtQEHaSOj6o7quymGlN32PlHvIs6S
LjaFnYOG9AYSXj2jfddVswseTRrHQw4nZ0jOV6M+MMAjhckGLxzvk/HzimCJ5Ydz
pskuy0jMYajHFRpM9CLQBHkimdLqsvoZlBHQ99O2RdTak+/s/Use65P1sVrBTNtS
BbuHnmtvcQSu6xnpXeeSXundy70lJZDiHq9RJsqNCs34kZ9qG1evu889HUJdT7E4
Y/IDSIl7BGzeTpvkCDqPtsw3jIoUIqhwDGxMDLOcZLlmoH9iEG8kSJWX4F5o07TW
N1u7dUITKB/lJetpE0roOou8GQnVzP8AfRnsPNXiG+7wpmv+TSoNn/GuGbqfMtZh
Pyksv3RyNwWBMmdMvrolQg/bknD2QW0ctIz30tA0e5DWRNrG49LNCHbSZW2FuDoh
/+WTF4/5lqgS5oTGS4E1UUG0g+5O/vMptflZNMuLZggXSPU80gKZFfvPGjIMQqxK
b2lcVRa/M7tV+JExFOBusuP033ep9pxXhATqC7H5+eX7+JMvJYkpTKcSgXdOUnCP
Sj13TRVv5SebpwyXf93EM5M3ttlDwPVguavvBz0XJQCp//mEmLXBU1UcW1PKy6H0
rj/xZzgBw7NK1msktGQXr7w1huzubOaUiuKJ3o9EBKSHG3BpQWJecV27soqLdpYt
yLyx7IP4sRY5SCE37ukso2JzjvAYqrLzdAM4A8LVHNTVY+cvza8pmE8Y+axhQOXO
+oG33Y0/REmeomE+PBqk5g7XMtbaeJ2cXi9rZehN2U8+XM7zTEVfCl9ryqX9tqQb
kCkJakzvtI5POiVX/nuxL2mpfOku3objq/3ncCwEw7xig/WduA6CkV1nohqVJwKB
Rj43s4p+PBfFwDQOFSbNYWK/8OEZeTUPQbFWtQuMYVCfTV0RyoL1Vdm04v0KyooR
EDmAe0XxC5H+uWhLtUVxFvmWr5+paB6RGsv3zI5RHJm/SeizUphSijj3x2f/hWDe
77HG4NKOg7QZ641uyNolEmBcQ+gbpTvgr8rFhrcHEKWVWnYBSGT6wjMsJSFX3gdz
t2uCVYKewJFn0s/y/DoLf6GxfMp4qTJdeIz5nvgiz6nxE9KujEAXUecHiZApKzKo
5wgP5MzbIdWPSE882AT1mSoI+NNHGwyoDV7oceWRyTU63q2gXE7D/bPDbl5H7xGg
0JG824P29CdBPUvm0Wg5IA0YzWu4wXUtgX8nYi3aOv5felmg2vWMl4QdCXBnJc+W
vpklXwXFLpPXvLT2phRfwfRr8XGEhWOttmEZmYVH6NlgVTZiz1vqhLmYxPTRRD6A
mHvkLJzoVSmWZlHr3VH9GyTAXpXZXqUDiE/6hod2bztAuc2BmTaFmdi/jOZpLeU8
WrNZ/N/5v6vc+7PTopyWRLnmPWh2J2k8kY3Bl2yclur5rRSG8zEfLjceAFtaAnrK
MuLnN88Ra5HUQ0k8SUbsmZ5QXWgd3yKcYqz/bgFP2ZVsxfk6kBMik/qy+jFgHdc4
IeBvUZ/NGfEIyCLHNO2yHt8Hy4sFPRIl1LbvXauoakn6nF828SfcmyFTFZ8FHxym
4932ZVlxn/Ee7Krsp7J68+CdD7o8BaqBsv292rfkeo4CQqYRY/J0Ebr8MOhpjF5A
dQ+9yFor14Vw4EciOBR56Mc16JHIiQEJEqQJL8Gto6Ym6GxC2jIAPp9F7nGNa7TE
B2jBxXtE+MaWo1H9vKdyjiGQ7LLx8EblM9PHVrgT2G6SoubNVnPFyJ29w20EJGSD
imC9hY9odvO1e+sHLngjreWbNxmAvp+5wspg8YOkBA7nHFv9jgbKNuBP4gL/ErRH
7CKQ734LzDvRPnk5wgPCxqPrt2s/xim24Ncpw6eR/Zh30fQkFjmydko7CyP2C/WE
AXE6W2MlEi5yhqzhyVcxX0NAV5f8k3tNTtGmFJ/Lg47CVDDDz8lKP1jIR8HEoxcF
90KRClH8qJZogz0doM4LLvx029eKi9mm5Als3ZHseDZJvWb6L1JyBwp7MZUVze95
zG+AMIPcNkcecxwvDTUKvJ4dZQyaL8HDvH2JOA9pzkDlGFTzD6HRpobjvmSOjAAj
d08Maty7Gsa5n75GRweCtJQ3T0ZFbXaRdOu8pWzcO9Vb7c9RNSe+P7Xx0Fed3ye5
DIwd6k4bwWRueNwFzbcbwL7DKjl7JB+z98KQ7Q/hrsm2/E3rvFeUDcasfPIZkgw5
qMsUpqIGfN8KKXYC8ti0UxRFvSdJpsxxYhyz/5+bLWs4t2xLbpd1HDcNrYBnhroJ
TROr4CBTa2/tuWlbth5bGuYgjZ2SycCgHd8mugtGbwD4rXr1uhpaF4bLU+MrIeRC
zpC4nIMXDn9fogAeN6G3HXLlXdIcSJx3C9KcCTjsjGjenAqkH0ZLM6xSR8Sw6/ic
lXLhbLh4VXjwbRUzQHONCaduAOXl40xtrBLPtedX1vcmVoAoO+evAWFeNdr5Rk11
2kApsgIlZZ1tfUPNuOIuam2Ig2tP3DJNDh5GYcpArY0CV+BZY2505DJdnYxGmSZl
MWqu1eFKzeR0vCkZZld9wcciZwD5uEp/d3ag++DE+Gn69MjNx+umcxTyeJguaQoP
Kc5JF/qOXVuM1EyGvTjYvnOixzLdGm2oyj9JFU5uvAd4DN+HyZuBvqeJ6YAsKxiM
Vzm2fwzVyrCV6GNhyEbSC+wqQd0sYRyfYPr2oS6XAg6Xrgg66dZHN5ltf88/Ciaf
lDbgRuJlBUPqWzg7SMjbwLA/6n0KzvzgV3Z1EDsUZYL5c3MNieRzlhwhyN19ZK0j
zcgWyn6p5A7K0//EHuqUjlSF5IBettgseu6j3H50LVDrYKRfIdsl2VS2LSiiKri/
uxrQdYizpKFiQisMQJbDpUVW5MEZ/IL206Zy/y7hZpjmsNrTjSzXOmUPCyLASkeB
SUXf5ms4K6tej5SdjwnuCS6fF7wE3LMyJK+T3+b+j5C3lyDuIeViMTfG3vjpCvZH
1SMf+1JfDrgS8gKw8QyOfgNQ4b7LB8kvgiPi5hBlP3ZDmI9kS/D8AF/bihd68v95
a2QVlHLxxa0On1SBVCawBhtg6tCUDsDSPqYj20gBJYay3XjOn+c4KnX0zyYsn7oa
F3QQtL69xNR22mET++c0FnnaqSztEdyM5hQa72osocZOHczH8qUOA4wmaCzWGs/e
FEJaaOuAq8ozfDto+lusOoi7wPbu0Gaf3TQSI/1pB7UWlZiDwCiUf7jTm0wPe8ni
xF+TcnjR9R+qIvY/7JzvMRqQn5A81f/6rAr5kQYIdw/hZOX7VWO8vSCmlM90rJap
CdL6WbAy4t9hzAEQj/YRu1azas6DrgNXkbtKvvxfT5iwVoB26ROSsn+bVnY3wfUM
aoKBziFvZbOm3aS9K+HFqr3+Cxs8Rz40sr6LJNVR8Xb/9AeW8pQRn9VV7gWb3bJQ
QS0BaIe8rzdDdOoeQugdrITogoDnYY7xwuR6e0UdfwTRA1EAyBUFLIDGvQgRtKD3
n9O6WJ0+MI7E7BFDahWTFQeI9b+Kq0T5FgAiFsvcpxzRU4pATZDvXVYG5Stfa+2j
54A2C49H8GimYf5i78RNbkGwizpgmSMVZr7wxeZ0uxwqbzNLSCbL4Q+oyNT67tHl
6ojyI1CEykuSQFVdmZe3rIoTSnbr093/LFj2LfQYYMNkbiRogz5+ivqCZVJpRJlW
7rvX6wfKSI7rEMp8FRepFRw1Wpk0VkznMWrup3OnpcEzHBTk1ds+a2LUDVOXFgOY
Ds+n9yj0hT0CmlNFPDxTTxQWSMwMr8fvviySvRmnDOL/IQYjyMUv7OyPSWwF+Z4v
4Zz5WPSLtOoG3YlV7KXeBqJpz6de6q8FG7Z/Z2nINc/0d8bjNa7OAy2fu87fJK7K
FsAAocb39Qhd+BjP9yhpGt+hTvT3qPqLJ4tdbLyfAevanxxAxmSOdolhaHZUyJJb
SNs4emrESpVv2IO3RNGsNYKrxllkipLGTnUGeTf0C1i0uTaOm3Dl6V8UtgiF0/vf
sKSWMZ+2zWjS1ki7ASqHgIh6RihDgvOJFOCZtknB0CK/Kg+u9dz+G6Wl5bEUCxj5
evYriXg7HhsWCAK1pzfF7Q02Bai4RAgoflVIFh14nqX+XU+G1ztOMJIhaoqy2MQJ
hA5rzg9NcwTWMSR0ccXKkOJ4YR44QtFpa8Q58LY2/yCDcw77NWL081EyIrLh+k0A
o3gXcz88Unr6wvam/nhHZ4NfAamPucs8fK62o0g+T2HUg+hiokaqRrcREtmGNYAP
hveGagxwT8uhXp8f+8usQ8vTB18Ut+YFJFQCugXhIpdM3HB22eGt2UBFQGy+PaMN
rI2uW/Vx9HRkrG9IqTwrcSaMrq6Z+0mkrPP7nGGblf4m5gDRJ3QFC5Kypxz78dNi
fxNYWXNI7ehT7aK2jD9BQERHh2abTV1iRJgPSojsePvsF+AXQOKwBekeMKR+2APE
y6nRJmW+QkQdencrXHvDv1sGO1tRluwMetQ2n8IGP2gVwgpdYSYYVf35AHE8xM0l
L23oxzdvBZczpTvMmjhsM1OzrLZn/H+N0LXouaDQ2zRlLCUzMyscCgPWx2S3zkr/
nhOELN556GYMiK1iYftw+Zm6bgxRTMaENUSmYb3HcC3q+ZYMcwyrBibonVw9Ph7P
KjjkByDf26huWTC1+GVoZUsr4z7r/5GAzpzj6W8ENLct0l/E5L/UMQJCQcad1bVB
tg5m+k8GQTyvWsOUe0Jxxn1X1/1HS90+2PNP1omSSfK5MmixE8EiE1zMt6kI1QgL
1hoaIBQhtdIMrxG0/GTG/CQOzu8R4hL8q65meu2XEr6zF0S9vsIAB64H2Jh5Otls
2kieGlfydzyt5MBsymqvBdr67bVsHg/ZawrpxnZA500AXGLwnFvN0s8izLtpomtd
kjoA8YHbtnFx0CYmDEv361eOPlftTkbo1mkubl0izltETy/YB++ngPVmQ8pig4ko
AX3+p2I+hsDSFo+xDQNLqWYVRx2NAm6KowXvThDzkKPXDn5DRAdcdUsVN+mWJOae
njs4Yk+WYcdPX2DlZFc30qKWk59KQVNWFlKLhVBSjCyV8RqsaqHmWOguFj7plWkT
+WN2hmiOz5I/q6pc3GiLR+uQdsx5LrzI/qTgWMX5UCccfsbc+O5Y4V6NTzCBBzOZ
8zdcIhhVFHWdPZbArdSlrdSTlbEH1JypFe4TxZEqWYgOQlv03VM1RN80/P8O71KI
bhTM7vwmipToIur3PZs6ySXllKToyIWhBc56yoVzDRvbjcsEnxcb0SqEmOMGPSok
mruAmPJv/+y4USQ8CnReA9D6TEmY2pT5Shz5/2soTYQwn983qs45af7kg/Dgwnd3
MItV6cZ+ABxBdrXLaLxDSe+BK8MXmp3DMA/p0xRMUdzx+y/Omq2XkGsbrgh68n+U
8AE4WkvdUEfGcXgxp0MFaMzNrDv0YkD00H5kq3JRhLhmXGVEk9cdPvIJli4+X0k7
/gi0Zt0ZnIp2vE/X/HtiNoGicxJ8xMzb3COSfpGbOyzK4cSxpBJ1ZkuHlquTCUyZ
KA0RMGSlCl5fMwnX0epGBRAC3a0zT/L5iQJ726C+2BjKUM94G3RQ4Re5sSHGLyla
moHaiOm5EkuXw9ue7udSvKSNayIPY6OfL75qXg0DY+B7SL8b4mAQfr8oxJiAdgZQ
X0hI997dR5BLVoTQzlkWUG1gTiRNUy0cPTVHUGRJBp5a3mmI+/yfsDoUOyzrUtOH
XGsEN/3AMZA9R0x/5cB6apks7MRViOX5BIeA/wFpp/oc2bxjThHa71uQMczVXU/e
o/FLOlgLvJilW27VCIBfP49zKp+h6Jfz53/n1IrWQqx/bgV4ZT9WeFIrgXthLAyq
u35hJ3kS44hE0tXJ/v3TprZEbHuSWgDxeZsCQQRmfk3VtDW+g8TLfKGHx5iVUVvl
hpqEEo8rJKy9G5WnZmMKmtOhvVLKrT5LGNnVQvzvyC3bibuCArvpQ+Na97AzxoPX
BqASBT1/2dn1SzlepfE4xNHHs9ADZLKsovUca85meLlugwNj8BqNqGV6RZuR9jsM
bP8zx+Wiqy2M8Y48eQNSjK4ZZPbFQrcDVIS6YULOGnxznkzFQMl0gfMnIl53bhaH
QP2hEjmcic5pGPvV/tN8DPjUjI+F/T2gLbSLND2PdgAFHBlfthAkOY4f1Pu+tZYc
2Kn2LURAGNN2t28xq6x60glwsm6lqygL0X9FL7zBs85wp9Q0PZUt2H6F1zfW/jiR
Pn8VlaT36S7y1+M1wDOwaNsegUyEP7FWKRH6C0BHkJEvyHLqWcJNgEASBO98Dxu5
cY8zTtPCzXBortlUGkv3850zf4cvqObtaHCGx6XG08m3g388naJJxYhDxlK6Ntj+
o5jHfeAtQSYgDk7eElQ2Zk3XrYzg0VmAtNar/ksayRSGhIhaNkt2GTGRl9dOj6nO
znelC/9RP90OUu6r4smDA/klqOE1NIvX3JgN+PaAlvQwIkFykcFUtJn8oaTaRe0v
VAlR34zGPTDmZhbz0AjvrMRjMXixwPMvorvYMTKHq1w4Scl/FDpGj72rQTAyOfsI
xhGra3rndrg0+AoGZdSfmOnpNYfjmbnwSwXy8TA2iTgPmGKU0E778XyoTWwcLQPL
QUoUHNcnlr8z/K7lmeyrJqzYoeYgARhURyzakoeCob/t7wblM52n8Z0zkt8bjcNW
R8coIdRx3PJACs4ZSol2udhNz0fkpHrV6FI8mOYQWEKOa6kSeV7e/ktwQjkzoNS2
4lsj2V5Vr8vWY+WpKacSHOaegkAif7+qG8pW1+vK6vIQDv0Jt9KIV0qQuJVbiX5u
S2jqYura6/8083rbG/C7AY2RCpU7w4XHXCrL51TtLU4nvsU5T18CCP69F22NXsuG
xBV0+ksolir+g74Uw0xaSOW+W6eFaZhjBlyN/n2JdcttWAOPq+nPa6g7xcl0wVg4
hy1wc6il6xp2blXV5ViF0Cqv+2qZCBlR0oWs9N3+qlRYGq3c4Qr8vpRVzHS4OT61
D4vRSDd6G1+ZdoljLNWVfQrB1aTx3AkCE/gvjIwatLlrb2hjZzoPx41ldKkyhFam
u55p8D0Bi+agcRuv8lN2NFHYaRVu5MX43fhaPghp/NNydS6ArE7vBI9IJGERlQQw
lamgA90zYjBcz7TONKinhfEBVNL/JOkAIWvVdQ+piN1XTAu6OnWegVknQFvFpsPg
qUbASNm9jDOWsfrto6JAaydNyQ9vDbmjrQYj3YkE0++6o6sXiK6WCJzMfSf6Gm+g
fO6kdIQpORQnNviYKQKAMJUkvAblHXqMXQO93Ju4In77+dYuv9H839vAswGqJddB
FL2ZEK0E62QEHlWPguP4yGe4ib87uh7JsPcU2J43+aWoXWekQ1ti55eXT6Cyfbap
XvsAiTSstlg2VRZ0/eyQVTc09CadC8AHapuk5pvGEFR2pXfD5zmc7+uHpoIBLNKm
sa6YFAAt4kizFIaxhYvFeOsH3BRCRMkXxcT+wjhH/svUlhsKfFyZ7MnUw8zCX26Z
nhmgq+eJQHy26kZvlAy/zelZHQW4D6XjAXRrqYNmuthLXQgl3qx545+3Xx5Sjzb7
BtsYuTT5SM/Ym15h2mzRsAWQsiOMmc+ZnLD9h+LeJOVci+lbxVfSaNTk/Bp+aep5
R7eMUdbWu64gah0CwRYeH84QSGSU20maheWrv5WVm0m0/Kk2fR9j8XBW0Wff6/qN
Ln5FZ3OiErUIb6bqnnM2k1YrbyoLRt13GN0o6xdYhGDaaq6/4h53kHydtcFkbXNA
KlUR8Y9A3aazKuh5y5Be5p8FpSs9pg7f+MU4J/M5xaT4HPflxhE67AgkylL9rUr4
z6Ku1O26eQ/pe1UpZ2z1oWmoh6BZg2lnwuLyhKlD5+2r/XNGO7qmAba6bJQ3WLMb
4BSWlVmRaEvIuiu5aS9L9gEUhCIqU6VQGHC083KQJ/5dHjZ7ynEFRHppPUaU6Ua6
NsUfFJPYuhqqqkbfUjtZmu6eMVOpPzrw9ywACFDXduGfSm0DR4sCEV0YP2q8pXbQ
XfOdJaUWae/nnjCRZcQhDkT+b3/J7OJM3qllGLPxlApl30j1oF34mnEHFUYARHVZ
9vQ9B3ZGA6DJB95QI+XmtCxUQ2MxpNjHeJp+jYdrC21Ss8yQSstOf6u3vtGH2Mkh
xIDmHJv1LX00UepC6BihwPK7LF8gjNlkvGij7Yg+07xublidkzrb2G/S5LhQpjiz
U++52tR0xkPUal6cYZaPQ0kc/08e5QRqacM8c2Bnm9dn7JLaV0YhbVgHMgrKJeDR
wVChvFxOghFAj6yHquykQVqDu0JpEZYtCYtuXaLF8jSlkO2qys8dDGAoj4Ty4vxZ
YW9dLauMDVMaAYNsxOOyDA5c7sqxsNRr+WBJBEdmTvC6BabtEkq3BtSF4knrF5d4
x/mBg27rm/hfxlVNf07sQZ6E3YYLh5FRCigOqy/BGb8c9EBrjkWUkUSvqmYHCHj0
aD5xoJS1TB/+Pv7OB4T9txvk5TibdHkz+S7yjQwqEWFVMwuyiTQJdV2Olu7+RlF8
mORZzjh9LzwRiLjS9JvdHqBr0wgG4fv4VoU7CRJo3nkTP6TtUvXJEhQFMZ2MgGJa
TG+6rZ0pBhQNXu215aa831UB3tg9hsW/oLt+OFNS4w++C4kqhyfpKJq8MFpiHPGS
s/33cT2mylflZmUNjGPWxo+uekycWOCqBscCGh87hMV3r/RBEgKmbkH2r8tGoGSS
PHhXAoJ823/4liHaVSJYWgtkVvzEpPSDCK3NcncJ6StDBZ0u0brdKkh3+kgiGpIK
LqZcJ66nXcWxbueqZq+FOwaA12U0aBawGzdqJmbXR17Uq4wyMfl2UIoQsN01324n
uyaHRF/WRBqseE5S3kutRlsZADMbmq8goS6tRW0K9ra5gzD6tkcmJmGqvOBygiy+
cqOTwrlYwKwF3UHFxeXIb2rxK2MMxlQT3KIAUeHKeHBBAxeFfe/W6xqUWCJcEHod
ULt59Zcnb7jkQKYFmKjAGPb6N7DMpWUehbR981t9WNiWcInRZxzKG2xEqmfUhssr
EPx0DFXNOLhuvbA9cSjCaiK4CVNc2TZ1rrVEbH8kGLocKyEHE15pmg/X3uGyUxQV
yS8UmNgxHw9z7f1ETanSlxZUo0N9lGOTqzRJ/BgoJFqU7MZ9A8a/ZqR7hJRxGJk1
bbE274XC6FKorouYyg4TuV/QUQ6be8e4Eb1HIMtx7SiQ4VkdwyvgdHpWqlfZWZar
GNRLpSq9PfFXPB1JB7B54H9Zzd7VarsI596pslM8qbmb+lzd5yqwgSkM+hZrtrwo
k4TRrWNV48NvTDpm9io0bAr1U/0SDGOdcDca+Hm7pFKxrFw7uz2nMUXpvY7nUyhy
zTk2ynh0hGWxYYet6OMOpw0WZgQYjL99B2cPz8PMUe8QblxKxUrKf6JTyVfB93cC
kf9ajrjl484iLwY7kNLmVZnU7zD7uvIjsm8TCoOZekZErPrbVWKIxpOEPVGi2owT
xJg6IFTvK+ZeTJzBpVZFoBzf7KCszWF4IBGP8+M3/mM6iVUiGfanjHcUlKaAP576
ycfXwQBWvV3bUbsZDszmSasaO0YN7Ov/wmAiSNaGytJU7dXpc8Z591tl77LzPjZU
IK3Iz87vU3/gQqF0TGY6Wt10giAV4f5xzL8MCJTN59dY845exznhrj2F8fqsSq+/
HtyGiAPTIvkorkllzu8hMFLcT0YZcCXeI5zpsPKuJu6eE9cG6oN3yA/cbgPN6s7z
Fpyh9Zs66gzJOQaSwVxBNsbvq1GQJVRcvIP9pPKsRJnd6DAm9Vh1V07lB8eZzboh
EJXTguPf1OlGpzlJgES7AO+YuAsbgV+qr1sXh1sP4QvAPG7L2R72D91sCPHRvwQ1
zn90rO2Vp5Y9945HLFkWa00nk1Q33c/RB4w779P6eOQapdTRtOnRjHuvL7fJ0fGG
HYD97SuE8E9qiW6j3yEES88btmXoC2pWIsu2lnnU9K77YJGAufBJkXZzSqSo4HKr
rwYMl4zOORFRX/OLz3x0meUP14EfuTpsx6SHqY0dspOjGmW231SjIReVanEFHlQM
+tFsVANZlgNoafEPFG3/NPkpR9rO4iIFIbJdEkQE/EU7DgVTaSyAe/8IdVZDpO80
PRSep/psWlbWG4idMmZY/O7Vzg9gu9Bi/t6oyzOzDFpR21vemZKHcZmF6F2Fxl7/
Qpy0Y3sJUgKXZtbYI5Nmu3s/2Ba3afVhnORE8Q8l3vLhBDr+Oq/h+eCOFWtLN8kM
849LjkGBYYlVzuTbkTj41i5SzH1pfa6b+xdZIfSCMrguTMa6eJ9MV990rvdT2Os0
D8AORa4ID1zFCcZ3zdnZVYhTzpqd1y+LxKSk/k9ECsC6mJM0ziXmCbRDL422YYqz
lkDoMCynfmBEdM5ZUCPA1dqMFplmsgvP/pC/HzOxgnFEInRENnNtTCmHyVcwCbcG
pe6DCdDSLCw9i1v0Yv9n0hv9cbOKDf+AeGamEmUM0/AEsoEKnvJkjJ7pibm9E4Cr
MFly9NkuzQKJMNB1AZDzuNvLEF7BaYi9l7l1Oh/x4xguo6rJKxdYARh3cWLON1WM
7/dZM6Zzo71/sHUEL9gHYRbCpyUH1ayYrODjcLoQywpfb1Bb6TzNQSTgoev888Yo
8i/Tx3xinId5WVCEhr/0y6Sugkhsqde/+ceNCVcSokuh76QcpxbxT22A1Fknw33i
0SY3svRoXfDvW3aFyXsNkHmDrkBilBAqG9GwmXj3MrHYseOBjt95ZSV7NxA+2Msf
mH3+0Ehv4m+2gIlx8n2LDozRI2MJS39rmGOfq8f2TX65Fp7i+rmkn0VHC2xp1Zzi
5RmP4aNNqntG0HtUykf5aoLefMZ5u+n5/qHVG8kWVi3OdjB6yqhR2HMOBBZNgu47
bStxOqDYxUgnkNuZDZFIwQHGeMxTXSH1nmEti08XOcaGJXfAcr86rP+xbE6UdGpY
TF8+QCYlnOFx/IS4nLLT6+7b/lghBUOompleMaCxIRqqNygFkGouvEDOTIJs0bph
jj4M6smPyY771MPMT6LwaySL8APPDIhlnYrCLBYcRmozNWR7JR/k/QG0+JoIUTE1
j/Ykvtkt+arxnutvVYz8YgX/Ta4X0rxojDsF75hHFCGoM/pPkrPx8qRL0zSsW1d7
zl/op7KDERkVhE6jSV1wDuXWO3SWiFoy9vb5kPzV8ciNWj9HH6pKkwqrssaFAbo+
IcLnfJffnoGV56Bw6pum+Vga75552VuGNrT1bdH2LnPjShtwqreQMSV7zw1EKnnW
6XTpcGOer0ZDpbVwf7dCYQoiiMwAqJfBQA7HVQfNXbsEozhzVkb5a3JUAUcn1+Gs
Yzig2jpttKDEp8YbPTiW6Cv7T7KUPY41w2q1G8F70Rqy0RzWQuJdKaHEJcIt/HKB
7SrfTSqeq24buYUZMXjOQS/utq5Kat2K7otePvdKLAjmylWYrd49t6eRA4qW0koj
juTk7xetCe54V5atuvmy4esFsgwH/QuGfixFJH2AqD19/TLq8oM2dqnAJpjqk4e1
M/qAPpnX2I6EMmmeIFHyDdmwDo0eiMGwD34Xaj2TMhOCkqyUL6DtxhE/M15rU7Zs
lRUNczXJ8KnRVEbZz7ErtXUkFUCR7zEfyxJlok7LpTlMhCbws3akD3HxoXheNyZD
v3trhRl7DGhGS+sHlC+/rLC6gyMC1viIf3ULLJUZ8eLG3sS2Bx59zxRJtKhsO1S9
f+vuGXmpljCXBZqfecChQnJxm/MgOhVF0d79w2bgGTesLTEzFSXeOtmMV+mJW0PK
Ds35N/74CzTymy0EHTsA4NyFLnEiQdwCKKZzXWW+0OuzU3vmWga2TNZDXbgYOajo
CVuxjsyVwoqTXI/7mbDEV0L9uSxd9kNAPcmRB61oSSqzDvYDU4lEbTo130oB3a9e
17Q4CgUHNg9gz4s3dsd7zWX9m56MPySx22756PBPe4Im8SFhYlST4bYwbgeEsgjC
ijnm7Oov7OskXVfWB2A3s9/SFJTF7LG1oIVp0hCSfy/NmjWbA9Viygy+8cI+0QGK
QzzgJMVEyM/K/6jgjBN75ZxmAcqp/SVH8kNx7qIvrot+/YPOXXLPImEPoK0BOtHj
fzob5qKBQtVJEf+HlPuVLYkjsYVMofOFJST2eQR7ijWvJO71YuSUKxHFGPQ760QN
6Eu6M8DTgjfY0OsHMqh9ELmjKHuxq1aBFM7bawIytRKt2pj6JL8+8WqZk1mHynjn
MWAtrhFWv+qW3Pb8rX8MyTKohgTvz3ymSIUKkdGskAZWKp8O56M+CTh5ZFuxiWLz
rG+ntW89ycOlV/18FnlgiS63tq+yTZAgNqe41aF1xCh4MyP6Zf79eJL3VhgJrrT3
yx9mJ3hDi9kw2X724AcuOQLiAPgOC40lYnrGlBWixWTCbb1nmxjnzybmZYj7kT1i
JQNmoI3q2urR2FKXxooo9djQufzcDMMPmgM6wQd5HABf8JyYKfs+v+NHUVFQwkj3
r1tbjgsNiFuPaEwCVD49mdHObF5YxcF7QyNRBUvhLcHyTCFE/JPre+PckOQo3Q03
jzPQhdrXCaOk6z7MTZPu+rfUDi7VYBm2ic2l8K3B3pjs6iQVInkzORWUl6TR22OG
kuOf5463rqlKr0c5Xf+VZAz3OcFMnCUZcjfMnbtmmxiO4GZWoeLdn3Ilj2wsdEzB
NCNRclfzprR2DAi8XJv1dpsyB8UV67+K5uPNzyHWEpKeBX9YdUjR78znKq8+4uMW
T55890aa6JZlaEe7pi7J/Ct4M6abjIqaR9jdDmBiAYrBmQSD834At7NJYsUvFSow
HjfsmgPazA2fExoCd4w/GuD3ufrh4Ou3f9iI7fR7VlQEAP704hAB1mY5+oV4xkdQ
1NLvo0nIo80kJbV9fjFx+qEmTUDkZdVVEourbiHUWGX1uQDGm9xjXyWtioUg8l0h
5LygZM60aqUcSjd1lR6s8s8ztvLv7/t1eGTFWcr65ENhmpuo+laGaw1cuhglnQmy
IztSc0AVIAD0t9yv+PzXN6a+Ys/1YusgxjjS33qiLWk6NP51tspFlnLz7EcJYF9S
iiCPQ+S3lYZZxZ0/WnRhC4eitRxhXeEIyI1Gxhd+FcR4nrPsYlmWsHa5xkYpb1tq
fH6wVAaHvKkp7KHmQdZb1f/MUP7OSoOOxRx/CJf7ib6xqsnBfwgseMQ3ugbpefEj
GGdDoKHgUQ4J73NGWuwaq+q9mLp48a4A/bFSTtC1HLfR0/uhm2cKMasnmWTm5thE
SqdYilbofLoA68nrIikukrjLEOHcyhca61lHOvjL8LZhnNc3yjzyn6aB41zUXhJq
tRxSQ3LyWbSeKig3vw9iin8oLcvvdZCPeHK40t0atEtC/fAVCTzjwGMOdWqrekt6
3Hgk7vpoRJZF+WM7igcAodS1WiL8ZriFMfBHRjA/zVRCqZmdQdHasKGqsWIXcMjw
DlBM3fVU/SevncgYFiISGlTPRN1gzyxu8rxtm6fDcAM1o7sL0SAnVtcxjFzh+Nx9
rIU+2bKR1TZzIhPkON+0l6pcxX9gOcXRyC99+pVJJhkTtSoRXHp0xl5uos4wW0J4
JOjLa0rteR6+0ekLv/hXaVYWX9845ZWXxRMlmhz/GP3gD7P+cDg+TM6uwKznscdL
QGUJgD2T+hDxNkQNT8EDVJL4YocenbMLjINUcErQv+FG82XnqCToqR25jJGaUlkc
ogI3+4m5UyTzz/lEJjqRis2J7yqw2C1vRwyJn9OqZxAvaHJZLzMHgxaq5+D6vj8i
+1OpRO/MZvnPmE6/PkEXEN8jJoVbl80a0Rlm5XmNc3/TjjIcUvPbCvvZnOQIDBb/
24ru4lCMoyJ6WT2PQ+Wt3veD16elTluSGtgN0F82vZxv/nwf+t9O0pXrxaTzcRpu
ZumPjNkmc3v5O3SE93n/houYQih+/Z/3bsKG/CEyNxLQUDolpWTfEoYJpDSzJF34
r5zEx0bOvsSneM21Ig43SnxE2B8fBavtr4SI1nbYC0Vp8ibI4d/LRm3f1VEVXzoS
Jdfw8aFV3gNMbmTE8vU+5tBrOqlfXS8gf6ynM3yhpx9I5DSeO9nG0/i/FhiC7Vfe
8RU3zTcdxRXpOruyjEmnktQZUlrYckfHoJZfiFJXNpI6BNEospH/K5wkSHtSbyN/
IOcTDFLBVsX5V5RI8newm3bhBBqbEmEDW4m6hMY0EROofDjGZqrgijkArQSMEUlC
SMFsFVVgNxrnRvT8Asdu1KEGCHUpTv3WhYRxQqaRWysuW7G5fRSbzGWJPHQwoTf6
hr2/grsqQjwJQIZ+0gleQ0jQPJCL4PdHHeFxTtEgVuhMYTxcZYKnCG2IzpLd6DlL
l4sdWwNG3JHSH+9CZ9NlVMAFVcnfHcUEL4KHNmwJcui9g34c1kxsBXUlPKjiKEyi
ydBmREhakSuBzANggRihe+sgyURcArxIKmheO2a3JnSufIT/z6jAi9qvKjRLjT1L
W47pgd8hHOjsnzItz0qbylc0MwKNo+lWoWsbpSQuZUVOqLhJGkO5EjoMvZZRRu1w
WPvMnOBV0ms4cDnR5KPbn9rrIKtWQqJXjer5ImOqbK1SvSIfNVOJUOebN4cKzCI3
T4YddaxpuC+XQ8VA3AeS4Tu4ySd9twl8SfUp0Nbf32bx9UljNlQ6cozN6G2+DUwi
xZyG/zCaI/G1NwC3YZsNtxSYHYng8NZAoX3TnfSM0Avvpofk/OASQWAbx2fAfAV3
zdyCwqYyTZFSaalfYRNAT6xvKoGuowrYH6b2VjO0vZUydsm3qqNWL4h2wOzjn5xb
/liQaAIFVGTG4WTfB+4u1Dp5DPZCMkeoKHPF1UU6PbehqKS+wmpUesKyCnuplOM2
0DYwRyrkHdq828tIaYZGiPoVsbemI9b9ibOWYaLvvqLJuY8tJ9HoJ5NSomQZzp7w
hXccHVxXoiHbLTVz34FT5fhioDVAX2hGSTXEHN+E3MPEPtg/m5DVkFanR8Gy8vVN
yxJosR5vO8a/jqm35nH5vLUqA0VTNMap1N2wmdNJTPbDtWtFT2ch59BaG6DyoeJU
zjqX/uZjtELbZhdbxubyBAAn/rZSVpkev81F83Efi87HSS/X9YUkKtmqB8Hf4MGp
BjcEGRW2Gks/ISsbApL4yPlCEO/IkldDKSribAFwDHAn7EzNoZ5kdf9fPtPT1PB+
f7GGE+PeaRhH/Ph9ih9PvGi2fdiDMazmC7YgZ7DN8i7kKpQPVxOpoSxhVG0rJzHD
W9S23pFBuzI3W+Ya2Cy3RFeENfiq8Zw8WrLd98MUneyBOLY4eVOLWWpaV6qXeF08
D+vKHBQU3pcnJTqBd2LjeAUWPwPRV7/XBYt7JgzP9Kvu1f8g3lyZMS3L3+KxfKC/
f1Dp9D+kO0ksI92QmPtujJHCbABjeR0cFTEV3afeCBdSsWoROSfMDh4zlkr8lUVS
Z/LcEyzEdlq0LuLv42l1qLXNWKR5tFGGv3jPpYXp0B5s8ox9aZuOXUR2t+9qCZrw
tELbhv1ZXgSWH7UyRey/f4ZIznUp1X0sLOHZEbPFPMfDFRi/L2sfr5v/JacamVqM
KYDFlMU1ninNV77BOCidrEQYdNY7IamH6C0apjshlJ+5bUACRp3W84GkCoZ9TB4G
c9k+ANuNw9Idw4HqQoO7XKRt4YdVgzHYcVXwNNsnKbUcVvX5Fgx0BX26FbWsd9NZ
njQx0G2wRbX/LjnW3CjKPiUWWT4Mq6pmxZkLBrerXpe8gjQg6I6bsPvnYem7mekF
MqfTwyG21YGbRhczHRf1JDi4ZbMDrngl6j/4aBNtGVGTaNgnsU2Mw8BGEr/O9THb
EX7vtMWpyKNFKuIWyyflVmKfL1An8QLmMSH8hK6PaEHzkPKqycTZbR9FTisi9yDj
SnXnwkaWxunc12OLnXFgC+AnqjH6lQZtEs9yoHhKcYNJ/sD5L9NltodcCUYQxTRe
P2jv3vDPuCZTryFmZ1w8IGKmhGgTncqZzk+Zv4UGo0kp/395zUIfnp7ZHSfRnB8g
5RnqXFlrrIPAx78cbRYZfxqqvcdhsPerqECmyikknlFEfuTv2g7NKyWrUdoNKCpn
UEtyI1KjvkSnyLMiNtpuNb3f7IXndNy/MJX4b7fQdyFqz2kSkHMGlnYpeccB+EKd
v0ZuTGcyJAFS8y/VNFZo9OxQrrL3kE4PuMJ/yV4lCahcww9TBfAAj+dmOsJkkCr2
s/L+MtQZEv/9dzjnIjbgw5GpPbMt8535KPA+e+FCv01BzzChzQVkMJv4NVfc9aQu
h1ZCf9rupsYKOFrO66Tu67hbn+TZqnadxyw6jYELZOo/hS2vTr2wYgPd66JOFSyq
sob2g4hGfRHmk/vidkxDxN6EvraDE4ZLNQAPrciwceNI17+D6E4kPDeuX6t9rzK2
D6x7478LqPZ4Ue8/L1lxXWbVVnQJfp8oB3o6Ikinvbzo2ODSrL709zwUNzPFJn+B
bq4R5gBD2/H36PSF4l0wUByce93ZW6zli5iMIhAKnTmoSbjkrCEBWHQvvTbxndyp
j2r84Ii2bpssNTbK9alyO77537PmL6ALRDEfoqa7N1cdNGHJnNRKDIhj9uXFYWxb
B4yedTRYOe8Thndi1EIZn1/6ZBEPtPjsmZYsvXLi8Q4UdVTG3N5/fVdqkaHiYYRN
5JopnlJAc67diIo26phwcgcJmsExu1mY5ZRWmfogR//aYanbJqXfQ7wfP3hAOJyR
LhaALTUpmPJarsjf6ReTB8UZPwLo2zDA4rJF7lZC4yulmsskmH42wEBHDlztjfGq
KIP3f8d25lUhwYcgy/le+DohnSsacrJKd3/69pS8ai/arvy3njNb0P1vG4J4jzpJ
UnAgGGyyXdoTMcYMJyl0+oIn7HPgSKKxOp7rQTXyEjUa4Put1rMI6bvUxH1ktlyT
bk4WkGBMUiYZX1IEvO+l8/o37i0q1cXBqzLzsZWRP0n/Q1t8PvRe/0Xk4lybZXaC
OnN4eG04sz1vWfwAsirJtEE3ktRHY0fq1sX3w/GDNSrsxPRU3H8RoPc3G4ylXqUS
tafbOZFLlyAfA//ynDJOKJyflH7liBXzniPri6r5JrEaPG6N+ktjvvHob65rhTuy
3BEHVTYV1GuAaKL9T3fsemCSPmXfYT9leRl2kTcVa13ME/CCGpm9dp2dy6WVvk29
Od8TmbxpPvzG8TCsNSh0kgPuTkkMjcrtxTb0zYbzX7f96iUnCWos9p51MTKIsATg
vzrdTKP2leIcvVq94iPcW7aExdELFHeFDBDpdWmlAPh41QrIYwahFa+kbWb561f+
DaDr6Qfex6+D6+B8GCwT2uOwwsIHJ2+s9AqtRBJGmpvLfijD9Z8o71V/xaDWQZtb
Q+lEFFI3GyuIOqoHEhPGvnLMYkVa3dZwV8rr0RT1VRJHKRDdp4XIwWkyaPM+u9op
f/2BJGHdp3NfECVufwFiyKtXhXOUKE9B9xsHaRAgK7U6BODfTZrsyDovx8hwe6OS
rg5cYRtNrDnbTAo890OXechXGZ33N/Fn1nq2HnApWpa9BZne8zC//IdKFEbMIMhd
Y9dT4zwfZQ0hhqMKrhTLyp3mgGZeURvoQXcOG7b6M06T5qvNhs7o7bnmMlCJCn6M
4G+a6rJEA8p5Tq9rX7vYbA3lR2WfM1ZUeZLEUxlLIZ+L60O7W1j+Ust3YahCWK2q
FKRd6nuVmQP9xVH7PUIOrdAvNFaJPjZ7Rzs+zksaI9SqZSEWwv6SNnrTuSpW2tzX
QLYcdd9luRqFHNE35qhqGey8olx1ZdYuGkHuJtGkfiHIl0k72gOMOqJKmISxYxGs
2k3oTIdxQKBW+vLtS0cllZXTGdBOeUOx40a4P7GNSwSOkeJieDYmv3pA8V2FjC49
sgxCTXX33IuY0KtWR/VfZ/b2VQNAUF+o4w4OBEYq1VFFgzRP0DTrMyfxgct9ZCE6
YS3TVg0OAKqpHt/PZDiFVfe/FRUVQgNpCbLjoKF3hkTDLn3oezb100WiZFZs8B4R
RgdUzZ4foVwaXWV/gUGSJhk8e7G7buqMVfNTtEnbWH3KPPgvuAnvoM6n6kyPAHDZ
5dei60d42CblmWxB7LI4dUw4vvAGoVtZQUATKFms36UcQ+BODaa965zUUqaPZNBX
cTyArAirvY6uEUHhhDH0jIUcQCb+fXaGzLZmqQat6lyV5g3PMUqC/yw1EK44viV2
EBuPlg8z3Pav/zqj8dTZ8cgsrUffG8vviaiuNTykyijix9n+aXRSxMZKIM4KlSbh
suaodWwdH8FS8cR24jZTwzbC2MkTVJpcf1zXNlAS2WOsuRbeZElzSNI5f9CTuMSO
1ySXV/uINjYG1rjZGbH3BCPmVcLfzUquqlFNiNgrs8qi4TJVd8yyOBtfZ5Vz/Vxb
U37aAgY0Ti3DIykTG+MxDI6EJgcrKcaUcWKEYut1zVa2iLBJ6iWmZ/2SPRpD0GR0
X0Q+aKtpkXIXsw757XYk0ATOEKEpfnVoQAfYWZHypd7qAOE0RPf1DdB1APTll0r5
hXh+mF+UCqGdYrOmZ9nca9I5vuc89SpRi/Vr36x5Hdyld4Mem6lmXx0WBU6/UiCA
7HrlKAtWbVrBjZRuYuom6Ym0Tbegm0tpNIVdxYh7TMLkCuFbHKfHQpAUutowsO0q
3P9kz1ZWSVFpZd9mmfU2iRcT77BiRqgGipQ8c2+0rLRJjnPSe0I2Z8ulDQR92Ey8
dQ3ZqTy7BmQunlP2ivcTZz+NBbzbVKC+hVTu7+jEmYS254gzd48O7JobvVuTTqQA
jF2NL9J/fiQC5RmYyXnMduyDkmuFP3S5An7UGEOyKUb11RPx0b9eI49dFdVeYKPF
fIDnFK6TyJLQyXoLFG7w29A0lC+NbEWCljQ8vVBbCKcXsMLydDnZ3EAu0GKc7QbA
XNm2FinYGQ87dtKpq9OsRVRfPM2ancOy33tYv3YZyaUEKeQOGb6fOXl/U5rFsxQT
9Yymc6hHY3pSkmw6p9OqMUwMXUTDqFriGlJBe/3Ynwox5KJJbBJYzEdagXectChB
8sRloUeAebLsC/OYwhWH5TOfEpupfK/m854MBcepBOLsAjB+k05b3InDbqZJB7Op
Fw30lJ5ZE7HV+Jj22+CELoDFuX1Ke2Dj8O1zF9Yij0fhvEzsywHLQwSRSK56q35R
OsStIu/4ufpoiOld1KNPd+BsfVmSeUp9fc6kfSXfMDfU8wPwyzh8yXmBtzdSqMnN
c1yY7kg95LZgoQaG0oWVWL0REp+5QT/1uLdLhy9Egwm35ogdIokWUiDsGbr2zMeQ
svX+F9/F7EawOEUZ8wUohczLl5S81/va5IazjrOOt3cUg6Ar0QTinSKOhLWVTuld
sm+QEAZOA/hdOX42/3880zfSde/i91l68T7dtSo2o7OfEAHntpDtUDSz2RHQD3lm
XocHZ54x7eTgub5A8kW0f7uOVYbYtrYrKnZl0h0ytqVii/ASPftsr0iL3BDwjVL9
yxVzA0JSl0ArI6xhhHaaUsmb3HXDoKTwXuiVTT6kh8mD+a8OW2WRGS4wzsaaD8H6
//khhMc81KV//aVmiZl5FNwY4r6zIzyoSKs0qqtyYEF6KQ009DvxIpwxJbCBkoNk
/yhvO5vlZiPiTLZN+eMVUsnzBtByISYHYqWqMuX1dNNXBCH2n/xyiYpNg/9tiNYG
DNhEzOsxcwZwr7KspRJyR5um2vMlPex3dKOoopvihIJ85+c/8rh83A1TBeBeSUgh
fnsH1SL8VsXbE2Isnm9HY4nZHYelwofDXIYnrgp898D3uESZ4PWb2L5I0q3aG2Uj
DUAx9IQmF0tMmdD3CPrO4gMakwDj54pdw/41lUxvMRzYy8KHsMHWracLyH8j715v
S0siDzmPP1QMTyZBae31n1DqFiulm4OlwTYXHta0nTAv71qyauV5YngzoxbvGdji
uz9i6fUyjJYQNvTZVbUFgatubsx16yobRvKtHQui3zL4l19RjWEYPE7bzLAcJI0U
qP0xXjEf9Jif7ZYkPHpLrY/GBudrFNENsgWw6nTVIWw/cYTwDU/W6JqIzLm8wt6U
b9RqWtvzy4c2oBJEN9s08IHY4PJWwlHmB6F/3Ad4UIEgvY92t1VEn+Y7mRY6snJf
j09qfZ/EBddyE7oJ58iNAilbrofwfQ+b8AGJMPNTPy4qSXJ8PfyShncCRWAXJqw2
hn4AF75yC/XhnLMibOtfO/xLdJscccCg5vdZ2Cr6mHIqJay0YLxNhGfOdxkjtsMY
wnXGzqpesO335OoT09q3w7fblUDloOS7T/d1BbsFP1FMeeilLFgT0t2kUMAzhxkf
4MRbECs2kCd8futDd+MgXngPiYUN9U5N8j1TNnJNJT9Krpa3/qmd++8Gj+BlDho8
GSQFaZq204Q24KyzPo6uuKTQ41IqCucZTnb9ZOOz9bEJbdGSFPDCoIV01F4mir/I
BH5xh2aXlYE6quhVmghu2/4H+eXIxXI0Jyu2mjpHCMObEXzbWCra6KzMKGfXGeBz
qZLjCJ4pDQ21HDoCSM8FKvrf2iCrgQ0+5HdVyk2aSBiFvd1ZdfkN6vajpTEICZ/G
w5DLrKrbYPNcRa1dWzcnRfPSz6KKrjYUWsCM+f7qdMjDCvL3lzxQpusb/mfel7Wz
+7S0n7TPcag+l/0wePHJcv73ABm4SwHK6qSVdBGvDmMAvZ7GpFRkLAFkCpYIjlXw
OYxqPHJkzbpW5+krocsessIn9dhpLp4cc07D9XtDF0wmpUVkOzRWTQCRgNHvtJNU
+jV/ljBu15u4mey7FePqBaykjMJWOiqpXxhCsMsAsIde7s6DUG3o7qH98fm48r9o
wOksM50A92SHp7Jl8YSnaMa2Yh8xGtVDr8us6ZGPQf3HV8Y1FPgiazvxAIEheU7t
PIkgtHa/X6K4HCZf2o5K057VqfGYYDHGvtYqENpuv6G0kbfHgBvdT1rMLgp/n0xH
iLKFi8Un83biEBX7lmQOgAZ3lIUBpjp9aTKTfhngqt3HAVfHAWmXlTLuYAriolUy
E++F+wn+PlvAIviLerdwbSGsG6GBibhD8EBQTfr9bdpNvg7cC6qrTfkowhU3VVwY
xBTCm973X4Fn35oFPQvTK6kHjbY+Fedi1J3J68Ge5k35jsx0m1CWK4N9Hg8mmX7C
um9bWfKhqco/WQbczXCEX5B+eMe7tTlxm6GrrgG1cZuRwxm3XBFOOL2uSH50PsfY
rpC5m6ON2m6ZVncq8Z3D3pUVEZePDRV916v8m54u6q8xbRsLNcwKkjTPTNMOZeE/
4v/EG2A4Ot0eyTr7BF9zYNcyyyz19r+KOJLs1XaHhBPR7BdZEwVbjkEWID9R8s5W
DIoQ7vNaowwr+E2p+KChf7AixkjeTKZdXC8e0z4dHjK+zJasKm0L+ndxru6+iJ3c
UiE6Gx0bsFPPljy/oIwPpHLOs3VvSC3pnqgFqrW9UuU2yDzfSzGXaCzVtIb983Ae
xkkMX/G7dagM+xZZv88HWc+gB1O6vZxBfaYZjDsf/+h2Cc6Waz3hIByz2R+Qnfrw
xiaKwSiBDQuspMv7GiZdjj2NNbBs9/KQUk5CPuXQTc00f2iQEgpTZfTmj6/BBRpw
fBzwJFYHBqX1xFDqs6NrVgrwnKuAn+46jA/o+glGamLOyMiSnw/K/50mn5X+GBeT
X9tT7yltFDDZEEVEB7NfLTn2HypcPfQtH9zrwFNO1fTrbbgxVtkAnl4g9fBlcTJ6
PyS08k65qKJ6DlSqM4jewupjIUL7/PNYT84Fa/+bjL2qPJ31w0Q+uxa5/70da/RX
JuEkmMCKaSnqJq1XJs20C1X+HNe/PNO/VB0ysV2YFBfuG9zEJWQ97veeUT6FnUCE
zNyAbTOA9hHowOa7AGVKMcGCReRTNAWTEwtzFkNpW/OisCrPNjf2SVEKaGu5ZBR9
Fbw7/3P/BWcf2noBH0GaW8N3F5kBi8BAeymK3Tb22yWqtR1A3CoqVB2dQGNMCSLq
UlJtRPbyNLJulgUlKAC+6AuLv0JGAsiH84bngvnJ1Taws/OcFbg6PyLJ2jHqrUpT
GSATFJH4BJyA4daMZBK4XZ8BH3QayCpVSdTwvaqDFI8njowI5VOytGoviQSsHl2h
Qci/MmfzURwDSR6ZFurudJQutY6+BS1RjdUJKS8bLG5w9RfbxNUle0/KMTDkW6J4
rWXj0tfaPS9ci+M5InIQIHzNRcYbPTRLEY4YTff1A6hm/U8iIE0GDGgriBRb2HiJ
7dNk1GFQxLc82rSH6Sp6g/sND20j2jCarLQ/+J0zoowYFAwb4jHp744SG205Sbhl
FcaKPA44pPxqlo8LZTgFYj1K1I2vzVM0thgC/QcveWTrWkSlo/1nxfLh0BwUyVti
B7E7Q7OuQOgOepqYoVcqjhSGXUo+T4tFad/Ppgr6pRx7c9M+4RM/HwlpWwjVcROJ
QPvKg8We3L+fAmfz7jf+2Yx4aH6UzVd4M7u2DA790EjEoIVpq3WmIejKaPcHkbr/
UwOXSkqpp9dGZv5j6SJLPeOeMmfdfdqhnAsYN8KBjgwEtjdWU4jYhZ0BzmayvbXC
us9VmSXqcR6exhLN4Un86NvdWjghQguwgOf+MyUxzsJwFrvPeB9IwZ6FiujEThNa
/3w2fhG/cPsa8jLl678jyc2Et5rQX38Aclyyug6IiRYLE+CGMw+rDXb2/BQTmTM/
+LDJjKZQ6H/QJvin1D1jgbk3vUQxdMv1RUyQQ7JIfl+qT6EaKE/pq83nE4bbYwFk
Xh+3MShbtrQoOIeLKa1uaRlZrh2wv2E/t4tyy386y2PKqcm+uDfJrJS+jxqlXczE
0o321VTrnudYbkBIAKDMULyX6xBzP+M81Ktx4jsadR/7OYzPpCqPOCW+EWdUv9hb
ZCrBUsnGKJaIQ4H6ytCMWB1aYw2G4/1f/OfpLU5o3gUabp9nsXdF9YGtTU/+GfFA
mOO4jHrGKA0BDUKku00yW0f+XWlNVKBYQGY+g5aTslXCzVCzCOxMUjMQaahcB7YR
m/O0zr8Thh0WJcJjBqkVz5OjcQYOUWDua+asSIIPzMuwRG1JjoCq4m5QnsnuNWqb
lHsHdz7TYSX1RrYciHf4uk2EWHZwAvMjQJrTPlmIHZdrRvqaJ1PdUhkLsfjma1ia
b94ssu1/RAqGmb0Yb8y62KLu+fhnTp1OwoZitXWjYuMZVT/5scoTwpYCdC7ToJv9
pvrHQ5rllltbhYZvGZ8MbRbIN+AOA3tuRk9LluwM10wKuUkvFHd8IV4j5fRLeYi/
LWlvA+sPh0p6Ke2BwioVOlbI6ZY+ZmLSfkZ87kvh4t43EneS7d2B2DljJrmSJ4M7
98jv29Ur4bdrnlctsIV4uZjF+0S4v83ObHjlHif6fGrGNnCRDDttnlx2diWpu4R0
s+chfa18UQUl8QMicpy6Hzz3wpnnutbNMQF6j33yRw+rAr3AbRms5dk/JwoyIvg1
3xgSoJPeDSs1dZpupK/+IMgIa67usI1KX22fXsmjc0QfEnZHCjjV5dUqqAWmB2ls
vfQXe5xK4y4sv7iAmJ+HvfaLFW1sCzWjFl4xhOviFKCwnGGT8PX67d3lsTpou/Yu
JVUBDNMitUlpoM7fVOgP6qNG5oHWSLGPBssp8PW/gKbONwsDI+6NdBKMtMoRo4gA
1Yh2seXBbIFzDLSYB9tdXCr+jXrtUazRKaqP+R8BsioLNfjNBlDIbmGhX5ujwK5u
nXaAZWSyP3T1k4BeDtLkW+aw3RePlz4DpEHmU90OtS8XJZvehw3q6ZvXdryqG57G
UUQqXtKd0K00V097YwNB3JdAIndUOlT27u3OVl9iqPZVoOvZSpp8mW+5TLY34jo0
HD8rVFdftMKF+75/8Rr8/Z6LwgljueffthIqfH6dUCWt7yaiduAOVdd6f7XY4+6Z
VeTC/cyqOn4Id8zFzrG4hAPAgZSp7iSpgINpwAdtUBmTiBqjfz4TllFMqDIPhRWz
+i9TlZ7Qt0se9JVSyb494Y/aBIZUqkCYqiEpq3qdaYFqvmq01F5IXmQeaQtkI+BL
0RhW0zI66n3Gdld/1TGBcWRk5IXD/smXwCMvZLfs/MKwtUV4fvH+aLEFligaBu+M
W2wH9Nr+tGd4dvN9zRyZS+L2RZEtMxutFcbnrfwISLdG5Wt1agjIzPBufcnUy4Gf
ggMXxWCUGhi2eMwTz0BekEg2BVt2W74eOZXLf2Fs8i4nKq28CFBGafH6cEOB0kdR
W/ZMmjOyVGbi7frzinkZTSmkyXwHH9/MyR2wEwzIkvnPA0GGhfehfudtj6pX76qc
5NilNiMgcB2b6QaqqSH0gvf2HBbvMj2vu5pizaaW3ASR8RTHK+9JhCzHlxjnkxQt
nnOztT4IpQX4sjvmHoBZoXrG4+HIzXaocsZmdUrYZYkKPPMKPgThr7ZZlnQY6vdh
UU0bJWof4CIKmI6IgPaSS61qI1Ze9k8v3F2kQ9qYb8qNB/p6SlyQ68drWH2yy1c2
9871ik2bhyCT7X3d11DlAFixKarjptioVY/ka+YnkvrKCb4iHjFdqx5bBpzxXeub
AKJzbWWbqoAyebnsijnQ8GI4qI0WG3k42NZJAdcemR/Ti4MawQYwhOiGTZPBQaF3
btU75WJs9uBHsBVQF2wutIynsL2kSsUz7KDLOAoeLgViKRoRbwlbYW1+A6oIVMRn
ZZCYB8ENaUz1QF7IFohHkxtpMN0hOPXVA89/QlZZ21Gg6x26ue/JFdR8uu3LsXtW
F0+vkEKeTc4NYjRQhOmxmGVoTktDZlwwywfN39RdwJYqp+uSK051ndZtJhxhsNfo
M9nbJPia8oxWgkOWfd6doxVHjLnQsNdcFjkvzTxDVorz1EzFqxRkwIhzrk1h6D/z
n9uQxF64OkmoGz2cnq51h+qlsbnAYa/YTqbiH9uFeXTsONaPsgZZlii2fUYVuNmp
4Kv2b4zNG0O4yVp6dNQPEM38wgSlPEczeXi5tWP9J63suB5guxvm2XG3tqTfUauF
8dKm6/+9RRF4r7/zd1Q5cyQvixmoeKj8wzYNOoXSTRrp1cpgzT8/qYpRbkK4kIl8
2yJGXDBID+PCffVpCHh18pqlq4J8wYaAKhLaJ7dbSOFe4keafLx/+clAB5Lxd1SC
S2v4ZGd+Y7kwZX2wCAQ0iihOLtCAbe28qk4t/5O4A8G81OJC5JN6UxUXEOFs0ARw
uKMovQznOQ4WlVNzaPPEydINDbmOVUjwSTooy1oSUKZpfpPaID2KTKnhlTM4Meea
p/9kKVPgTvVhBKrGIVKezFidgZySvi0iqL9RKnw/FHGOZts3bLF/EOePyOr7nhG+
pW/oJxsNAGzLJgQE19YS4TedVlO0a0BW0yDViXtlPnFJb3pe9EdCiuQswCQ02Xif
zwbS2SQTITJXTgu7PDIHzusdBpFBStU/gGFbc88aU4wr41jkWg5JDq3tJ73dkkE2
LxTLRE8pUWCB8QFpcd8BZaDOXbe7Y/Ux/4exYB6wYSi4X9FVvV5tIJv4n7K9vkX/
XEn7nnFHJw35uin9udie7MZh33GYTxz3FKCNsgk/FD4IOTA/JDpYDw8Zb3t8uz5L
/vB7hLZzEpLWtERWUWg9qJR41FKgPx7hlmtEwJjMjdasR1c2fKMoyEWLxaB6wi2a
1iv3F/4gre4AyGKgyYH/nS/QmHo4UkOqninQtP6toEligAapLxJyOoL6oTZW7hHD
Dy8ZPgO+fg4bToWn7oc3Nna3j+V2MAyBpn6WdN9nVVdmZz52wIIsWhXRSukBh2K5
UdpM8p8tdl5goEup+X1eFi1U8sfcQLbVxOzDxyUqeFpomrwDmw2PxxUJvjr/QEAy
7PCeNfrzeDisMXPp4A6c6z1V3KlbhyQRIeE39T3SRRNNUzc9Rka7PMgCTtKH1IGh
huDG3xHJzOEvp1AQuoqErIdi9hvg0tGnTxwGNAjwitmCgGHuzan4bzspgOHhVbH+
ZghuuXn+LLsIT10IwmWFaQflCok1/WQ135uCDfWgnO0A0MktV1QSgEVivC4tQktd
bnaEupb3VLVqImh/nYvo0L7NGy5y9bdCmrRLqokJHZytnD83X/s83xntX8/t3CqP
yLstXBisUEV2lxXYINLpQX3W8KMa1WZyjXg5iE3tBPwMIg9TeSFlBhggRXZWH9wG
Cvi241pUXjmiSIvZ5+7vzUoKX/zyf1YkjPnUHwoTmSBrckN24wtwDZE8+HHjD0/g
AR7Ery8OLfnxDFxSoJrgbprn9aaqWiJKLOnW3+TWigAjtVBdKwiR2s4rfYzisLCd
pUT76twb+FzzDyxHNRl8z13vcy7d0Xxk3TUBaF/dPBtOchO5MRnc7/8Ai+TS+Lkh
hQ6AUT99txuQYZDlqyvHeYVRkLnMYT83YZXl282YzC9STF1Yr8xTzUiEyxYtR6WN
UfEzloNhWMWJBLK9E+OtH21vfKwiBVFZBOYyzKUhs4mzgHSBElg5G9LbN5e2Y7SQ
u8bMjcvRfAyaPjVTELqIkT0YJk9pRxyYVNlqILScH+mIA4HH56oY2gW9Uuh5wEYJ
BzzsfnMOxQkm7J0zFc7i+CTD4Ive/eP7DsCkvaaEOQuALKDT3ZwmrivsAWPAeF2E
aY0JoRm5GMgJVztkUJLJu0rnIVoGqqDMe8JNbqN0sLjcOIAZSsT6p8LzO9rE9ckx
9zMAloKacG83VnAEkUjK4e0dHTJOqxZsixlPSrP6/iMvl4pixgG7vtXQJu+16kS+
drksbBmFG8fCbuKEEiDKL87y6LUIfqCIUD7Ra5QbNrixafp7fqXJ/Vv+LxyrJtbn
UBibHCArPhvJ0MN9cmUq854JFwHxi5GMn8OZ6m3Jsoj4zQNbceI3ge0WOmVTmiWG
NMRs/+KGDw2dY3ljB8NBivCHgU7HQRK0vNrRkrh+RsVd0pUksGw3+SNnUbvNJzSI
W80p5VT1156ZWM8lVmmda0iY9FzVZ8ZRnzLY42uwrnmymkyhNZmVdRCVKldqHtyP
+qOE6VCZf+mvclF90Inq+dzIVKh+i4+LRlZql9LmEQw4n4pXNjmHp2eL3qdy+S58
6hAObVSc1qkQihNGuUm1AVM3EwocvXe0tL7cVvEz0eNF8D2TyE5R8N26ae0hu40I
vpYvHvbLsnwA+qJ2IlAzswZBjAb4FuhV+i+8Q3dePjSgONfaf8Eh8Vl29XOBVPS+
lK0AsPesrnD3n2oA/UpZEWe06r2YbhQsVQnlyP/fBY0VG4pe4CJoiXFkjB/Bzl6P
dx2mDAsOHsqQrGcPc9pBtGXq4ZNY4P4HfIIV3SseFuWLwlI4hdftzqZfiAFRBL3G
RahqiK/vdsThbVS9xMSmrSwxRUi06rSGTD16hu0g2oxrH0a+1UYasEnNx/R002J/
7edIpr/WGr0Y1IaTU4rul72oYWyKti/qFd6xDKivnWlePaZmRKixsoj7YvfM9Qsu
TeOJZxDy7JPcWiL51q5FZo1ML8Wr/LRmVRbU2/FHMxaV5CgrVcj9LRYypjRkixIC
ZVfP+au3G0sUqeEpHjm8mtj9j3IlV5FBQbunhqY0ZFvQWak1eVMBnoPrGo8QBILp
pEKVXflY36XBmNRYvNQcftmpWAn25RbizhX/TY/OZaMnkhqSQ3ICqnU/Uls0JSCD
++ISz9WrdgiKg/DsedL47jT+1CCLQ4Qtwep/mOk8cEnP4UqvINgnrpxoTpW7nnY8
hb3C5Ovi3r2gQN7XSAQrKFXskWx+WHOazaZ8Z0+WKCF6aJ6uKpi7FJDnn0ab2ORq
nBS29omtHbJTePTPmTbtj+AXtn0es1kAJkXVbt2hw5bMA+zz4TjcfHDxX2zE5kB7
jyC+oTcCVy0Bd26YG2xfhxrXLMG1fkkazixpgcJ06TLlDRSwrxMJQWINrK+o2LWz
XYUo196AwQkcm3qKhAPEwxKqU+AV4Lgu9QI5xKQTZ1ldyxvCO88uS7IMajiSBLoc
pS0+y3BnVFvttG5hcu1Djic1xA4QJ/20+j1MoNmuivp6Y0LhZ1z5ftdaLXNzt3E5
ZgFGKP7tu17B5anstNz2CxAMgJWCdcKnEesJ9yUWaHoIsWanIZPVIkYBJavH1B3t
XIrYmx3eRWZiAgLgTaGucHRZAsyX17p+egVqfOHNPg+bFUCzQb29/A1lNccu9N2f
jPcq6ic99+UXpUE/OmTImLtfEXk8Tv2MWV7PrReBEkD2g5P/liT1eOTzjDtbpXY7
cenOMtkYZ8YPA9EynldoW62kJrVLYtfGkm1qrcRH37kee8FcybBbhZY/BEpg/qz3
YDydPHxGUxJD+B+h8g6P9nmqSDyHqcC5aElJQLh6lUtoltScQzCGmXftpFNmTZEt
8CfE8ztCdLb/t8aB+wuhQtDdDrToaK9DwdOfnw+S/252Fi5RJlhW9RDlxa0TJL6/
hXlBGaERmCu0C0+7ryE9cHqSqAjGSr4J4DgVyEu/xo8AYuFLGmX4B8WOWPZHDfe6
M7KUHkTsmEBHCmX/bkwfKwxuH0AmUYfSj9wqhTdZLPkSzO3k7SqioKITGjx77+oh
F3D5Ioxp8hEjJBW6rDM53Xh4T03dmRji94zBNOgGQbToGdfz1QbzQucQAjWG4tFz
IXtq0/EPGXrFv4On+ErPtLO+6lzOGGDLKWgfL04tRcIb72PvQe/NwnoksTbu9Ss1
ajQFjqOo1Fmcp5pcaWZgZwasFU29kCeJDGiNQ1AgcUgpeazEaXcn/faEriFKIEog
j82ULzutkEqrsnlSbOiEDxXTR8w7QE8QjiwNtSTMvrSVp76WTB8gXYQOt2nN2LzO
iwhht095a2dei7IsBk6jp0B91YSAhUDOkiGk/W48kCWCT3GTbaKr2zOOPCUkT+Vp
s+6vWd1xwRe3OIF2owibWYQUIXne8/1US3EbVrXm9TWUyf0qlDdZsBEBSuqmbwdO
+EMVqF8rSUgqCjezRbJxQCo3YHYjQchxQidrD4esQq0PhSbQttfxeome9G9CysnN
gGiEeBmr414Hbzhs4J2fpSoasZGY/W9CxIZOF+N37XVfO7UOPoBYWc6y4hgxrRpk
IAkcceM+5/dL0PI7wiH71VvUveZozK9t/9+ZQQwiHpvBPhX2fQKdwRxCaRtcFxlo
5CLDOtJSm/nk5jL4y0n8UZyypwyYQohAha091dexchhOhqP+yClKaXyhJT+rplG5
3McchW6UZGGLAKxzfFHnUjLlEVEWuq/wmTqs3mW5BLtYhovXgFm6XN0fgMxDRONq
aTXHaKf0cIgwfcazgmZYjHBNt09LdyeWShyuJ+l7HnA+UksZxliG1/DNd+z/5Ep8
kRCIvrdKEr9kPTKJYh+t/6zflpntgVorqbQ53i7YuhyIFDMOCgo6ZO1+pdedRbKy
Jf+r4rWOAFmxYZRO0Hc3ih7Xc2bUXSPrfmmvYJKZNGyPysfFII9ImBCtK8TF0veJ
x/h+L5vXEgjKW6PUSUtsIEoWScARF1q63CeY9xqz5wqMS0I8LiZCI8euK5S6QRJV
7p/yYuMDBl4r708pmoj+69sUcge62au/+WT6+WR2/Ze2LEWQktMw+QbkI0s+6UFX
MSpH5bOW9fVG3XS5JltevDSPWfHvMcWhqT3WATHg1sYVCNd3g/xQrriwVZfDREPO
gJMW5KmpBTKlnHtK3e1kLrJqIgWmIncRyXpS5P7fG43HXVWS7j4DxN1mSY2kK6/q
DXtUiXWGnNuPzqlfRh609l/Fi9QJjFA+EKQoWTzcfp+yCGKlTLtXq4gulY0y0j0O
InSMCsfq+rGBmF1rYzOKpXC/B0GbC0ATrTgvzRBz7EtSoUtfPF/jD0IqOPCGJVVe
Q7eVyARLXvMNqtzB/kq1C5qKDGRLd/DbnMSh2eUXjh9zf2novO87n14iLRfyKcTX
LNam/Lz7gFwTODVuZ3tmWOOyjWY2ld1gq6VVro8Q5uNYxIw/Q07bweiQWzS2nXya
ki25840tuPjce72tFThzFzPFndu0SMPl/sIP1gCMoyA+Cl+HJpKJpyQhI03eFyYG
YGC2fJx7vwi+QwJ9KPT/fOgYN4irzQPlAAGTKmkrW9xfR22BJ9aBiStEABV8tSo2
1vBklh5OOu3N3FItMrDkGCItSN//ZYMX7Rfzseplsdd1WhdoZEOWv0xxR1+MLUi3
gimSP0nsXY6pH5rTp4p7KunhPjoy0XRtTgqi8xKYgJdEUsI/rj6lTUltTMIgiN+o
7p/+GUjiNfrznAC8GkJOZvQ3KontcPBoSswpl/dAshFhoMYkNuKaX1N6HvZg38u3
l0Ms7ZTO9PYkWRSn0DPphpvW3EJD6X/zfiozQSxuAtLAt15mWgiZLujxWn6V+PqM
k8KNfcdTz7FiHup04P0WchPy0DQPrtiWAxyECocFiekClJrUCwZvGr6TP0II69Iy
fH62YAVriKB7iatScfyveVdrieyTCZD4JgNxy7mY7EmIgkLqFdwn4M11/VtMZeio
NyEcdq6G0kZluUFR3cPM4+jkBRMD3BfcWyubgXX7oxsLN0Bx1P17VIjEDDelgukc
qevVJ6beq4WzqUeAKBwYOsU8h9FbqnFDZTIt8fYqRwtiibGf+8KvT60SV4Y8yY3V
pTS9WzITkond+2KKvM4BFfIgm+S2v0kL3UFLujXpU8Pfgqyp9hW3EOUgcEdvNsod
D69lbX8bhQqaUdbmwAXqHMuO3fBiXpTWqRfzLDpzpUSsoIE1Rw/IS6KFVHi1WnNR
hew3aHOmPKBuGg2sGQ00mqucixAtqnDvhc+CqWtQH4K7RtEndpwS+aNW8bXbBkCT
/FpueYtK1DsbK6HedgCGJH23LtCae9p17XdJjMnuiriyyX+1SV5U2y2CobLF6Ztv
o3R/lfk8Tk0c0sCSkB+z8P5hKchmCZ+yjCgM2zrI0/OzShC4pQCJC6nWfyE1v00W
s9pTpzFFyPfe3JiIJy8u2F6p/XNcSerynFwLlbjhcC9JznJTnlzRQDWYcp6qzhso
bKoURVwVN4v0WkIEQq210oYdI/d2UfY0A4WecT3zayQSS8fRqux+l6F/1uAoQNkT
C7RmlFZM4RgINDZY4afY2B7zidvgS4a5hoG7e9uUjCPoXh/8Rtq33Xj9QynIdfR/
Z4snYiz8a4XP1GTmn6Sw5go+BWUOrC6YxhWybWWnVEB5sGQlK7etHQmmxCNSaSD3
P0Jt2fDUUBlmag8esYezf8/AoveBapp1MgC1+rbh6xaI2Wa5tc81Kdu9emDmHvKH
EwLlJIDAoLNdO1CxGf5zgsYtbNnvzuYZeE5or23tvtxnIoIB/YpODpjAKLZwWqld
wyrY1Uq/qqn6MhlWQO3fZcCtJiqfdXjAHKnsNMjuxsdt/ahQ7wRtBR1sNYsADMaL
7xKuBu6GcAugSAGDDkPdfII21ULp3+kEKtFuaLIC1OfTCD/YKgOy0QC5xorOgBXZ
M8yN5NEsBe5Y2t5QSbj+IFVRDrOo0xk+ofog68lgzDCWF9j5t8gYbBOCTbbOhnfH
oaMG3rOstAhMz+VbR5BrIdSNPg5lNjqm4C/yJfot6uMdKDcSGrR3YkBrt9kjZQVM
JUvDL/qIYYFvQGB4WpmLbLg04lt4om7rUeh+s4KLVNbY3vhtbJJkTneneNIDc7eo
95vfKvfmJ9fSWOVIFokpHy8oPdAjbaHtlFD8pWwEO0nhTNgM4Agz+ok9ZPgtYEsT
LiwvNwHfSWJtOKEmqdmAp29mJT4Q+HEfcloh68OGg2wGTRB3LYMLI5LE4kSLPz/Z
rWaWkHMPRK6rifYmg2YIEzJaCstulgp7A/H8x0IMwmCiRZ4JRjDB27DDRcBDXD2Q
//Jkci0styyr1/XE9I2lpRnLW8G9Ilw7vBJc4D8c7WhwbszmU49Sgh7iYgwZuaPB
sZ0149yQQs4egJjQfLSZTthe1Bk8FXsa5e2a/LS1cn43oJKRSe5PL/tQeJRQBAfD
Eda7mBeSILo9eGDUm98EL425ZBDyGnQnaUSX9iT2AL73ypt610TQqTCy1tEMM+Wb
ilb8x7fX2dIfJrSUvjPsQV6q+jk0Fyp3LHsmw/dy+wtnOA4gjrbaAovXGhlSiCBx
OeLMWQYWYGXJMQ61ocYtlqWCGCY8N6mRG9ATLfvfE8lhq4fh07s15dt18v8WHLdz
C7alMCEsk1L8YJIrjUF370yA95F3FWJzocNoCN2/k286eQSZPyFnvsLJyqUnMNea
Z1eaXkgFPzHJJnWquq7GhTGLKdJUlNBRnQt8MR5s8FWwjeG3F4XhYQJy5BnkScm5
tXDt5FQZpibRlOq3vzPQH8/2grGsKRbbuRmKqzULwA83ehGfdcXNSBHmb7jzjFWq
4yhSqM1d6YUJVCWxMm2786JeVBnKDOJc4fETMSnwepRC8ft9gAIy3a1o12QOZtOv
c51fNgklt1OMXnRSfAxsLE5EvS+ZtyGaJQg2s45OlB/h83AbpzOvn60z1BOZEKpn
UieodRAX4Br3nCCBqVjg3MW6rHZMkV6kim5st3QjF7Raeb+Y9GDv1Pi94NeyRrYH
Xdu/PBTplJjsHEOr8KV1XdTbzwHIIcbVBUJgTDXKshzyhGz9U/e/rnVUwp4sjL4u
S7Ci25PVLw8y69Iwk4vs5aTgBICXk9RqEWKYuwdkFqOhf79GjVp+T8H/8qC8K+WT
PwrNvxUKPmKNCaeu05AqidoGZdsqACGb7NGvb+epXINHuuPW1X5dWIMR5RPJQKE3
cfe5dMBvx3Zkg59md2t5IilB4Cy7ZANsB3DB5/coSTvNBqab95PpzpROTHDh8cR2
rkyYoYGhGvILBOJ1+Q9DCOQOTBObRjWfYpvBBPaL4IOpoSX5Ldk2O4hzeWltOn2y
97jkfVE3mgtUIcVK6+3FGsD3bvjMXBGcCaBGNoXD1GGBzr/I+L24pL/KSugD6YLO
i4f1DTsvHAbyDb84SeIzGJztzUnQgUXacbE5aUPP0qQ9eLpoeV0FnezNAnrDwVRk
ZAxc/H7PoJjbYOtv68W4VCSOBUCpuYDDfLdWer5QMa327I4IB3ughmV+BebREz6W
nWK0KrkFSmXuuffSOzAjuxIRL22KwccjrjaMoTjOAVF8JiteiF9CPvbOksEc8NFP
vONHqkbjB15mPB/OsPIcpM/xU7kHMaCowa8NgMqHcD/V2dJlfmDUR9TgXBbINyI8
JrNtuqCtZub/7VqxjLnNNG4W+SC7cHQVr0rKv8jzorbesMXTncav41sjzjUJlLuV
ikUnujj1yaRoUq9DAQyGVm1DWZ75OtZdl3VJdWxpOmeVixZHMSAM/hFbaU+8uHV3
I3wRxTjqFYpj3fIwcbUGzDhRftatKjVSYLCOVUmGGrHsk9+tQYoVgW8bk606Xs8r
pT6JGIDQHZkLq+kjL5naK+pzm7mOKJlk2aBna+sdpgJirWRpZU4JFw8ZVzWjerT2
PL2k6P3MybmdfW5785JLplm26/yzqMLiadp4HC8/bToRkkHKabR5sE80m3+LC/Bn
70IIFR2msEJMz/PtyLrOzoXuud0NhMmqiZhSWQM1t3OvFmEaaV/eDcXo4GkjuMXv
sFLYalOMBNN9p2xquyqLUjIdXkML6dHMaNzXQbbv7BPGpc9IdYMMNIF/O1JMN2wW
fumSj53+dJwEiMFFDdbSP5xXr4DMlOhyAHedKHet9j43fCutmhjXRZWdeQX4tEO9
TWHqY3z0f5/FjMC6w9do7V4JuWXS24g3Q/WSJrGjWvs+Ocg+gFANDNeo3ygqmOoZ
8SaqYNvH3RErlzAnNX4pvVVjWdtVF6PNdEmKe1jez9wBnaADVElQyFl0wZ6QNqN+
ct6Y+Pcq5Xiow3fvKObSJ2bs4kWWc/npLtpR61xP+w3ls5mj7+QdJihGwtetbix1
pRyFJu5d5yJ77Z72VxSVKvxKV0OxIml8CiumZQDKvshFb++npUteVKCqYw2pJ31C
D+5ym61pOSIFC0rY8lirsJskJ59mQCvd9wsCcChoOxvfvCgowqtxNDxGZu8b2d1M
EjMz/NkgjHvbX924rQXMLOAK3H2mUs9ddlI1JazBhcUboxLSmuA6dhC7q2Ar1c+t
csULi49DkxDj//88G3yf8vnIFmfXVE4i9zKkMVKE+lyRx4dscxgbtPfKGgOwxqk9
51M7XVeFNeWDqlLG4zreckI9ZK8GBHmj9Be8kMUOnkPlCNaZQbRNuT+2d3SxGBUm
Vb7Ldbmwatct+QhsDzM01R9cwKkC80U3ArhfhDAfa8/+falmg2IE16q8V9sDaq+u
0HmWa3lQq42oboM/XP5lq7zTlBpgxtUtXZbd4d4znrWJiQzePXV50KjouDpS+0dW
FKfA0Vybsu1NMpkr0xCvRouwDJ9+kXmuJ02ZQiHw8Ya7CmlpIBRLoLOwIcVL7vvL
4YxHqkpA2Des287HXo+CrV2hOhTqhH1yEouhrj3qbRZmt3prarCFhXcr2j4cu6bn
bKfmviXtlatVNZpo4mZKGxw+BLtfr3JD5Pzv9VJWJbyhMxxO0wnX63Rmh/pepS/C
h5riHgbObeYys0gRzBOqyBKjGpLCWbpUrY5yKmgvMgSK0cBx3l+BmgKc7bwIVJ7u
SmsM33uS3sxySukxWOvD+E2HLR03uB/7dNtlLIohfxCQfE1KeaCItNzVYgWYZL9S
nzvMsxZuCuA/YiTXEvIPIv2r/qk4PTN8Y6vFB++AjjVUDazzgDi7jJz4yDE69nrT
zNQPVI7nmdsPnamh5KVuUpfISu36a7vDdc9aCQYu8ZLmlmEySkTHIr5ERzS7U722
uj8/9NRaQhPVYW0sQ33/mMrMxqayLPRKLzd2aVaSSm1mnozgFWnGu/pchQpgs5rs
461prYawNx6a7sPkNbd54UmMi1w2+CkTZ1oCSP9MyPQQb5wSaPd8YkXvupwXUt3g
kETFq7YsfcuCk5I4WZjeLZ/yZ/cQjcpmKxQbPEV68OLDZiXwN8Yki2JVg/632zF1
vyi7RRi4V1vhJAo45U68SnGLZejJwPQK8iClv/6n1uiA7L9XAdbOFoHAIxK06MJD
g6GAlJIb5w+7e+w55CpUBqZ9WFmk8xmyxDvMa//h7kJIJRNNBIcTbBA7KXxH1qTH
6bkboJV4NeYqGSKLLl55eO8DOfdqaVI2km3QZXZhf6EEUFBSJOi81NnpaBOJzhca
uzy0h1rAam2dRlUhNmkrLJd4RHjOLyKpsiXp6gqP9Sqoq066yJm2lFt3pfPlBmhl
ZlwtEiWNVPef2e4vAORPdY8RutxcSmVz1fcInbRDxvHveRfJYyuyEDEX/V21tgd1
jEyrUjSD9ARJv6PPE0b4zWjPW9x97KRH3yZyyO6Uoji1/+yv5jd2T/GAO3EZkavL
/7A6e+YbWj4wsNozV1MPiNT7Au8ZwZPvPy9t6MalNPYuny3/+Lg26EQQiN6v0Wsz
U8GePqO/m9CSqWk0uFDz0Bj079fJlEaD2AVRqLtxlq2bbVCXLlXEt9qSmrmutnAe
55h4HEwDu5zd2lB10u02tnoxvl7Zqm0RRq8NV5jqb2ALOz2Sm/CfCERsFWMhd4TC
4q9hJgNJBobobPRPafv0Qs6bOHVMO/JqQk+AIEoH4Lc59L2rC/4ntXf1LPCu3dNH
wk5gt1JdxWtoMl7Oc57pTCG+8rbtPEMwQA4vzrVA3ZDF8Cu+Bm7D5JUYfJnx+z9G
gLQ9eqHFSjAjLSeHM0Llba8GeBIboKeinp1BIG5tdv0tncJGizq2mhwfuvsb/jf/
15586FL54BOZx6xEcEmTHzzktRkiccvS5IOnOL3aGq0+Gp8c4oGc2/QRdjlSGzq3
0yAHegveLNcL+UXrKYnKveaXavBQNUzAOrxtTuxmtNYwy5M0acP+iBKXM5SnZ1Dl
SFFGgck+9S7fkLa9pfELw6Ad6YnlxtDbT9FsOqtJruacwzcQpDiG/1Hy75X7vft3
JF7BMMBSvZLHy7ari1xmRzdYBMGJJoSESndEgGtfYhM4DJpjqpykxhIORBVa1wp/
IURpfpPjkcDw7/360PC0eHyFgh7M3HtKIHJnLOxvj2Hw9bk1r0+ui75AINKpfKTR
xBg7UM+Avt371wfiRk7P9I0q7+Wbb9D6UIzHpTwQbkEqfJ2WVHOeD0DpbrDMeKUm
BIMAaRxRgW7OOBgo042Cn1L42mb+eLUwxstdML7UrGrvLoupgcQ8FmVXOIfUldGw
cz5CdfkqG11612UqfdWwK2n7S+n1OPgQ2BbR4P1tTGeo/eSVKohEywU30UWqfau1
CWlM9xw22Yr0WJWKpqfOzFu5XNknnglvA3/HjKV9/UmIoEZazWv0dK4fkZC3Diet
3ik2pXYAlbC473cQkP54FRIkLOhoZdu96c+vq163k5hHAdCx9+bwv5PEWwQYCVVT
lgVj8TFdXqmy2kpmpZRvt5wVQ87P+GUITOAyf7pEN4I7ghFySxm9zgVL2iNsQqsX
K3D3cpQbb/FJUw6cRP6FWaCVa5ZTX0l2mYnFF0fEWqZSr3MzBoUD6MpgQh2AwnyY
9UPIXF/Y3JO4U8e2BmbfeCA1iI1kADFLoU67m7RC6mkozjwq6TYxoahTt5bB/Z0G
cd5fgqYbxQwllD9yHraA7yCYvXLEtHQ6oTPDnal2iY0sT6nEvM6Nq60q7st1Ms72
5hdT2pgq3L2/lR0rQh+4kqDckZjD2+XJTxjV+H2ug/Nn+sE4Bmjwz46Ge8LMmOiN
YTFge2pkc609YdWgMZgV2meGJhTuaXZsMpd2f8a371dCnyAA/B/kLvZSK60vcrnu
K5J6ZSWluHVg2Q+C86aD4CoKYd7peDWPeZBe5n5VHqvSGUrKRn3P1AyYeRoEsUAD
/TnmFSVkLZVXZrC7BhN0Pjfi50VWzcWx/y1HLa+8C7x86rob3m0ZE4IRg7RoG05H
o2RRaDDruhz8W12TDawrwoMOO/pudVJoggLxF7PU7KYVDy4lX4gaSPuVPTAByAf1
/eauTbEDO0imDcX4/KCTjisg/r/EeqPgDdtb0q0yBfRu7sQO+hRo5VIls2LwFnrc
bMJtxM15kzLu5KpJ+IxaRRZ+BPFsF1ogyC61UeXkLqxk91P7FPmyePSIMSn5fwFK
yh1ZEgVx9ps/aSpxQ9mh9s2a5vFPBSZXbgtLRvNlqFyBiUp7sDx3eYHhcOjf0OqC
dILlRqJ7K7DyStA6eNCt0x2QVPZrdGqjbj/UOT0fvYQA+4nIzSwbv5wT6tyY3itJ
RhSOnKqoxnldFwf920UfzI/TyFLSQLfIuZDgKwOASeErMqTGAkhBdHb4CgBr7B3g
fkFGrwZZeFn0rOOrPegiF7fA4xCrF8ni7Etbx2FmOkwvWJyya/7TZS32XCplWcbg
KRcpUJriNSv1F0z4caCrtoCwnhVcT+DmYDPPN9sXG7HeT36lLU/KZ8VUxBu6lx06
NQRP1LK7/WFTFGHgY375gs9ctAPkv3zcVs5tVjdHlNHNfxODpn/SZoyrGpuMLvOX
KKkdHoxuU/N3N9QN/BaVR9Rvfl7J4e6Gm9UQsAPmk59Y0YmMzUcERW6sIZ4+4PFc
2CLLsHCJt68cm5ZjcY9jaFcTABsIxJjRgKPz8kr4k9oz907GT9Am2pgps862720u
b8jA7hMqK3J6Xm+8PUxGHUbIL945cJ6YXZT7FjTBhM8ah2weiefLMZ/IupToQ/Bj
f0REdB/GSGglg7LmZWZGG2jsLG57UTgZTYOpFTJFCFCgMwURkBF4HX8X+LARitFV
b5SOckFh0nyN2BD/HTyUtzKim8656/PA2bhTULmjw5UHfvvxGxjRZ4N5bqHN03S/
F18YDyPmyr9a1eKhNH6ZNlLDH0Nif/EmFEE7EWNeodAvsnXRG4zBrb8xjNcNkBgr
sMKYNhasP24kwdTCVb2eJi3W2Dyr6v5FL5vXrbYr3Rp2C4GMBElAK1B8i+mqbb1P
ZCsSgWrgXiv7SM1KVVCTPRUbbw0t7FNHrkIX/LOP1WnVH6lHv5qpKqUsoOoEtIkx
OkJW8lqI3u+f4I0M8SsuGs4vk13i82aNaOGpYt7wkrqCJ6SISXFcDYQ9cCaqSK1U
Wtxwh5PBE6RrWq7F0WnRYuJ2aqu7XwtamumxD3BHYSHvAw/yS2jAqeKXGJWYOMvO
PHMD51QlGxF3GpIPRq8eMQMlVpZwOfyI6jrWuwwU4wDKeq7N4Vdmg2AxCC5mdOq2
5kgrA50LZs9EDpl/7J//yOt00MQwVXQ0I35y0LTUVi4Quzjbq9oyDTaw3fy2MrcB
hh3NYIs7tcoW4CyG6ZJV/VVMLGNFd5Jby5nTx13OIE6ugTj57v40hpCCt8B0WaF7
NZu0o3Be2Ggq2hpyr1dDAZ6AWb04kYhMuCKSTeXMViO3e9TnzNrE0DiuSPWUPV8i
uWJQT5Rc34f9lAfWfNDy0zeK5F6xPK6QYXJ36s8ESGRBUDRsidpRirb9d76GnRFi
nZrFG7dlVlgB/EX31mGM4Xb2ZHsDAvOW++SIhSw3+2yASxpkXbxoGRKswzc/ucZF
lG6tPsvN1GGF8PhIjYfxaJNtW2j9xdbBfbrGyw/40BhKXb8I5i+7u6fhYV/ah8LC
+85dP6Ki5DSIzeqjv8y6Qw9eNw7TTczFKHJGFQYla+x8jsF+2vuyCUabCBZ7j1z7
14X9KRqPbdixW4eUtw0fiRdybWhJZVxYv4AcJUbzUmY3QNJpcqnLo+oT55BATZFT
5pZhpUoUI6QUxi4d4MFk8QXZB7qKAltTXJDRgNPckkCJsiWG7/etFBCb/nUq+jQF
N312GHE8Z4Y7kUB3m0nSQd2P+nH/fMsuq5VQXfEvfPJl3LrWJe/fKMyAeEEQ7aYI
G3MidrPp+nWz1m8AsLRpuTGZMz0Eik5oUWluXaQC5lC0SeSSUlHbIoLt96I/YTO1
3rkcfHDhUpYsxBvLsYzECA1JvXiXnXVc+/O3Ldouz2y7yuF5KmR4uzpgevSxR1Rp
evV8gztN6p44sDLu7+lDOlrIdJMETPQo3/gvLJ4C9tOc7hZJjxqioY4A3haE67j0
dwJaS/6TC0XcqjeoKMK/pW/NxVw9Spm/uPQum60tI8UVDnOhuFl29IkHZ7j6fof3
iZPr5SrEBNLQ9FJG9VCXhEAf34cALMxpRotv/Bl6xxrZKZ2fQ5pNhGZM8z/eTbni
tb3av+BQ569RbDrXwFjLcyMeoiwMqZeyoexXtC2JeLWBcbVAusOJBEIpLuchjvrS
eyBP4leQESO5n587jY6D0+pfpJ/9A30kJAaYE/pRWh1cGy9r2sAygjrzpA8Fa6Vi
KMdWht5/oKukbTvylhDCARZ54lb2O3PjgWyggftzRloSqa+FG8SsZRNwfpS3fe80
h6pC5r2wnKGOllrtujuw8v9DBWq8gsd58DcIG+vldexvYrvO0zRg7UyVwdhmk4Kb
1/WE0uX9YxUG2nNd0CNFbwidg3WbKAPFwV5PSWIbjFx4IRz93KcBuieQVbXv1d8c
kYL9zAE27upOLb5zjbooHDbqLQN3ntRzL72zehbOBNeA2LfkdDIMYgB+5DCzG6wU
QwhR7Com8TfcKcgow7H/NfUIqKHhy6GgsetcL63+x/euJRAL8SM9lx7Z1tGJvdSr
lYbUSHWGwAuQfjmbMARQnCIECttd0TcyohGcncGQN5rUEVQmQk/CoNfgpaQas3nI
Hrzx6CeM71Bx2b9ylyC8XiJ6CNa9F9gH4Twb24Dmr39JNOtoo4oC2VmJAVPbbGcq
CT21WA1y4CRCdbE769aBy1Dmb2GPnB1V2OSRGZBL/gdDjQ2tGUNNwcvujwd8RCZV
UHmoKGc/iPpuJkx61CF5XyT9YAVqvPtSswT7VnFY/NzU3/TrGt0tk7GxvfAoneu+
cqHQ2OoLWNv9nQIpYKM3mIM8XDqeqF+Vhou6mgUPLpzdNaQHhje1jdYSl4j/9BMi
MTt9whaRfFMQlF4p+jaHUEZ7e4y0RBS1KutlrS3qn7JLmwrpcLfcnmHzbLQj5YhM
mS7JlRwX+rW/qf9FeWLavruApxKmogfjjXUHt3U2oV7ZHThCPp77ZU848kqC/wom
URgvoMWEg7nMLYwtTT/1Z6ZCUv7WfB+DtiBqKd0AKTAeqkqygHsSzJcxihQTUmwe
FzhshOkExmBHdcL5AZpHFEnHbazYMQvXH4Vp5xHshoNxxzovJYJSfxH8ddy9fYs9
HkrEHVMuNjU3BrrgWBUAHqlX89rqyo/l6yZZ4sPqx5DPHC5CDs5V3L2gQ9jl7TPr
L118XlM/R3kCiJ8zRopbOXDyLS24iwS7C+sFHv5Xz81YeovH5hi4TgV0UbyljyJ9
hH0IbvuqapiV4EGoAlk2wDus7G9SWQVG16CtI2sREHems2Bz8kUBrxleKp7WwIOj
BfG6QnVE9ujxLOsQhr7cCWh6LgvQzRbJeUVUgFb/eAf7Qeyw21neS2zkUX6ZI0it
hNw9irjpftYoboXPL+edLdjT+Fq7PFwmOaZpD34y9IqjHLWhvUUvn4m6xKpZxQPR
cntCWHaDXPJKi5+tTVDOhmpWZ1d54S9ShdikIFzTU/I5e5Wgyz/VxOwfvPAo3XLI
HF0j9dyjstWX/C/sfxmYRWTmElqS6aka+p4ODSd2C905enGcRAeaQWAYBitka34s
hk/ugFzpf2QETU6RUR9THixJ81Rait80x23UkZRhAQ1hJNwSrq4rchC1butytT2l
jEIx0nRStONwA7woBIKrByoPk9lAqouW4AUwqX3bwIr9807xdaGLmmiGV766RGu/
nYkQPDFxW5EuUBRpbX7kfxXxG6bmBJPjZU45vQpxOUCAWDfAdIWgijfKEech5CWA
f+Cz6Udaec25Py7xw1nIIzG5V+YpZeKc/64BOSpTLf3c5MQfJvHI/rJZYulVmW/0
HNtant8100FlNm2yXlYbf4fcVaDhmUQb6afjMGk6P68f1Izlu5aXL5IhYpzpdlPk
TULISBS0syBGXPUx8yEzNUg2SQhw9ykBKNBtkoeFfcLy3qw12+vq9jEL+zM2erov
X70KxtH645VzCGmcnKPKCaor6xTvH1brVdDdiuRaGaH/eu/ALveXTAk1+SKf5A8W
p7rOP65ItF38DDqav/sa9nHzRU/5A8+LJc0SNCzrpqTYyBqSykua1qDR9VRPXFfS
MTN2gvVFEmyMPJJcZ6DRyl59c+GTkbwNpZDEKdYKySRel4Fa1rMDy/or12r3HYuM
96kQkD14alXnbBt54weQMnOjXqemK8dpZkHG0qq/cZoc7zUWGG1wsIzBYN19odYL
8LLhz094GWYiJTbQrcnbYXl6UWB0vpyzxjH2Mxs+mtdmD/gBCgZ/nt9YLzabIFrh
Ey9H4MzHUua+J+XurGDJqvguLJ29ME+wVfdM8njzrd4jjdFCcMQzbs8qlDtFjZfT
xqCB8vp15wXHTtCWSI55MCe2EPCohIB0dshrn11r7KD1Yci9NZZPTWe7PgFXn91k
IvdN1qDwI4VtgG5g7RwMDRSb8vh5YHWBS3FCYlR0VVFDXB2oynyw4HNkkkZCFy3X
5+pCywAV6OkIlNASvPP/cxvPUpGzB5DJLN/OUc9rXWJvqvijacLkamkSdRnra09R
DCrCxyZ8SN2VexenPmVd/WBjw6kJrbg3K2YIF2Dec9JvR3Qsm1zizDp/Wu+wq7l+
HO9WHKHdZbGcOiCFNyvT8PvItfpuDp3BtJQeZoLvPZeNswfJbMF50UotdsBm0IIQ
AhSjqlD96A/YdfwlPhWhNJs8PGizyd6S882x/q7VGYrPuK8/7sD8ynpi4oQ2IBHv
JYRadboppQm/Kj4RTXyD3kIX4Dln0AnOoHfiKNZo5dlsI7SQV6GTHCDT9oz2+/bF
VKoRfKm1OhXkTmaWLt+GDTLlK9WQySPpbblBu+qtk5BYNCSP9Of692hoLKlBqLoH
jcpg0lhOF2ejywXUW35XIvmU7uJu3CrDwBgL1rv4F83vIEd8TSo39oKth+7+Ye4t
v1soP/wvvOOGW3vo3if0P71Up9xs3AUqzy0tNkx6Wk5i6YA3m7QDpEpByefS2MMT
fF1x2k0iSHXp5cUAt/m+/82yWI1FnbYEL/RdLPBXsQxIuW5JBcAYn4qTfCKj481e
w6K62uYhvOBGC94XNuHaw/mAMdkqWYEhftLKiUQ9bIOtuG3H8AUgDcQVV5nwxRVo
9iEvKQFY4RDQrY+Hv7PVzGTRq3zNmXJS2IuiIDYrvD/7bfYTQhy4SIFPl9b9T3PT
yGjbK+Gx1BAAMMBSCpRCvDmeUlU6VWa/ugIl+1CEKm16ndiWSZ5asmjqZwcbIzs3
6OOTY2IFnXaTbyU/9u/gRG6FHXxIDA+hCKpnpjLlcj0QKEKol6JzCIHyLuBPHJTs
FfNTFrZxlT0NgsFDEiIpdlXNvAOcyrHDN1gZscyIxWxKw+8UYQTv1FMH7nIUEoxZ
7yGtR7Xo8iZSdjSPi4appJEwlZ/oy5gFYyKV9ODQK7fVRVAuLL5iMiFZrCsk63KV
hotitbDV/hEsZ5o6dcIif8m2Nti3Gwb7i1la/fZpUH39f2yVf6PF5Jml/0hxkzzO
sh7p9r8UEG/923hCPz1GRp9vYAdiTwkSb/V0gsQqz3iTixf6FJWejkcdXyeg0M98
+b8Oy88qbOGQWgWeaMLrMM1L7wrqkQFkMOdbFaYwybSTUktXAAXFszX95x5oU/Ol
uIA7ZLCj3BEXh8qgfmmrebE04UXPAYQbOzJOTy5ox3lT2C5ppD4YK30WiTXFcpKM
vhthnwFHJn5KD4/3qUB3iWRGLQf8VEvnISGptvcT3EvMl+3yfq3QxYrWvoi0OMk6
6z3+OFNUZaP6B7fgk3hO7Rz+O67iA0kXAQOISyFvFf+jJWGV+g8bwqCAR1iSiqci
OkVB92HCKThRfJj5MxF7chJxF+zjDm+m3+rISFizcLyl278lQxOc8n2G5unImXQs
yyuHpiBxoplTyqeNrbjIlHmCoF6Lq6GAVqO0RlhGI+zyw1qu87mZ8QvJ2VUQi1wY
cSYVTelTvExVgbu7QHvR2g9FuRBouk9z5/2UMQIFiYO1lQp6+YvqYRl9vCp6P8Kc
q2OCcRV+H4x5QhrBmBNwA2JtmjdMqxOPOgPaWIXQaMJeC8VEnfMYeB4NvadA1eTD
/gwuQolhdKS7N7rqofvHtqJqkVgU1Gje/c5JRQ6qKCLCwEDoYHPW0WyMG+nKn+br
IfwIpLnxXnzLcMfG6uewplPk883LvoCGOaai/j4xDu0ghfp5T5NLNvcCjXgVqSNd
cBjN4b/35eNoyB47/Tq5dW04Jv2tP6NJPVaurBac4pfMq4fVogwW8yaIrOubD+P4
+qgsDv6p5tLaeuwanrU1CsQ+9PGwJyp+T/MK5/1JV/yWnEyf2Ri/Uf62wG+BfNuI
AAj+daucQq9m7zSeAnTD3ecqNjcGa/SjxNq1JPtp4K6jQtXj0aTRv8lGK8GSKrhU
3Vu9vRXNZl98ikQX3jdkRbt1+0wwDwvCIOMyjrk+SjZyjp4MrGnlebTbwzSHuNRU
JVSfJ3jP0rqNzwMlmnAPL5j/FJ0IILhysNl1mJ90R5o58VPNKs8MwaP+dg2be2fm
hdvcmfUEM6qKRRhwLvbbmqXhD6Nax0mGmFwF+wrBbKatm0SN4u7r2cBMvlamzZNe
AUwVnsp9YSwS02ReaOqGMlAuR1gXZ3MX6HxE1mb6QJQCz1fxljnG9EysZv6E7aBC
K2f8TvD7OGAq5uiqTH+Kzk6OYlwsld/+0h9gyv80RjyHdve7D4t3eqaaq42nRTvM
y1RrHctVqMEqwLZvN6CKdJvb4JuixZELkXcBIYVFHZK5HYKo7Hl1vIksaMPkqeiq
eBPPI9ylLUyDwMUt2nJ1f2wQdJDQ68cqFjDAQz3kykviwwY9uesRF+KjTS9pdGBE
0Wq9EE9nj0JWevhhiGw42SoS0geI84Pmw4W/pGcZcZeFkbIPXuYjRZAai4xVJvV5
9cM6q6tYO6OpPqay+Q5A3fCEZZZGUX5niQ8RqvR/5of3RsTOXm3W3yVUfCwrlvao
/tfoSQUJljw0p88rSZLnciZbTV3z++iprE2N6AAX+mDxhZ0+qTFdwf8lqNBlJt4t
MaH5R02TiHs9arzv0jRzxi1b1mRLyFcgueXcRYtDXxpxfUC30MHKki8oPrUzfUH9
YnyOKquB+SqEiDfz1N5iiOysBbCqNDABZGKy87Q98wwrtfac3vK+BiEIfn4BV7eW
hwKqGnYrmlCc+F29jDtFB8gEyeTzGANBlEb8imOvzMgzKR2/Ga5Vt6Dpq79+GLWw
orPSPBrRnGOIrxkLt7igNB8qM40d+ZK/ojSUHOqi2X5Vp3+PreQgYpnKUHHKDPj5
mJb6SHQ6riuFxngpUfkeXQVBgDOeIjnYBBJ0r676+8IX4QXVKhRLyFOv6T2COfFy
Vh2bSXo5TWpyVZQ551RQjGNbpkTGfsyxcAiqokTDhFf2BKB0gT0EDah79lUGD4ur
ohmNpFE2O2HPibSysQ7dY9e3beJZyhqm+BS7Cyy0YtXpWwcyKBX5K7mUfhsxrZfr
Fwf2LAQUCOho2FJfWFYb6V4qVqDPObB8Cnh20DGaQ0C1mStNlJD9/kdQla7nKtv/
EGDql1dGIh34qsSjGjktvIzPATZLCN8rbBHvnyGGhmp5kqD2GaYBmBVxuJwI5MwX
nxqUrSSEKr129LSxaq/Xa6p+XGfBs8IU0s5Iv6LsH22l++GpbZXuPB2QieOMZ0Io
RF91clCetTDxe+Bg+3tpkJq/YhwvRN+XsiQwQRk6CWPFEHf7KlT1NCB8RLIrSjVf
5NnTg6vLj3kn916jveWJurvcxF0INmmWD27AosC29wkr7V7BpF7Stnh8fwMUv/7V
2FeU1Zumr2Ot+8hJpkJ7O2bjCvDMVJGJ5dIcGqDXBmTebGKF4rEC6+m/QgRtF0Ka
LgSDkTJ7EQhgsNCsIVQdCtIQdWL3OaKRtquRkHmXSQYGAnb3I3uOMLiP4fngEdgq
gUmdkWpYoOoUMUw47QGk1CYgXLRq75ZC4t7sVkWPCfl9CrAL2KS57F2F8l0srNUz
BcU3iiZUDBibG0kaMlBeP2uzQBvTaqrFioJc1rFNC6BBc3MNj0x2cV3kjU+QzM++
YOIjvZJFHJeeax5Q6gGboFNMuwNF9KJJYkO1OpWdt7z9ruOI8McH3Z0yrTTH762n
ZEWGloXtJ4mKxd2eqdED78Y6Kr5xb/JAK1HmfXILsbHfot5YH0w0nIjxB2NNriAH
WnSsf2WNvU/oKxahIFYsTqw64QkxT4t2kD5lMM3QZxFHHl3MMQJQu+HZaPSsUNqL
YTvPPrMcxdp1NlT6r0oVWokiat1oVrsccSqrzRQbxZKbxbKPN0oYNY8ghPzvCLdd
k8uPpxyHT3MAn7/B+7Zmau0bO/YTzuy+E+ocRUM3Gxd8Wqn7+gV6DnPos+22fAm3
VjULbaC8Qib3p928Y4EPiyfeM8j9bc+YXTgvgkRU27mdVvlkjdA97Wvh/VbUr++y
56YmEZ1TUapSvL84awtlZtlTjRpBzYsZ+0RoUlltkum94/9j0zXeUnN1ymIi3rO0
fEHw5//qFORq5hBipZDqwVACaeegN0INimSU2j82hB/C9SHqSOoicTOJ1Y1ykn5i
uNWvYmNeYxMVyxhN6p2aOmuuNjSO0YJGvG84epzTZ20M0nIdcad72F5wo94t5DyL
dY8GCJ2BOlgpo77J+A9qAaftx5AOrf+C4DCLS4adURGqaTH6NAhg0Y8l6ATTLCym
TM5w9DGnJtga6kUnMuHjCzu9iLH9dUxMhT+tTs1VzAt4b7QQ3ciBmSCJhV+pA1IA
0/yy3oFdCp0HIkiR9VdKXmkh8Xv90+2GJxIdtcVutqgzVqgj1WTzr0J+yQz9F9ei
D2siVlQI3BxR4vc6IzsGJJDPoHjNejB2rTTcnd0ZCBHGP1/iFcTLZNZ0baqTSKz3
5k2ojkdzm5+Hj85Xs4FkjgJulTCwDB6EpFrT5ZD0j0oMLiUcx/NwAA2sPZk36UG+
0+pAp5F067QsqJzT+Q8juEDcCbVMmFrs9WuDT0qvk4co31mAb6YeipSC+jQUqt0b
YGihGQI+sRH+kqwSkQZ2RdcuNNWd7b7qqSGa+8zARxAU06yQkWSRuJytQAb6Hqxu
Y6WwzrSSeNc4CjgLYlf2w5VN8dVKBQApfpWKv2li3GnuQipLFTl7a3uvIcqgbIK5
TMDpy05HbGFdQ+7eX3WTRyeNxKVyPhZsdME4CAgVNtSR4N+BT3fc4/uwuSSi3UMf
S1IfyGCIKNsF64Lq8gh3f9e6TuOuiFqDEBWlWEDFKyNeVCFSctJuo1a3vcVYG96R
oxMPaBccJvvOy5IooRtMzCJjuKDuJCdzUE8iPNDsO9FndPBuLpYD04BC14oligKc
YIcFX2NGES36Z+bZm+si7vlyIVtZFDuPV807CFn30dKZ645R7GZtVPdzIcGvoh2x
L+s3tQUGuxngboO9kd6W6l2zR5LKybKWXU6bWD0T3jFAA4+XYndWSV3sWjHrVjYV
5IOpFvOZc2Pjufq4xt4Vi9wEDM0LmchoWfpcAZbxUIvvJ1evnfdLcZn8R8570USL
BciLmcZMfgvXNdYQBEFPbHm+0W9gk5DRSRYc0zVa7wC06jLs2vTh7OZwIPQW1lxI
mCbdtqb26AGiDZRPBYWnPgN9Lo3x0xwH5SgbF+8XdbWBigVONbwUh0/ushN+twFU
lrT7Jsh5zwvR6xhzCiSfaLx9e170CzaSmSUwu1OluJ8yKrQ8lmSPLYvi9dl4yJGN
iA7hZGBgz3jDUuQC0PVQmLNfiMneevAxcvb5qUQ/H64xWd596gK7GUco0nRL44YT
r5jMQ2uNYTbyHL4eXd8vc9UrgxZgBox4MRv4zqJQpnGsScffGxn3sh4CTIjk9znQ
Y2W7bhL4PFu1z7oTrmnlDnVYO3g0si9wYeYM3UkaFqBKwMVe7CdsnlJFjLwgrrLn
0lrP5DXPbZ5tujzyXincF0sfWP2c24VTGwhfjN6O8bKTtNqleH/X+Mtw79Y/OQLr
23GNqIbNYj95ylUF+RDdGvo/rw9j7ycoji3USq/CQQ1yiqtO33y5c6J5f1qBLjjl
mpl1booBznoxf/3JhHDnDmUuGNf0stgqQgKR5HrKoa+DxpZ35WwatikK9ysQY14w
+iRLfFg7hJ400QPv13PKmzasIOsyEU1jolIyQRQiJebfHYUw30H33NfZeDY1mRq+
bTLGIIjNMcE6m+NUfVuzMMLZtwA+oSaAFDOfEHI4mA57Q+0l/Yc4qLgznt77mM10
Ftm6qjeeNCdveb1VEIB6IOvzWNTnXtSYrG+I3pxeiRJT2wd5/PHRXc9BeEau1kfH
bye/yTPcsSNyHIA0QU3i4yhC7f1Cm6WkeCsB/awQ7K+vG2FP7VCmfJgXZywlgO37
ntK2Nxq9IfMQLNXhL6os8xCtPIeJs6d8ByrVQNqjfZ5czg6yYIg7owZGrN1pvF54
rPHXpE5YE8ALtT+qzmrX3riY3M8JpGXzhs5R20TxUtMSQ/asaDQv9JBx9IUBaEPD
ZNl3AlICJ3Za+erIrFAYaERBjnxQBBH0EOHILqi5rwaQHyzNQsbZCtnulYft9Hnn
5GkqrfDbBGp9DLG9zgE326loPUS3Sr9E8UXZuGYx0EG6bdA142uj/j6K9+Tj2xOy
PXOq+kDZfRFNrZA/PpGIOCNq9T4c870+MmhiggL26WTh+MLenUQp7S41ts0geTAI
ESWSEEdLWPYJ+X/fhMCkTt+R7taY9jPY4PTbLQZvoyZpCanvMym8oMsOzDS9jFwU
+FDKaQjNRbED6b1/ejQnhqY/Pc/dHN+nhIwkWkVYLfuv9q7K573VOw8A9NZWY+J7
4vXC0ftxqMoBbEkya/xj3BHgVWy59jzUVRkZforsVTsCPpbIknZecWCDf2Z/Th/X
pnItwouUE30ymiZMkECpycpwu0+SfafbBz+RXPaEZaA76r3JPrCjODjd7fJzsVYS
JqN5FbR1PnKPFuO40zZw21Pur/NPkMbbkTw7SHS2pv9IZJ5mvfPsma7TCquUuU5q
FC0PK8hRDaLFMGqzWCehUVynqpH9diEoEguzNYWmCgDiRCk4V9sPmtBMUh3DsOpD
jJZKcOhwV6wLP8xo0uw7iLJeHI9BRnOvmjeMIRPtGdsoVya6RyMDX43q+2loVSH4
IiOGeL0jnADVb9JqiZAD8OJKD5pZgSzFcEEZWyHEINYVSHZTmCSJs0+poeFJNsWc
M1C3133MCS50duQDWw4pPQxwyUmljWzeA134GCcuAGrP8YKyfHG0+vvYfKkLqrH0
6Nzal31y8vUpZO6SOlFwM8UMpH7WX79c1vIreAEIxq2GlyvRBxv5P1JL2eKlu0lF
0eAd+L1nm1Mps+pxqa9kLwJkfuJlIhDgO7X9aAbFSV5Kxq74pHx92MkrrEq8Q6Ki
iDeTLILTXCaeBR+aw/D2gKCVwxFVwH6zk/S+eSPE676gY4pxd/2gUCjPnbnt0PNy
hzL7fflQlrgf4lV/+/PDY5sQ//4X1ey83o52g3MMsup+kil2EKnHyEmEJ6IHfm0L
h2hxsYvyXC88q+u0lpXtmw2VKy3vTeZUDWeG0q28pb/e8aYCcllKUqLlF1q/1Q/v
JzxicX399ZeDzCpPw8ja2eYIfUPUmRjA1OF0Eqby6D2XRnGHRZIjjAgBz7ElhFdA
YACY+gzOdoZ0krS15fAjvUt+wK74J0B2bzPyDt21WmOTt36HWMBJ0grmgSzwOWMe
9PKbAXnVnxrvka0v5X80Tyw4hAZu5/n3rgR25okOK1Q1+XkTj9MIV0zM21kr5U7R
9hRI9bRTQLVFa2t/VzEqD/74jGUbhughlKxu1jI3CqsqeivW771T57+ZkSCoGG/3
eNQI2+RblA5rpBZqBaNnqLw45DCSzgpVrb5L6QJnjGJwX/f4Lg29kXSaxxfqunb+
4ZnISoX+uNDlL3llqsV28lXetJLJjeIUj2YXbokOxT0CSirDJp8PuXRwfoOMwlU2
5C6PCVkRaYizIFakjXTBfaRyganDA8gP0Hwsnmep1zSQjt3+Fb5yUlwtAz7OfZ4N
EXhtkuH1JE0/KUWBlGSd4JQC0uRFabIqLyM6nwds6p3yTw11sGwyhAZkoZbvtE5E
pooEqL6QVsCi48z1C8JcRPYnxyqR/6wonhDHvbHE1q1Eym6QlXgLxydOOwzDPzFS
GygGgGvSB/ui5HkJhAfuJ1qMfPcSmaRFSzPDj6BgofA8TvJIQEmjIe2DIemGzxkx
ZAULvWpobFZSlSv24PDyRNfsvimqGaHlttQw2jcxEBuieOtNtnNZFQ2m6v9WCqWs
w1bKWHmKckOKNAa/Fggqd2TolgHwmFyd/K/kROzBB6klyvn4uOlyOkbGgT7jyQiZ
LtOCAT2HIAECFuC/52bmflaOYj+hE2PlvcdY7Q4PV+g3et/UFvv3TKisy16fj6Yi
UXYct2IRrisaktLj4ih39fZ0kQw6NRS4OHfvW5zhrmLlM3Qvu5X7BEIKqABi1Nc/
5VpSIL9FJTfXUz9G9G4CQOtMWwzV6h/491Eeza11INCw8qu8PrLB119avD1fv0Hl
0/Rpqc/jtkSPhX+hOla/kjh1fxVh4VT8akSnEmBCvcbjN3Ko00cIPuFXECBUGzFS
/f60x7MPyC5yeWsdlotqrGvX1ofpCa6OjpgK2ikqb7f+5boAkQX4CHhmXJXrxEoE
emEJWtCuG6S9T7fYmbObvHS+DrScB75Dcqy+AcopOZUax4IvC1dpa2H6ECFjCv2I
cQh1/ho8PNzylHANOcGN/Ec+/+W1JD0m/I/3wgw/eoCh9Jq+dJy26Xs7qll6HRZ4
5/57fSnYEGKfTzKka8T1uL0xE/LowIjs8TX5D4YLFrbrsYMHsGot2wi533XcTs4f
8YSMrOrGD1bHiUNuAfm1IQKH9KEm2SzfTCt/AeywfYsgtZx+KyWYY39aLVdNIymQ
g8dePcKfEwYYAPtwH5i5iJN62d01W6CrRIJ/XjLoYCM1xeXVzQlBfcbCU11lKTlA
cpRG7cg6Ua/PgLacbwkPWTbalq+knTjC0oE3b07bVe3URjwksM324oraM2FW6a1d
r3uunI4pwlBDXmRVXXN9SL9v4+f1+yk2qcOLCqw9v9D3f6Z4vR+k44ZddVM4oKja
7S4arezyUDiwnUBOTKhkj+lQk3H9vhXTHuNZrZzVoT38qFx5bUEiPy0zWK+FVbAV
KIjz891ROHtUmSsfkme1/ZEPaDkt7E/dRiOJjJuPdUSyyqb+hXXjLf89W3lioGwi
MI5NL7pgkxxu/ykPx20Z/hKv1pX5Baswr3YGTqdQyR2Nf68oG960BVPJpDcPX/TB
4VOi91PP8HeqlVPTQ6T8jEvcHWjFr6XZrYH2sZGSJkz7/aFW5F69KMh4ENWnKx7A
godOW18L34KYGMWRJuYd//xYn663u96bEhSwJwmyDBTZD9RlMawMGv1qGCU4DYNG
4JPUdtLwFbEej+BQQR2hu7PqsYrCh2g55rtI6bjKGOh5B19N/o+SmT+IR9hIc7Qa
uJGzIITEu5ZYaQPCzlHw6DMxEAMSlbCR1hdtIBu1UADkqXMB6G/X1P1Z5L3EaKMr
XkMzgkWXc+KFXoXZxx5Z6IpLakFRH0sIXSy10WlDcRsJX2I5tFOzArZJ+o2yUo0E
9a/NX9aoR/qEQy30Y1eus5CC9z5hjz3GQzVeDfTkpzFBgm9mGJQYvKmd5UEUZfTN
2zzPR4cAkdVst++TgePv5dal5L03idlk50kYuRHKoNtM15mI2HpURY3DDX5NLDMh
KPQ/ZO4F6dXiEPka4mYGAOsK0hYx4aY5GHZ4mWFluu3iB/VR4wwcvUwGz9v/7l7v
mWyB5VnGXgSTNJ+dObyCdazOvCBukUPMmmyOCIb4i1bR9Q1Iq01XkDaCspJlbTCy
pd8ndXe5bR4RGBw6AAz2x3JS1YAswFjr0odwZu6ZkI2GHdp18fVBQcqgiNXjtNku
x+3sA4r8qkc7FVNcs6KzcPR5XqYkLK4fy1EiOhzv6Dtf/ygZc1mwoaq6+Ngp+xcb
6fdylaMvr6eMCjXt93DmV/jHEnO9lIEKh4alISMyiCBh8yOnmB9Qunvrf0VQ/ug1
Gl4VoVwJvSBzf1oOdTZtez/Esl640NsAFDir8shQ4Sgeo28rtxwfxZ0h3kQl8Nut
2gjWpqbRcEOLuRdljRH9TLlCvsLgJlqF/9rITQdJx8TnEQjQ3h6SXhSrZsw9bnBw
SjNN+n69dgPkdJZFhzDFWzcElCTj/hFbK2489aTJkJ3qLvCnaawW8GrzQ2IxBwYL
dvJRhJ5oOx1z40nx27k+L8kOxJ8sbw0vyLcASihsLukZUsR63lb9hVyHdy7Su7c4
vqlyrvy83iayMpyh+6DTo+4lZcQRT/bpq6JrvRGKjt4hi/6hIYPQsfQb6hP4hg2/
DmzF7wjAaTjKWhv9V++WSUFqAiMA8hB+Tb3WxXNll5qt8BuIVZ1n/Q8cFhwK1WgO
ELfMgfASJMmJyVnJgY37BPPhcA0diVhDEdrt72/mw5wsEJq3Hhedx9rB5ZAF22/b
CO3HnoyKysZZlUcobr6rfJS1eO2XGWrfY4WtYfMl/9t4NNpVqyS1VIgMwR24ndem
Lr4uKZR5t8c0TdMmo20VwEchXPBb12GCur/sd3NJZJAlg7kE1FP+9+DVQrivZ3Ip
MEl4LN50d6iD5fBpc+amVWdItzVskO8/+xLq4PGQOXcDS/Jo8dCu97+8fU0PBcdk
W0SW6gtmSqTSYfBrlizW5ySEWq5IcBhWhKQwDusBdOoQta/VSn9+bA2F5xP6hVKM
12bXoPG8JtAR53S2gXRyqgtTPVZoobjxDQCDlnTsXb6QRDsUOEhTeQKdkZWYMqov
bFJCk3u169bDFeTLw+YMY2UOeGahEO64dq99hUZsFT9fbwYvSSaCVTebrnf0fDK+
dCae9XIYHIDLxXzBNWcLO0vb9WiO0kG8/jVEs4YfCTPJxzsJZ8v7hzhBfFlQshGz
2JJEKbSsRKes4oY+y5pC1iXosEEbMc0FWzxePbpDHpMAI4DHwVxh39irN7AByaSJ
A0BQFQShQ427yc9hybm8bvJyraaR82gSyw/6EkYDbb6qcLEEN5ZUnfeJ6BcRWTLV
DOn8pLPa0qhyFUpR30HpJXUgOMjt5WV7atg4+Lv26p3xtU2wIyeOv38tX6VY6eyE
CHKpW9uaClwqa3noqzPawRXT/CH3gjXZ95Pe+6uFQXR1wCmd16tWjQ5vcusfMpxV
XvIo3jf2C7Zg0aXOPD0rcS7DLIZhtPi+J32/I8DuIS9aHXMJSkMRAe08LKQhP8eh
NqBjOuJ3NE9D1S0Dz3oFaSKUiu8QJhHhjRb3FzwnGiqJ0IW/a4FYAV6gt6/s0lko
xot4Yz1FvPU6ZgnC+jZBfOAHZsSzS4mbbnpBAFfGxX6xEpIWOWB7IhuKhaaNuID+
pAS4+66EuWauztm47bMGBPQil96QfnOOmXpKBcaLfylN5J5vgQn4gL8oDKsTFYnd
7gXsTA4dO+di7gRY7GuCPsYERAiaH+rmLpLEAnRriDMo33HvqbnxmIbQUP3w8JJ2
vPK5VHpH6JByJf6oJzXWR698Zqn4yiwghHyAQILrgOKMYfVGqNAzJiUfG395uVSp
hgcw9gaTgjENnV4HvHIpeaGd6XGjGupuq2BykkMwq2ZVhbeeSJGrF39x4YH9OciX
VoUYbB1WLjcCuB5j/bRMJC12HvVZIXFsGNcuOImesCtKBwU8HsfgCXSOe7ChqIJc
LQ8KTAtFnyrOMmng2X9Mu7iQ83nkbqDcEJ4iSSRsZW888iJKm/nhY29z+gtXIQW0
tOu5bhKJeX60X6bSh9Oi9oxORk3MP4QzI16f1q9OnC2O38lWCOC6d3hR9jJwh9+y
UmdurXL9yEiaYMt4M5xHJcG3M8EwfVuctRRdn/JXkg1yZPNfBhqusYwXPpuGA6ix
6/2WplKgAW13T3/DsQTNWMF+ZaqX5HgEuItlb6gE7+Jj4JS5WOk/5j51DeVpjtGd
HDO8YfAep6Oa06XsCe7bcV/Hur4gaQD6JpkV/BpahvySTrENGxHcdS6Hkbq4M2DU
L/Kqmxr8+FmRb458ujNyBAcHwltsaIfEZ2FFX+CNqlNfnTgA0QvqhC8wogvHE4A9
gQ6nh/5QnHvp+KQg5N0IybmJBffl9aK3cDVZLJbQPnuixVwXVXb9M5otRJYL6rzF
SVx4kOc/gixXdx7mU4QhAzwon7btdbltueMgL0FZvrk3taB3NXeA/LEIdnQtt+X7
rCxKhKW+kqrN0OxcSCTY4TtvzA9gJv5dwhPOnyCcREijiuMk+llw9ovHv1sIbSbX
uOV+dZLGcJYuniQq5zk9AnCXMTuoqzxvP6eK/CT9JgBWQGMyNm/e6tumtzbRixrD
9cqFD00NgfqeSGCUQLQ/2zvHp+bNwketWZOCUl/Wkoudhx2Qxqsv09p+T7DIpBSV
SWZFI6w5YHvPkFu93UtKDyR/2m/e1jpyEXy38SWdUs3MwkZqlgE5Ng+1zKPl7eLj
yYtaTvgVQ8cHqr2PxaSBN+HL+8W/MIX0/IWKf39lbcrjz+2RO/Pf6mNnfMtaP0wZ
ZD4Y6k5IUSM5aRKDQtvKxiTkxyf4LB4U8D6MY3VWSR0Gfy7zxxC5KxSKgVHd5Flt
aRpFaT64SpoilvGllN85kJHhpuVwDxQmK21JtdOz1rsOuZFWHN7kSsYg2CgmtWnS
bQFXFJMxM11JVusFs0UcSZGzx0xzUEjsHZ8mGBpHo7cVehSqLuC0LJVVgHNV+CG4
SV9qGl3sGvOEoj2HcI3QPPDwz95imPXyAO7ZjsCY6wdZRmA/nlGVB1p6Odn34AA/
SENsIF0CBOK026DSggjZo13FmD3Vx0QGcwIj+pdiaIxEeXbc6AeinBhZR7Xf9SL7
vlYWFo0yoJy8nyapzbaGcScIdxIjys4jM83sEdoBtZTBby9Hy/EdFFHR93rb7oFP
77lQ9/hF9Fbv5Jk1D64Q3xhbsAE5Ytn7osNLv64K9I01eNJ+QwFSI7XBt7pgaAlV
BJaEfDDZPEYrvFWfTe4kq5L01fmOYFI5n8G1sazk58GsUNPmsDhV0V5maKwoX7kw
JkcH2JLp/dXh6f/QUUNFhifOZVsw2SLjGioCGctQrwpFUDRR5v/oK68/vdvkQ91a
A3FcvvcQF62sSQMyMeEgA5V7WRNlqrr/XHCMTBMPv+jJcRECW4RN3SlfcHFtgrpQ
EtpxOY34s/jE5TcZK0jYt9xr2kTkUwqm1TRenBFSFtbL87ImYLh/RiB7BEcjuFOk
D4kfBK0L3x/f2tiSLvMQyD3r0rxj4IfdWjFmN9SmNoRY9+BXueKiZDNe9We8P3v4
WYowsHmAEorpt0b8Br5wISRSGBPUp5usCd9xymcCv2I4U9C83yNgN+eXNv8jzxRs
KH1LOgPxba8K0pGHVsVkonYIoByi1+xNNXDl35dV55pnDhc1WDHXunpRxk3V7GwB
VTxyUdL5Ge6Szx8t8dVmyQe+Uy1q7uwORFvZ3RZAAaWmTSMcIG+17YnzrmFCfCCM
e1gGXKE6yomKWlR2WaYgXNf3TICpD2p/JaTmycJy/nviNNih7kjAFx4bEOqLsTFi
MDPNGeEXoMDjlcf5Ki/q050it/La5OSyVBNlXsACJFYjxKH0zTgdxzupetBhi13D
mE2p/BR4XTdsL9slBv9yMjeptuS7Uon12w+b3tmsfa+iOmWxminbOjiMLRHCZM7G
lvnUraDV2+/g1DXK71gXwTIilBjN85Kes0sliwF5EwlW5/LEoBgbBOdwSXkcqSV2
8Ku5yBZgAYJer/KESzMElY+qwk3UkqyYVK8E0DNhtoL/SRCIdFw8Z0EqfWMi23ty
e1+/IHZDWdt6n16NFGB/7sNoXMKzNpSBrLpoG/uaiQh5y/yUQ4SFKihFSXxnokq1
sTbV6A/XND+czf8MXyjPGKmQ9aRU7HoH0ZESo9lX7bQEJa/ZmefyUs5eaSIClj7S
J+2gtggmBCc1Kw1R7q/h61dGRrr3sB8htqQsOj+MRAw9iVqmlIc0nUT9xPVt/fg6
JIXX6NyV3tk+iF0Fj88nsYkMi9UKi9Rt3Mn+/jfAHrlWUUg13rk6kpBWKznrZkY+
zsPUpvICKMe1ciaVR+zsoKUwfpTD5kDELjRmarriSMTQGs5FHCw28gzN/cRAZo8S
1A503sPDlxc5HcXs/dcz2hKdahDzWw7DgHwisvjx4DC9i5MaQstLhvxOUgqGDUjW
WwV4l3vUOWbjDns5Nz+sAozWp9UlxuEY/yi2uokAP+Fi7FH+TenSbe+dt25UEVcm
2rBtYq6IQAzlw/axfjJoIn2F0ikEh/30G0F6shGfvQurx1xw1STS0jBor6bmOL1K
gYJTZN7cErQ4aEbTw5aqOYdEcRRQskfPcnJwAJoCVa2LIrxAql+3QlkDEUVOdMB4
ObjYzRyvDUPtGsujttZJYtsvLXDop8qYTW9CkBxpRpmssrCrLDehvKbQPEmX4KpC
9eJWksImMIZPCfHFO3gvN954bH4GHtgjboLm3S2kE6sSmqUoUcq2TeKapAf/vO2Y
6fTyhUfEA+WnxXsFNwiDd+uj34LKj4Ky0pHynCZBlKmkhLz+g73jxjHEWo6u71vl
tHneE2j7+SJsGqgMfcEb9KJGOaG9zcm/8pIpAoVMbhSzASH92DKeZlNHBv2Cdeyw
TBccPZgUnMAZ1QuLio96yixxrP3B09JHnvXqSRqVtHuVDKR+3/jIMecHTfzF20T7
7rfmpRAwEHRk4B2DTLlzcP/YmhfGgDtQdlgVhW35gt/Sx+42mMAq28k5Gfj00ehE
ZVnGHR0SdN5aLsdWNItZUwlCEJXeqW8hoRbgspnglJsdT8bdfNdYXtMLWzgobmSF
YYWa6hzSd1ZPGizUjv8VYtUnVREO7xytlfc66lQnQyeHFQCJKtIA4cNZvjIogx4p
KdQ6GohzQWAqyq7Gu5ixIJJGJhMnoF8/yqt6iWK16eKPABUqLWbcKtP5VC+6Xcin
eCGH4gTP3M07i8spfUJchBtkUR2R4uZTzrkH+IKV88p1cE9U+xSahx2qtEWxtoBi
nkesxU2D3dNuUoEI9jEaZYH71hjEFaXSSvn86UGQDvKeIeT4BWqpOdCMW1+9INsB
e+65805RPC6V9RURz1oRGtV/CfevmPPHZjlXEmnIP9X53wbvHosKT1ILTamdjsph
rgxdDx1tOFoU3S5SYGXIljf+zDQ1L6HghgkwoKfF+B35Fz0ALf9iK7pmo8xj2KWI
JBdxL9HfxIqFT5Ppu3DH27FE1ZJmoY8aTBMnAfuMtc8dZ0zepJtnGEMMqMRKnjlx
G+kwac+dC2iaRKwsDTTmvT669OtNrKQXNdaUl7bQSS2rD9tqEJImQS6wpXkevs66
PCGnFs8rAG9Or3QcSl00PeFshJCvpPCEQe5/hBBAG10uUaFPyz9accDCJBeYSs83
VLjBVLgsyQ3BKw3mj35VWLRAAbfXcJjV3qVXDjfz2jiDZyQ1NnXebZAfiDWEJQg1
99jvb4fKQgVlQOGJHxVVsJcC8LnV3jwUJYoApMdOtj8lcqK8D1q9BlvzI2kxOW5Q
GLi8pDWUg1CWDogkgWXFIANkVbqZWzQYBy5Pb9HufMCaZGhdqIJh/wT+BJd7bMSf
GEAAWsrXeDge5RQLXL36v/oYKer1gc0fxKsyb6qmurTNvAVwVP0+3v6G+LzBeS/S
z4HhToG+Mpl36Wd3f7hAhkJSkKlXT5sbSIM8kf2WOtbeGlSwRMTeZnNoTuteAk1h
D5BMoOu//fJOq03HyAgrk3l2ABcc8YP3V3Y/jDy4tORBRVz/FQPyrMQAYkfEjamC
NqxUf9gWK+Lxaq5p0GnBNp6kYoqHr+TEM8oGm2ZdrMEm1i17TwjNLjqtv25rpekB
CieFnzBawn8w63anYRVPcVAGl19bqOUmGciCC6bvttvxQfGNIkCD0ZfOOOXhZLsX
Aw1Lzh46VD2l/sPutIWJahMmX33ulF5P+cmZztXdgr2WPrMd1cEkKcPp8l59VE8u
heWqHBTE94LjyBZAbyfFIeGqVdjrlxG3MBSzCj9lIwCRKGc6jEtS3kH0qTRWBuon
R+6sDvwPN+7X3aIbJREzh4sWv3Yl/21nYTq9ZnV60Dm5WTGGovZjOTQEgcodlSds
sLvrGu3QWYsPOMGP+jGEvbLq2GPONX8+yc2pPn7w1uEfVZeSLnb7asLIxRuQf93q
3KLLmqvs3jZ1bqzG5/fJJ06EDRv8u4SWb0RlJpKCucioy4Xll0Zf53OKr381JDs5
AonTKy1pKBMiALzgZrJro/H8bP/tlHMyh6r0IazMMAF2zej1TdnIcvCTDhYybj/2
5CKE2Xg6ATkKFEbx8r7Lo3TEADOY/I8kU1JGuu4HXA5lbMze/0dYpQPKi4poolcG
RL/A2akL0MRbdGyUHGoEE7sO4BCCu7KAIaocA/PTVeYxwqI5E4y3S2i6EaNJht/i
hv57lmJVY17aptS9clZIqb3AmES4c82AgsZlykXRhkC5ywyKG38FaZyVNIykUCb5
MoiIYqYCEpU3KaPT9PcOozzwZVvu7uui9kLF9PxeI6ZW1LSW4jOv0Y/ow6J5xXxa
5d+OZ+6RSZOAdv5X0ENroGrgM3SO1SFjXeATUyWM/7SGgzSfI/P3AKKdOePs21/g
723GIWG830P1Jsy5aDSfk0mw4uv3XrvLMsl1TM8UFJp8cZoZn3QXGw3zIYCv093e
BZxMTKXRkQj/tnmwlRKe47z5Zu6+2A7tcbmZpNlAZTUfYG3E4nWjaz/KzNOLTjj8
m34SCg0gnGB+TCfc4+sEnhM/YOyK4TRD4uyKk3Fc8zNbbn0A7h2lEGEOE+tUEl6/
eCV3e+jdFYm+WiAG1BQ0cFQ4yY0ntbgHZkYgg2OEmhA/P+16zBo7cK7shobK5K2H
s1dZVboQkluTAN+m9XOsjhUY2iR1mJYGgq82BZxwroOTtJ8HbYwAjtcd69YiFcx4
iox3iWKE6Hqv1SONYVv833i6urB8/3MXFwz998N/k/Hz09aOAt/leG4p2PnI4KhP
Ve/S03fKgwmVD8LhEIkk+bH1Eo8LxpITck+lzI9eRTfTvFDiNHntFNVfsrAm4+EP
UxsNofqRNngXbA2MPCYYwAVnbSSkELUyOq97tqeE4nH108TiL+C2kEL7AF/y/pJa
rrf03lR3LZiA+jU/P1MZ1ivMt7E3Pv8u0pa4m77LBfIHDxOF2Aa9+2FoFrSp1oEK
wIJ5CjVmfMotG05lakpskAF34EjWOQtT5y7cCM7EYNyTO1sH3/XlOF3Woh0zH6rn
UANAVvT0or9HFqL6LnSEhvJbO1Wd2FakWdvIeCaZAm7vOMjcgXTvGlFeHO5Hp0q/
VsowrNpgAZJes87PLTFfWvKRCS34YXSFI4hT/Dx5Dt2KxCUVgXN6BnZrwj/msbS5
vwN8iSYHiFK93NX3Xw/PURURnHzrka+hlkidRsdz9w5JdUBv+NnwzWRDXxN92oDJ
yW2OwhkB3Vb4Li7GOgPmTeMNuKOKh3esza/bpQDK/T5AU09sqMzb5+9wpQ78Y+fr
wHoQMvxKzvu7CP6cWcs0sIbXkfcW3EkbQEbJQXD9lR+LvPv2+NNWbkISiFxDzNrW
z5O9CgDPl7GxP4RXSHS7QgMAlcGmJY91yQ4Ma8iyx+j3vKkaQNtuhhQv2DXPA4Av
GA19rlu/UgdKQN0/bnS+P3hBN4JTX6pzkACjUVVA+IdKBoDrtzH0tk18q5zlFIyI
AY9Sbmu1Bp5xGFK359Y/4L12IW//wa7exGO/t2ysTuGH7ZgNV8DHkKgLx3yvhNOD
JiS1TOyGp1sIDoluFAXT5+2n7pfCaWWN2zN9eQkXIME+0knYLFhfuurXgzr+taPE
HhnpbTQjV4I8B0kQKoSxWQLbNGIgW7zh3/n4B/t8oSU9LXodu+TuNgh8PV6OJCLv
mda2oaPhB+dVtynvk989UgaIv+9TTxaLPgz1Ng2U974+/oR2hUcAM+2fqMURo6tE
iuKCo0XRqMbgXbm/HXaXXyh18s4xbFIF4NihJqE+NACCvKmpUfB416AAn16MTE5Q
FmVOJT3+m3izV8M5PoM4UA9TClI88EPwY8TSbWBKh4V4QNK6Ha3fpFQC9GY0rpRz
WzBYQVf3NOSIU7AXxzP37mQGICTrMzGux2AiJh4fWIB9vectC9lcQ9NQwnVvR+OU
+X93QJfVFYLxRyHsgQJnDHSKD1SZ53CfAGJ9QZOipdj4ZnbkV3arQEA//kfA5KkK
NjtZsCGLvzdM3Mj+Q9ze5WkA2kZiCftFQqent+5juwj0InGuFqus/WIQM0IhUpQq
0zv3H+2puQoHa2kxfQc4RlR4vR5MGzUVa2S4QAlfG3xM6ej323C4QOFoAtjLDaQB
3dk1sVpG5zr/b58xDGQjsnHvHBMWvOA2Ce/aJpziMpSsU+80WJOF0q+rIJbiXV3q
B3QrvVB/vVVw/rQCBSA5meBD+prAMOs+hWNNkVSULE85DEfQYXeQjgEnYI3C3Pb0
YhafDd9pawZyfbu0mu9GkxqnQP6Lr6kPadvTuK7K7BrneX1L3oskM2LyVS3huort
kDiQZcwcZnQEtP8WdUNhm8VFtc1GTR3ydTAT8lbtSwERvf3pGMSKf/PRw8gkOFXr
nf8VJ6lp4Glb8pd5yWZs6rq/Io5TaIQ8DzXUdjiBGy2OKtNcj4MuHyRtzARFZRsc
MwiolawaZpDfFhd1c+gUAfxojP3IyQWO5vLxVNjkBIEuDjyw2PhliYHmlovRhBA+
eOwrscThFd7SV5NYdHO15G8G7GNHJRNGDOVfZHcISuC/Na712uMu7ajpZYre1jsO
G+t3yUFi/+7dV2NR5hkpUlhsMqxl5ZBoURU44sg/wr8/j5cUMa7yDdQl0F2ImKYK
lFMabIF/H5YA1rqWBWpPsHgL/NRxMMINSGRHwEUezf6x0XU0F6xK6iZuzKQnEYMJ
8xIZhn1+cLxEeJq9WounCydzBRx0g5lLDE1RhvTvkP8vf/WCEguC/BWLafLHYTzZ
2RBPPr9EAz7s87HRLEGiLL/SR5UdNxRCr96+I67lmIQH6lKcJKk+YT9xX/RAdc1E
tdwGx304mjVuGotmx4BzkC+cMSofyfzu4q6gnS4zZhzp8Jtrr1BrzeVvqsQ1/YGW
V3ISUvgeCHDNZ/NlpX3ZBUxgIbizQoSX873WdCsETHI++KAo4fkjj51wifn1gQsB
ZPjWT0/2C2Wr/Xbu3Q89jGyj+qNreswKsBs2wjNMKZmDK1MJbIUIac42l54E4Kn6
86z620FWKAGt0GdewZ+w9UxperlZ1seBHp60RE4zDSGNh1amk+HzWo9qil47cbDm
wvUWyXXlx06vCXZamQwtG0vQamQ74D2DvR4pOWm2airY7l5E8cOPEUzUppQ9dV1f
ZYD5ss6omHSt8XOOQEH/XNyefSmTrfGGJ5nEQaZUpL37o11T27Sr+FGe0LIdYthv
zlHqQ+e4x5VJiVPXsvPFlR0v+Dnzn2sGsfIf5tYXrYwRMsq/PHNT1TP14a14loBI
q1b7x/zMJB0GRWuIzyVOAKmqzAM1nb8S0WtFeJT1iPTsS1BT9cYJp5Y8K7Das7Eh
gE5GmbL1srT3yqqfM+W5ND1FKLRXY943kq2jbrlABU/t9/tqxTVmTLbznave+9tR
RAo4QUdyn4M2J3btERetDTBl6URuKZ0AA75xtxGRYTW709LPdpoTBK86oFg7S/Yx
B3qtwlzWYbaNYOYZNdtlgGTMpVx9mCpoHgzl4/fasvis97Mo2LkueMWo6E1/3FSM
zmukNEBThlBudXbkVUbLdm2Neiz5BbDtC6WF8xYcV9739/DeZSl9CWDw3qC/xtO+
FmSnvqW7RW8WIe5pOVskYeE4gdhAlMMvgwGD1B5JcOF6SKFibK1mtZBOjGBE7Kp5
Gx6PBHkHyQS5SmJQHpqvztKLm7nur30IVDpfunuHPMgobPzUXdq4XLHWaSaOjYd6
ksAf7XsKjs5YBzSoLW17iLMX8GlBzLixJDFVIHNgIFdxMmOE3OZJOTr48SNTwCY/
JpHInMCYmeosiK15Dd/SFDj4JehFhnP/1fwOQSUXRTVeMnPyp4h4JYtn8/xcvKcg
t6XRH/f9KSnf70p4z+2EzKjgeLuBJmccVBEVFdj66M5t2wdzXf+NhRN07Dd676zs
/e1CHxsTB+xKjm9BYKWsa/ihu9zTwnaIboqol0rbS5Z+LZQNHIJmtvWEjsQnE1+n
YMEY2l0hlOUMPDKUp4i6jBux9LHeN9EctUNi/q/OxRm1sfZpyOHrqMIg3H3S3Ov1
MlJTFl4lVmXXX/l3HZPwMoAatAupbQ6DnJUm4yrUQAVsR8vtjlmj6E6OfpO8BWwr
NKW5iWkHubqAwZzryUh/h5/XkUFc3pYrMzlysAPoOxJFy8bJ9OFWVBYgvETZalB1
F/SfhvLwIQedsl08mAiZnt2x2XLyJp7wW6lOmywrvkGe4rjCtYYidhKnRK2Y17R8
tVelHH0W3HmbwzoauncXfoycb/Bs2+XO+2lygFIwbs2yKsTCPxXSh+F5tY6zrbSY
nXJ9lhiezvw6r3DDz/VzHUIysjMWfrSzNdGInin/4Qd7CVJmW5lef5AcnP6mqx9r
yOiawLAzGoArM/cIwU2016GcSjzPt0q2g4o1MA2NkoQspV0XXTOF/z7BnZbvvYaj
05HC6rwYmrg9D0Kg1HPWJRSUhSnmOaJswhWTCjlBhImTXZBkAcupIb6ztWt6x20n
ea3JG64jFv44P4fNs56Bt2AwAMc98b8ZIXYsK5X+yW9OHDlZ9jqbIskzeEInvRDB
a1KFkl3EftlIyqvVl7xaca/spGstO+UmSzYNgqg2abAnd88GdFQu+wtBecA3I0Dj
WLFsV0KPf8ctSy1cBzAKntQOtSY7fCBMtm3r8VbY4gY20w++vqxYMF1ARJMfh7VE
9x+8nnQW+l2ZUazKlp18dFlRcBhfqJvLCE+e46KlQtBrBE4Y+USAj9uZaFQx5/79
+9pz1VNLWLrzUCKwybF02DipccwCVgJBgoJKsGBm+ooHRqOdiZriwAFwlG1e9odw
6ySCUn7rF6v5GdPxw+nu1dBUdk9jKaLEWMnvKcdH9VKZRovteYnLCauYfwUmj5QS
BbTvAOpcapmwQ8RZyaq3ceNLl/mNSykSS3pvjkQn80FlFmO4Tqr1Pnm0dNkQTcbV
tmuF6kDwLD0SA1hPMf7aedsgz5pqCYgkuiYU4+7Z8gLtCLwZrE58kKTGxIMPAYcM
swYVHfwIBX3Cr1UC6whXnvS5xTuw0C9WDHcN+V7k56GdHK0Um1SMg67q1kTQfjf/
Y6D9ZuWa5eONlktQEA5zeJ1W/Ee8ekTjQ2KfeyASrfqeJFUYh7JbEdh9aL14ivcJ
fNQzxDC//qOpCSsa40yIKe0fzlLzAv5I6e3ADx2/nutB3vJnTxXuqINO8Jex5tcN
Bwlol9fszg6mTUwgOV7nDa3CPIPV4X8YPF9FuYL43Ue+rl1ktb2uRZtMz0s5h6yA
gMTEVdYr+mQT6fWJiu3hfmARzZgDMcvSsmbD6lZT+7dkmo5VrOltYHl3baFYzkRX
fGeHFHX7g+2wrDBfU3GTxLz3JH1dfGnuk2VRLZdanLsNzVI7vko2EO4rMViNxSLP
MdVCHMZRE0AsOoc5riMq1LfyQDMfAgQxOX+HceFygZLvD9xqQZxpWMNlzfOjJq4c
E5fo9C02nm4dpQwcqTDaO5G/cgn0cPYKxpcAM6tz4m8x15d+iP+UTs0aoyjLl/s0
/rur0qkR2FhqG8YyMepq//4YJPKSuU73bRPLJT4h20Y60lhH0dPmfeU4pjwk/H7F
Hfgyx2qda4ysX9Ai6h8C+LLSH0uXRwj1NxtDQhB0W2iS4twBkLGNttYfV/UioQNg
xOOlSQYrvxTwZhq8JEjLP7jDFn0WYBIjosIHsr/kWLkikJu4y2YhF4xngdgCwcbI
MGsHOyUQlBVvetQ4i5WXV+m8zDItzd5L1SdKPQP14Yvzqdyi5qFsO0/sbTQftlny
P01+dzo/oYa/Ha/Jft3u597Lwj59tFyxiohb9IRWgzfOhfAV3UGfFlg4Rs2rgcDx
kUaSsHZVp6GLNHJjxzl3jUIOeuCDzm3pnq2gWkzOQw8FDL0osyR1GtXeQzAg5SmD
KP7Zm6TnhEsiEoqxx7YEJ4CiIJXqYEq++ImOG5kgZ3m49ijWaJdqXWcMmU3l82O3
HMg09ZzIx+hsd5KO78MDzEsFMHNgSyIj23zMYH60ubLxAMqa3zz52xUbJh4waph7
z0ns4mFALJo0VKCpHnPWPYA/Y37Xoi14eO4CqNt78WwjOrU/sIZJ6vN+tRVPbFVU
BuXLFgTFl4zlMWEAoO28ertZmXB10UXa+96cf2Z3Tylazw4Cvb4ToNy9/4xeuV2B
XAZghgu5ypvxP20UKN4KVQgDTAsJoAw1VZUoWSBkLyl7et2EWvJkHYpvQetxZAtE
kjk1Pnv5uBTCVW+Us9XDPD/oPegBzpeqoro9CFMeyX7QP5G+IKY6qJDKsNec8Glo
yP2+Vg5oNQIsO3VMCy6wLE03WXQ6xHoAIG+GjlBlVto0Oh3sm86CMLWyHlYkck5D
RBZkO0Gzowm/lv5e6/tiV3oZjKqBi6aQ7Rl+rDyAD4h/yh3jPI00EYgXYYaUulNF
hYM49cPlGwmh77KeuSVWJMWk7j6KW48HP0kc4kfpR9l46Om6ohPPxux7DquJVMQs
/pj/W5oNRmF7doZqyuiNuhNp7KCTl2H/8O+YauUVW23czAKT7IabYyppAqbe8GdV
9kAHdD/dyEvFoaL3tF91hvoa68ZxiphrcpSLiYkOkGivsnoO2ITSs6ACyrQeoKRI
1jMdMoR9YDxLFu0iSjk/C7i4/7pNKaovzkaLJp15cLjK4ebe9KWS13Rk0MM09R1V
oJRqfV7Wyy6A8++DPgskcRt3eJ6Bv3Qfqa4yR5Sm6DCXtW22PNuT1TnPGbIJxOZp
VV9lR1rZaV9dFPoOQ77kSKvhflz8qw9dvUmp0dI/oaIV4gxYufKfPSL2xP+eMm3e
W5Hh5C7Ze9C9pB2bqetqb6/zigGGUmI3hIICBQ06ziY72Ai2TUlKW6kj1rbm25wC
+R6yDF+vi+/ax53Cx0wxtw/0RHXlUs3b0ZaMriLQWsvfB7ZFb303u0HssYV1J+LG
R+JUPr12p4dYRphXukM2Zs7N9CZl2wZ7Mz6kiFG0G2Wn06nPkoBQq9gZJrNhpCx+
KsOnpMZlbyQEArKr+raR5sam+W/ZsZi96b9jngNgRCCQTWkAbZxZpX51o89TBuHB
UZfaNVt9bd7xb1jdwVIKrHCRN7sQ8VEo5Ttf5vPVC24nSwWeTMRNNaVHR2lD2yYR
u++/Mii9ql0ofe4f5CHYk5KXs8a8Js3WC1mKs8486Ju77ksjU3XENdnLAoeRFK/w
2rZkPSAe2pE+M1A/F3UjOaawuILXR3DTQmWhXq9h5dT0SVziBjWI67oSfLAFPd7w
jBvf3KpZ+G9KkEWhlBkqA/3a+1nxkR6YJh9TXXuVsSKWCL7UxYKULrvpY9miRAL3
B0XMAwNSfyRVJrovnTY6po4ke38j0sgbNVPIgDrC+jzgPGsmZkxEV3tUL5krNo2M
S+lpy43YEk8ifk6vn7YCgoH43LZyDpNYumexNjSDIXACncIJzsIbQH0V3hjHzKuw
hzGpOp3UzBdMl6gsB9hPdhnFyNRgX9b4BHETIBJN/AIZYfDGyVKm49BM6KpDmBv8
SoPtIYBCqbsO1ZlAywEnqvzaQw0KrJc8ojsa8FInp/9tWTeUqOfgoV1WvDwMNhEf
ILhVstifUl4cohPUeK97qrRRFHbl/uDKQrzLcAEQkeNS1uDxrrGE/7a9zi3i6QE6
dGDm0bMZKznwSbypzAxhhMmA8iQVD3RQuWw4TgnvPTFpduILjrXSQCUa+WVapRWP
FMdP7WP6a5m9kDrqKei+0Udl8QD15YteoKZgimb3UK4P27jLiqUqgwp/Ko3ZZx1F
rWDbzR4JlhcIRY2+qySdKqo7ltfEq3xqKVa3E7u2S6S07XsiDsWSIP0sGgl/FVlz
ZWkz5Vbo92kaz3IHZi3dm5+775qDDIYW4wunNBE7bKyNx/H4M1lOe3LYb+LLENVi
d15BlnNNSovAXAkqCDxLXFcZ2ryid4q6B5kUvCqFiSdhRVpEUNZA3RRGxgPqnlo+
dITvHe1MPE4WjtM1izojDHtAmGf9LOfiBJq13RrQGXDIGDlD3Bh+LtapTOjM0xqS
SV6oFrBapBigCzaSVoXkyvVuDd1SXexth1x9VSX4hK/W4agyL4b3R25jjDVR34t8
0OSXK6q/YBK46UzXlvy38nftkiSMYDMyBfMl8+xwHmSnbiTfM5eyJmHEz5io8DdQ
BSDBq8Y9IHqZd8yGzIQ9hRI7oIVI/+/haK5rX9wWXMvGQFWQ0rL6GxG05HMcLXlB
ARZZeEPaDcnpJP9U/S1TISyz2z4BiFnUa9pgr7UbUt1iSd9IeMIwfwEf2EAlB2QI
9Fr6Macymnu1HSq7la7LJW13/jBWZWE5EW9CpP1yHgEuyW6AfAXLKzcS6g2ZFyZk
iXbCWBNhv+H0woq34k3LV+rLPGsQQFEmFnitIRVjKXK7qepruQpcpHzqXtgtmiYm
HgcV+N9o0n38GIp4+2k9Mvi14TLIN7O3dAObVrrD9QdblTMBFs++dW/suCTZD6VH
dcZNQtQNjqXsG19Zmd80vkjo9YopI3tCAQZCYpJyoHtaZrUHTgG6Q4s4lKq1yhqZ
7KBtstTVcyvjUA9ZWqYVF3vdqGnHUWWlgJKO1IzWLu9w4u1XRt4y9McqwW3neX2I
eHsU8M0lCPd58/M2ndfomCUDCup88ufvm3uTQFZasx+xg8Umgupe/74xi0LW8Oob
RZIAo30i/wcOUY611wXJY3lkw4A3PA4YwDJhH2pvvLYUMLRSoass2ByswcZiY20y
IVshEPj1v0MKOMjEnPIJrNwAtX0f191/5OW6XNCY1k21cPKeg+F8zIcubr4rG8kw
PmDByl8V7EzAFK2dUmT0z39wj3HB3We/OTNn4B0RkU2TaYgrjm++uwypLBcdAQID
OS7rhiINHTmDFgtUydGVymcAaOry5YlFzZMDvmLQ52kXNVMRacGWTuyLjey9koyZ
d20L41aemaPDn+JDeRiLVqta/9jbgK9qw65k9gsEG3XWwYwDQcUfFe3bFHNiKZEM
TFf1GkZGFOyiccJcMDCj0oxxG3oxkkPFL+nnVOrDaHwaDQA+jKpJapiBr9t0Omcr
o5Ki2s6+359tNUu47HlPX/4zqs7eJ5v0TfrauWiC4T0CIbNMSk617/F6ird52hHx
bm81vFq84b/EGuneOsdPyYAk48zXAOtHXs9vv7UCctVtUMA/roC1ZfA2lixxIPpd
YHXIi6bRsFXlKSIUr4ugJSxgUCjGZ+JRm354J8RGs6bCOCZDFuovT7yTEwO+8nTG
aC2QW0NrgYWxpwqA8uisNcpm70wyLnwM255gAQrADdvYi3igQig7qEqXOmqb4Qbg
nyRlvowXMPcjotrunR8xSZ4PZ5U4vd0aAoXpEOqy9Z/IrViHjxzocuTntLgRW8S+
jT5AbtJyXQykzctYVsXisGarkVKBasrLeYsSNBgUX7R5bYkSr9lj2LiepG8UMAoh
aaXSDor9rm7rIK4xqx4zlSD5veRIog4fjZmuxrM28NoIDUgxbwQlEsQc5QNyhznb
o/uEtCXNCCdOgpiTPeMHAnTVp32CmWgR1kca12SB9ksl2d8fZUap4tK4qzOg8JdM
8ve7RBnxz848+bStv9yG+c8Uy21sRDT11Nw5lZtNNbsrVCtlqvNQdZTF4e+rwHIz
jot70vYzHQkGbk7xKMS93O4dlX5PnmV4zVlL5xlfcnjDf/kcDK2Sh3CFFKXYpPsq
xtKoLNrEPHeSlwQAhi6GR4x4SSFuBkt52Tbj7LuIEMkiDi2szQG2+geRcFdjszJG
pP+mVtjgaaQtEWpCvM00yLciby3r8hv4/S2tL7i69E3evIs8KN486QEcOT1nupKw
jY2WanwrX6+t7FblBSH7kxgqMtmCdiYxAYi4ZA5hZroBjs7inY3EIQOGZif8h/4b
A6BDUSVvNumxtAArAZYcQ2/VFSD7tuTNLmpFraUqIUAQEcPZ/z87KqT/s7QsfSny
Z/MAMBgD+blVbfEUAots4aEa/1UnNx/QSqInhbMzodz92w/Fv/CqJq96LTXj2Nku
yGF7x7eHkxoZLgpypeFi85eDF1VUIgFo93ldnk/2Eqd5evIHuMwq+k53RRSHz+y/
5FZZFjlyT8rs7EJmTAi8oMnpcssRmxDckqMGDTPs6VU41nIBjiCs2TJaxEQdYrMU
tDaiebCIPsSnNyx2lhe2pRRdAQVaKXa/6CGotPseQac4eCQEuoNm86iXAaeLNWRa
fuqyVvisyqvXSg3w+VUx/gotBc4Ivu5dlbJg4ntJN4+LaabvWuF7LjzHsFblsjU9
NzXvhRcFK5T3IDAEeWzdOnW8aTX17kRTl0y/VP+2b+nxIDMbm7BjQcSXvwejdT5G
Y0+lHy8e6us173JwOG1mebjl/66rt4o/rUBfz6zzAxg6J55taN/x5LFmdEQ2gEy+
5FE/YOtLNTvfZPtfPt8m44kQk7uHujqV57tBJuza+Od6Lb0+BDmOtk1Pf8HfN/ut
Pc2/U50iCDP7ZL1F2SJ/GxwyIDioAo/ZckCJM3cqO/TLugFHLmM+DZrMSapYLZ3E
luOCU0qt3VNzFbTnMTMec+G/GpNCnGrqIJZbld36NgLogWs+gOEScr6bwTGzKLGA
JxbrdQDf5r9EUfh7Y0XNv2x3ZiJN36kU2i8vROf7akbtkK1weERce7iyih/M69Kt
Syr/oVGiLb1brNcVaQwZmpgIR/dnpS9i9f+uGHdrzdxvviTOiku8nEdiuMJxeSCw
XZnfvCPCM1z06ThakUDzDFg32Y4z8r6ADPOt1EBjNR8IXMPXxPewOj+bHwONIAXJ
FtfLfXDZmoMdebU4rgZMw0vboDEE8A4XbRlOGcpLjM1yOKteIWBcHrdoJ3PvoUwJ
XhpFyZTTSq4pEH82mmXiRo+mQHaDdKQz7wANv2oBgAwuIw59OLCyotpfseUtMTyQ
ZBlZyhVHQqMKWUZrtjqSzuZHIUCO5Skr4nhvx4OcUjR3UvsLW8A1fznlLmHdFhJO
5FJu7h/DWUDyX0WCqoqKU4TG94il/xbUrFPeqzGNSXXVtVmHBSsu0jO/NcFNngQH
klyvlmRgnzAa1EMlyQz+MAyxK8TzIourVGcouBOtqNxFUqUzwxR50dsp3BUFQORC
vW4gcpZk9i36MLooF1bAU2qNES+nUPixkgW2diOBAup/YqRXY4sIxxgNx3APNMI8
zW0yya66AN7Ia1I1Rk/zBvkhpq1nSYOIhdGzPQkgVhinP+RkelVNRm9N+ezpE/UE
OL47IH8O4KwMepdYVLovs8ISvWrO56vl6tPMFbAIMZGHdHQPKaL+l7NzB8vm5TzC
FwN+vCaNynN5yiP0dBCnIqn1KW6j7IBhNHFPpvZiCE905df3VsqGGPlgcXYBTxX1
DjfjSUlCXfwrqeLazo8dY4+puLjVO0cMzx7Myak23OrDqD/2bU9M0AWH2yDJIrtS
GrHIrCE3DI6A7faAhCLUv5OuC78PZtjT7AoWCsM9oTMflF+4R+5gr9U8YU7FryKI
DVCPQU5F6zJFr40ujEPQMPbx+AovAKPwG7lKYlXgueIokmiOPYgK/6Ryi+HA/Pem
Q4HCiEAXl6hYn4yehp+kKBG5lSXHT/d0d6ja0Fm3J+kNwin5XBTZcA5bR0eNTtCQ
MYKpKA2Mp980+KO/74epIsS2QbQk3yo9HnCFJxv1VTzbsyTImHiAsjoWTBCUyE/A
1YMju7qJEFNkxwQqMZxPa9iHL+iDoU0+kHmnrIHz5ObBVTjt0BrWCbwS5A7v1kU6
z2kHoiUTXnhe63qRIMyknTEBHznN62bJxDoOwtv7ye6SH5jFOaBdQhv/y+amq4fz
LZ/5MEkTB3RqdQFECdyWrzFYcrQo91XL7I1/TZ6CzUgYiDlF8SqXnT8SvkdM9+ur
Wc1g3N96niUijjIgOzJn0/HjH8Cvd39vMszuXbS2VOQ+Q6+MFvc9YjkIz+6jwFi0
ZLR3WvTZxA51jS1gIfUOqR9bzdStu/aqzIf2+P6jJEUVcRkMUVwQmmXkPiPEbwNE
xDdIWF8xk/6s6l65xQ0RoUeBcedKsMi3HMk4jOu9Vv6kg3HkVsKLIWDXoe6UoaIq
7cDxGTtwIv/pwVbBa2Yl02PPoOImfquoPceyFbEHf0tPmT7tHn6UGS82GniZXOok
Jzdi2iXrXettCeireZgyS683EZfOGLZlcBun4zC9KqqUbrkXijSkS7yqgf3ufgdf
FLMw+s/+YYbIQrnbBXsNqeBCDVMcnCzP/yYuI8ocxPOQ7Q4wXEawp2BO0Cy8WwJZ
JuciM49lWwtvesVC1KfWvFhmM9U/cFpuBGM3uDX4eCErqPWBsN/oT0JL85iaK+hA
FyoLY8sWP6t6uRCe830YPiI+4mH5kHJAYFiQJrRJ0MjHRchfrqbps3RX1tj/JoIz
k+e/MtbqdJz1+DtUOz/yVd5Zlc8GdHJVEezHq+u/wgrih+sqWiRYNWt27TIrRZjt
Jani4s7GFZdya2ihfOSvysZekuHSib7VW974rmlsa9b3MKAK9LYEp2lzcuk31bnr
jN+ZXHj4WuftFVgEWeXpMklaES9aJMs9AMlBxRgXcTxYnSwqBXiUhrY0DscRBYym
M4FKggliwWBwRZUMq7J/TjeWwBr+SVTU5mCfEbcAG9iTqhuc34uNLD8u2k6jG9Ba
n+GhzYh5DyvN/hz/NcBEQK1eLbSd6SgL+/kxe+WDbYbGMAp9/S4qMkNJwVxr0b0U
CL0TZ9s/j6qTgS7s3kAHoHuW5ThImBGkIVwq0iMBKQlyr39uvMq617fIfXAdM1cZ
8CqTPwtQdEsQDI4NwK6hrAkk3vH3jtui0AvSfFT2J5CKdAc1YqP0lEFFGxn8HyUN
InOz5NWCu8XcVCWFxYvcKjHumror/d1RAQ77sEDkugrl/eZLiljsHpmXSqv881J2
xKqNe4LTiL63V0iYzLUNrDac/OxlcOs9oZfsQ0jS3XVF7KBSur0bxLDQgMdXi4Jq
75TX4qTix9RGMuMT9KoCzwQzn2ZdG00njlxXso08Y+jhijXDiiYadInpadNN95lU
EBVVZiNF5wW0VzDy0j7ywgXFjF+P2KIyLzimnFcv4kVtAGSX1lKKd11tmXsPnknR
Mb0baPrdMgj6kGu+FzNjx+/RFv00UrxV18nxJOWjYK0FoGkiLITiwuCcDQvPfJuo
gY9u3kcIxKmAH9Lwsi9XZIQLBq+WCpY9sLra9PpS6x6VYF8eOViSpCV1OnFI6q9J
+kIOQf6196ZndHcd+MkAno8Sws6FaEsAyEY8H5t2ULwKABI2VfVU8zBKiEGgqT7P
fFIGEqS9dxMgnY8A6aHVKzvrjwR/rVJx5KTPjqZmwh+HfY/seT3FUan7nq69e2+n
B6nToD8XblKu8dSxGSs7xxZP0t91C2zkA+VRAAA3Ubhae1JiPKA/66xzVTD8DyVY
CVOBiINHBf3NkIWJkNiKz++jZ/Xk4GvnSthHFBBumpR1CYbMpyv/ukEaS/r1Rt98
/9tzq2nvdwEzSTgLKHy4kBVfZ6ViXCsMt7l8SYUH0MOAUQK5ZZ2DiRr9pNwUMg+F
47ddeJli7c5LEtEuiLGJfNn6XP38QQstjUhThEHc2IPk6rfrzf+6/ivuEb9huN9G
x1SUOfEmQYWh0PzMqzdW3kIiXv73Ys3AoWrAiiyqr1Kwquc6C2hZw7PxqhMFlrpe
vI4xksatNVcn/ptQBcRTApwMbikbpn0hppCw+ZLENS0sJkQTNNkHY10D6uuf/JkE
VnfofPD19BmSt6MUBYeIL6McPgVSKrjbEQnO/VP6a5s5p1y7XFWxFq6YVPtuCc5a
17jeOF7FSuV1ad2l71tISnl+BkYc6DrHSE7udvni0AVgXIOsBMBwBMxlz0vCpelz
FgVVUF7pnb1cCjS36dgVb6BMIep7GlM/kjw3U19TEZ9ILg85n2ewCIZ2Tza0GmD9
7LcrylM55fLo4gW0Hyg1/o0+3t/KFtdfWlnDihOut37uVAXHSthSEzfGAOyks3+x
sGaDiqLk6k7H1WXWJ4m/93sjx6nyUR2OhXO2JbddN+8CBCrrt/gJFtODLf39LKsE
B1OW0Vrm9W8+l2NFFOXsUUKFAiRGQxy7+C1NlUMFT17mvHkYIrQ3KvV70hvktbnF
RYHzOn7Zh6qn2PViErP7p7YG5pRGa41bqPMg85M10dZsr4jGofwNqGtRtOqlzGIq
Gfc2wNuz7TLedk2ANMgIaBhsSxSKHflfwfuRT6kuX3eyy7T6Y+2i5Iq93M9RqpJj
vaVZvLQAPoSzoY4qP+mSVjiYbJ8v1qxXj2ELEfiMbMM8MD7EGGR5HDt6gbtw5ryg
9vu1rmJzH2ko8nErAIdf2xidG38PpXZv3ie+SobROTJ2ejklL/O8qOoiVFcJOmQG
zh0aaBdZPvqGzOrPHl/br2DCV1dDQX+s2s1Sfp/h8KJMiC6PGeK68uh1lbPl5U9j
s6yJBMDMG1/Rsxf7HylplQFxtj0HpJLsiF0PENxm+6cH5Dqzf5n50XOrBIKPU7Ej
CImVCmDValh/1QiZLw2w9pRJR/gNwYd9XGKqVZpFjMr8+VUPYSigxkSoGHOtVsoA
0PXA50osx2Ll/pdho8dcdU5tD8FcGLPD1GdmMXQb0eDDEzRE9dSWPwma7cZaWwQG
/0JOBAEVjTL0Uu/7TeYQFE3r5cHnjAmw+wnkqpdFIKqCN+v5tNJbnMfZfIjbs/5y
+1md5PvnGHWvRgXw66qbBGfUaU+gypOGbDAuV4lYuo+B321OIy6LsREbJIbjfae+
GScsShg6vgfbu1otwT1kF4luY50Gk0xiigpIJYXsMpPaha9jxmS+2tv/VQpSUTe6
iWYsXckFz5VCk5R6jLxF1HUfkys6vOULYXNmwjE2CGV32QhkxGHlrgankkC5Nogm
xoU7yDrP+zYJSu30qa1SXsApkaOakMEXnJiYo9TPZEIi++TuLHUBEs2GN0SYBbb7
2SgGBhUauDQpReIR2hGRB/U6UwAmKWWLyTXTf6q574qLX4TUioU/vL5d19kwm4Yl
f9KV4hp5ddfJrLP53IPQduy9Vy+RPVzJCJNYMmKnIUD5IuqgxSq0wg0DKtNVsMFv
onOwtbwjyfXNF9PORCh010YF5WP19e8FJ3BzMZm3swg/x2iOxiZagUz5eARL7IKH
WO1QiKQG5G/8eQ5dDcGmYeHL8TZc+FCoA1gbynkjFt4CU/lgGOB58/sDj/orwfKI
lqZ5jbAld67u+DpA0edaaYpXHfg+wBjUqWRlwx07SgDCNV8TuzT/T/7FR0R8V2Da
y93GRrjLgZENG7TS9ZXZr3aAXql9ond7aCtq9NCcTkhE2QX8Anmg12qOY7KNOCiS
808vAHsjuvBnymJ91MZRJ3Wd/r1+EO3TiRE/DUWkh0/vLYiSwPTkruU9b+JUkWm8
YqeZiYNG5ZFadE07NqbPIDbJirSx8uqurMUEKCESRL0u3siyUtWii4kM3pPNAYCV
K9k0bdBFZ8r6c02Rnfs8ng6rbE4E7q2HJpkI/e9sDBagxSyiOH4iU+YKWlPziyMH
TFAIhqURRJpwA+rA+VeKK70L23R4AQ39B7ymY6l6S5vfO+h3w0X9rXbLkwp4J69u
Evi1CaS+nRdLcGAebyikQPA0ii73HNWE4U/9WTwyiOgWGGWTvNAhCQGxbnwBqY6t
LsShnFnIpmsreyU5JwBlXOBp1i9zxNpVsPxYQNIYBoHW+Tj7HjQwWLv9JsKx6C27
8zqLS6Visv1ZhQAorKS0LQYLYn+/7qyPAfjkQ0q44D2B8gbGwFBSZuM9sf+o4Wc7
JJs6KH4JQC4XluvVyT4GWM5M/ZpSVd1/6fr3AACtTPFVs9knErRtT6Gci0Zq4/0b
brLC4TKhAjFs0oy2LlooaAF3HPHQWoZH/q67YnVrwgOzhj/iPaFtgpogEmAzfZ+Q
bAGM68L3/gSqWuFxzYSOSXV9JjYheMzjdJFLgptIcQmODtrnU1HF8auZ34+6oX47
olH1cDEuv856Qf5pYH29NhtffUKx/XJzeKOV7KKkknHHvF+5xAbSLJoSX7qcZ0UP
v1N/YS/DRi0BmfY5Luq2uQ/cBOCcBxQ8QI+DMMW1xwfWiVmhIgWdzHSsXywGol+M
dBBSbw00hs7QbZ2lVIX0SrwANG2GP5sLYrw4hE1jqWiRTxSwmkNrIjcx3bjCPElg
t/ESYFSwi8kdz7fJkdjm/DVmMtzm68E4DU+6NGHy0rsFKMUTA7BrFe/OhEvJ/EDp
h6GzkZR7wBfIy3ZWLZN1P17423K4FVVWzc4xJ3Xw+pFkQGM+vzFH0cUYwY0BorKm
TUGE2h93ygFEcGIc01ssVPwld3WYfKJfj4bKRvAFzPZ4HrsC5OkuFovzfG/ZHFNk
hf8CAFAYwgFuT9VKGEw+pTcqzjcWZriz14SiEqE99ToXTwTo64ficxZKkhfilevk
eduwgNO+/cZN0zW0VywbWapoItwjo0RckbFIyntjUg/736wJO1Z0+qTKk13Nwjna
935VZW8qVCognqzdQQdQKFUrLI/56+j0wX5NSJVCzEM8WiKdxCVhMGG584IRqPI3
E3CSncnXgmfD5tVZPBf5ijHHQFoN8/Q1s2Q/a59nHTTJ08larEjHmGWA7766+uCU
dqpBc1ZRU3ZLFskOzRi0Jecy521Eqz+B+epN0TPnOD2CbB5Zkk4pZFkaToNDvWD1
JQ36Ej71Y9tARi4jYjQiy40nG1B8sWYeuzHE94csYQiXVOQ7UvydofFGe97OoAcv
END4nGu9I2b0649Eyaa2c0ItP3RnTrR5eWxBdyOlB+HLAqfitveBRR3cjoIjIhwJ
nZTUhp1MN4nt7OBEeO/pHk7ulpWpxmZ+AsMelq4GyIkjSAPTFjCZ7qYvn9H48+TB
cJgkgVONIluNyevU96nDSWOihuo48cahUTNUBwcvf1fZRNQeAJJkbf85a5Cuxe5P
OXHlC8tcgpNs4hwvPtX9O30ivUnUFmEUxK5nnC9ClECf+S6NnHL7gUuPezNQmRm8
8xLGLLUTlZQ1pDgVZxA6NDv+sAWVxnOM/+Jc1ZiJ6kIJMfdgcXDryiF5+VXWT3qS
7ytlQshaA9oLtQorCAoTPBmxSCYRbtBsttXcDitYfUMkO6sxqZYWCq0hz4ZfBunz
a7FBtQH49KSqaXMjfCqMR4eOdAw5Xp537Q7S+Q25ylLK0owYrXvnnT1cQ2pFZHhl
Nt0vFtIpuosE82sfnULd/wFSVbrQvmtYhMhIEKf4COIdPB6PsGfvTJ3xD7WZhkSb
8LvqW7eOuqv/xQpbA3/cFQeoLNW9+KTwkoyNNOBgH4lyWqcnGn5nYA0U8gqeX320
C6AIHPWPwzKKHCA0AJ6tWj87m/8pSo0gflmgoLQ6rP5zKUW1gh/l9qamGWe7/ZW2
wSl54VlFGEjgehZZ4ld9C/yE8OJRya8jPn2SmKXDE0CVMvuq55II/eefTFgs4mNI
DctHMkawXNgPD2pa54PnGqR7KOKOmKbyA5wrusVJydNFzJDZ2MCsaU8f5ij9yA+7
rCIMEvp7E+G8byzrE4dNKLekrX+7uF3lfu1/t1NzzQiBzAXKEMN22CtBrt2z/eOc
qxwQ8+8N88/mLfmHR2Vkr0HqNj98mws2r/hnZHAPurTwcmJCvaF67u996KT0yjO5
NA3lj4SmhVzCyykaxH8yBt816rvGNYIRGrAA/T+ZHH5Vwe/00FGSTAm7qmhNrwoq
+QRbJP6mnyr7YpsCDt96thbT4HMjbFfbZ9RxeDsyakLd8bsZQ0VyOOeY+rs1I/sM
8RU770FQ+Xry3SlAnL+KBUUq9Aedd1ce6JRW02+EsHAfQGiPv960TS498Jsks6eh
ivnxA/erx4/9wySJ/MIs3MBvLKchiYm6DtF48clXxd84YgiUAsntAFcmniI3nNTG
MFNkYaWW8WrbtdrFIusT9Eh5dYgUFeWN+DcIMy0dY7T42fnqOz7rRJu5IjVOJoee
ix2S21qK7rMVUlJeZ+gKEBaKuXLE+c03Kd0CPAUB5KgX8P1pp/1pUp3PI8whntuV
AnOoDVIv1gvjQuQSL80dlv1ALHry4dJb1+vvwGr+gMA+lK9J2u2uAcxZjK3Kp+18
6EAMSFrPFke7+y9S1Dm+Ob8t+8+lgSDwyZ/fvWK0Eqq1u4b4CES61yDVTtR4PQia
ehu/fW738UQrd0EfuXLfcAgPxJ0auvyK4o7C1hYjNrgi3ZAgbDMx3GfhulrMIG29
L+5O99s7AnVCYnR+rez5+j8p1944ht3MvhfcpMXHDtQl1P+amKVq6RzOzrzKjbgw
4wK6F3TNK6rBs8WZAFewGAdTjMjKqdyOcpFvWOloiSUdS3RFRSuYSQz6rBR2aTe1
EMa8n0U3FGnSCPXI1j+CjUTqC651tjgJPkr9PfBK2T+Z2r9vMl3eZcu8/pixoUUI
KEuxBKBghL/O2s6tOWQeboRoYMR2z6pk49pDzdCeHD6T+k7tyOwZpeRwUACWE4gA
GKV1/b37MwZbFFx69mbHB4iWTHcEQQ2Jk6eU9YCiDZe/yOtY1X+BfSr2tKPqHVfC
ioYo0jQVYBvk0I2VD83cn+DvF7CpkxBkZmSMYFBQC/2D8kRfYVW9vkwioviIVdBB
u+2+vBsrBdrmT8kEGZU6TbVAHFw+4LIi5b2wCjnF1D8oLDJBBhA2ANOEuTdZ8FNc
NDQFa5YzNGFpjAhOWhi977cpJZbokG5ooZZvUQ7v2rqQszDdpTVOpbKKxAT5bv8g
MAvNIHDLqTyIosXDb8GS4FHzzkiLVoI67uGNRnx9aqiwpMXlRoIN1jEY1zdTKHX4
PMIaGM72R0ymsDsL0zNOiGtxlwnVn16ua9OfDYEHbkIKeV3GOEU2wLKmolHwvqe2
6OWDaLmUwo3I3LpeaF0fVVgjJisP1ak0QZyiU0pkB76JXOIRLWkXPep+Bhw2dZvd
r/tTFrj9/KDjIGj/TBrF1zqY8KmvF0gSX38bofpznvKE7CiAb7OgfE5jHFNehTGf
E/LHKyfGN9J+Q64DZ7/9e+RN1UpC+8hPxi4M6Nhq/hPS4uxmIiId+0ToI7tjD6Tu
AVXo0YhbjDgJIXdpsSStWEeM9Sin1XOY2XS/IXMehgmnfQVHw2fVRZBnkXZb1IUw
6oZZMebTFvC8TIrN0UZAeQrtFKt9jp49/dRv7ej7SqJLtS8j6KXkm1mP3bvqd69J
1qacG8DzIO++h1c0ya+3R3sbQdT3tzRejzivApyDE8jQ6vR6Rl6MnqhDDBxPvdEz
mWiPAiDHU446aGf7jG+WyTjy0NRssAyseqLiG6UKKWy0pO8WKMWDOM7UHLmS+dF5
2hb0QFBe/gx28j7HkBF7ali7/XmBniif7Yegr4aldzY+6MV+6FTJP2PmuVEcU3zx
mtivn32WsUsBuAlCKFiXeqVGg7HctK4fNic4ON13RaHPSQtOFKTA8ybtX11M5BoL
WLgbTKyRbe2XtjaySekQ8+8QOXAsbMj6mGe+boW7hkU8pfSxZ/JHzj4N9iIZAhGn
3r05WjfQvgkiIxw2vz7gDW6C4vaUY8VrNe0IkP+mHeRU3HNvO7s7fkoyq/MZYy6F
T7s00mFdGYox4+oXTF/h31xHQAP0fY7sW0YGZ+mH2h9ENGajlvSsBoespb/5q+R/
bE3DYFL0nKpehufbBIBg36BbCdbEclVdKyxpmNnMQQObOP3Tbcm075MZbTT2recm
3UJV1RLO4oTdYMqu5WTFrm5UXJ+r9iWwStgXd03AZA4AMpB7k5Hbc4K6YzZRUa9W
u5BP9NL+KywuFFrJh0COgyVJpt7ACus62o1tc6QF1T+d+YNuvWqMu9mq/0qwad9g
z2aWvjxGUwbuy0yCDpqGH/oISoXPO/HvGwtZFB3vrivWka1fXq6ioRsr5irh3qLf
eII9TJZINoJJVnvU5F8OtnAbUQ1rQyDv1lnRzeMouES+JqtbgmDvSplSRz9aTT2P
ncQzFT3wS6uJ6DnYNpSpOMFVCvavahvDyXtD9rNpfpu/xot1QYaqpZbcbNBa9bjX
k3PhP35ys4MS/J4+iaosLTOsjrm5y1gxlYuHYkAYatLPHjPo2tEA784o30o5dQUF
oRbP5pVw8ze2TMZloAKA0gSr81Ts6j7eOryufTYCV6WXvCDJym3LFjPR6y0U/tTU
FSsf896rSZJ58qchW1JvoHQxCGF6K9Zh552BHSMw+qQoXqEQ5lesN0B/ZF4Ajzv3
aI6manSt9VdYfnA/ytb9R/d0bN+a0YN2sr+SapcsOAAochRfLwIzWsbD+/Yyy3fm
XuFwJ+109EmycWTpqT3UZGLhp6bgNBOirLa9wJrBu5PxCm085mDXip0LS7WKUMb/
xMgq2jSS1W7hcz6/bIDsGJE6g2Z12hhuLLfo3l+/n+YeYhfwXt20jpvQgHEH3cQz
o41W8UBjaBT+ZtRtUw7R6iURZxo55ll8AQgI+879N9F4HQpgLKY1LSfGax1jrIvD
oSF+eaQbZNV6OxeCCM3yQda7ArixckkQtQtNOXoyqphbUwh6lQkP3xT6VsCw38C2
8Y+xgei402DTC9BUQbRBU19/sMhkKgLOkjaTKHt5lb5lMm7c/JOeEisQ2yLOKLgx
TVi7ul9VLbH6dbOIMQAaCTTxhM8GLbtKpProFvoBZcZBwUIgSoz55CUelCVd3ybX
szF1B40uHXWL/m94gmqX2kHWiJ0lKQa3s6JL6UuVgprBecve+16w7AGq5RtrMIzD
cSEfX/X2N0Cp4yKEY5TaI2Bs0iKedO/Grc9GuAo0FIwYIIJ8OJULYpRAeeh9fD0g
Q40/FFcdCS9N7EPR9I0Dz1NCFMifbWFGeZ14FK7hP2kEvqjbxgXvjwd3IpblQdiR
T9FuVfz4vJUY4/WmJJpKc4oikJ7Di5CUGOrrC+1VTzBKoqON+ncwCJFKgdX8USHu
FKCptDaXhBTkh7m+wk4HDMnL/g4F3MV9L6va25JotKFK0D78P5orUyYmvyMoJ+kT
IC8bw7erszCbTSuPp0pa5C4dxF9pS9fIJSz5hvFPC20OMc91QpSLF1PSzPbboky2
Ntdh314k7Sd6ZrVvmm0K+z7BvBBg4CTJBuQ6Siwuk9ajMRkV0vd2ZobiTSxO8E03
g/oYNw03NiOVXJbpLq+krR2BIfLL4TEtDXCxeBoVTAwZGe6an0GxctzKFaqw8ROj
AKIXchkQqmUCrVUOPrCTtcRhi4DdVrFrdDCyg63nSnjYHbDW0yD1r6GsjM6UshmK
8w76Fy5WxJsBY54Lyp4vTA0p1+KozTehQvMSfQpJTRh+4TbzjmGuW5uv2E3Q0XbM
SSkrUwWYUz3rhHnbEKahldINa34XYxNsA6rM6KhBW1RQbZ7e8dpDOBgGmZEcJN2U
+LoBkkDRAWm7MAtF94kIVx2BXZ1/tcsrRdAlI3Gd0SSD1INT7RqpFxok9DB5yxlL
KfqxbANICpZDCmQGUlAWGJkgcALex9zzahPKW1+/k2mGBDBcImJ/5Itc0/kwORea
Bv1sPHI9UkT5D87nc0fzt17maxHIlwdUBzD6T8aSHg15WNVMDLXo8hYGwHFEFfIC
nwSHJ8DM21W9raDCSk9POGePVi7sXe4Ojz4Hu7who70QdmCDeT+84JR/UZLHHJbs
4pHSAd+/wmgNn0RFs+R3dVCtQP5vAcLQonhV7PEPm2TJsPvVjT7hdNSWmCrFpmbJ
gUMYNWlaiYnTpQcfYRdQKQoRwJitC9M6oR73xtO46HyWBNiI0nYal1/E2qPPhMh+
8byS19YdjVLGKf5WA6jdlUFwYF1M39EDjEIm8kFlgCMWQXL6nc76ycwFCkvCAw0I
iqQqI6UN6KB8IEjhiDPILtsQorJbSA0hrB8xOGmSsig2+ku7iVrWP+vQJfyOtsUd
YIwdM4T9HeppxGEegpSwLpHBPWrhozlmx41WtTQpzJ/YXQBNsYN5pQRXcEz5MFj3
QEz+JHjaA+YsRYK4sCaQmUO39krLZD/Z1s4aXH9IxTRXG2JDuHNzid6ngupDQ012
SwOCo/Lf6I+/jl6rdx7JzTATQmnKQiEk4/hVDAbGAA3E7ere9sKetZQ8BciYpR/1
qr7eMjadkbGqHJrIbTPqYBKbuLsIdEed635LgFZL5MZ1DXFX9BsrqarRuXTs50RQ
eg+txFl5D9bHuX7PHqpd7Jwjz9HDuuhxf1wwPJOYAbrDVGtEEpnJsElZBhXSs2f6
jdBGoLNxBzcdAZ9Cv3JKIWV4dajsRoQ+9iW+jqwau2BxjdA2AuI7J19hlL/ijoGU
B2Nt09uOpbBcIl3vWKUV44SAya14HpnwMYPen8TqghwfVaU+G1HPTF3x72EQSfei
+d7M3ef2ovRkCWJWEz6Bz+qcSBMuGNr1MTXANLSUsIUBlXc2zH81ZnR3EoK0n/c0
i5/KH7nNLojvvblDPHodhzESm8yXw3hyT9Jx6aMtjkWb+FlVI5dPmSAsJaMBVPdF
9nTzWbfHt+gELYdpjW9MICSlPodkhputpsYm9iM4ZDd/+qcelDeOJoMolsglPHSe
M1Na2AtBOAJrth+nud2n/dUxIKA/ZacBELpNB+K2WjGnP0mJl221ljWc2L8XeWl0
3XDaX3Pbgle293pgZ7plURIiFmLiMtTrAnLXmOLryzwHFZcfBr0RNBgDg8DshFLk
UYZjRy5AHAeIRosowCBNSEqBFuhjOjcKNJHB5KpE2ExDyvqmKk9irPoTtHMv54Dq
dkYyvHs0nj/s9ciSKemuJ6Tdq2FjSsxt814ap9ru+sO85HVl+6y1UUkj043vd9Tc
OEdx23Li0vnI2p0CJ8t+0Y58PHFtNZYGHk5Yz+wOcRpnx9dL9vSDbGX9kLzu7m1P
y8Iaz4VN3+4NkV5ct7Bam93lMXztJFcJS7utmyVWCi/b/QpUfO+bdAwa4EQdQDtW
yHF1ekFHNnzshzZjQhDmumv5HB5bbmotgb1jeM8XEncIMFDNaUg7d1UBKsd6HEmp
Rqhq6vVb/UBKcqgHPZW+mIZQuP/746r6eO6WZnyfp2DfQ8oNOc3d15GV3v19tg3z
Zm6BO8DUyVV7ApCDfY1NMUXwNssxoAX2Z6ypOubObqK+YpcZPmh+in4cgSJmyCFN
l+tx2rJ2LvB9MkjSLdrLeYK1FGOkjf19VhmRZ4gI/SGtCcAbd5B47zXZlBz6Qml4
16QsQkhmOhnzWcezLjcDa25pQTguoFqCkU/MU3DR3HWiLpogQhXQxfqlRODFYesg
kRmfnY/zG5EpE/chjVB0LhirQWi5MBbBsQYaoA2v2HgcQewgdDerUf/aYroC0lyJ
g1dlh9FcXQE4zrnDSwT4+QOVpzMGu9sL4RA93j9TdWexSSxfgXXVWvnrkF0Wj3g7
t1q1v6jzpOlDb9v+Dxc6WTISq9BriO+tsErAMYM6/uvPXG9KvLjTqcxd6JIubm1S
sknWTGmu3KjUO3Kg9rA1kg==
`pragma protect end_protected
