// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
C77v31TTASfIZAPhlvma2tkw7He34Gd+MFhr0emp35ljP09bowGLynz723rb9N6i
bk/YC+dovT30kKWNhevbW7eVJ5cCTSPpQrWCiK3KhfV6pofB6ytgabLueBejjK/s
dxQMIvTzUu/lsj9VIICqfOa42cQKXV2OP6G98i5k0BU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 61504)
39qXYhew4pS4ckO5ZSi6z1hrmrRpKb0vUX+1qDGRmMt+ZpOo1KKW381piuJZq81E
s9ozuRlVgvfSS353NjSazQXDLmU3pu/uFkNSUl8KHk0vArPymGO9WueHhNtebzgT
OI9XSO+hgY2Be2324ASJTWkjfw60FKG5nJTMR07C4OFNtkQ75FwY5o5M4WxBgoyW
qIfykkkg2CJ+8wpxXte/3Gw6uS9zEWhjrM6W2TmdQ/V5XtDpPZjw6X2jIB/pmBy4
zWDrj44RhciXbPeAkQWSaKAYtiG6Jv/KADzUmdgAITQqK48TiTHZhDDS/H98lXg6
HLZlT/oUpC5UdIhb2kR2mxM8RNOawrk9KuBgo61iSo1rbIx9i4roPIRYybjpNpf2
2E4Zkz5m8stVHZQKsDiFaoqNRfrWIceFUc0TGm5ACbJ3NNFzMs5YxeA5F3uF7gqq
SsvXojFR/upForMtcCybhkMgUzaP++X/a3pUw5XBIQykvQKjD6nrNdrXUbVlp+Yu
oxxQDnZ+bRkdqCyQtsAi+lVVfnsgU7Y71s3vS17ECvHVo1QY2s5IkxqUR12R7NWQ
+GzJHQENlbY4usn+4IDdK9yyGTCeMDS2Xr2+iEDSCdjsTeYAdRrVoHsBW307Uqno
A8QiCiiU51F96q23hyaPiiYRVw7QMWnBKBM6g+AcwMiHb8DIKEv7uqdYFPmveExD
R45jTLp6gjd9rsElqVXDbW/bfcS9vGcTcbUBSL61XZ++tvcsoqSl+CL2nunKC8OM
vXdKXRRC6qN6x4LoRtFc736aAbkxAfTFOj4k7ZdlnMdgNXFgHc1pDsTornw5CEY3
8ZdqqzLifwcCfJMJjjmKDJa1Vhg8uSRF4ShM2J4PFPIWBfa7QntzcV3WTJ72nj52
blavdYBzKeq5y/Dti8WFUOjI3urtSO47GaR7JaGjd9v1LkxzGCOi4Y50bOiZWsj4
sLrSTUd+/STkOL9X1uFyQD9WuyQ8ZgEq143M1iFiUU/NqrK8nF0Rvy8ltHDU8YsO
jFadYjAjyALkLa6hmvuI5gBpDU+rCnNotEtkZ+i03ZoseA88e2M+oEWOr4tuwlo0
CIYtCiXTQx0qr+q51Zv48okMAEHkcTJo3e3HOm5JbU1KbHboodTgKddf9dBWznvh
ON7NRoITyc6Epvaw1gv55S8Th3AyJrDP9JXdudnwtSqbFnPpgGd+Dn4b4kHLu1WO
tZA+5jnv7LiZ1+CBwfG6PWRRr2NKKlRwhYqQ2q8RgSPN0usivVKDfSlyBbxHajrj
4sM5KTH+EtFlIS/q8SjjRpF3keI5U1q6pZ7bLV3lMZ++uu29Dmm8NTLJlJJ4xcWT
mx47eBC6TRJagZTpU2qkC2h5sAjWilvMGaJgUE1MsLGeGkziZ/jCubieQProvr5w
K0+XZG/J0w6gMvmSrSeNDClihmCvYWpBcPGWUdrJhupZWLoA9Z5qKXiSFvHBUisy
1pZhQDTiT9xFRwTrSuG+8xY4rOkMR36Z95EZU0PUvHzzLlhNEE63isZU8XkgYA8k
7fEtdPokLIFyBqy3JcwKP/OOesapg2wPclNevXQvAWi5uoxNoC2f0FV0RF+IFnFm
I3zgfedULabhsrZBKFlc2qNZDHFmiJm8SLO/Aa0hdub/ouZ1qOVkOdGZ6iOHGO7i
+QKAyFjArn+952j/1vPETriVu/U8URXsQUnn8zk1+61489tRRSPYErWKPXxmsQ++
AYIMgp5vfQCf/vOhyDgCGProX7ZRDgWJl1lIGiCOqkfPWmDCOK4ORtgZRCNY3xNf
OTgtoEt641mX0QPEjBgTe8h8IFa/ALz9C5ns0KRAKk+6DG0xZut67pKCW55+PWXO
ZJTUVfpKLrtD2ZMe+p2N+UnxUPYVmMd54+Qb47JIci0aCM0RUVg/XPfVUYTNjHlS
4WP0CoBHtXA1ZJ6rM470/uLYDdMc0J1rY+2WfJYRruPmFMcX9DaREooAx7qj7HKr
6RT9tgKiWXBBJF9D2cKVeExCqV9RTdBzb5hSBwSGWJWlWQTwGaqtZZaXF+gVFwKF
AMxwRtECl1Jny0Xfgb2U3DGW0qwjnN/7LzoEXdgDnTV9iJJMtnA/aBmjzCA7315r
77sLVf6+wgSDe7OXMPqzQWyUfD5V8FmJYboiax6RnznzBFiNQwlQi1PyRz1NOQfF
kO64Cxf73YC4Wyve0wgbzFCAMJy7AgCr23gZr50zrFjncGUh7P9icJWtQpg7X6MX
WKTQmXPrLlgScKdogc7m17Z4Nh1novkG5JybJmf23uW9kB7PuwHqOGltJnulanMW
6Qr+mC6trN+fLHQhVqYnAgRtJfMYkRnDaCJFjqymYBrwmdW9rdh6ECpSAFqRjS3H
Hh1VzkOi5oa6gqKbb44F+/DXzn/MWmhe02B4K90U9l5tupsgh9BHDC7bBB4Ussj9
2L9H7fxZE8Hgglj8Sil+lMIfh+zoVxrftFoS+BTyEN75zuj0t9PWZfPcCwLjJmyL
CutCOQ3jzfzbXJqecneCoh4tCHKlN4ztttVvwqYgfuHCwCBYPQYKAkimb1no607T
6KQI35SUGu3v1eT3whsKT9yRe6y+xHBLirLbFQK1NQ+6dg08udtoVu442cLu2s0K
bFaa0kWUJfTK3x4axSTYHk36yhhJaD2NsXeyGomb7QDL381yLgFErOtkqlnBBraU
gsEbPoBdGo3sOvm0sq1iqg85hNIyNIncCpiwfncSREPL8n3u8ES9Ipu52gWaEsL/
5SsftaXtGowIiZeyAKeDtDEVudFdyd6tGq0760iEED6yQNng30bNW4IIjTXZEs57
aImbuAi0tE6HClMwjGOvubq8jTedBmQ3TzdmsbC3Q7fbI+DjA4aiM5XgmqX35B6p
ysm82xnMq+1lkWyalrcxpbwJWOlr9V5I+p1IGal3pgCWPpYTP9dgACB9C7/kvTcF
oFzk2gXWz7R5EXS08yLeQw7g+gPntD4NFSAmTGfplNfqvaUEFd3mUMLsKadPf9Q8
ib5gotwN8kNawTOm6vSH6SxXnl2HXfYN44eUvAKMil133elS0fZKrexzAwCFT8Ba
hQy9HSi1TLjcjINd7JnJGuWWvBxDBFTnOsIIFZcJk5f6808ukmnT+tNTxAtbml29
bcE/KsOG18NozIdTE/spoQenwE1kChNe5+b+Yo9aqwCXw4yca/OoP18WAUn7nhoZ
1QD3qFoXiP0heALyuF71bgnTebqO0f/Czytl2FEWPZ73gO6B1foxsPxrVqqwylhI
RGAQL6Y9D8kuSO9ZjbuEyA2fSJMOKFnfjbXHzWxoICW0tKZwODRplKtotXtCAVJD
mPbVPkitzUjQBf1DIJTI1g00pNne3qmrVks5HnSN5JOcVDwZF5Dw8cx/2LFKDgXz
Ll23T3FcWFUti7YYRakHLv+KIJhkDiOTrckfgda+0DdyAuy/APDL7A1epRfR4odt
WDAvueJYydJJ6ZTJDvcwqn/YjY3aCddcdcV8Qb9+kGyJ2aOfT/D6O6ZNFi4nHMfv
OJAu6RSkktcjC28A5wGJPGTUtbnJjhplga0lQ03nUS7HxdrdnuYx0rB87AaGj5Nj
qkjBq95ROu6K2zbeKOXpPxc6jKDkLEqPG24J2P5LSl0wL8DpCaezIge+hwwI2EL0
v1n/NddxXf/tD+0rL0yDmtjof8Z9UMF3QW/kBzkFqjtiXv74DhzL7LVwbXu/97wg
NC2UN5hiR560N6S4bc8wVYii6OEt5uU5Te0e3/s3gb81r2bc1ebcRzySIXLOczd9
be2fI7kX5Gmnxb+StBG8rXoyvMG7fQ1Sg2xRgp9n+5RRLRr4/knyAx0cE1WmMRkL
wZrf9MK1lBUFtFjVlEPLeTEEt2iuuqmnm24rfwOZcvbkB1Mv5vjL2f69WelPCH9L
OSnC0x9y5m631yQWVe1gLT/7/odxd1WnuV6OgzE1ffeOYfcyvqybeiceZgD8saHa
i6xOv5tN0JlEI53s+Gn8kSvWOOuht9dawdZ6oaFqiGSpjGQohrVpX4pBG7jED8cm
1YVPqn+lj9tJZKp9GcRnorpxRfXGvxzPnTFRalG2u16vTqRshXITncbHr64SG/ft
+OQgOy35hDb2SoewX8uCnP1o+klgb09Jzd6bB7YQxpMUjcplDoXePaDDHN4ruVdK
Oa54P1tLJEcXMlZiuwMiz0IsITVaqK2Z2aJU5EwQMMx5uIvFTn0etKodr6ramSmw
OjkIOQfoHkcArlBWg9K/fgbetAbhY9/vjgMa9+kS/xvnjBfYgPbWLaye5muiA4WN
SkHpuVPi4+uv0cmen/GpWc1jZc8RRvpE2INej7vZWFgrNHFxN4ynNu62ZIwcAIk1
iznLLmAxliQnbkXjLT7sLEe/bRq18rti4khHm74okZsvJHH2AWFToBImWkmjnqeC
vnlXJQpR5DNaGPF0FL+rcvRXilfLe5a0I+yF1TGI3hwKr0pEVWUKD3Cjij/flsvP
ZSG2le8vlibKi/xyifROKkbBNYBHWDKpYWdXg7iwaKc35l07RHBLgWWf2vQpVOux
EsaLldrW/vRaB1lawL7IZsmvHqAR7ARkLp5tu0TlUDKpX5FzmefZEARERPErrW6H
lYHUXB9vYa0b4kThSxFo8ju45Hp5H3IKZuw5zFYGb1iOs4Sfp6pTOJYiho9d6P3R
AIemphAS98dBQz6yZygZcJqYkAIrfCwyBdKoLU1U0HnicfEhrrEFfwFlIDSi35C7
Gr8EKWoZ8Wuwq1OYFhwhKWfWpJAZikkc2FbAi/D2DFw670Qjo6H1tG1ye+js1M5m
gJIKFmx2qS/AP/2UBNxt7Akr7Jb8ijOvJyiC4E0iQwhpWk8OyF968Zs2/5xY5xl3
tTa2U8nVJ1gDjknP3o38O7ylCJmt/BcRgupKu2KMS/Lg3ly23UyHE0Hk6wfGjBhP
1W9kuozeYybIFJoz/D18iO/N/hb0Loqju0Ez8ESjQdqPaqeHHPHHEmXMEH4pkMLH
YKtQsTjdloYYIDqG4zRoTj4q3uo61re/SOyGjf98+MXY3oNAGxdAiSxMpg/VMndp
uZ3KUV9OTRG9gcywmNlMN9QcRddMvfHjbqYUTAUsbErLLjxNjvbO7Q3EPWzaX5Zz
NEKV38hxDjCcXFNWgqPFxUkNMDojOOZ25L0PwbSpcMe9xDw+c7HbrDpiLvUeKmfc
Io12bxOo46Mp01kc1phImY7VATyY5OXl0iBJDr0mnjDXr3sB07PU6uRYxu8sM0hC
PSD89lvSaKU6nJyAHvScIoQ4A8MHzngg4+zNqj1XAbhKvYAVp0F8RuFqtSQViczx
QJFn9LPbYYK9jlR6Pr3MvR400PB495roS9LzK02tkVUgtCQcK1b8i3LOPhniWDoO
OdZUzceWa9I4mes9aVpOuQSzeuPsNvl7NrUgeLcr1+bvCT0znzwCBUMb6AVhH+/c
cGq9jZ+WYjYSPYHnkUf2/fGLxjUbDVQrSgLr4N0IbIYUKUOFV89Qt0AToPq+h/ay
0KN9nR4lsnX5hLTW69hQYVEFe6kcLD1rq6Bv/42nsM3Ds7Zpt5viYY+m4OiYc79K
uACoCc/F+nbhYGzdQZRdqCLXN1Ae98gIaUn3ykw2nXhJ737vtCPUgATL+ZP57x7f
ByYq6Pw9onzc3o2fz4IOeQE4iOPe4tOc2RNMXMO+nmwDvCaP2wN0pJ0IilLUyiRm
9VPgmjR0VA+xNFtHVPQKs4AREavhUIchE9uSobswnxhoE/lL/Coz8ELvbmiE4VEY
0rBYq5I0dGuLFJjpYZpkQIdlECpCrNtcTowvNhnWhH1X0+Uk8NiuzAaZpTi4PFNe
QXFmajiq8HPLfeQRaFMRY6z9j9C6mzM7K9lYwROYZSTlDXe/eGcog848lrBB8oIY
tyZ+lbhQGDpgd6d+N0etAmvJ2uFIn5PiK4k/Z01cb+KNjrMet545+d65KFScRfXu
fUGzjJxpWQ3fybygHDEdmH9uLq5ERrJKBxicdmtW1w5XHpClQdbLRzSQR7RjtjhR
+zSB64JXfVLuELN6kqLEFKbJqqk/zPP82UelpMrqXeWcg0HkP2Yi6ay8qv7zPT9x
VDo+aYK/1Kq+sdEaExZzvz1jMa0hR4jBtLeVtGw1gkRCA9ERr5ecrB3II9J1+LpC
wt4HGHuMiDJZz2HnWkLA1Cx0RAV/Fl6TaHnthZnNcJ/foqFwgnvQKQQdfUoUClhg
/FXan5sA1Q/P/+WSu3YgGHcUG5+Nri7trOjHyldjmR5q56x+VLE+BkjjyLeOVV9n
TxXvfw2RrOgM/0YEuUfmQagPJuxwCRyMumltPW+PnbIVc6c5DK8UuCzln9NauNGl
Pi/rOQosZqJwbENCDCLYtqdtRIyW3/83uQbmDZE3jgJwRImfn8BGrO6SvkXeZPEI
cv830jAbzUSq5VA3CJPGRjPsnE/FChVca9k3vYAvJSXcdOzhO+ijN7k0giI5UAjz
lDYPomk989WUggE1LO4maXukI5w6zesmV/OD8px5MaT0w62fcox2t05iMVLfH+6S
xAj+AvdXoZqpqxb9T4xEswzveszIzZtX1I/ZKXZWNtcBaDKzZNKT9Uc4U1EGSIGn
ypaMTbF81cHVAjTiShT8l19WfkrGLlYMvIsoeYmj8ZPrSSrh3vcdJ/H+vEZMZxLo
YE7ds1wPqQ5qEPz6rNF54VNgZuFmrWyLU3CKSbtmFn8uiwd8cuSiqqyvgRL01zG5
qCTfuwQUTenMhRHqaKsJIWD6htTKNlsfbpjyCv9LvScS+PHSoAb7ktyg2nMMDkzs
LJnsvv+VpZEQskHMwV5v9ezFHvekgjOOW6GVNoPHr42d/chl8dc8pT4vii2OqZZN
m88IoknE4pG4ZeXVTN6osaf7BEpsTjcpmT+LtYGgwjRNoTCwxFG1712iCXZpC84U
sWx93JoE2n0L+51gelEiDjlQ+Mxn/RfV2labuz+nZgbwurpJIG+EXlsBYYrQxIAg
m/3yNhyNBZ7m4Z/nCFp18HoLIKTv0ZprJvZ0WIqu+/WxFj2kc/wVCjKgLECAx9Dn
+ENC81qtxmaVE4M94IyTN7qPLvpTcw20U5OLG4s/PBEguvnCQ9Eu+7EI4gRU3XU7
I//7Aku0rbiSQcPVjzIosLTbpivqDjkssxKAA19G3w6UtwLihUUqelOO+2SWUi8v
ysWOSlrfkRgURg9944/2KZau6CMG5tyGv+51I0RQ7vg8V0dJZQ2Vnsxsu8vuMT/t
pgTepc50HO1FlLfGiHUVt+K8OzDguCspxtl4/Iih+iyH0Y+6mfIuPJHFcbDaGF7q
3GBQuYqRXXwSOE4WXW9XkDWMIe0RyVDcqkkNp+I7YM1MuRKD0F5ulETu2kMnIhn9
wWtC6M3XJ9B8Zar7KxmnzqwCqvgsmJQavCBAfnJPFTulhCcoEZGGTzrkohGvk5wk
IgHWVXIFbzWkG4H6/zPUTlgfP2PUj+x4yHERb2IwM85goeccaYvc4BW1Ne3ufSfM
P11aGRN6Plp6TbGbB8k058fTfmawa10Npj1mrkAvJKdhWVgbdGyvh+5GKLLuzWZ/
7z9izWs9pLQIepRq7MsCSMTHE46/d9CkBjb1dhbtoxI0eK5yGV5Fx9IUeU8fqBpe
kAZzTmEYxtR5rnFfnXsVY/TWKkvinLxF+r1OcY7rujLQHFMtBysd45SjhC1xHZyp
ZGMXtB8Obrx9bEPhkUHVnZS5qClV4zc6oRKYrWqfNVhPsvcIXGh7vihj/tL5UwLe
DO1yoGifqp7MwOezMy6fynkKqGFOQCw1uLTktMBt0tvzJPqxewKi0Mo2fukp4fmt
cH3EPsr/6I2qlBGGTAD2gS1Ut0KOmTY25RXlsmP6ZzviRAcLqimnHt+ycDH8QNs7
V0hdL5ifzqnV1/3ymVkY+hmtWoiWXL/zXt8ccpuUKKYwQzsY+FnYzHlFsgVOKyrs
hur8vJ2gJuDCy5B+e+hCYhvLWig23BUTLUZoWuySpQbpjEjcOL/gkD+is19cp4kK
MGUjq6UiZYDr8v94Km8H20X/NuUvgWtS/Quf9TI3QeBHMXrXndGLtEUAwNF6rxEN
n2K1m6/RrJ1B+fmUElLElnod76kMGGXsHG1L9SALNoynAw7LwPPrQGQ44MpLRS9g
qy98KsutAOfTUN7vY2AmZrTjXsf/GT0r9gFiwTQrqyQPiMYGiHP6hMf6UYFLZS1p
z74QL5HHESAITmeNM7zgFmazbS9FKUTYuisMEpZhVdUiKYi9/PTWks4kF4MMg8TK
5RxbdmT5Gt8kHyAX7OK5LC+AmQvD2SHQq6CqK8H/wlez84ZRLBRkKqGNNwYAqfdi
w6yuWO8iJoQv+m9D0ZTP7l1dvdvS+WZYzJEIeKC6NRYdEln8hc1VxAXEkoWP1LQQ
NTMBLIMdUkUPkRo3BpYhwZ4nVuJQJzBkBo42P/crnKjLXw2zUEfW1UshSLx+UWfG
RkJY7B0I4JHTqL+Au4YhnWcihLJRxsXb1B36G4Keoaq7ItkmnuZVq0bakOLzNCIG
UetL7RBYfSSnN7AZ3TXDnEJNQ5+8+M8fUldcrCab+3nAAbaxS3Fnj9JdI08DjjtM
vk+pCG9hAiDPTPOh3rEFto1ZwG8/S2KIo2iiQ33lBCcfQbdwmABvZiENsTJURhVS
T6zOk78DdQaHZo8AYY6uhVm+nlTmV4e0ItQex9XQHP1zzmDIpJDQ+VoSKz4L0fzp
8WWI0qeJQG6wthXKM6Z0xlDGbDX3UQhaRk9Q+gtDRtp44IBZlqBdX9DwWattTMNP
qR1sI454LIgDU/ECxTGAZI4utwV9rCOI7kp7XPS+SYLQkIRpxtfHffVimLGGGWU9
fRnDutSACjoOmjFNTVMGmdnxbVNHxdlFkUPW1S7KGatNQR37v7734mh/+OM1qhvS
VQRYYxNhfjmnZGug+miEBNZed65SWjHodOJTl+WGbUL965qAYbSyQUx3JnLm5p1L
OaDo8R8LkmgUPNEoE8XiTNik82eb7hjJgvfdsy8iaF+WJcQiN6BR7pU1+mWiYouJ
YghySoxyzNq4fZcqJFekCgKZo5dLy5FuszSmYU9jebqYcX6Gw4YiYrrKnpj9Hheh
wbaPrxtjgOV5fs8uwarFnydAEsxs9Ya7z46uw+9PnkebCPkN4l91ad0DX/mwVosA
m7vr+/rKmix7D3QB5vvqNrQXG1/KVsYta7qrtfMUKyHe7ORl7xgCL07CXPYMARCG
nK8+bHKPemKmJoX7+CiiDD4fWyNZpl1kci6LuXSsfMOmYWO89rC4rr0mQkMVHE20
LkLYIn3iTYGIi4gipAa72vO73LqW1lKPuNGgHiP3sVdSJwmbS2S1cuoTe5p1n4dE
hWXtuks/t1fomY+kld/de/jejelbtjEPXjvgEDR1vUOvijHFh1c2rb8tToUj43dB
mLTnqqYhSlsZLvdDEc9Nxy4VAw7dTlte8mntHmnxWRPIQiRuszYLmSGsV5YjDCfX
Q9oK2n+KTJ/yptTi/Vf78/7LgxRrBXO4TNsh5BHQtSl5erGxF28d8u3wAhd8nKA8
a+yAd7g0XfO4A6D1sM/CgkKmdld0AEL0JXsfdkUnwCo+lBJEdHGYGa8C3EMu/zSm
RJAj1CweQCg5K2nWu5vw2007BRf0Tk+gREqVyKnH8K3EF67bE1gWb96/IK0ibdzZ
bru2sp0y3/agf/JhyqgRuLP7sAO9/9VoD6AYZEtYPRMatqITVdPYD3tZ0dJ8yWWm
cnNN3uwjSrvf+Ahc66EGguJhJCdQKaBLRqC8i05PC+mJEKm+PYH2KflMmATw6ihQ
kE3hcv145uJNQ8Eq84H3P1hCOGApgn6P5WbWBdd2wgfg3AaHjJmFYKW9rjuCHx5K
n88qt+ucr4wl7tWaAszDx2xr5WhW61PEZ2tHi3mm9w1s2D2dhcnz+wYKDFIqOWKr
HBPu8Ra/Itvm6KWxYdQaJwE/L+OKMWU7btKz3TtePTHryQD6ievvzHlx2qHxCgCV
k4PboOcBg6zwfhUI/dMv0GtmAsBC5i5mrd2+lVRXSdPwr4mp4Q2rWNZkYYRAmtlU
gGq2RCjrC7+9V+4CDny9UGZvR1bo+unetEkjscSwSdJbTAP1SU++A3vH+dDK++TI
7Blwoq6eiaxUNrNgRPkNlmd1PNL6Xlr4LhYnsznOvKIpwVdH9mKDZVg62VEPkUr5
naeOj71jqxjCv+7tCOwtffRfxAOPVFP2GodesS87tsmM6TL2DTS4VwS8ivrMpgyg
yYOYoNmwKEEWDneUcRAWOlhnuBYnIxYF/KwsGCbiky/WqK3ROZca6CDHZCrTdGf1
TvfUmIGg4uP32PXMc34cM34O2ZubuAaCl9VAULKIsKaSrz/t1/lYRHvKDdU+iiGK
39DPrj0xG/xm/OJcc424cVSvWjM3EDsrodcaN6H8UBwlIexXvXnzyVAMNZ1h4+S+
9hMoYe9czrPvr4ZE3qRuugoobrm8JfVzdcDp6QO27/SMM+2CAkUiwW3PLdKlRE/B
qj821R74aLZul2qZWJJNSfcBGgpdB1j+VC9iO6OUmC1L/E2ZyiJAMpOoLbWKFngA
EC1rVzjGLN6GhGyHdC7jrvlcBSp+UTIlMShAliJUAssDE05AyintPegvHllOM7Kk
XN0RC/ikRuWLTaSHNsx+HzpqRTaG8oKyTPw/ncsWW8sky+1kd+8ifIEjYzmFo9Zd
5yMs1zyKvLaPIDBdKFtPellZTVXmDuYTuX5QBfGbFdArJbazCwFDKcOdnNwAzjVp
Lupwuht54C2dqI5KXm6rTtF4gFUu2/QxPcm9Nj/BYX41ZseYybHdk9cXtAPufo1L
ncTJH6y470Pg3XUwtAkNwrguzZE0JoFPBxMEHigea6/5/wgS4DTAXWoo4s7PaTpa
5i4zf/lXm5tfUaTwi98J0Kgbr3IpesvqFGRVsP3ttzpM7zOboea1gNXOeZWvTPoB
SbZJv97C1J+LBdEGdISApJrnPMJRG3lYdjHL5h9r5QusKgF8VyMAodAp3rdBy3oj
QuyZ2xJkVsPx4jGvJJNIQgBbIuq0c9UI/TB6DcTbP2t596r+zlOummh3UkGAIzPR
XVgzrr3cIoHecUFG7E2dp3eFVAsCSyzdkQMghY6/0zc2xQxzbVBWwoYBKt2u/nX9
VjqFx4lN2NZuCDvT/r6zvbNIDHmIDtGXJYYjTea63haXTjnCMo+OBwEW+oHhKLX+
2ECTaQOLrvx/szyKWdiha0u9jobjSClA5Rr3aiXrFtLPZotlQZlSHqC955MiSufR
BbkGcYOBBbLM9rdFs7BsXoSE8bbyATai/2fGvLnu3kyvXp1HjqCt/Qx8ne63qDvS
FuPQGovnXtsSNp0r0ytYGL/ZEQywmAiv4N9Pz07aWhEwAFinZcqTCHIuKEV8Gm6L
iU17bHhT0ZrzNi16wfcKLvpwhxPYxD+Q+vfxw5vihAJmhTdov+KVYpxv8KWGohtR
8XCkSESTjOrb1z0EDdFapd6I7Oto6CQV2Qg7V9FGr4czgMbU13COU3DVD1FuEbdG
fmOMjBqtet3Hgr5pdhZrr+PoatJsSH2S0OidLvqW4GyDmnlZXHcet5g8rRWKBZxV
JmpXnedCeBkXr75ueRZ+37bGiMmV7NpX8xOVXMAZR9v2TlK5Hz+asAjHVizRx0RE
/HnaPsj9nXuPkt1yKG5f3Osej5WdV2B2OY0ST0XPh4FVbdgQNnxlR0uUgXeA9iLD
1exNmh03F1agYP+wMjkzKwiuxRKWDthIrh7eB9VAklpiok5n5a67Ia1jpOCUwKqA
C9g9nh4nCRBHkAD5zQtrAYAK6vwjfpRq5Fxjw9nfYC40mpVPbwm/+EJiEncFVs0z
BMZdw8pkJ3prkrb5kkLiUExrxZVE5YLwzYx5laO8KmtKatO5TwS4KuDgST7mGFjh
h6Mt0dwxCHzWg8goKVwfhdDWYPLZO3/B5bF/slqrY+F5o3Nfq2ezmZAXQrFfgyKj
GhbbFjjbWWf/FM5VICwTSj3yJhmx0Z78hNzB3apSgVTd5PogP1MTDSYW5PaxlcBq
xi4O7tV1oI4v0syuw7hs6GwDd7LlF0JP+G0UibyoFoNbQtOoarASf7gKysR+WRCQ
O4xJC68JwrHL0JuSZe2TLGZS3xJTsYCRsAsdpOwuxjzGEgi1F736AJglAGWhkWMM
DxxRI6VA0SwMYqcJh2OUfsayQHUk/4OiJtO8gjCRhaigVxWKYE7vwaFJtTtow1fk
CZDVKgJ66UP6DqeayoJ0Q/ItE6Z3DfD70lbiX9wxmRHKEUmbg72Uze1X+E3Xc7dr
V5Y0iQfKbFUWPAmUrckO0hZd0Mgh7olxvoGtbKkUwrOTEcB7MUQ8fbe0c/8pmk4z
V1eRRxmaViK8mo5+b7KQbxViLJFE1qiAe3HAahKcLbc8oSvqka27Zk9KJ4xRzHTx
hDVMToCxgOuNaKBESu7nX+51Se/EXtYwg6lqnfWyTrADsY6TKK3B1oqMRXyjWpR8
ZsCKDaDj+zdydwMO4+Lc9uQRMM40foyT+Nm36UXBPK/Zsi1ztR/HKpbhPfkDCSLm
sat3vwbt9wj5hFjtnn5ap/1JO3w1F48q+ftxpDpoZOZMrI0CgxsX2LpknuDxP2fP
Ame5aojadcUAlDRRyVi919cokWDNCShcpZk4mn+Tb7zaqA3CUPGf6XvOoevu9+Nu
mONoW/M2YgDdNCoi2fshb8d4DSjXY8DfZYHnJiD7IVK2M96DB2YOyK+/JP1irkiZ
P1Inugqh1bwUbT1TQpXwKfSbQqJSufY0hPQC6XCjw/CXZa/k4wBk5ulgVsQhjEru
G1X/7OE51nF+GJ9j9X0DAUdIJggyWiQ1oIefnybNfpruFa0FtkTPQNQRJwnE6PTl
hiYTTsHukdH71rz+O4r+EQfrMC8G3Kx0yBBA9IWz0aZx1WKYm0883h0Rf9ElDyBa
ygr1Qhjy2SqtytB9nrjkwuXOXC8JoyHnuK4D0eKgb4JAlBd+Orty3B5B1gftPAGw
QUwEGdaWolrQvVLxoFKNTRRLU+aiQtHIMVMwpUPH2kWLC8bvvMEbQyHeIetRjgZQ
KlLXgIvTzI++AZqIepVDI60JdAloKdsimRdC/l6USJ/CpQjHC3ZjbBhncERHky7T
tGqSCbsg/E0CNAIbdPbxjoBHKFtBWdYbfVRX/xI/PNQQ8JeFEtm6A7ZSwkUpatK7
A6EWZStR8VbPjKGvCZXIeFapUg2ClWJabGatBEjU7MDFAvtqxBJefNQjvgNdGqSx
qDwE9/wK0yaoTZW+cCOj42VClZtVqmjhcXzoGg679UbI8SnfZfPv4EWzvGroebHQ
oFDrsOlIX0mlXb3WRk/dWB/xBhaaK1mt5Mrin6VE8Kt7j1t6KVvS4e41Q5RPRL+X
qiOSFpk0W9SVgHjl7ChXpqnu/N0ouFJ4ffgy7tbN9AHHxNWCHFeOn9koMBR6eRhP
ZgGk0ra20eJus2tbzDY8bOAboE1dl+Mzv0xNE+f71SXn4BivZ/1Cthew2SHJ4sx6
DAqCYXnu7VDMRYkkRYo3uS7jlASvHhcZkxH5Q46nbT1aXlJZCrDUsYUCd8gfdOVG
91F3rZVdOnQGgsXhCAYYwcgcw1uFVxo35FSeibJ9uwGEjNbh3k3ST6qPiyG+4qhS
TcVlJwpTHQN+3jxE/b6U5vpJoUAloyFVPM9QHMIHWvPXOKDwsnBGF7EXd06q2sEB
rZAeOJ+U3s8UhAxnDdSJK1Ac0/JiE5aupR10dkh0HGD4ypKuzCZ7Ul2UpAitz3N0
69OyCBDDyE6y0Ccmimge9whB4ak6MjUG3sQRD6MlSEZvIH7b6F7lO9lfMRLzLnR/
BkxNXXL7sfCNTtpm/RDxr2gJK5vIISzcj7Ho0Luu0ULwUUY3hB1pC9ms1WI8rpel
T9cM6UJvpzPlVwcTGQ/vJK2/3p+0c8+oidW0ndM5zZD/xYUm35poL2BULjefybUE
SDZJiX4tWk7za5Ue4FlQ0lZZu3NM1YBqJr8oUecSDNzJQyK+p5eq8+0a2Kw5oNo2
Pml0PxFSofCjjMrDBshFJnU8Lv8dBixNvedqeWeRkafxMertGfF4Qg2mXHNG/pXV
H8iCZZwW6s5fQdhsa+ADau4M1VYcwh7wDnFaM9CjVGumWlqzq4RQu5s0AOPreN+r
xoCC+/pQEgeCCOLO9kufL0oA4A3HeRpwglbmTnN9FtoMQrWQDoTJXvhmOy0HOK0w
JfU+cz+x0PEQuf1iGBNHHi/qTxUobqTyb7ZiLe246vLdmPZe0WcjBeJ5P+21VxNB
uSMX4bnV8Lw2dkEiEUihd3NSAekDwjGghqAr3tWKBL/7PX+J2LEWeaEx8U8/KQBe
HJXsj/yIXAbCKfxOCIW/L22IAMY3YaMLjBAOmhDeUw0WI7avAezxsMgO+fooN6Sq
whfe8ZDd9aAN/5FsJDPfpmdBC5W4ALss17kuSKGtM0gUUPpcNhiMqC0T+yp6rIiO
JxlVY/qhjJdalF35ZqdCP75QbXwEwzOyXk3f3jINzCUV75OPLfIf30fGo9TmyBbL
h4zIwF2OTm6l0j6z3IxxDwSLAbpTsaDfzjP4ALomGQNg/wck9/e9yuh7d99C25JP
/lKV/48oDSf3bHB/B9LwNorFmApA6cEGjGeZXGJPKHGn2eZwoAlEH5tlxIahdKLO
ia+Kei8EFZ/3OT3SHjbCKCyL8mnm4Jp5k+66lKPsuaQMpjWp9TLb7JukjAnWo/3b
oqc7DkNzT7YP5+Gvqs8Rd0Zx21Vo/x/LS2yIg0UgD5vUnN+GZoJOPkDjYq8pqLHN
awb4WfivyAmfpR++ZWS6XUC2ULa5YWPJnSg4rKV7po5hvV+zyW91DkhPhf8KS77q
LZLf6rtOrV9iekPng3yrB6GGlDbNKNMxSKsZWZL6hfBZolhRbU3nZLvZcAwvuM5E
gM3oiCxCz/KrqwIM6Has7oLKzfnHLVrMhQBg9bcaIrEzT7wd4PAO8kgRWeLoJe4Y
CWY9VUZ4Vsa3YHJK9NLZ2KUw1vzv3kW7ndkgY59zZwe7xfVNhjbMMwwzaIsdfN8t
jS17v/PYt973bJK3ZIKiDqJh313wmoG57muajm31nM0hPt0h5jBfhIu5R11KIAvQ
bRkl3gvq9ClqTeBolAQiiCYX0++1N5qzc8lkCuWmAbyRDUG77MuJvJx2Vwn9N3Ja
LCmdoQyh8YBRb7LEtJoMQeX5t20LID9SR4vy9R7eNft/IsTTr3htRbZwE4O9bnQv
yO4qUjFEcYAPQ7AtSPEW6+YpljPNOPpn7w+W5F/i5cW5sStGPZ1MKTrQtEiFJeS7
orai4rqKPzR90xacZmQoO8OCQ7ASaInZuSYNzxF1KN2NXG+Ik6Dhym9yJ2rrdPfb
FF3LFvJMrsPT6c8rA9O9EwyUS+NHJyvVcbw6lcYKMpIwLxj0IGU3SeNOFVRIlspn
cwMSZ7WJQG1uaCU5wjliOHV7Dgw+t/XsC6kJXdKbg4Oy+qNxac0OEU69Gk0sGgRj
WHe+cyxj0h21pAlwNyanRLaXZYHvLEmpF/FZrhDBTQDEaKJ/CQtRzFRKT7kBUicK
uVAHqNDZht7wsRuSEVz8075baXeLN8Sn1AoXKdBetWHXyoSpmpxNzv3eFTL+jBBP
CRTUn3tTDK+dYqIfJleeb0JZxpGjupZ7aZsjZM42KfithHQaMfMiUycbiCho6VdR
24Eiktml1eQFNgHPacezMb5x5mZR80DWBCdiSOsp72+cJUYgXmgQTzdJoeAaatR0
lLLrVm3yx9FJcVT3hIrfb0MAD7XHXLrtFnQiKr6cHj3pY3sKXIWewqrUiMQGE2BP
qjbil2o8WQHisbsf31WnttUiEjzjqQyujzjdST3bZ4CWrL6FgtN7YpqcA5wqfSNd
vAOVRCcG7l9RXBcAGm5N9Nt/bylPmQOsqKHX38nbzazbNU6aVqmfw+0KPUZStrw1
AT74Oi98kcwQMNWhSk56RDgWNP2/cedgatYHqSZEkT7ljVV+XbzDuwLNVQxZKron
0OMBU2N9ear3835o0EggK27Fti30OsW3e/XdFW2guPM/nLwXeq9Rxr77z1JPVVET
uiLN2yQmRfQDT5fs8lCbIj+BpFdn/82CfzaPgwQnkBcloHruy8B7CYPgGRxLk1tQ
XflE49w91cuUaHiyc/eKEYw6oe5ZfSLBuBhephUk/RLe3NmdYmkcHYHCtA0EXYMq
OmOJz1wLXgZ2HEXd7Gb5HY5HIaR+Rgs052DLtSFh4joyTYLC2Tw4xPrnMwF9aIvO
AbXDFrPKNto5a8CmSvO9qgNCrvO7Tof7LW10ws2rSTHQaljnvwenH06ob0zPOGmX
P83yKELfQ4IHciqw2M5M89A8kKUvOwgSQa5HpYBOaWRGsBL2Mwd9duDqioJ9D9On
f9xjDiHOZjaixMTgmo+M+mc0yNp8vgu2cbGRDW4guSFdkTb2smYgB0tAKApsdLsW
FTOTPzGXkcpEy1aFsQucsjYihtP8nqAuqne5DCbBoc7mbM3JzhDyKJHFAya0JwS6
hoZCn2ZKYT4KymrJqmAOVW2ZTwyx4miMwaN60frDZjIaGc2t3G1KUoimNcWYbWwh
zDdmzpkgNWFjcEO3vCZEzVmM6qfvvUFuCP4TH324Q3ILoy/RBkhKsNhcX/Y5bafR
l5LBi8934uDt53SLUUdCsBmFB1uGYmd7oMrtPxC1DRjNDd9SV01z8OET/0izV/5v
hFnp/aI38ohlQ0XQ7PTQpXCr3nU9uIy2BmSUyJ1BQ2OPXZ/M/r63K35dbmVu5CPK
/DQs41Z9DL5Fx7+pwvE6+gYIGl9ErGVR6W+itY2MW1z9NxrWmCvjL0c2OucqPhaK
bxUUpwAcXCOe6YGpejD19d8WO0byxgKY2ZHcZrTci/52iSKURp4fzRaA8vN7Kbik
2nMYV7GBQtlWFtInVhvNkS0Q32E5PWBG61efzEjRnK+VgnyAE4GEy281SDgcbYow
1CTv6OZSONmv4BPL+66Dob7uO4ya+uvpmzHvKEtIjJ10sAFwOg+tcT+7Qiv+ixl/
IkPpSUq5Wvfum1MuY38aP+J62zMomYZ7vZd/IRRChYnDXwJ7a2tBGsYr2gf0Y5s+
GZ/SjRFuhdES+Jprf39aJ2hn8GojUptizLvYyX/o5Ebk7pI/dMi4y201VWYc9d5/
wiVyq2A7Eo42e4muP+AUkS7k7r//ArQMZswN47ugYeiDvar+Y8Y3uv6yC5TU9B7I
VGMaUg7MVaTEA0/QVisOgsOPOXNcOSOaeaM9ErzIW40khL5Yyqg0p4+TbvAHk29r
dsSRv5YDK09Tf+qr5eB8uA8a86yKvSKY0Qa1DelGO1LEdp5aUmfin2ovs6AOJh0/
H5yCUM/DZYGFu2HpZ3fN4ZK4PhMoA94T2rt/t4ds59L54pB03mwLyYxyC0UeK60M
aJv3npcaLAUIh6f6WKQ+8+i4SoKdSw75sTmF/7pJgXxctWpgpodOfFeww0XMxXr/
PWXsI96Btci4z5m1uDHVtXbR1qt5qgpZsW7fvF6o9siUb0LRA7LSqTdY7UfeIRUo
Q0YHLt+2eT8CDJT7hnjPm3iSIIQiyBqC6dqSG46Nkz1xHLLg6O6LIySA9McZonn0
kxlZ/MdTZAn5kvfTpSuVX59zsv8trV+xQbjkpVcCfrHdQrpMrcV/bspFe5NdCaQ7
sWWo2Y2ilNn8svtnu1b8DS2qAm7CK1MKZr7ObBorTV+Z5pNo9sZfdqREBlm2E64Y
V4hebEHeOwYe7uQy6a8kJf8RhbBsm5z5GUjNk3iZfaHAFs7+9htrw66evdT1b4O+
tXNzm0doEi9XFiqVBwUj1hq6mg1xmHb8g6fuB+R7hiy+qMFOXaQjD/iMi1/Pjo83
FFlb33ZCn7f8Zk6buSrMUj+3GW4OP7BkmWX5oUf/Dx9PIlT8QYI9Zb4V+fZ8AXNY
IyLpgTmjsntf4grrITEDCPQwjJ85+SRHLQ6AJVJtI+d3hwCzYd5T/IMoBiuboGdy
YKzbv71w8QvOezbmx+izPcxyiAezNzEGDG41auWdUJ3YUHBjjtsspKMJD/o7cI0g
Db/jF5mB/heMTvS9DmekNw2UAADT/GyEeCgraZxRj2HBsDQxjIwL4i/Yjl3vjFdu
j5Cf+a8DsGM6R9ySOOlN+O6+9jtUzVNihX1/X8c0pe4a4iP7V3LSGcTPZ2epBbkY
+oL8NohpBDVhkPJFKzf1sRRXZm5CKdy7f4wByqyyGeEoaixWuZzhbcM+GsHysF9h
nXRVa8RxzohDwYErh3zeStqLkA0CIgRtFXsbP3MxX52BkkdBICo1R1nC77IthGgd
f7iQhKrmlHNjEdnW2ULt11Q56GZfi2wDbL3eX0t9eeLIS10UOHIsJjTN0t60XO+s
CjSUNJXQ5rE2alA2oIJJrWIDTODeE/tzHuU94nq71VntDV/HreNlaQ+UO5yqMupH
Qu8YVsaDcKOHhn1c30NuyAJCvrne7In4h3/0VJoEQnG/bGLOQf1kDuYQVs1A04mO
pfyCmnQkqeJz8basELJUGXr2CW4T1lSkcwU6HCRRYkDxnqO/TZv8b7quYaXBdLJ1
ONdiI2Sup70ItsXKUg1fusbDxv8rXSmGJJnoIIWFdluhLRyyXG3oywIGZPdLzwV9
MaVTMDkSbDFFF+y+c/au4atUny91kYJj+25VU7ih2x904BBd7A0B2gtZmu5BdEoN
6gwvFwMcS9M6fTPQa8qXSbHbzt035F7WSpmr4EIZb5lf5zoiJDBNpfAZWVqtcUA2
EclV/G38s852cp3JYps+1VrELnYrpqeFrkGNt1b6GZAnOG9DkAsfKhDdXW2lhz+i
V5iFF67MenVkz/5WPyekAwmemiA+DrWyBwaNPFAj7cean2Lp7y/4YneNEkwM1hYV
VMEwlP2y9HUEDl41KUh1HnsAuO7lWx9jo7/5s02INdRT24UNG7B8yJy3h933P/cE
z/0NbIZ38DMFvCqdmayxj57QOKmdhe6ooCYDs1KE143WV8TMvc3BeLRby3EuF5XU
4pjf8RTAlcE8EUlJz7AfsSggFu7B2Dih4Z+052RCBEaHgU4iRsDJohQrHI9IAgoT
ovlAslA86QaIlYyxETPSHzHVWIRNzMbXT20WQJAxfg1LxrsTHUDFzMUec9fExjH9
Glz0R33knLyfBtBRkf6ia4AEQy+7A9DkaDU8gRbRZx7hLXQ2ruytZaM2ElqjxDWV
yKdP4tC5dP6cfbUa9EDaYco4oG+9/J/3Dm57EdAbxwF8gZggSX/beOkEvheWm7Or
gosyojdKnDzmirTKSSPvhX9rTRrEsUKRbUHge3elSXG/btUnMVObsJfF2kM4fmCg
3Yuf/Xtwrq1GdxmCgn8xvg/t0akLnIcXj5dDExmvfq/JLJxwsnXlvKuJ8SpxSBPq
t7bSh9BF16gifeuf16CUmnVReYezO79mGXldFhqqLM+zNj9ZrOjOos5FCIOykZxj
kdW+d45BenV1k9gwVPC7CiWIEpHu82KFGq40mI3ecf1+tCYyPtZITWdBnrlx3V6m
2FAumtnredR3ruRPyPBPWZWr0VLx8tOFnEYVlpo1TigRE5/g47DeRs3E6nQ1c/cu
VlMuUTBLDo1Owq4TaTTgnqwJ5WRObIxa+tMF2c6YneeihkO6i7Lf4o367UEhRuaK
YlKB0ZXIgGsejWg+ZJtNsH5WRJII4SHF57WzzvKvKzbiDIjDU7njWTXKcDUGxLXr
nRm3Qsy+MxJLnBSfTqtZm4Syf3xpjJAK62sUgK23M/y9XANEOV3u/ujHEl4xE+Fo
nR/GckyUQl5usH1hIpQpMK4+Xbpsho5Wv0fnEelflLmMbt9LLo4OTliu1uSHnkK4
/5OU4t85wjQAJ7XX2Hb6OYQTyCZuZikO62eTxTWVBNL5kcC72cafd+hGVYxK5dE4
lXp4wEozfTAK3cMGkwmDy607WvxeFQtHkHORbnQn/55CU9tCw73HBArnt18a4m5V
WWGjo4GN9opSEsQkCIVBV5Pwy4uMURK4hOiAYaivfXDdypBsfwQWymRfm9yTOJts
ep/Tp4QD07l0BYBcrPoSUMjErUjNoM8V5mGkdodKtQkWqtoWI+VaOXEPou9zoeKQ
ge2Yvvqe2EnvVMnRJw1rT6BhI69KYSfvS/JGfpMI+1U+YKOQEnGHqAk9LpYBV4Ca
jZPOtjBhWrp6kkWYgWxBDcZInl4Ggh/0cyVSXun+1BujRWyQDuEq/52YWa8Na0lU
LX7lvjzDSIK+4s+8uYBt2080Omlnkk/Wge/OAKJWRcJ83rrfs4LrVtgHufryWqZw
Zhmew20MwRKhGCfCiHQj6N4auNOAubH+kbYPqBwkJbu6C3BgBWVDq4PQBmi5AaF6
1v0OB1Fglsi9u+gjLN5WMUizZ85GTpWDdUeHSgD8FtvwKs+2YwYPJN/bXNHvAFyV
K3upsgYwigybp/sF3dVDiWQnFx5DLdzn7ctpA5oGdL2YNaiGMsJSCufs8v1p31bH
wak6junCMYLYr816DnnR71Jjs+3Q4oc4h/mQ/peRkxOfaoIHUom79yaUcLOsvWzL
nuUdt4jzOfaFrNj5SIS8ickST3oHf4JPQtoP8fhzGT3VVy8N4g9w29gIWTruWF7t
Ei9ttm6+KENYb9PwFl36t5eYVdZaZSTOJqoT+am8VZitIC0evCyK/53de+AeGmT0
8EuUv1uD+oyjoBKT7r1yNMh5ERLNkCfpKAbd58w3XDPPY8oBgQGCNPojZZxTtfKT
T4BYV6WwwXvNFH+M1d0pA5r2VDTLka1AQDy3blf49carHu9hwsoUvdr+PCw5ycX+
mAtcQYCAJ/GGa+jtv0KfCv5avz39IlAneZJqZYofw3mCiSlP1fYoqntAH4yL+Tip
lxdCz8ZoB2hww3C/eM8u4dZPPfGB6lnkqgONS/4ZqGDL02KGqMhlnBX4Epe64Ryn
6L3INkKo7U/7jOx2PBYFDI17LI8Id7tru/eH7v1IjJl6DJEQhpL+f/iFhH/bWgRo
pekNSNX1gJgRTCmlUsrJi6nRVeoUA3XOO6hWBog6ab6Jr5VeRJTaPBv0Az1iMKIu
oRfP1V5PgzwrxwEvPhGtq3cY8O78Fdl24235RTlicdbZH/r86xA7xDynQpN7FnMQ
F14Kokg2m7qwjivAgY2bqn2xW/feUodfRF988M/ypvhEhTl3AU+2sewk3Di+Jc4e
FjS1SHvCH+aJlnSwRa9NlkPNiwJzoHBqSEJgNW9TLFXjAl4zc4Pc0r3g8PpVRUhR
dMMHPFwsX0CeubJCaOB1we6wDqabtPEYgcoDHkbjToxmLVZ/HayFtjd8nW0oWrv2
wk77q+9146dUWwg5SXA1200EWkqKQZUWtzKNiWHz5NLAfALBq2r/HEBHof14WmcW
aqbmHpp3e0DXO792iMr182mClN0xEQNTTD/wn9MQ4py2gPKYZEp7wFI71HDTtcEq
S0abGw8PyeJHZL8XXHFRuAG7lx5CVRWEvFGuOeNpGmFKBcM5rfHDo26Ik16iC1u5
f0MIYsUbx1eyVUzwbVFig4rmRUChz8GjOtJ63cDn8KjYAxQ1Q2wL93hHMb+XQzpR
Yi9cOkaIFrAVaH0+XXsToKOnJp7uzkDGTpp59MziLio5b2IKSQqX1JEVZVbk6zHP
7gjqwZwq2pOpnKE9RzfxUu9D6YhJ/ESE+8mDPkpO6q/HXJNcYfO+KBucF9hzox1+
nsMgEXtzseDxzGICWdH4DdFJXwoG0bJGv/+rMyc3Ie3TGglChsuuXlPzwh5W4cXB
der0DrUq+/mpJnCObPA1Cys/1ddiVnZfXb6U6htS+4A3r8RYXscS8kiIkApYmTkF
zvGiw54QXiUnJZ7Zpn+NikbRNSpQ1OfuVA4pWIck9dba9uJgXBsyIaLFoR2rlyxD
0mx3eATFMTHLal467ldHFYrmredIStsUyXNzcPA2hyExtkIa7Y+RoO0ITNiXlwZp
Y2/qgEbtHHg24FyU4TF3OSqpLmhu+czaUAe58uvOlGZdFreGLFZiYGfCGBkvGsFY
gdlbRRtL/H30BPLUdCY8cmdZVk9lmfzLEzmViLf9Gv9ZTtMYXKu+R+vPw9GtiabE
XzHMil3hxzGP7JFG1s6BKqyQMHZIZrKpsgRwWKcGgnqn+Zw4d+yvicxU6F1KD/+H
xLs6yXXyKcnX0Iv+Y+6p9eWPz/wJc0HtLiRN7fHf9FZVot/NQGUa56P6smLU9+pe
J1Q2Qt/Tj21evrlaG6a08stf5MKRUU15h7EcOwsvvhvNF6r0yu3k7g4aUz2biA1x
RkLQobhAnsTRCJaq5Flzr606GMYgtTa3R9S2JT5xHqyZWM66fjqTgw/6XFnO/bWc
pZST6jj0TcNEj3SXhOlOj9OThl749Ntv1djLkHfwLvQqQYj6vpY14W7PTAumX1ra
rfLqfkf1NVSWX2GdseOYAv2YaAFXWVQiHh4iG1r1p2UGtzHGq2wAkIaDiwZO+lm7
95J2vIphOo3AViMJTveJnOqMtcSDN5oHeVEefztulom2GwsRT3lLyi9BZszedOL2
fFIaxHzWCovn+aez2tPxu6zfsM+xKo0Y/4GTCvmPHR0wePPamiVR/VnZzfE2KZVn
8REG/PggHvS+HMFJrv8Is6a82+NLwjy/SPJE1v5HlUoB8GUyrxCrPpP03Qb3MOO9
BdXjUs9nfgOV4p0bT64at3/YeLfUWow9EmVP+l6qu0Ls1d/gAEfUDWeVLsmM9ZVE
82gsaUNIsYAI9tsM/YiChHCRDO81kfk2AgSy5IylOGG2CA5UASYZfwWXplyx1JvQ
fOwpblIJjQgwOfQQ7ZQ+GDwt+L3m4Eg7HXtIMXYOhgUpvgR5JQlNPnyDwx8qhLnn
ywtyf84jAujLEDSSbrxZ2foUpy9gUYgjbOI91IselDrLsURMWPE95qJa5lFCzMl7
CcYWNSkhVSgr5Zcd1ds9NY9LvNw7HOA63Hi8VwZbvg98i61ywevbU3uCSy0B0Tjd
yn85+Lsj2Vf6h9szGYgAinarVGq2n+JxGXtGF5dHf1vg2CcNkdWIjNTC3RTTBzsX
nNM8u8mQiPpOF+/4viv0n9IGzdsbcheUgJGz3A/k216c4iF1MPZ0i6ozl6trD9kt
EKFdctCTLIvO3+/mORQoIQI2gubmmaEExgqRP8EAnk5Xfe0SEWKnKYGBAXCMWZTH
BEKTj9G1rE1jWexSG/FN7WdnnnjBRLJu+q3A1tblCZR/ppASzxdt2ywR847X7j9h
L/CSREYKRHLhpmmXKF8LP7dJNqwmlT9nMp0ZQFZCB3XZG8NNvlnXFw9u7JQrMTdm
PWISqrHy6JWiVc2YQ9aAUvw6+3aExNVBsGbqf+ACVP53c1PDzmPXp0ILX+Xl0lTR
4nNOPmnzT+c+v6NWoWMjk0T/ILgOMqBUb+Cl7DxzeDdx6sqp1Fgc6JPlq5+Jq38N
Frfb8noRpznA8syer9ori9cUxp4qsXgUOrf9chpMyU2Q8hbUEGtzeybIJ4tJxuy/
6WfPz8A+fwFc7sLAlpQia/e9Pq5BI0vh5A+LRN+xjLV6kCPl4LzMDE8EQCV2ujIO
RPtcygT2lZeWzpSmyTboBh+Jnn8itlozbK4cbRjnKvdxDZPlytAu4XZJnW9zCI73
rUyzGIdNEl0L04jGuh/8ZmnGAAxd6yjLpkiWclmpLUfN/9cvA4tm44fUMKBPbVAS
uzTDWeoGGmFxt2lYkFlfEYH2aAsiNHG+WSw22GjPjCU33z0IEsHeztJlfUvECOqQ
51RG0LtjwoTO6Z4d1xN0sBpLbs8rXZ2ILqb45EctgLBGEYVc4a3PNj3C7R9EX7Q/
S5/8gqJ1Hx363ZjlsMQIWhSafQOa0quSHLjGwdYW4ieDuPATsveRCC9rCt+Io608
nciRv352cVefA1SpUZWyudvBA6qo94plD8SYOOq9SWV8MSQQaTCeGubZyHege++1
9DCatLJmLR6INIcUZI7UirCy0JQl73OedpB4Gc3yvNw+Hfl6zb+IA41aNESjt7lp
ZWLy17L9P0pRUZkYadvx3vi6cgTmBqXKe+rUxCiM0UrP6ttutHZAPbhlM/WhZCkd
GPFGGKpSWk4HpuKgzIRuq+eEtbXMr78Dy0Uwhi+dFcTecV+cs+fOHqqr1Zkg/bcl
mIhDHQiVadpQjXgY6QNpWQVPgGdc+HFrddZ/WcudivXKp98KeIcgL2VANzTe7khJ
6jZ1kT0jCcTLSo/202iwmfA8c0h63imfn21GfiX26+Dw8q/o6UhqEifIj7mru7VO
0hn1iIJuVAsCEaRHXWziSdHcrCQ2z+eY8ZuLGRhVF0YKXZ6wEMD/inBImwvfTtVf
/BhcLZ3lH7CJeB8U+DM5WbnPM9YIol1XpTgy1UGuSumFCXPJilu0snL6owQN6Jq2
fQk23Qt5DoGllHAxjv0q3IhbUG/cIXAIV8B5FI7/FPO8QuDymYK7MRiGiX/d1mZs
ctrn8Tz8D6PoZD/BgtqTd70EfLJgw+ahaCg5StucvTtcxpOrv9KeqtOno9Lp8Usa
m+/TWsfJ0I8LzfhAWphJhvWRuzauE8GgGkXH3SNgO1ym8j2rSfHnDQkAEoXbm0c4
31ZoEpm4migOWbBs3o+qRjN+lXHIu98CITyT+aXJrm13MQd4Ya328cUFIF9+8oRW
/ZE2FD1zcpDVF5XrqPhZRex4h4KBavWkUKhpFpCAxwrxM/63ivIfBsuYyhharQbK
HaBRE7cWzz+O+up1LQJA+cPBojMK5bKz2ru3HBvogWGOhbguqg91Vk8aTtwCBfy7
2BOK+2qqXcUfnOFrOu/1ErsezNPvbjAzgdLn2i/g95wEnpaoQAhyncgGOxhsxQxr
H13UET39ELYLCe+j3CdjTQBwcbKOqj4BW2xvoQGZw9LFlO/J56vdLozEblp5DrDw
3MMMUo5F6OngE3Py+BMaZPjXtOQXu7nRlvUgW5yfpMqgN9OGSuPzjJQSouVddhB1
VE3jtE0ZIuQb1Qoa4EtIZkntgYSLFkB5B9NS+35MtqqGRkNVXazVYty/5Xzrtxfg
ciqmvVidpJ+94Fq43qL5eiaepZ0Sr4ICDm2/kg1E3fExQyxhlDbCFTldatyEINls
o4UCQSWE801IC7ZH4MfmakWC9sfmvZ/EM+S/d+4gSkoZubJ3ISWufx7UT3AFyYhI
X4Q+D/ZW6UkItLcicckET98F/IhcK3fSQNXPz15EozNMHUwQ9V1/847XgGvc9Y68
RIa0kC8dadkqYzXdwUj8A+UibWOD9MYJA+dSeZxYa9DqQY8e6bHfR8nEu1rCFzn/
JyKhTS5hNQJi+w48+l3wG24ADaX823NE0eYUVmG/PNG+HvQpw3uSykc59r3f0TxG
YcoIInI+5u/l4K8NZTY8jsfJbnwRO1qxeL0kv5ohhC8auV7hEKwFetf+qQSnxcv4
U5kx/Yi6/6trlpgy4LdBpoRvDaDCgLC/3HC0qCwjPkKk9M4YXUhI9RB+MiO4gc/d
hqMsbBVZP+SYbAxv5xGFLMb9k+FKzmEtNE/RoZneM0u7QL7iL4vb2ts+ZdWvvFk9
t/w3+JyPkboBDZSFTxdf7738AhuxC3IbTEsNGxV/fecYCttwb6DrcvydXmIwTAmH
aiIizOrFAXwRG+IZyxGIejrJcfujoJ1tE11aqcU1EziA1ejAKNJ2Im+EV7b+bJJz
aWYVf9Vr3aE6/xMHyOsbAbFlzxXELh+N4pAme+0PH897SJyj7KyuZaEMr7jKDGqV
LyIBfbbMdmGhx2j2Zvqw9ueOvB+vKNzcqrbClY/JhLVADQaj4r2IqT+m1TFR2hS4
y7BAwFZeZkiN+j9rfYpc48Qf7C4STju9xbwkJtkYKRd6YXu9l525zh8T2cz/kD/L
Vilt63OzlOqDF7gcRXfydXhOxU04O66bCGo5/ksV/RzX4uiOWB+XcMR3Z1TH2Vvx
K3TJ16t1iY+AVgzfzkXdS0/esBA+m4qWjCkGL6p2u9lzrEj8RYlbTnglwubqSNZC
7WgMLTPjVLCByjquVRqRq0IPnyI04UVcs1gqOfeAVxNKSWPt3juytMEiH/1QuEAg
PxxClrrbbBULWiI0I4hjd9wOKvvzMGu/lUJg5j2IZCWlDaoTYDp5us9snsHKo8fM
StD97FuYO0PgylgshGWai1gpyjJMamhy+LuIe1xp1GpNqNL1vSSJWYmp8tVgsUYB
I+T1Ii9IuMyUutV9ylo+BHTbPaYul0ePQEq1TTvixOVNao7IXDh0+Qyrue+kOPsX
LNUXYAVPr3tw/80Vq6UT1FvNDbtD4mn1Kx1yFPYw4dIpgV1XtLJf5j30lhqYzbEI
0hEFHjQctxJTsHoAnXazsxYPtjlYtq/ZiCI5J1Tf6jeZK4V0myCoFw+LBcep7ljg
B1MmbYi4o/EC2ZOyQRYBG1apuDdWDCUn4jKt29Wd1u+HNqkAJCs5/tkJNJDe10Zt
HmNzJEzBtQWQzij9UmFclZPQi06Dd7h/a0SibjA92IHBvpvrhvr+H1Ug798HP3wh
e/o+/rjjqfqOyVYDXh254dhoq8xxy6EV17gcJjl1K9VPuG+fqyFGB5jPpQh/C3Ea
nDdMYxyvhsH1pMK7ICL734gnZXiDf+LOV7jKs+a1nPupzFEmUYCFF4ZU79x3553R
4TvYa2CHy8Q4n3sZmh18f9lSUOBkVY+GRuzDs1nf8ci7M8XA7xrRU/v9kYpoaeDk
MTXpQSsHULuxqC+XmboNppquo17cY6EHaQ1Rl4PrF8UbxjPiXvzVlKBKhYQ0VBvn
c70zk0hokWhJWaYO8nWTOaXRDWyUWTmZ/CpWxGG3nmQVCYRcuuEmpzCjdg3yC6ol
xOUMaq+TElfnkM2uKcIiQfTiWWjyu4x67WbFHZ2i+sC93iRzbf5vPH5/PHeFJWb8
I3pFfCvi0rLO7etN/QHUQj6u0WRhkaJ7c7OGKQPt3hsARpQ/XCYb8EWyXMDnD8q3
oOSsCPgC9DksSUJeVZcle0/1MmXn259SxSsF/ypx+1O9bLXGBWYVOGqHigy3XvHU
9Q4OdgIBmFgORYct5H8fMFbfNDT9Od/P+Y+eIJJSLoBjkjC4he5R/q1BjVSbtY19
IEazhd+PaIamHRK2B1wlFwLJCT6jcVz9pUqe4j2P+1YFJMYNbQ9gLbkiq1O7Rrl2
/yuzBhvWpVjzvpUcuu1aPOvWVfYjv4iLV7x7cM2+/eD8jIhFE0GnRNumO58cOvzr
kGoAPfiSsYHFWHjnTs7hfd5VupPDzS8N7XmDBx6Rkh3a9lfcg1mjLZPV7JZk3Y/n
5URQWdtYbMEWAv7Ul7Wl0xVizfL6BFONdQHHH23NTTjXgVxYzpc16ALOgs/d/efu
dtLvyaZ/vf/MJXHCm17Nk6TiyCXfcPzBS3KulDGUsFL4Pl2xj/bJHJoFeAM4hzLS
g8ChG8h+wSyuBAKxtgxvkxpAfbqAGBRv5zfYtrn5aSxc+CIaK0Oxuv81/qoZ1n3U
hy4F94O0jQRcouNmO6Erg+3VSwkiTk9syl0GzMcMC40gzFiJRSDAHVFUGjAmjpDe
bYWVAAq7Zy/kJ9sKaE9GSJrcyh0AOi5j6I1ScoCWg0hF7e9UmblSlRWZ15Qvme9N
sBIKmFxxvIgH0NKs7/oXI7e2RJvkAbmvuzJ/d5ctne3ULSSAZ7Ns2PRblckAvm99
dBWIkI3Sm11FK6G1LN5iMeIyQhUILgLYSgcnIvfEdkK7FsV6fhmlx1Oy9B2kBuIl
NHaYocO1wYNiF7istzyTrZ8oO4a+JT3+wYTxsm04mIwBL5bLFOP/ZsaNJVUpLwto
VirTZY7faYEBhmSTV15Gtzqivqu+zhduqETaGjAxZ0DCEr73fMBghoxCU7rMwjI2
sFFj5gqFjEIUqH4Pt6d2AJjjRrB5ECPPNfMcS+w/337+jDliHEXZLjPvffJ02Jza
lLdgwqL96X6wdId+C1U4QCKyAEYyduPVR4WqtxTDulFHk7X7QFbGqMIfaa+laj4N
uTKGP2/xCblDf1iV9JJKkBZP13eTb5XgkZlLwVWa6eXGA+4gFqlI8pFV369RUYsc
ynjibWO5n3yJjbFghAdTYtduNDeBFA0TLfj0Hi82zKsG+2n/ZIE4X9IJ00Pogqqz
SFe0c8ccQQDBG1CT6/qCI0LcjPMTunz1S2MnpQ/B/3Oyd/Qd+hC5QooAf6M0rPqP
usDg/UrSUVxT9rIPok4JP5oAUfjhcpk6GPtC1FRgEK/MXlj2yQu5FdmaOxZkRUFv
OTn87wo0P3r5PY8yc89kC1CdNePTYoGNwOZ0fgxHyvouWTL6i4T2cW5kCgsliu6a
YaCm5UzQfFw6xXYCrBGZYxd2j04GBBlrfyb8EmL/xaAwlqg8RCq67eT7uItaovlj
mcxElxOwunjIBNI57CIbRB3ggkT9cU5PRO3ybJ317Td2GgujaPzSA1mDm/O6xx1P
DwIXsz0Una0N4BOYaZVcK07tqqTNM3ctEFybswqd6TFP50ugl8cyn+QBZfhfce8U
SC0VABBMb2DzMm7MX5ibeh6IMN7wK00TwqFNOHMeAia42eS6dY3ravEOAh2VyTDN
zgyezSFg0KFZnPlPBD2KzyJx9QFfdLbIJ8KSQPUwU4aVzIv6nSd1dyw6OeEQlInF
PEJLi2Q7UWzItrybp64nSExF8awqXJ+Q35irXm2b5c/ZWm4vxOzYPTWqyeYoFctJ
7juMUop2L3tItLYdHzg4T3ZIYXoKz0HFKJGt7AcfIxn9lBL/LNYfPCUH50FKGbPm
eR9A4GOdv9GelLjn85hjU8UvFPRIlxsXZpxboU/wBNzntoXArjUsuBr5WsGflSWH
By+j0tIn9OSUpQd8Kupsz0xlXCauAwC/JLsIOrTN0qmO2n2mm5iG1MFum2TOUi1u
ha5lzkdYFBevw68SK9kQyclSv/dRAVU6A8TU/5uWEcLaGACNSMVf2aTlzgk4YsfW
W3u2Pl8Pz5NzmR/QNGeJ2h12p/a2LvKEob8ipVA6FTutTDAKKHnvkD2hvQpwCEZB
UEFaQqiyyWZrv9y+TaUewvG/sD6O3uQ0SIgc12YAP04ma0zlZk1esfKy+3TNuDId
zvbWBX9Ipi+Q5IU+eMymXf5BeWnwKF1h6KcWuoVQjoX3JuzJndFUf9LGUV9gYrXx
kmggGQJ+Sl1CazcrQO9BVTIpGq5k0Q1PJepozGPQmv2WCTisqB7mqtWvG9eSt6+M
N3lUjw3fhNngqhsnEcoJHwYMCzMmsn5pN5/+XsK5yhlaaeszqM6xBUM9Eha8vD/3
m2LEXJpKcwr+zEFTpC60c7TDL4+G1uyGNwqEqheGLWSML/VKeN+3Q9iguyxuDJzR
LrblyDDCQAwPQNSIJteugyOagyQpJXtMlN1uLyNWmUqNwZyjJ52dFYMk0IMR9R72
JxUo7GmfhxxfJIGn/hHKrxL/dwcNOUGmdgixreRTivVJgTZv0rZKg6cQrTocr0WU
ZY6EgWSOCYtH0+ReZsnsfJWDb3Afdem6Y118sKggDyzSJjsF8lR/owL6pob0kJLy
NFwEE8VTr95y44f4zv3lmpZtaVSfXI7sTQZKBJd9WHKu5+FqqnIETo2eAZEpK9Qm
RL1k16eSQdiSi6QuNiFm/8JqDvFZAhGhm+hrsI1hNNlnKURE/BPwJjL4c54RAiNC
/EwauIFj2MqOwAbhT6tO1Vs1VwX+GBnJomrDvLVUkJLMnIsuE8zqaK79v1ab8wDt
7DVOzclyHXus7wL5fijB2M/mDlMoz+2Sfo1yXMTPd79zVz3n7X4o5Mt9cEEboHJp
u5eVdpJwcmd53AP74XJXySA145ukXmrPRmuIi01DScjAsDbQTwdl6y31ZqRBg9X6
9c1BvCHAAmbRJFFtgoHxtBUUEkjKP2qdenZtFWmJWRHpl66+kqDKtZuJmkl0VORd
em41fMP2r1oCbEzZF53/ed0CuiIiWBwPInF9NXzzRyidpv4oaQpn8B+VuT5GizMw
O550H2u8IXu9Ih7+ihG+9IGN56P3Rr71CLRYxYvCgBXPdM6GW/XwBEitrLRtiNyt
zhGYQWE7fNG5Rj7ba5DudhiAD8JfUMNWDVN3U2H2N4oxO3ZK+0YQkzB1Z/+fNQc1
8ZPsk7Ho4FwHzaCwl7OFNjW1rjpK3OCv00+Y4jeOZ950l67HDiIeOaZE2Y88FbVM
LDQxm8JN86sfCtQ09x3haZTqLGAfkJ3Rp14V1lCEwbBshDa6cOJblLn8EZD3BBfF
sqNMLfQqza0lyIjlw+E6QXt+ANvhNnz5J3H2G4bixGTcaGATw9QjJ/P981At4ziq
rzR705jm0nAXZb3+nI7cLkoeNk/KzehAL6gPPr1VqdrnYiPM8HqYlyqizDDtoOIq
9EZG4QFJLlJq4CLAl0UvOqnweW5tLD/YX2BTXqXVyPRMfX/5KUygWJIqYIMUcXwZ
iYx1OH3yaSV/klvE3qJ3H1gIBTGRGQGYhpHmr+PSbbygcCuPbihj1mYk1r3k2lXf
khqNgqKSZmUdlWGWZo32G0fEv4P8MIEgJVKjnVt5hwM6dMBon4xRzxzNjJDqUngR
FKEZ8lliS/p7h68qICOvdGg43aHCFcqjH2mRJl9R6ulvPLepICRHgXrWgRTkhRO/
zQrojT2skfiH4m6dwHu/SMCGwMlMAAOCvGV+a7XrAJla6M3nFnLiHt5tVdgj/oPR
Ar6+YNCYWJQA7b4G6RT2/jPtujko1dnuoQWvw9MHZWv5FkxFn41wF295RNaGnZWS
oH4TqS6RlZ725tBKXydDcvEJUVqvNY7KQDgxpq4LpY/k2o4+Gd2EMvXkKVpOt1Om
D2ztW5bQOqWLVP4kZk2cpQ4KhfJBiLDImLFI16mEzEW+MeXhshPSUKaBi+WKII2c
7pcKRMuwnWjbp8HkCFgn7fnR/u4eBAP4kkv+8eJJeqas97NXoQot5vj5OvKyPwlx
9X+U9GbTJhULltZQTIlnjkUM3jXGTz79+SGYsrKqfdkf3uHQjPIfXdrR+LSejRmj
4TuLnRb4Es0MoNXJOWRjuymKyIv//IrXDtZbjXJcijThMo0gQish3slVK2ezL/lD
0A6yt0vdXtDfSU96MdzLvJWsC1teDtjcmNxa/t80WGHOj8cJNGuTRPr3zpuYkaAV
PF6TdYKrE9SWOF0iujEDSZ4eP1yrb7zBb4oS7eCtKb6GJA8qkO4VScU/GJT+jGkO
u2pvsJgqxJIwlAjVc/tAcPgS7M6umdFr+0bgLb8mNehZaIj04K6KKzW+1GQgQZ2I
j1s/U373V9Ptrj6DopGqpaZab/EZ13DYmhC1s6Dm11eyvK+Fj1RfNdaEJgAFunWW
3GusaI6yUhZpPW3VQ96aMRaEteFCqp8UA5P68KIPb7J8m305g/Y+Naf64xuVxgeU
RN0y75MjmmFcGo3l03YmP4kh2Bg23eHtOoQV3tNz4PWjzJLT7lGeGDXIDmi1j3ex
QYsyJjKbXpZ5Hw6Gn84ntVLd5FmAEr2NfD3+mthGH/gcjK4YZx9lrEUN38gGnFqv
jSTYuUa7+COFzewCZI3CPXUXuUS+kdezfMfm+2knRKD0mtTRXCLjuBfWWUPJ0N0Q
CjYDSYsSdJDC0n+fUhX4lSu4CkuoCYYFi0aM+qnHFXjoTPHXh+xhJ1oSxSu9jkBo
TfC423/VpBnef0sQ4h/GQ0rLVMfZb5DBX3BR3UueH7gtImV3LzhSlgGRuFTM++5M
ZmKOB3R6+0pWo3DTW5Pw63xlMihjhUU8q+jQg+vjt/xwwPH7ZqDk4eyMByawPnE/
3pdmGowgm1zS+BEHsJzXnCeUgASVgT4eSzc2N3JRGihQiNH8bGE05gLpAhNU5Cyk
l8rAUXhgQCf5SwfO8idvYa0rufMSnThgHswdXSmLSVGItD2EaagJuNeUOZgXLvNT
jaUdvdz5I8uYXXgB3nMbMb37IjIXDUDoUsqyqpI5xJe9t/bFMrwVFDyK0Nbxc6XS
B76XF9h8Nu4Y6a5E8/1aPA7zsASwGpOnw+fqcj3pINil2ORoekvaKpna/A7IbNPk
TKt/4aGwAfPTWafs29F5rWZIpsBVM+rc0zZi3/z6hLzx8CHJ49QiTG7bylH4peHp
pkRgkytXHLSUrE2FaGx5z/ktsALBgs1uzBjxTn1vKiwTTUhwvmuxSJTJJQ9SQjDZ
WterbFUZ58wBJpIKyQ0GJJlsQL8M44jvZ0PwFc4Ofw/HRW20h7qHN3gKrwIkIxz+
UlLYUBhuYFP8qe5DmrbADsKoGxjhR8XbDbQbDcrbMYXVS7fUkoFLtwdmw7bE3/eH
5zs3oIm804IBGWpSyd57IAFCF9XfVdJPF+C1tjKpbo329AgWizGc6oB5qGHXoMvG
pmfI11rXARpzWFDK2TqDBB2r7kW8LiHxRwojU0ehOQ/HxnY2fzQauL9MC7YNFez0
OAFFdOIOu1R8Y7q6XdCSR77nlZDsUwwdPHfX8XGng/lcLqn9FWzYt3uaqe5w66NF
yKzNIq69wKaBCSMVW+Pbb7V8NjwpeNmTDWq9AW5BiNzVJVOns9gO2hsO40/ESHJ2
PYVR2uHNC1lBcsL6FG34U0OdQUlj44C3nAe5QSPNsOGppnoy4OvHgyvooS9cNT9X
t0daa3q6Fmd58JQSNDTiVUDni8NxxE1Nim0azkx29hXOiHDXPXZTgjc7l2/dwczs
iBnX1whqys4MUs1vPweQM83WNGKwTp3UoMWb1Wdao+eRzDGlDf4vz3NuP/43XIxj
Sb0MIIRGBqNyCMWuVavjvXVU/h78TS8psQLFpU+OkX1OGd+BCuBqssQTenxjdjgk
jN95PaiyJMqG29SOf6LODBUjp7CYN5jeqLLLkbtJdtBSAt19UIGrcKtYsidQ4gQK
32+mavO3+vu3mEuUtVKP414afUadb9kq+2dorzVLDqOcwZgBnPMiuIQeSwncP2pK
VXHLmuD2aYFWse/KSM0du9QDEhsOvnTiAKGj3mO5/7w+lSXjfyt0YWFHJyJf4xSo
nzFuRSnVSqxqLWcpu8kTPKp0qG1lp4/ECyV/ZIe6uu83lP9dMNwfeq1FSHvHzfpR
CrqjbZD2TgeOHBShRxPCtkj0TcShnfNB3IFWu60lwTPs3O12LMyKJtpp0i2s1KdV
aW3IxowJQWXu5lAgpxDZMBVIcLCmRG/5r8LZBoNQFo439cMzbjuQp5EXe8zQa8rp
QrSiBxpSeZo02zJc0RNkgLRzgBcsKoGgHUwfckdgXnSAXl/pi5P3RWgO6YxOJgFK
tFCJjoq9vEMtAVSJiauTS0u+DpeazB0WtZ37qmFzCALCqpvY0aa1vQtm83s9DlP/
KDVkKx7NhiSSqAaMNetIfJjaQLzUJ+Anei+ExR7tVYtfTAsyjP3nK1EXL80XM3y4
SsX/j8tJrpkwTVjYkohM1cexyrY4SL3Mg5686UkR+JvhVape4qrz8HiSsrjzaoIy
Wwui/2l9Ghgy0z23nhxyLJ0ozXRkl+lpVrU4c3tb3tlt+XzNNgnhnlhkH15Z4rhN
Ql7app8sHSFWEH4LI8JMBBQZMfL+MhfaRympwbXWE8UIB4BSvlIT2V4lRUAIVHMv
UV6HQVa5d9NV7RN+e77XD9WDKtZuvRjmKv1lt/q8MGNPsN5Vqtbnvxo4mNUlz0ta
AmvfGH8MCjvOEqdkvoxrTAb7fJ2CD/WGCYM+5ZE94giOAWdY3OtxM/hAXwwP7yBn
NxFk5ILpt37XHGfaI5Z5vcv9/7U++pfIRtPD28jLyLhzucITVa31RRj9sAWkrG4C
r6qxuj/10BR/++kO82AxDCBx5thPbsdmxpg0o6ZFIF62cj6hfNg9dTFrykTHDHTH
UhT0R6xcJnrBIaoakDKKs38Ooi0gpQE9Y869ajW/duCXuMO37Zxah6AOcQedz4Qi
8Ut/+eGmpnc/uJnNzBZ7GOa/KeFP14dOfplpxgUfAwx1Cut1jjYHq27uslzCCVsX
Gn3AEHTPgXEEcuc5oc14vvolZE2Mfc+fLhmFBgh1VsrO96OqrvtetCGnx+l/AMcj
tXqKAHuN1YzrMXVpRjqCfnfDHYruszqS/9sIYs8vsHoiSVz4pE5o2SIL5caEHncc
njp9PvzfmI7CujWNaDnWvQcGRmvW02PXe14aJ1qRCbQ6BIIQm40dAh1fvXsRlSVk
zuYmKzGzKRS/0sMAt1fIxUAMvD49wNFrPFf4z2Z6rcuF1KiM4wDQY+AHYlZm+z29
LsP0+h6c08uzAz8ArA7bcJRoaE6HXqtsdSoBFnbx72GwvrFsDuvsPTc86xfTdiTi
V4hq4yAA2Almp5txoWNqg07X0eDe9QGppdk48uaBCtRuYljQxeCFjdvQrMFDCprr
3m4VnE9bhONfk50fqimoOU5aldPUnVg/BtjW2EpGpNNjkKM1/wF+i7FzQzorAkjW
XYXPN2X6oOSWxvz7CFS6jnDtCGBai+932hC+gJwkC6SmVHkgogAuhQZlZKaW74vU
5zziHOliAt+ZvGUO2W7p05iNlwjmW2LLhl1VyKAuBJ5E8B4ZuDMqnJtxBaNj0XoH
fSDPZPlsRRMR2ClRV7s4oUaKzp0l1nNTuGIeEroibieRoJpr0NkFGktSu2R4d4vc
FeF4VdXU2KlTxt3g8GuOElHrca7ncmXoNfVb61+kD4EqajxB+iZmGdFffTBmY7io
/ysJ+T7XUqGdansrXH9KCSBmrk2vjGQEYq/JtL0OzNU9qonmSebmHVi7sy9fRS+I
SeiH61YDHsXH6C0/0eadyRB5yU3jfhJzxuU7RoOYGiIEdUz3EOflO5+jbgEl+zMw
2ftTEYju52FRZrv6VHf4vCqkIfTImZQFOMDFpJFG4ZEyWU6faT8mGrGZ42OTMa8Y
VhUqgp8k5gl9tb5Ex5OKeK3c8uugxoeGsjgqH+kRHqap2YecxtWvw7NHhjblLJ8F
VBbES+O6q4QhG+E0/QrygT3iCDSoZ3NZV6BXUDqHM9mfS2tik7EKMetyRWzDcDeo
5vCs8jQeCKfl8afwiDlPZqmRgK6981LlHVjDK9rKcG+l0Ft+4Yx+B6xZRzhCwTkw
YusU+wXdsh8IzPOUI2bMFuxo+fv9C7qd5N9WEXp/b/mIgZ051ZbPD8lBsHqI3/bg
VGJ+FA68Sn+coJdoOn4GJy9gSFWfwImD6C+zqGSG2DbnMuB87nxY3gRF284oOq9M
8GbHBpePRiiXkGdar7FZB4spjXkzPxq30OHpdmjUyiuLxRI3X/x9XABnPfimVPVB
DR/+QhT7JB3DVG5q9OUMiW+L6HBiRbV+8ChsIWdP+8scDQ7SQ5G3BhX+V0qvnCA6
zmlHD74z5nT5lmHT2CNS04aNodxPyXUORyIekF5QrFUt2sjtJPvwzm0Qtf04msm/
V0YCVJE6eu3L/PC2fodHRCjnMO5OMUGFw7CffRDzaWavgQfAribhnHH8Xdy/ASeM
IRyxnexlkipycsA2l3FK5WegIL8d78KirZUdgCFJICTfR7MrR2LpdkE/M8/2F02u
j1SP14ej+5QI5cUpOazykpskB1EB4NC+RmNS95txL1xz1ihFCz+1PcNzmMobKKGf
jPQEsi2iNtCayt/3DaldhasAgElaKq2nHLnLGW6Hxex9nelOQT99vmYZ3DSWBY/w
YPH+/UJ47jcpr04NdwCJPt0qE86iwYtUMKmuxWR0FxXmbWxaqIu3Wz6RWMUjGv1Y
dybSpqmIYGr/jIcCmB8KFnkzaQAr7TxNUYpsZ0gKuKF24SF20xJL1lr+M1nq1ttN
UVFBt0gr+WaqMAE02Ft2/bKnGkaMRT+tasUsHE83XPzEut+0ZYmRhaTArdbHp02D
ALxJfJRgXROtQepmO5eCnpIWhqIyKnr+qARChTQRUgzyf7/JjhhOyA8igBHEkRVz
Kf7iDA1XAXP6+KulCdD5k0FQrQ4e6siBiTUbOMSGOW5ctxgqxQuX1CU5qNXDLTpn
RMLjkLA5afCIfJOUpgI8G8BN3v2y9b9x24otO1wCEu7zYKAGe1TWefBwBpXONBg1
DUIbpAeTygUkNOA0+bONffRGfXJAg3CRZ2MMVIB5wvd18lDUOLOVKZTSuk2fh53Z
73IWvrbH9I1VLOLwmJ+Nbdjuhky1DjzU1aQif7XFq4GT9idm1FyopBl1K0Pyu8xg
GmXCiVnljxxmPPFKRQCbHjA6iubbf28MWcyyVaxtWZ2QcgflR2j4t7AxW6hoXvWv
3tNazlb9js47j7dIEYg4/nypTfyBWYeV8tUg7dDe5q8pmbCBFIGMGyyq9vX7Lnkh
VpzvVjazGB0ZNdULLqhaC3JF9o99cGOQ6xAqlYPugenBA9buqMtMKbg04TiKvrBB
55PA+o7r7MWwmtulDs4T2kHET9vOMq5BL1BnE4URyU8cHgDsPr9bWUBxq8Q7jmN0
2kD68+Ks13PsUa1wG+ztspSkM8Z8XRDNcT0elsMQOXvK/5eq/Iq1WgdchZsSr5Su
DsEX01ZdJgwgpAFTSxkBrxJkfxvcYAGO4UARqAvSEFeSy0ySe4cMgDzPBe8MvD+n
u5WoTwPaL3DFaGSxSvHu3QLlGV0supfai01UJWD4dQwKCM3MZM7vb26s0Dkucvqh
QKvO6TVxBAs3ENgzQE3hACy1ayKcfnxxnOfjGlsb4/5xSP8DR4ZcVsDFm0LXOyB/
JjXEB2rhix9ut+218zauEY9V2nec4Tyn25oTOuOTZZARNPrFcc1oadLRWuLYmfWj
L/9eIw/7k9cgZ/Uym/IlXEgh0hc+viBwcT98SpcZI+MmkLlowN0rQzoBwJer5i9C
k/MP+v0AZSDTfAUdViOHOLYaWJTYztcETg4k35vj/a3FILjOBfE4/abJ+dO/4BrL
F7fjwa0WX0VZJGsbBwT8Sczl1MVVA5Pr7ZkAbhsPWPaHuRCx72+9KUA+yLcMzZWi
eki+Kw7qp+r8KLhspGNo4Y/GfEoj8Agv6qsjjMAQTtZCZ8wQOCrUqTWPHeDsj1B4
5NIXJTimKCCkvjlhP3EyPZ4WlP1emFcOVdQhsxYsDi6cxHK9816TzNrWZvJvwbqL
ZsxxTPmtJD31dC+mpx47myVrDVeCtrmXbm5euFGT/Lt4nxcbK7r6ts1dT6J6Onpm
ttQm/QHIzXjIcdlrcAb/AoBeaREhg2l17QA6pVo35n3nFno10ZvlYoIkg3yB02jD
M92ZwiCWbtf6AMLkKSd0UvdQcjUND5BK8m/rGY91fke375CVSGuQaiI1MskuhLUd
oWOjwjZc5U0nd7tceu61V9pNsRpcwCzASVTCT4AuvrUCxa8KRoWrfLNrkHea+xgq
YbvsMYV4IqM7t8FsXGVBU6EG2WuD0t9b1+IpyZJEcIb1HT3pzqv9OquTZVI6RChk
k6RV77iKgwWmJzsLnNHqWkm/vMylfeXXg13bVmlORqlxzbSAuJbjgnzwD7MU97qk
gfM1w2sqdkTrB6BL0pN0tJMQ6gYkQeUmkel+lhLLhpqgf/twyQV6H4EUTQJXKQ7S
4NGMX6n+aaAuKsZZVwqI/4VX700IDMboYmpw8cNeMTP2CfgjxKGkm7dHbPn9EpuN
jwXPlcIYrVQiL4vKYO7ztJrLnLhsgYwm72tOXDRkasPkAvpvXXI7dD7dnOu2LPER
XjQ52zc+U9y2GPgQb+O53iE1JZR3FxE3dpud3qOG1dBZpqqrYtJfgTvMQTQkBZXJ
0c8yeqmIYCI+zi9qWSJ7bh2xPON9vabU9JT5VWH8jYPyL6WylqDE/B64OPldZ9Jx
RE/H0oWeqqF3H7MYfCT+AgiE6milZoY3a8Nl2LfcFI0gzi8snvryIha5cTPmDC/S
d3HhQepyN8EYrkcWS92jWFdqmzrHg+U4BcugHnmRENtLfsq/omo/zceSlQmRC0jH
RMLTF7OShgavfnxiMc7aqa1PHTGBSDfq51bQtgVE600htds8Fml7IA2a5nKew+gT
LRGHGGsYK2G1N2Te75pwb/dmSum1Ljw0yE/lDQoSp1q07gqRCfDU22wLk+wyxq/j
tBPIWQ1oq/iKMUykHjCoDGFfo2y2GKrq3oI3k2mxPVzXDXviCzwUBM2TZnKGgaTM
SmYvPN+DFGnA7qC5U05HYlmbqfunjdCF3ohGfr7s0FOZhh+s+hvRTCDsnCKv5ER5
/xd5v3V94Ah1xLIcPpTaqUJd4gw5HwIGXbfgMrIoTby8e4nM+4iheTjA4ZT9HimJ
fDYSPk1CUz17iT628wexauFlUzC3+689QjqBSfi9C9vFl0lmPpMg3JHph77ogMp0
Ov6ku8xmGddkUw6TUFn+GKfqlJjH7HDM6dlzDC4JKaGvvcZ03Fbu8sd62FUJ6uiK
p4SfHIV94l80ycFX89h15QFon6Mok7/1Qk7LDtD+JUdSc70gdoojlbMWRk4nM8it
vGQb2zLJczLFSALAPDYbyd6/GIDeKRAFYGd1e+AV9L8bca0hkB4mJCWID+nIoUWW
72z8jobrOWDm8fv+i63lHqJYT9P6Re47GTKcyBJoDE8PlHV6C6KMVbLfg7DmH9VV
z9WXpAksFx7vsYKLFkxKnKZ2+GuSSGL0mNXax505JHJ6SqKkAqsjVCyB5oAfMPkv
dS1ENpiqBMxK/EynOujEtS2nChJD9yRwCsRLlkO9aZFB6ql0dEwZatLfctOr4c+1
HA9KMMC6AWdFNiSADhGhi/3afBGHuTakQZQ3+mZHQsZ0C+B15UZgleY2vdhoipg8
MPJDTbVVBBsWlcf2ejv2jS/DvQPv2lLgBuP9xSTYwf2/UG1M29yFsHmjMsiCYLQY
gj7mNvet8+6QC/GHO/Kld/59Cdb9rBGK1Y8TdDnvsI9ZU812LBKKZxTGBWW3BpXZ
pJ7yE03vWlQvoo4or66h3zMnBqYsX9LNuKcfMZCgwA/TrEO/zq/wR7ID880KWzuK
ubnQbBl04masXao4zUDfVhp6/AzBLSCKcTvXh4dArsBZYwptLnBy8XikNzFO6BFs
HEhEMTqcu3TLPzFubMkfJMajNj0ytqrwpF6F3keEE2CLM8P6RVLoqDANUl8D1WIO
46WsW8pra4BQ93mbpE9inPgkZ/T9FL+lmMRcn3tR5qhXFk+Hgt9FEFMUE85weG/k
1RxJoHLqOuSvEVN+ohDOJ2RLD+jXnFbPfBMwUZKBH9EFko2rMxcPEm07gAjGKtrd
ZbNLjQUF262VmOPd6haCk5SDxWPUaU7Q/SnahAt1yOk2Ljk/GKG0oYeeV5cnLjdD
gjfcCoTh6P3/Gd2YE3YFANQTJ4Yunxoln7Ccm6pE7lvaLZSqmj4WHgE5vqwI7LTu
lDMiptkdu28y08pX1caIpETuTf+9G71pWj0ipJ3TWSSrUXP78+7+//GKtFpogP/D
lZpcf1qgYuHGKvOQL2zRT0n+YYCG+4CqsIPlUzFZGglV7zoKJJL/p0rodHfPB6Iq
Mg0P0nRz3IJgLh/GFF3KOPUJ/Nhqbubuf8FQUwxh8P+F4qGcSkfm3RRQa15UKalf
dgS2KE9Bd9ftCr+F5ysk1ZwvketWjn18FnbUPiJ6xZlwoLZZxZFaqAQidDX4180t
1pxyXrzHSJWNIVngtZrwP+b2C6MGMmqn5fhqMOWb2nj1lTDiv08rza7Rn3PoYVW9
0I/d+tYzrWEhGItUbJ0bnqnpWGBG/pbeW427jv8ewcqQVLUKg0pfzOgA0K4/SlCY
PPGhf+sDtxGJsG3K/cEKR3Ns4bSQjlqnTjmUGp4mLgA5iAR8iBLIuh9nynEkvC1+
gWSBMuifhg0CB5QSlXQJJyrNdLMtzWCXc0ZCajt4BfUV9BFIejaiW5y1MbzieXA5
J2v6G6dJK25pO7EFIN3TOZpl0NQfyG1vYeiw0LqwQsCcmTOVshBW2j+bzPxbahJh
PmwH+sqrFWC6jty0AhUSUzyuaLpLLTDsJ1fbqNMhvbFECVfQHaSV7sYr+IVU8g7U
zo1WAGaerqe/NBZFYwru+49dnOsLH/lvzzMkfrfHKqNTW3n3D1UkDJAUXvKqUyOz
bAsZxc80oNg/DSsq5XNPhL7ELwtlhKoQMe6A39lmBmpGTtVOQohdZflvi39fvvla
w+d5MOuqTGSCYD8s5N/VQ17CkwHiV9j4S/VuSS+qemvQLzN3Usa/qcJgXhZIIZ2Z
zK1cnNfAs8GDkAc4j2Qozbav+WrccjLRyufEADmOhhR//qrsExP46/oW70tE/HVo
18Cey5gRWP+qKnxeI+xi3Xjra2rG5IVqxFrEROucpecGS8nPNp9b6aYU2cS5sHdH
rClcIj91CPUM2W0D3u/LwgxJ+bUKojqLeDJoqd9asqHwJvIvVZ7oMnJO/ZDclpHy
xF+jzMhilzCohUBo0IVNVRArko1WUJftx1bqIZF6hnD72TWOlMX2VR3RyknMtZ/e
OiURRENFhupkZ7JBDh62i8Xw4TCizhatjkuTPNpRWZftdUd1PN/12km0PIHfAGTY
FE+nNwLO1m8L1rC3M3hqE28uCeo96YWF3naPwUel2mpUXS7domDLW2BX70xlK65V
kExECFVs+CDPkomAYGOuoZL+Qiuhn1MyHHpo1P1hT/+hnlDc6Gm+UeJwIuS9z/N8
EsJup9QbrhmxUVCf6XF/UjOzt7K8FA/NASNpdErljAVZt518wF0nDigPesoDxWFi
zNfQdi1fOGYQMyavir4i75PosXXDlh/dEsjqDxm94Eq1zU1rYeTrjqoXAD+na8Uc
68owc5E72kQqasUGxHmGN47yCEX3o3oC/BoBvIpEqRoPJ53eTD6mOlQl55NP3pN0
ty/GC7/wdPSBaQRG2HoW63OIK4WBhU4PsCNstzDtwrMyp85Uv+IgbpT9gyJbRWdz
X+QTTZT0rYQJJBR3K8Ez+JWP9HfgQMKKFJnxckKxZfCXVhi2QsEh04wZGSVZQtZT
n3z5JYvuttunPDACkfMPmnoJMYrs/PsoW5Qsv6dtav3aMjplzgNO9q+dNrFpudlU
ho6/xjIuL4zueUcpopZjcVPVqUhPBILSj540getBwYQzyfKilUXBujc9KWLz40et
jG6+JXjpI42E1iPr133/hsKnYYeVChpmjrLTE8kkAD8snWKdrQxitt7r8pOfbQx8
Tfbc5KN2AAiVQysTxxfE10A/8mLEGSSmd1H5I0caaCg+xYPQNDyCoWwRnTVr5she
cSQRdIJCNiy+zOtSskhTDu+kMPar3T/Ckn7yfMBQrh1qodfFsjFqwBcY4O93nXsk
epXhbOFJt+E3xhLvw2JCZQ7JwKX/3anSMSGhgq30L6yKQDhPufPm/pe7vMp9Whd4
qJqaMIT5HvBK29WE0pRGvOBWsRBobB/xmhdPreh1H1kfW5o8FqlE8Xd3kKENcNy3
ijkKJC2+Y4F0r3VsqqBl+lnjvM8aAw60gVy/NlWoJ8ry5Ax3USj2Gr3f/yNqbA+K
zn1OoKPfjYYXOJKCTyDU2acgHci09mQjM2X0vupmpp99pNNLkJHZuQFaipUmz0Ku
G5Ut3K8/EOqyyFc9Sjmim16Rl/cWZXgk/yaq8uotdoM1plL//Tt2gyo5+lRvm1Su
Pc59vUPNW1N6XId8+ebtZxEp8Qx6av8QIiC/liyFAG9IKW+DsPJpEQhQwyCZWB2g
XgznmGc3+CyHrIKcTMkavTPU5lDwDs2J6wIFWLtR+YIuyEL0b17ydgBiANJbKW0k
AzwKTFABWuTU6b7+uu47y79YHuOZmn5wpUIWrw6y7a4wIb4erG8sx1xXN7fjPd+7
s0yFeSwvyxbv7PC4YMR54YXnMmVrcFRZX5h9060g9g0o35bm2sifvWzlXZHGD5C+
FIwAXRklx94Bw++vrSfmuezCIeO5BNFyaLEwr0TDaKUduM3QZo8mWQXQ33i1jBuB
Bj4UDKX5/+p2Z7g36haYTfa/uf1CnJBEhxFYyp7ZJhZfD72YdHZAHaGTA+06BzYK
Ar1skXgvA9flDh7kudvxBo3yJDAdP0CbtnzGXp2xS6saYXR2Dm/bRfYFyX8LcDz7
HZRhpGj33MjK5lVtoSxfSlhjJHcZeah8C0zzBLWpNclsG5398j4rx23TbWsOCyV1
1hYp0QDuwnfYq1TyW82jp+HPEooO/Y25Prm1KS9hy89+S845jM44XZVrpdywFrrd
CB91VbOYoTar/V4x/ghE9zEYF4qmL2rh0MYDJrjBoPBmufXzpQA+g4UfYsNMzppH
GljzxO0HW8cvxHaXceixWVEz4OENjGAylH5Cg5nPps+oLOma+FJTlKFpBP7klTE5
mKbyzSjymdFoAJn8sqYbA+ub1oX9g6NaInTF7R11acq3lxajx9351wpiRlfGWLFd
v1PL1FlymGP3xj+HHYg1Bz8kUeE9As5aZu6/bTwCwwT8i23P65wAOD2uWo5jThc4
N1RgNsM8b+4IeMw8VQvgtSMmB1xTzwOHNv4ajxlerLWWBGqAPUlFoBJp9gCexJaL
NscgCWNlQGbZDLpnWvCsi7JXL6QulkY93gyhbsGf/qMSrBgrk5W69M+wKysoAJwA
EESugQdF9srJbhtgy8U0oulrgE6qIV4qsFqwGC63vONQJzDpinSqnF7rWUwQlZSx
KzjIYl9ZBHGRXMzd1NWufEAuuN0Hh6qCE9EBMU9tKIbxNQ1XZPTWopVO7P4/Meyg
PQNHXN/GEsEsYEzSXal4ZYoytk6W/ML1vqV4BKJ4RxetUHkuaqUwqGCax7h55nr8
s/m7CkB7tLK5bBXnhx8/f5bzfHomk0wws5riMnIX02Jkih48lUxVF59fOUtye/o1
vENespBIzJZBLJa4M7lwzrwmSZ1oJwD4+4xK9nnaHn6QV3AfcPK9VGsPPwsLvT/B
OcMWWDj9FqV2XP+YsLV3NOmfVpu1WmlCw6x6T/KOFfUs9fTbyzLsC/MCB6qcjr92
/nfWtqqPnhBO9ax+hiSX24qKWmCfSgWYz6lcSRYLECCJhJxjd0K/ly9EFWTW86Sz
zPcfAeNrUGV6j7HQIxwN6jKkrfit3e9nB08I5ws8KUbc7j4BNTMtPgn4AKfaMHR+
3MjI6wChBt4+n1HBgGuN5x+ZQ+ZPbILTqj1u7GgbrLoLfCGQUE1b9mtS/hEtlvcn
iHO/1wvgqYsecNiOx2jZ+rGx/IxpQI1BjmOrCvzvwSLaORGgWkHI557kfZENB1FB
DeZYGv6qKjXkxxRG2CLhvNAClnXuc3jD6SZxot3UO04wELI+iE30l7g4YFQfpvI7
xot/YIkPU9dhax1JaKCNR6qsCOyISEi3TGr5+iq7Hj/7wW5G46Cj6zqLMn7Npbh/
x36kKoNERMzBB3l5vUkKHcFeGhE+A33VSBBxjdHc6NJUy0QrAoYp94FZvKVTX3/i
4r8JxoGtrtwMqJtHQca3sVjbkgbkBnpMPANI4ehP73EfJePi/ZfsRhSXKwBdX30N
Rf7sAPljQL7XBlDWRLRwB7I7MfmNCsDMZk620BoK8eTKDwRkpWi8/JS5YmOTfm+v
oO1aulVPc9v09Lywy0QQQzfn7T72O3kPsqkRwc3RnQEbpjDAvjAqR2SHiwyFYsLk
zj/XKmnpWJL+kx3JQJbK0BQZpMjggPUW6p80Ap82J+GQvsUgWckOkVWzMbhUpIXC
FI09UO4do6z++GWlfa1jxzeypWedWjNHFYY3asS7T4Dkt9dpdTKE3k1ObqktiiPp
veIJV7vHOoDVv3RTUfI2SdKZThqsDR24lNMbRFs+GUpLMgqBLn0wKfyRVARglHaw
/baSziKLiLnLLG8sD4O+NYvhak+Fz6PZZj7/fHtaJbwR+QV0hPA2ClleicNHDKMH
lpdVGWxgxQ1ll6aA/c49FgSDXgiTt6Ismgk/uGFFabSILAhZBlI9guMwtOgRgryP
dXMnhMgRlSeg1ah3oLsu+QGQ13nMgiGbOKsmfvdigvA+DrHnFnR0AS+y5Stm2dDX
Xzy8KbX4rz3Ik5VB8Qsete8dfFMHqmK2PVTYNB1RTCfIk+Zk4ihCf9KGAk0l+PuT
hpQpV/E4Ki91ShcWe1jK83FNNJtEvE14y5FXOVce/ahjojmG8tK1dHoEoTno1ctN
zwyHC9ckP1YcI5p+NskUCsHBQajaXqUTyCqx1wonViwL/KnXfr3QvULdr4FFtgBd
tJOd4OuVRNprX0VS/Vrglq1AkmKKBgh9fIqg/47VgF/gDyNayjajq+2MC/j268Uo
PHTM4LB6Dh+h3odAAwSThgmRzUU5nwcsggdcRgFs/zGZgjeqj4w09HHYw9hy+P27
PTQPzT+Nx55jyEmtv7Q6wJL/x5CP1X0AfIWfQkoRonSDYe+E0KU4lswssjXOJc77
51GAf+tj4JYsIwU2DRirONsa1wh6AuP6NNkx3VcdhAPU+um7+jQGIjso2PKKG1H5
uNqDIZtIggfHu78X4ubfWJMtwl8ny6Nk8ordIrYBac3Sg2Ppx9TizYGsXJXfdFoa
SM4TVS/s4NCD8jvy8C8nYjB8h+F0Eir9lpcyjUj5cvJA+yd5bqlGiDn1Cmdifart
WUnNaurugIQY/5rwdQ/brLkDwFun5NTXiyY1cxxg5EnHPui7J2yNO4c5jMdCVFPw
5qeSGd/cF80l+g5nGDqWEshYRACylHHZMcAYQnVSiQdhCXhEIoVF5BSJhcbw3MHD
K3T0qH4W9N9sqp8g51Cj65j4FQOz1f1DJSb/8ftGpZdNAg1F64l9+BCNh5E2GX4M
s4ZkaZL5f59R4W9XicVlyQ/PQ94KOXxccx6PuEz2Xdl2JdLiEY87jAR61J8tYRAl
v65GMb27CSyDgyvJ8StEwcT94Vtyo9QeJwIHd3frqbInywNJ+2Z/XnGuN+5Fkhuc
HcfkxBviqCGC2ObFN/YZ+aUF+o1n42z/1rQRC8G9T7OehMzLw2dSQo1MUt0RrsUw
tnRakTH0P1ARZRgH5sQqhJKc1xZf9j5gn5yGYimpil0I24k+9+znVv1PwNVDcZSR
ol+A1JAN0FarwezS2GeBwTLobhqk3MT/kbaYUfd96bcLQMSyFAk8+hGTnpZTP6I5
Bz41vQNO8OhetZ/fYq5L2A5qmnaQiSIiJjcKb04/+V6JV9QmgfDR/4i9pSBMHN9Z
TkV56i3xLsgYk9WFXROOKT8DauDwTLOhATnmEWUkeYsZViCyCySq7SdVgLLx8lCR
Id9WEvlx2ubNVtLxf/jfgjugRE/vZc52Z7DKQT1ihN64V//jMEH3ExmoAh9AhrKs
G8jJSrZ2tzT9fmsNcHi8l7p5HohHpfwTu6RN0D0cs7oIUz7ic3i0vfl1RoZOQoAu
BlljeJvnZQiZu94qPlJAKDqjsBRIjnaPP4KqLDewa7oGpdyOT9NxkVYf36ITnDi8
6MGuxBpSrgDn1G+5AN+JU6zNyrdLppe8nbcsmDAqb2A8YkUrdz9pC58YiuGD1Jby
dpchWHosviz8XDh7RXznIUOs95B/qg8lxhycCLu6m4D76goxWECsq0ME7CTkACtw
PRYggDzxO4lFOnl9pHiQ8R858nbXyKYIGxPMLXe+2eNcPGM2NUhQ6GyXi7gQXP/d
GiqMLjThAaJhedIEi3R0ZwJ+Jq7PU78I5MH1Vs4xXt3W9Zs3L35gvF8+c9gePEMz
I+5UYShfsprY78ubvtzHSFSQygWcFejr4OE45gw4akwTejBwtzT+hnRhv2hT9xPy
58t7L+fc8ykO1FswLh6Ufq3UYVzeJP5+M2OZiXPmWyHPhlPeNOy70wDKzKUsUHqZ
Zi4rFa7r8WUTyLHeZMa4vxTJ76NzdHIWWgKsxsdhT0P0pxGjJfnYxYCMiYMCrQRO
RGlJU3c/oDPSqb/2yKZHadtLZbaLGiEIFLdG+pHSGNwCdw2yy6wyps4fY4wb31eF
mv3VeEZSAaar/AeV3z5tH7L5fzIv9QKEJY5hgCtKUSOVRitT1Ss+0ugkaNopRQkp
DH0KsaCwoBv9rdDqORkFN4XRHVr/D0TZKi5y5S+l9+hF8pbplAqiSdApm0zU8YqK
+xIZT+4o7S6DMwAJpAAt6GylXggRowkFKIn+jFgVbf+iR0diWD1NQNSGuDAlV2wO
Ngs6yUcvLiL5vRilxwutKsQHFp/dKexKcGqUKjVi0y2A/E9cbRX+ncFA3HbIo5M2
JClUkozydFRnxIu7uMI/ege8Z1mciX6I8GrciEh8o4aOvHjlDDYrSpyxPPd9/D31
M4ddwAdWfONlF8yln67MMXvNzscOSgQvmXU2aQ3VKfsMJNOQN0H74AroiQNJiKLa
TsYXlIJgTgcN4nuqp7lALeLEbqlG1umew1KZsmIyh1h7YDi547GHxftDdBP+OOLi
yvjhhB1FDgRMBUybk/dPklTQugG/c/vbY0HPdsgWaJNhFMHtqrACfWbmHiq3spnQ
zz+tU6/uwZarrF/VSCaF4TGcHaHv7Oe+bJqt2LYg5O7r0VSPFW50B4TL6i5bee55
YfTQMBZmatBzqY1ZsjuJKteSMwYTjuFQVcPmtmV037NZFuAcvl5k6IiUW/1BdS40
9oKl5pKm3zE1S8gUd6t5TBu0kixCvHoWJtRioF4YKNePJGfqMVwxnzlEIySHMsNK
zdCXMUHkHEhAYQahDJLrW2mGuiYDfdZZaLlcbiBe3NruCItCP2XblOzZ5KDWX97o
HdnUwI5vSMo95f23VtFqEJf8+mpRgbJWEKpt9mm8fv0glM0vyXaB+y5s8sI4RBWq
c0NQ9o4wJpDPwWl0Uff6gL8+OY3iUVJmjlcwIXG5V4JWFFC5d2gMhUb9ocqaPiA2
SAnakoKk87/8zyISHukm2oOoVj3gNGsXgZk60XOkuBCuvxV8JcUs88xRR7o/revq
XkbdNRQ5ZXEk3nJ1TppEvMPOnCIxyAoRFw2JSYfPWLv5krRj+nb8YhhZUT+KSzoB
2BNvoxa0We5AR+x12FubxJkOlpqI+SZAm48sW/jkf7Suj5ojYzXoZe7v4KxDSoBV
4Fm5yP+VeNFGljO2a4FrWf1LwytU0VvxZEnQ2G5XjUnJhPtuBYGGNMW9oQO95kHC
BYbp3FvpxLV2SS7QOiOgU+5sUFROaLDdcBT3vq7mRCDyQ+eVNHAW4+UYmTYFFneY
bVyiiyywBiwmiM4LFSCYGXxcFikm8norj7kpaRxFQlY5cra/eQlsxx1CSEuvPgYP
qqoDJr20+pGDRDTWQESUBC+CCn4RH+kZEPhyy09CpcZqNJTtd33Z8y59BR06gBSg
ZPPBsndFbhVd+CYYP+MFnhpY/0S5AeyH/1xwUyc1/Lg7k7sJyUMPZuzqHvD/ABaY
LKL7ACWOXdB8oUi++TA6oxk6zmaVTqpv0QmdaAhNNGNsH2JX/7QzJa9Xgzj3RE3u
E0CBPiTvUYl0fgaI5KR59BtmQQZKrIM00nKD3KNXcaJN44wfWILG30lTMJFDv7N9
mx+JF+91P/5IUKGjADir4oPTPsD0F51DhcK644n6wEGFBeQwKdiTMLQtd9Qh3p75
bRUGldzadL5RxGytfJes/iUUBkZsoPMxC5phQpf+a5InqNyc0Dt5bx5Pzhjtm+9Q
7fqRvRapjPHJcu2+gCSI85q1/4YcXR6UONVsFTZ1FbIzvJeTWEcTD0QQ9m2NQbP7
OayvHiGi7/V3Loig7S3yHqo7mNQyCvwSo0hFRgdFy6Es3KKA3oGB56HuHq8ynB6y
9nEoU3qxFJ3nNLGnipfuz/P4Z3Ad2hmWBFblar3S0erjeO0Y1OSNGfnpwWxMkOxx
+/8nrU50Wc7vSrKy6RXvIx4XeHxEZ6Pe1nRXqYhHvsuy+dSrLNejQ8HsQAg9ksVf
95/LsYOJHVmIyiAdTzB00IpknlIzr6jLztIsvkVDU8AVrcNFvBVcLQjMxTxoZzyg
Nnfx8xBgwlkGoaL/2JTmOiXD0Je/nAnYKmKZFmNw17tUQzuirqBCeZqpzmneKWCu
HTVQysCjhuACw2q7Y2z2NViwE/iMnEzv5wvKhGadsvsdWrPnvVR4NFK40ZFGt5A/
vvKQtjLOPLg4qnPIe7YUQg6xU68YvO8FFzsGRXkhjwjZLEYfHpaTHBFf6Qd49R5a
+1ohRyB78RobddVGNDNw/XZtkShIk/uK7Lp2GOJtfQWVmN+1TBvxzRqO7O7+tbNz
UaMUsA3jkrTfvo5ns9OcgA5kszLbGWnIzMgY9T2kd89ReRwM7tzY7ZaPwjok7wD9
6bZP4a+rWKqzP4h59tjBp3GSSD24tViywRBB/lJScB6TowM1TB+Cc/MEjyfsl8t7
kH1qjJwFUTYYv51Du3WXwQWXK7MovgzulPEaEsIxLPXdp0s5ELasQKof0k48FGqJ
qkYvZf4lWgOpvcVH9kKOQOPm+8065kUEgeKcECOmd7/WUVXzPL8/NRP8oyHLmQ91
nIYgl8MOLZrUQUelKDhgmZ++DxEJY2iAE4AV/ReCMm6BxFHTYprSKlmOMxtK7k+g
L4FX0Cpn0O0IYMtt66nkmzDsyJKMeb+oVxYPgO0r5BZwTQupz+u30B2BxGFGIx0Q
jCqjOjxcHEsj7pUK+n8uEqNyGqrMdCjbCIEY54ht8sNcKV55B8qx9JSq9PXoKiib
YbSnbMKMZ3Jm7YONe/LUXu4s3L8AmTPfvldB/dyTuEq4UJXFOybYMCrO6+sXm8UQ
E8OcLX991Y2IKWuErHd6mxiwtEuPYB2EJw2EGwafSdSRkpxv0sxrMm/Gee4Rozgc
MZV7r3OkJfo97e9XtsduzjtvzcgXuuPaaP8tmgFkZNfI4UKGze5QrTwU5x4fYmrR
FiBe25is8unp6Th59RGfFvJ8YzwJSDf4vl8D5hgt8KqOra+hlM/kpqGzEfInlcM+
VG1J6Ky9RZG5kogNpZPva+bNV688VuJqrpMEuO+VpsWc+RGcDcdWbl2pajuKTicw
uzaRpLUtopMMzUhr8oG7jq+SxO1xZ2UmFwFO311tcMNyFIKiPaaZBM89TXS4gven
gvNL1x7LCjL176MlhZ7Fa47IeRRa13Izqoss/VRwN+yFbiFwNXC8+i7sMNnZkuyV
SYQlUxf4nKFdO1qRznwYPi7DR7bURPnE2+fvfy7eWResMZhhru5TiLM5F2DtRhQu
vRbBCx+1MiEutw0IvYbVzxHT8oKCOi+0rfpFV61dwtgYyohZxtHK5nIGH/2ctr1z
0+NQYkRtHXBbuziQP2piaOB+6FDdoicHFa7cN8n6LhyDyAqOGb7w8Sr/K2zWidMz
lFtJ43pvaQnW2FFVCNTX4h2vXjx4bl0U6RyPkqTa1gH7PJHHFijA8ncHxwJPp0ON
ANyAoU8wmTbxEFm1HHq2GrEzyfFe+SLuS1pswMPWr1pkJPq42qSqRr9dyD5C8iA7
v5MNOixXf+3VyqrR065x5poUh/0ScNWbc6NlOaMtwn/sCpEamrAAjLc8VbM6Gyqw
u7Oyckwf7HxrGYxY0gMpJXyvz9KMMH3C9Lwo34hoPP3/iLy4cO+LIsL8mfpWhq6h
mQfIZhDcxsmKyh2q9xXtkMvMVO0z7Ws0Pujf6Msmgx0SK26BQ4r+Vcn+2DdIyW2/
2p16eeQz7GAI5hNYU96BsjYi1brMSgLniHGlz2Qmp0m9cFzjccKlvBBYvVOskP26
2aJ+JcW4pxr2wYbRnmpTERh30fH6MIEVdY7kDbA9U1VBFwwqjiCpeQTfThv+thMK
SXIF+Xtg8ed4P2ItBi7Bvt88aoG6dY+PI0y8poPmtOqqHlVtf3SdLK2xIO+Dk3Gg
5QxtO7n36eio5H/+kqjvhn0MttQWVXw8rll6P0UcgZQdBj0xbnk/o0MnbsaUGsDW
QUgoJgyfR22CLH4eiTJKPP7gonOip4FvLRoJHYKxArWf1PEGC+AbPZYF5/UyD3b6
5WQwGYroPb5+7hfeclVDKd+k1MrfcdYPhAKoYrQP40NTFZ6AAxc0jY6LrEFHIWcn
E9Ne4jdY2Sp231yCihvxn0WnTetaDhbwOsrKRrDXrA/V3OXXvsUbA09qM96bSRKn
I0L0NPiLA6bgHcKAl8akUcudMiRaSNSSs2xSgj0kAy+74/MUTthC+ANBHfJzlPNk
IgDgl7vHAW+p7Dp1vkp/QgaPaNwOh2bUP0jCO6Ej7rx+GTlu/aRczcpYwmAEtCWS
x1mM8/EvErGWyVwLUXwh4xmYXl6veXUFlrVJ9Lz8eLcDGmmVq+6IuIWAN43hjDFH
HUM0HmnznZAJcPuPLsNPBXYVZ2yzlo5ZA7/vGpvOzI3kmvcPlvuUSRG804Ew3zDM
r2+HHYwCeQJfZMx5Q2j2dsFcSPbYo7kObhEGFPZ2CnvZrrPWb5kWJMQvBNNSbovy
MVricgfiPZ9UtG7Rd6+Ol/wX7b7FfPUGfqPxLNHtmwltm+ZdyF+XVqGGd9YP1mCs
fxH+urMHL0+QlLTYaevSDwxqBPsqfFPdf8UituiIfn3AJ624w6EKZXfAqjIepWh4
GA8d+WUsLk4m3BOvE6YAd9tdiOCgaY6+1Qwk5fIWkrZansJlN4mLktu/fkNtm2Fy
iWvgo678Oi7eEuNBmK/jhlg87Xc9/egOivNPHAHWcfbMVmZGBgl2OLA8GCVVfxK0
m9uZgwYCrD9rA6rS4+dN1Br/5OkZRA5/nVuB+W1O3oHaU4asYWksgvf7JTekI3cb
rM9V8Yf41vFN3PamzTaePvDOp6TN4upL50jSauA5tjJhW4Io3gT7Xo9uVSkxb2dK
qORemVIIuLW5u2L0iFODiJeJopVYBygXAslUgzuzxsPXJCTEDVcafIzX9q04LpAj
hmnx5jK9GQap92ScmVZ4WujCuyOd86HS9h6DqMu+YsfO9cGoJduPBr+IfQbb3jK4
oFpxt+aKls9A51RblufI87Bh7pvJWSz4OU0QxvuI940lrbMgUmzR0VhFAgroN6Pn
qIHPLe81aV5acq1DiXmrc/0OocwUE50e8DICmi/KRKWpFSrCOxUClcaqCmd8brZS
u6yj3bLn79R5cFqkQMwQN6CsNSfSRtJw5zT7dal3nlGi1YleZtpK6g5OHpdfcNeS
3F+fZEWjJ9nfXVNK5ZHx5pGNdsLhv8vrqhA+Ystzos6M2WowaxN3JsPDMqdTIpfx
T+ellp8iux1g6xeRuYDBxzYAQ+0FHv8bNm0bjYyt4wA5mwTiBsSrkWNQcZyYxmVD
0MNiGxoTFtADmLQ95EkH5kp3jFx9f+qWEfwS+tbA7dxaX6cIJmcxR3NhBLqXkasd
czJHsPxK4BE3x08UvGDMrBFXTdtqrfUXQR0bxWS8tKtwpXQTLL4uc46yog8WWrpK
VnfSuvHOiyCECPjO4ioHK4ld4RWPXxfRcIr9HMw9iNc1wHh/nNtIKXnpdgjYtWty
VhL0wymj0U5V8dtVawRo1VMVtpG3O3mCZ65euV08q/EcSei16nyZeVxbIeFEVDj6
9uhExspeVWs5jrkJsbD3lWYVfxDyJNnYDTdKp4hiqZi/3h93rmqXf8wKwJi4pVrX
ltD4XmJYCGV+mF8ae5qC/1p5uyjyynKU6THWPM3S0FpAljiAPtG/jtyOJ72MIpi3
gGOFHhK1fDmQPIvqvE+ddlBg2lcNqruzwdi5NnWR7lr19Befr6IxLxDLQc9wENQa
kgZR4c6ePxVPl10GUcBh1cneXN0bLG0U2K8hR8LZazmMk2sW/D64OD+YWRtBR0xp
VdD28SXN86OWdAndoC+Ql+GIZeW9hrSQv+51Zl7jQ5R3Fgk846UaZxWKLNLNJXis
U5gQ6VsvwEfz9hhSKKd29J7okY09o2e3jIZekEMQDooMPClZSepEHsNQdZojuQYa
8DEgS5vG/u7srdvRhLtK5JOtp0APKvoteGPjjFvMbGt1SAkyNJhrjlDY4YQTJoFl
RSiTht/VjpEbUQoHIuij+4WdD88Yg0dVkuJTCi7uCfFNNs/rzI+RH7Jquf3uQIm9
T4Wq6M6bk0YVBeAOCmaZaCdPx33dm1xLARKaaYXKylurK4ouK+cYt5sCnE2nlMRR
6yPU9R87bmcJSIjC/kJT+cfc1AGAwOf82Leiz1B83v6nqXl2hVWT+0ShAn9pj3By
k+ImDgJ4PrX5lU4ZvIgYMeW2GmRI518q1KRNtoxTOQ8D14W11LNn67fpK6wTFcpg
ffXThaUYYRgINZxO/CEDGRQLcYhVZNMI43w580MtZtj6HZJl0vsa7KMeeIbqUUkO
vYxN/Szwv9axDwi5RRfn0JPA3oPP0yQ4pGVHnKZy75jmRUv6bP+hjiudl1y0eqoV
r2P1jFmrCbNBTI2Su4qybOsX8EpUody7sBf8CXlc5NHVGiXsAwv7RDxRnJoFZpiJ
5iuAQaiDBFdj/Gld0CUZ2UNqOaLkGicVMUXgctPWdWXTtygca6nUnBD8hcf/YBVz
Hq3CpH6sWWaOS7xiMAJEwguufMpkgusB7r1Enf31WRiSOzr6L6gQOcqU8kTr2HW8
48naHz8HzmHM2JxpS/6Q1gUgsckxNjdf0AHzrrVI2Mia9ZIdXFVpFGBHBTA5k/4n
Ap0rEy92iSwibICXBoHrgUF/L+8uEXwusHIlAU/QZnE73Oz7E8/IOphxFbjYJAKS
HAPayu7glF3if/DUCbCVHWMSXDTzowUhJnxb5mwjXUNYlA9UxEbL+C1sQBUTz6Or
Y23rS57dmBRcVjE9d/Hl+ON5kfddMyW0Fi3F/sleQSa3IxjH6aDz/Hx8n92dWgET
oWyvOvp2H4cgqJT3OqZL6V06oYULre8pTJFT4A1Wqzmbn8C+zb7zkzrf+H44xyqi
Ybb+RIWjFdW+js3cPWujwq9BVMD8kidO50axR2bJbcEKr27MODTnaBWCrDIQ5BOF
gfp2QsLi9RABYYB5uOQvDFrXqbdjdjhVIK3pk8iv00ZKrxk59WMxsFdS3xQXg88g
QMSwtCPIKDEF3ZBD1DMmDCV5mz1BiKNNHnE7fDyb1sI6ixXz96W75mVd+F4NFSg9
vikktmN5n4U5r2nHXngZzdfCFsh6sMyZTITSyyEswSjc3BCUoLrpqDkb8Vnlftzx
rL8vV4rzi5207iAX9zA53Z0mA4+UY5CkDVTzNfOqsMRQ5MIq/Nhwa8zBVUNKlqi+
+yftFgczJ5ntyD16QcHhD/pxxDBtBcHj5dv3cASA3g/IQUNy8Mis5R5u7YXfkvue
fXPp2HSRrKk9ImZ9lY5CGhxr/RprLX/nOqdUhzklB/WXu6xNvIU/cFIeI8V0C5nr
igEqHLAFKwGy1eLy2k6Z/bY1RMRT1NV3dXoh1VtRjWD+/ItXoo0O4Z7vUcCwMGhr
tdDUZ7vOlGEhWvAQRDne0+IH0u/YoxNKZbEIryedWJXxEBYi9Ua3dSZgKiS7d9gq
xhnbzWhy114x8Ytnt33LXzZKisgQKgiutxc8JUcVx2H6kRop92sMhffL9ybI/fg/
JwJi5Utg6krzZ7pUCJ8g+p9jDylIDXfgR9AKJADOuRb01ulBkWFsB3z59XZ8PFou
FDCpWpHWbJ8NaXbR98603ofN6R4AfPGPJO9z/Ept/dGPIKgVK6LZO/V7TZ0tsa2f
VfFoNWr7O++YhHMLQoj97jOTkhUWudLL6DKKLW3PeoJhR6addWhGJMwEszd53cdu
/5peKJkCVSQg8LnbctOsgVlGt/20+dOPEH/pgui0V+jBXQw21NMy/n0biTWxa1U/
yQWoCp66U3sMSynz/a8/HnoPHhlbLrH2Mslglsrjpr2Q/5EQOUHxlBPl8fkYTGId
EiUHkdxA95gUykrxv++56UkETxaCvjyVaxyYTp9o+3Sb3EoOlEI/57R3w9CcZT9N
DyJ7k9RI+iZP04C3UqxMU56ftHVkMqG5DxiG4f97B/ht5E27NC/two4Y7rLSneQv
70gfwWHe9S/vdsFUSoz002/KTp1KQGy4FaOzXZYugyYdZeO4Hcft8oFip7lvqZLx
RvC0YsWt7Ot113EUCCxtHVZsW0+wJNOTervSqOc6kspg6cJx3VW1hcOLZEs1tIIJ
LTtdtAMtbBLMrniRf/sNSnr0kIVaHcfuM0ZcWWTjqzihsm3W8DTd3m7YIHvqIGI5
5EC/fpb1mVTz31tPKV6s+hrMIMPF1MFKRaVpWKmyd/57Tgevc3loEEu7gYTya42L
TJJcJDP2cKBtOJlt2b33aLrun0spcy1ZWFQLpQ0h4CgyNQ70XeMVMSwOdddaSdSy
1DW9+iGJOmljJoBtZcQXtXFNnfWgSMbdd6gpcMWQl1yKTT7H5MfUckLh4R64zwLt
OBNrGF2PGPr7YfqH/u84xC1NBz9du+kLwIpA47O7jO+BXAmecgte9QEHHLEIyQ6d
gN9PV+s2KrpNB1j1FFP1aCIZUUrOQztAbC40/p24uoeKnB/HCKQuiSUc55AW4omI
a+udoaP/ESkfmS9eUOsOK2NHrS/DrOcgKMxq9JfdpFzsLo2Cf8jAVh+fBFhvM9Ux
zGx865OeqPfjXKKH5YNC2Am+zdN+AtgHhJdwWYf3DMQyhNDbIY+loV/JrF/1Nr4w
il8aWQF1rDtxO61dlw+laCMPrGuXzjGB5hKahAMBjaqHax7VXjmxAo5IvpeoFnqw
tyTSxbOf4rIWcwnJFhH29Xool6HZKycDxvMIDkzplnQ4sq6K+ZZuKiMsBB20JSLy
PKd+ycO19/zMHO3Z3tqlUXcDfS2vMtgNAylWCRx5qjzH0B07St23Dk1G+r3UXl41
lKpigjgu4Ya4QY+GgrvHMq7GKWeAWqgBqGEZ8pvcEGnzZPck8C2AzdwJxrAjNbRo
SIxIdfo7zTUAvC/x0PyovebDQ22UcaapzSoezLvP/AHEB1y7ZHs1ow6IDRJuCgeA
97le+L70HmTIrRq7m9ChjjVY0S251OIGYhub2KxADzT+RdtmQtePGvjILowJ/lcx
0IuVGG/Jr6Ygm17fata4e7qpEK4axh4kWVBdV+2V0qf0hd6yGg2IaJJ9KB3Xjy6N
IbR1N6hfSNX2YF8eY5V7thMjeN9VbKS+7qEpHgzMsXt9FmWlxKUUAzDcd5b1MtJW
sTo5LDRgtsBdxJa7HTEw7DINbfjF4w3mOUkyvKasw9bZ0o9GUA3eOGWb6ZpVayck
kFgGvalwTSkeNM7NzhBxD5qg9Hozs7J9VZHld7lsO3TNkXCMxi9NdFVfCpgJuEGK
ZUHR9PuUnI5WtROIWS97yYkQwMGK+IQvUVhQSDO2LDYKfJoLqsunOE+mj0wG5Ap0
HM99nyBnC5/7nN+hLJIn8AyWr21jw/+wmSAelODya76qfWcvx1DEUsF7EH3aOu9b
gI95dx4hf/nI2zXGb8TUCwaFKTLi14NAssP4AEiVZMMHWdM3bAuPquD0qUMCFwLr
tKo8p3xlApGWl5ug6Y+G9laCeXZEkL98mH1zLE5b50VA2hDZHVe5f1YUmCbD8Mo8
RS9+5TwAdN3MwhBiNlBJQKysG0/IxUGq41xZ9tsaHuYFaZXcs1+yw+7/YgL4G11Z
28NmpvYfqTpCnDl1QYu0cfoWLn8ZBgXtuPpf9hLSeoDYk/Ay0qZEYItKa1Bxg5NY
sEh3APjEdqD81/USH7cEAD2NAK/dreomQDWYBI/aPKaBLsp8McGHUeuVqbZlK7A7
yIyKZDObVbqLHs1B56CC493GuSzH5GhviH0cxQ4piSVXPBAhptuqlJZtcuWXtpJm
OPXFNlImL+QyOo4P9EVG80DgpogYj9fsO05A3a6TSsVYYHRjnrQrXoBEym67J8Ns
90Cbo7vl+tJrrrl1ysX4H6DwP7Yfbh9Tku2fcJDoE9xSVdpscv089j7kbC7oQobc
fQx9g8Nda2pJyE8mPisOAf8xn8bCsBbvwPGtDom68Ll3R5ECWw+T3yJSJPWmaed9
QDs2JBWehC7ygDa6iO42QDSQvy+Q4vJ5Psv4W9CF9FYVjbQCzk1KzfDCzKdSAMx1
42DRaOAi104WZ1l16rdfm28Z5ajE9IgDKMe2MdVF4d3Ge86Ka0PhiDvxtA8a6vW1
e867eiE+A3IDbWG2HS/sGNmMs23hNHqKvSz5G3qx29LmWbEJn7HijzXhUhAtjjKV
bdTsgaj947KKaOIV/na/Ju0l97p1+ajxlzRkMBVfjCDjIxR7L1Lktl3aMJzAPYki
rXJvGh++hMHF+7ZJqm4hQP7SLYlqCoAPnqURFdODUr17Kws97D9zGrp77oahM3L1
spJy5KgGD6JflOTeVcW7Kt3CcbYejVjWwdq4i1xxiPt1YY9q70DqXjmNf7MquIT+
RgtUEQwXH5Ui0bOMl77PMPsiRSLVh7bbi58XSmbSHoTXc09zU8zcQL6/1G2SHFo6
Z6Snu4wqUnDl6YBk8t3AkEoq9OT0HHramsj9jo5GvGBmLT3L9kJhmfPR8P7TsO0h
T6h0OkelWxVekysBIYyzfUYxXgDPQVSVKyTblhIpcQcWnQ5P9nMAXa2NLE1D/98m
hMrLXPXkNNXNAO5bOcvSn8+ddjUNtp6GvepN/0WAOKS9JuIbDU4+eqphmZUdhSqN
cWkLxH/T2nqUyQVakOXSQutoUwJ+i8z6SizUQOq+ej2mbUekrOW2qfa68vC+hOX1
yTvdCazKTIa5F4VhEhRgY7Y4hSPIr/3lt7DadMB4tdLPpNrZh2y35nvKRuyJ+uwd
RkmladHIQ9s1l0e8vBIvMWDXnl6PZQ/bLU7l+MMeUgw/6PAoadlak+wafWQBDb9K
RNMpaWNbHIG10dh32YzFwoIdRtkYE+1XGBu9Q0+B11TufRMRj1q6f6qizN7yyIuS
n3zS8CqVKJs+95nMWd3puyhya7rlbz8igJbzJJWtXDVSpZ97XE9Cy6Mn/Q1Zee0k
dllrwhr6TCcekt8ZpI04GhNCQibG5rJqk0WgaZYDMyWi3iioKpFUvu9+Du+OlSld
Gnu5s0RCFzswPvLKoaqJLmu7QVkEyTciap5+Ynu5qXIHOfBEps8arBMlYB+GVFe4
fv5yJwlOeNyJP9X7aqM4h1aseFNo6vIkaZb01ISWm964fCLXHo7rHBo768PJZT5c
rZvEZkZ0uudj7WNB3SdRMauRjsQs73liwOQtx/wwp6sW0pMbWp2Jd1bW4YLFGNKo
sUOI8kM+uK46Bj9vaGO65xcr9iEh8wzkfWURYuCmj75e6i5qfEM9IarX2UxVBhru
0pSRFqjKgiAr9RxoUOnN0YK4DCEKu4lV0k6w9OLoAopFZjyCZVcOT5BVSsk2w8ia
NysOYJ3uxOP3ZLfSiuqGR3NllRZ67zy/CjGwYu9hUm/iYB8xRMMvfjLYepQMsetM
/+InhmlmB0Cvai/1z35YFY05aKz04azpdzwCSL7E3Nyii4Q84I2NGsYmcSVt8xwR
mvYnTymNnYnGywK21bBTN7eTNWItHhLpcNJptKm/mPxnAkBHr6tlnYBQ4B/tvT9h
JgxNx4OQuTr4QE3smMDEt3MSLKlytcKt0bXK7pNg+WRLSimWFLmhggAw3XdNVXtZ
lQc3EW1i33+m6TEpnUFeUmgrEafzEb6lixOu/qEpXSiRaCkKjD20lFXlniVvOXrB
L864DUGggPNGA09byc4mXkh58oiwfNLIEnL5RqsfGMX0Cs/62BQX2r9V8cVOLLw8
/ihl70NvSvb5LPMeMeD1GaXeTiHNOFJfZ9cbDEw8GRC+WdG4uwdGElQ3/9gMyRMZ
ChWPMUGeSVc+n2hxD7wTS4g5hwRNjdDaLr3kecIcc+KXYgFLcy8xYwyt8NfRy6pU
b6Tf8Bfpn2XBhZS/kYrr8VBuOcq4T/CeL8hkQv69iclzTSDP/hFV0uPDoSN99rlJ
IEZBy0Iw4ImQ6wK/2Tc03vRMVp6HWVWd5m9azHfUfX2QIgCfQaRZfwJeU3HGyLz6
yf9RWEZgDyKu6G63VTQc21aLyZNHPb9m3fWbqSsZ6kAgwmslBv4z1gdgKxhnuiws
Rccx/wwlQMCaaXpvMapOlDUS4Sw5YHhLF88Q2ePFyH2AXonjDDpH8DSCB6kq5MvI
Z3KJcuM8puFNfx2wOEbhgO4mD5Z9rbA0kn36f8oV9DUnZCLxC8iU0vdQNpsGFOgl
sfJGvv412Pt7mVhyvYgq7C87vqZuyM0TU/Lmbt2KeaNrj4HgECCsGziDbxOH+h4U
8KQpY0BvfIKcGYGY6tOUZClGuuJvIKPBUAxJQrI0z6nfpIdPSE/8msIod2EKOnVm
7+XzQI5R1WTKFSJdQAu2a3QnVrmRcvbikkBXTr13/d/+EpTg1LrbRVRNVneaj2Pq
L4RZ01qyHHnVYAH5ecB4EpUGUtme3lD/HUV4rYHrI4sVkENAFVM77yRVKL9q1+OP
S3uaeRgyJgEsxRGzEWr9+O77nOKf8UR6xWM9IsXX0tfgkkwS8RizOU5EIbA+p8hS
+aJ546doKnbByKoOmNrdsKjHO+iO2r+vcwtI72RAakAyoH3S2trm1L4N8sGbdtEo
WUsbL/HJjV9qU0PdulPZ5jyUgwkD/fgJoC45KbaMHfaRQCwqA0QwqRqmCttB9qC6
c3yCjuw/mi4l57kQs4FyLfwYSqaUYcrUDk+CN8pxyX31X1UOBbd5L5aMHFGFsp7u
DXG0LTjOCtDM2poMbx2jm+1cRWhEfsGERB9kUvWvikds+TF50zPQkNtwZMWZewrA
DhrRQ/Q32X6bxy93BrtzJ0nibI4/CWK4AiRrRPN8uHqOYz/iqbBizkpiSHFAwykw
iomUtQkYPbZdfg8camCMWb3viBAHtyM3bpgV+l9Q3tcPVQ2c14TN6RpxYXZBX74M
4o8Nezbf8yciDAfsua/+W2oxXyn/cJQH9GC9raBb6+ouwgl8+nMmZszMd05ho9Qh
4+y41k0Zqcbuq7LsEIjF4OOqNAL6Eze7r92Ng4x6eDM7wOXX+0g7GgzIJlQCekrb
RJFRP0lTksdKGM/6RlSuzSfHf+0wSqDu5ihwPfNdcaezl/lIfqxy0oa2y/qwEMqp
zn2KyZBoyShS0DnpDJFWcuDv6pWPsRlIwkzC8+OBnOn8kupm6IhS1m+SHnkvLaAr
N17VObcj7WLjN8+77SUM6/jnDhJmGsRUrIIJc0ANOk6Vgt4H+JMvl41O+youU51o
Vdmf5yLl50W/FTBgKtvLN+OTzMjPgdwO2QGaiWEMJ7bbcJUDfR/g7USXUVYyAwQ4
j7PoWJzFLcY+fGfGlyyHqAilb+AeN1Mn9dc2ln16XGn1iZivgtTkE5FY/qhgHVQE
osnRsZ1Hg57q7P7a3nJ1D2Be7vn80iA/pxXrnMjwR9Y8phd0CVbzlX9ItcsERTGV
zpS+QOZlErw+F5eFthyO+x0iDroePEQbOJt73z73Fs/V8V47Ckox3/eVtEW4oKw7
6mDoKA+hXg5ro6MldMeyPa4F9QvhbMcTAldjduii6FeC5OlsPUtcmeo2N5aBrL8A
+INtCbHDHEQqe8tFCgrrVtQ4s8ChZ2n6Rz5sJJmKewiVguTb79Dr3ff3mIT9H09h
jCWcNoT0MEruFIz+Jgeftqk0ClluFR1X9VO18tBu1NcF4HcxIlrcndrb1Y+ZN5+S
ooRE1naZ2X5nyFsS/5SSi4HhYENHvd9MuoThioM93rfMk4ZChk1VBS3tZpo0WfEG
+hUA9Z97eRFzyb+SfapAPWPLeIIXmfz6ywWra+7uC+3BNLsrHEPFnq5Qw8X1Qiuq
ryinza8ql3ipDrS8t6fEd9EVSadCEsdk547owk9lGoy0zK/RA81oEgZ6cba04/xi
K1aOm/WdwsAiT8362ohwCNgJaTQRYpyk/LUUTj8gdoE4YHFqqIarfFYq3/fj9DVh
0dEAkU+2QcWbLTQv55JB3EzbvqLU1PFTYHNPv9UpxjAKkKyZHVkTCOamyxwkwgGe
yKj7xRpFX5toOge3Lehkyqa28GC7Ibkloa+YSSkL65jS2iHHtxuDEsb4CwqZbrcs
+PBuwxQm8RSIspApSXGn/o6BZkMYs94iPGgk2spYqqX9OXcgGuEVgNDNlH/UTp8q
YVcBQS5KcOeu5jH52F5MDHvuTWGhvgi0chbn54P0soQS2Li9wPzC9nu/gSZ3HfL4
K6CK+/maMVm9NJyLMtp3/KA1nyHXch4MHgX89PKm4cyJth9hkcFPV1f00mK3715s
EzOT6KOYMKlmDnj7LMhp4PX8HZX+FLYdl99yPy2R2MWeKwhjsuWjyskS/TUYCUTH
Ce4qeqescIlMIG3MzXtCnDlPakcOwwq26KTNAochlHzrLYyhVvHxxU9nDKc3REfG
SEVEgVqsDE+oyj0rrBJ4lQxsKHdw3100u719gA7oePbi8jHv6frEho1cXDcd1X+9
FRT+qh5eh3hAzxynE1bikQJFo0U3+/tnvZ95UTZNMpjG00krmR03jK1Y9wS3lhcJ
60CBsCKkAkKcjUiCdhCRjq2f3A3jsLH6joY0SnT+W3kq2Wb0JegNZxfryyyvfuWf
fAL6D4kOLaNyLFtlajqFZbK/wRrM2AHDRnQdB4UyxuVyorhNEApH9gxMoj3g5qaQ
gdBGRkACwHi68QnxUcdyP8CvmY5TAG4Ww8IF4RzyQD1qZQySsK6fW4huNrksM2Xv
IGVg/D53JVML3YTldWQRtf00vHbxPtQuVMWJtfWqJbt7S3v9ndu1RESody8NJJCr
I+GRXBh3aoKVXZyicf4NhqOpSXB9J1bIxpIueq6ukZhFYDyHe2K1IrJPkksfsyvK
c18hHF7xA2pqzbZ9v/vdb0dlcz+2/7FFD79TNmr2GjIEn1pUvUZZ2tsIjLG5KPHn
g7exW/Ka0hhqFUD6lwbSx8Lw5zuNHEl4AhOq8QA2N85Gi5NnTaK2yLB6f1wmPuMP
m8UYsCJhnbC5UM4ihoKK6t3A4N/A9BWWe0J0EY2O8G1OySADgjt65AK6vZ2ODtMh
2L2LbEv0L/T/EP5L909sb+cxNsZQwxi9svrS+xvvc4mjpHjFLMqSEZP2v+3suRIe
ppEhKDU4sZ4iMvLvUhYzUB/z69s4uuJ9rH5i6aEzAlESU2JYLQP30jkkvNR1IHU/
oRExaE7tdql+HFca/85MYBi8dgeqc1AKzGVj2aeM+Fp7keOGvHBUypYMSQrVgFB+
hGVUVdHAsFxrezRcb7yLnTwp3Ry3sKE0lGDDXpUdBrlwpSVt5B+s36JOakAWWyvy
5cSHCN682m/knDT0FMIysnvG0Qac4nucUQ2FoFTgKT6Ve7ucW8bu1yeFuxdyDA33
9jl9Ht7OPaWUT1KjLIhXzk4fAjtpc+vTvzfhig31BkmH4ehsCxyzd/DORAD+TlYd
+Tj73gUti0QzkaqwMGSwDO+0mLvHI85YL0U4OuIK7yRXaKARrgdee6q2Yqe/+Yd7
xXTLoDgqyg5lCrUMgeqt9S6bpWQgdnvgl4/DUcQoNDa0SgzsyEO7iTinyWzHzUNU
Xf/beYejZ8KuV4DF0/335io8HJgpDe+CZM7ye6OuRuBNrETw77pBfeu2bUCmrovM
QT1QiYelld7k7wkfv5B/b0EsGZ1B+hKmHSxnIOOaEnq0chkt4uIdyrREz8mYK6/+
EX5yFkop7GVgGgRVSuTqIpdDsxIHWCl66/eG7jX5xH+0aIJP2XYZhNt7sW7CamS3
VockyaoJ3TYFfdJz+Jkx204q4fMTCeV0Bm78C0acFBlirfzrMBsa/PTRDTq0Ocgi
ihVfKVH6OyDl/McGFi+l8ggp+0dqeLk1QVJ4vf9Xm78B2ZR7xGrTX/oIB8xQMwc4
siZ3WYlgpBQnQjtXxwgYwWLV60qlVD7Ep25e8D27Egf/cwg3PxEQjNUuvE0/WM00
fcBClb7sOqq0bAL69V9ByaUfbce4iT7WFa/ZfcErmaLQAT6kv//vQxrvlocI1m8w
kyEgnAjAIvpkc6F4iwtz0xIofWBJEf7L5LYBr7pZ3mKE6oJrkDP6yh1OkWbCgJto
l3O8sD0isYhkA28xUwy2+ZTn2/T+3JIIGIKCzOritVzPaDNbbFMunWITD3FxdvwE
9wl+68lZ2BdESxOmFdvRl85JAuZJOf0dtrpuC0g0uTnvf8vCXyW47svtG3G68Nmb
QzoZgc8dF6N/55iYwFjbR3wZjmZ5OkEr89piXVeotnyu8LCPTPhCow/FICOGF7a0
xQNfkU4oeP2w6TRAoORUHDYI/q/wRtgfseJCrjMPxTMXhm861CtfEtBccqZRSfkf
SnSYrfa8p3saPcpNncmiJdH0kti4xH44FDV/OoQR6ID4QYMmUByB7TStls+k2dmi
UFlzog9GEtR05svgyj1Owy+GdwLiQbr1DYYohnRb+ruNaAZOxrrNfxv/+fsb+eIq
3s3UeNAnhdA0R1bfIskLwumqEwfVyE88X8kktxH5Vrad/vdp1e+c8kWbQCT5CsKK
ryymQy9dZqXTbkKnTzadJ5BrP8F3xjSU96PEipbn7Dg9NsK9PacYjl9X538jl8uJ
Q3GLwFn87KOabjWuiAAQYkqFr9ihVNvMMUwHNuaPbuOkhhEME4UvdeLkGDaJ9vjv
wOVofPH7wLKWyOjAM/xFamU7zpNgvM2RJq7kWjBPffojT1AYJbX+1hu/S6XB6aTV
RBzi6k9961eWPMTakhpUKIbEFFmHkUnArH8pV0fExbSHlueVwlt1iJEhai+alkSv
OH04c//HGVYYjdkh/cJ9Xc1TJ946ltGJ9GxbyRmkeyal9oCrrjZ3MCWjrlz/l8Wx
NH2EoEI5aElt3sGQnlso2llmOPX41Y6EgkLgUXMBYGvx3FXVn5sCN+eGgwSr2h5h
7Vo9iv5pIas3F5I8AtTYmRMVIG1w7PHcKbmdzZCQiYpIzj96WWNfE5SafzZCFavB
EoxGsG7VcjK/poPxzOVPfRrCe2tkrQ4g7sHS8+G45rSGlCus3hnct1hCeIoRXGbA
IFJ0EP/XzEH4K1ycnNu8YAdBNPOVMyeTGhXo7oGZXoJ0hZsDqx9yUlZljbglpSma
gmUthQv0OSAHjZNBmD8Touj9LwoHwUDgrWY5aD0qVpw90FS8TUAQnrcNhuk/+g1R
GKb/KNsinoYAVBFUnjrAvUoUg7++ASdNsx5K95fbScbFk2z4eXReCVWvhjaw0E4o
S9qit4m772YvDz+74s02g3XQQbJJNYlQKeEiI/gWL7WFGqNetyeAqqqTHr93maUq
6c24EbMDikFRP1JfECcVbin6Rh9SyaMII93BbytznhvhXmfILJkhsBK55T9xPVGA
0+4DNIXIZlMQ9DbDMDt/lJCwsG0J761269RrDSOTU3ifmMvhx1HkvHlYB7XInefL
0ApPXXijGYWyWjBcSCXFzDyYBkxyrqaxj0O/tTI29LzgyeMpwQgEmEP4Q14Mv9qO
jm/y+1121YXKDDjyjuTMxtPEVltn0v0fO6SbsJuAxJD9sJFVYoGIsVqY2AJLyknD
1HFPJGyEPSKWgxbeqIteFsh2GPqIS4/mch5wq29wCaly9Vb3JUP3TfLCBKRdvtSP
izV0qPgKLmMx3EyiljqvTbFFchCMmuqhQxlQjp+CgPcsbhpIwt+vCUkEPSHxYBV7
z0gwRFO4m7/75IyTfCZNznO6qy4HkpDLnArgnHOO3qhgYahZkSbERPeHHoTCJdKi
bkD1UOQH4PU/Zh7BSulc6K0SppGaNGJWy5ahT/cySINod3ViAcDe727av18ndiOl
Pf4rwJd0R/OJW3zEM6r5L9vdql/MkRk0zhBiF0c91DShTyj7nP6jjMAM/JmDNGru
CKmIEGJo+b4CZyTILFCa5ZSo/dnofEVggFZ1xqAye6zN+5mWXIfsQbQSfBKfgJuN
4hz75Lz1oFPT+1VlRo44x4Jki0R1GrrSW4P863BhvZ/wIpqW5x4tEEP3dHoVZ7RH
fIpiUEZuVQfIHLsl6ZrLHLduBVx/7pz6STpeIMwlot1oN4YwIYCI/7BFNY/taGeq
BC0/Wu2HTw0TnBdNacFUFkbHr1+K6qjwiO0Y6C9anyYeCwv4BjlwHaTkxGiackKo
NVUyn5GWDpDmKXBxj7zCmI1lT1XeDF6L9RPnwIJk6IHlrJAGLc0owmHu3dPIhrP7
AH2gZtaNMtC/qnNAuyA4pAivBYMBEyUMkHU7FwslOatj4+K9L0JoOPoB21ocD1Et
Fqdg3HbC5SNBDMYJF5AFQ96BJpJl6HrZHJ9wHasL0MhqIaxO+sDY9UFjCCdevv3y
P5Y1f0ka0XFtesPVn+6qMCNk3PUR1/blY3qRPjzTg6p9Fb0f2hnsYPQZB8Zv9PhS
hvyMF4L0jEgZkDp9tOGWJEx8X5yt2wSQAz0zpjQDlHVWOfPfNzqhiqeP5AxyWJkO
UfO21CijjSu0sertpZSsLsm3Qeg/kjjCDKLho04NkroRB7fp7MooFnU5hQEF9cZk
VY6N8/amRHl99vM1yfF/Q2Y9jZoLqvCF7R8Tz/8pBLixTy1FoE9gI3G+Or8do5Uf
XLeqzAAQVS/kr5SMJ0onHXvWjcpKtbxiWUoGLJ1lk9Z6SxiRO6+mnA+ujsTQrP6I
NJ7a5FNyW1e8DWrc8FWRO6r3chTBJueMGJLWCa2Ujxm3xibH0e3IKYEulzO+rjGJ
sgpQq92xsJjQKoHE0HFJCwmHbsTRw3B8c1nKe5tVk68hW9gh4Le94rJHx3D5MUTL
+Tv8r5kksEPPvsrMGNWle0xzCj/CnllRUrccR30r3REar9stzXGmZ9W6eMQmRY9K
kwSmDiaFS+34G01iGxpEf2gjSGRUuigOEw7niaW3BF3I9lLYfBo+zysEA/MdC0yR
HoqEZxShcyimoJqaXxeywk+oVS6onSxD+LridCXyWWQYB3clwBbNzRPKdfPb480V
QEVIIu1PFbB7fZJuEZQPjshbnPqR48tKQOz4FU0bMNHD6p5l26N2LcFVyeM1ojQe
i+PH7cI8Ju1tCbvVZSXu43NonQDA0fDNC7RTvK+jInqrUdmPu9uulsq6ZiH1f+3u
ZHpdgpsUoraKu3ujfY5eh41QCae1OZ++/ewiYObiHuTTQkZx8ZK88Rp8KCyk59qg
DGQhN7f7pLR0kpOUPIgOyc6f4KWOCu8p/UtWllAfsASSQnHj8TWqoygYccCWJQmG
l8cpzVJI4UiDIuKLECL777sz1tt3sKHnQIIwvKONq2erKpCTqwOLbn8sb/yq1C+U
UaqHHselJkYjy8DOUCzW9F3wNFZzBhuLeM+UXy8Kooo3Gntb0RqZ3MU3QkeudrNg
w4dBKUzh9A5Zgmy0LxrsrLrPyhtpMmtgsGuBPKacJPrXiNKiemSwNYO5h3VmTI/l
DGWjlp0+OeEVWnFiBsq6LiWsf/2vw3it1Ff+4bi/KBrMiTMGMbJhVgATnAVPGGcY
HF+O89SXXJZ5GYemOgs34xeWwc8KGJfghuqm6AgSuDQv/xdzfTh+GVItZUUA+MWb
Hy+WnvnwDfzjVGlRi3cDUXgCgEhMdiUuI6n7+i2tMEAzruNk7Da4PZpUrBtvu259
U09RmPnMaLUFGZzoAPDpQ/c3fyveCP0Gf29Em6LA6fBU72hnfUK5Qw3/2ZGASqEZ
PkdgH+8VukKYDO1RONdyqM7kUxLzqHg8Rg/vSEln9je/FuiINNZa0P0l1hMRQLZT
8ir6uvgdaDukxuYa0NudKZUam+BSpcnT4h7yXKZj+xK+QNGFfw3GRVsAGTFgekHr
jCU7LdTt3DK/BTk8adYFyaIehLPOf7yzzbkh2tMD9cin80GYejsM1+33XxSd9v6O
67pWXLSEix+itGW8Hh+2jZLCqdF1G2beO1+Lw2IZq+RYwzgF1iwB2rKri+wC66oO
tt5sqyzYgJvXnU5h6CafjN+0DqQx0f3/1aPH5T70IPY8WpGIPKvDjSnUApUs+X3s
+rCTXlNRJvR9sMsuMAvaKj/BB2rqfHykSwEU+N7yVaO6NjeEy/qSo/3rq2rF2+t1
1t3EiiUBUgq32Q6uAyRSob87UPAv+Mos6Z3NuPMKfijmhdOU/Nsc3gROjrpOLkAx
XhNekRzhNqd1nK19Fg6DRh4zRQq7rtZbhGu64Zh1cXK7D0Vqwpr1b4qbBN16c2UJ
0fBRP5NoesMvi028kdoaX2df4DMPEtmornbLNl9zk1qp0v+9Lujri8cWNyIatFdR
V+N5m4xwhYQvyH9+sYct0kIdhEohWFSmuN/S9ou4QNIUAusBXrzuIyg6QqXnneI4
saYLk2bpM96KCU1/nRSPLCprKdP1P5wt0gh4Z6vHJTCHy3SpAr7fuv4hnyFtl2O5
WGMV79ka8CJT5DFcG9ILy3E58gXp/g/28PuY66pUI6IKezKCS7eJLxRyEZxJRqKj
HGlBvR2ifZp/30FkXyCdBFGnjOvQDIyYuEZ8yzvVxou6nP3X6vHtynS/2mEq6xXn
glhm32tkP99oHogCIP33Y8n6tn9EtIbAlsoi802Auqh/zfYUkGtekk7fcmHmaffl
NJbHr6CsqHLi6H9kMqIeV9sWIe37KpZS/hiECSmZqi1BLd6pTX5T1uNVILz+5ISi
0LyMHeWm7/pVUygNrEPI8cB1dDOSd55jkleAztdbrz345V/m92vKbOgKMEth9Lba
jkaWmctvW4/UMRMovi3bLLjxDu/aBSIv07u/dSyCutT88+r/e6qvE1ij6tgkP1OZ
C5c8JYhCHNWZE3vt2dZ/Q5Z8WihhFP2SxTVWa3dLAqmStL5WXq3rNF808dEsuIp/
wgwI0xYXOnByIzAFX3XSgAh0AOY230l+837uhRjBB16wrMXK7Ge00KCHwKxjyyT6
H8S6tQ9IVyAT2kfpASsvyuXwBJq4B1r1mfFTekP3HK5DDxKlVEv9RVJ5a87bgAdL
CFSN8EkY9zh8KbDm8KD8Aef6dvd0+FNwMUcXz3PL40axYgcvIEjl70KsVL5QN8rn
ChOD+VOD3ptwM8F97cyTTrbMK4Rk6LdSfQivMTgn9drbhZ5GNV4wDWr+djUBe4UO
Jj8hHMlSH+i2vxtXpe29gZpI23L17baPwGXKetQvpbZk8MpsGntSqHUQ6+BxRIbx
B93Xteg/QW7GlWR/X5MkiwZHXDeEaN/9MYIzdWqIzHuoK4Ae8r4+BYEtNs7teY1T
DpI/F5DK5b0jrlUg+rkQg77HQG4dyliEOIpoIxwdGFMN2T6qKVlQ+aUd/OGzX4TB
N5ejsHiUKlhbwdw6U2qDFCGXqGy7/EYK/IL67D94cm7AlSPd3S9B6897tScHkwRT
tHPBHyTyNlok7Zi9utXY7hTvVNe/gX9nea8aX1tNQ+e8Je2wtTxyAnKHfYFJoAaN
iiKLTyYiq8jQXeCLThrqszaIuaLyCe5FNuG4YdMyR2dGyiedVcrRoQ4QXk/BLh2S
UuCED4Iyzo9oLp5zOeEnAok1/zYZgnqlDgaROvLftJwTOcPC7mxI8WBEeOwiCg2K
wZoBuqs+cUjjqwUGT4BMLVy8TLUejZMkPmKAn66Djz2/Gx7xuTvWa5A0QeYHB1yJ
X4CUOk+LYMEm1bhQVQMrpn0W4phM1LGru+qHemHZ/iHBHmnEThMgMuxKQM1jOVx7
KYhAc9hjmwRQxkScu4+SiiD/XuN09HVPsA4PFZvXisxGfdMV4rDlhaHKeIu+j0EQ
1wEQGJrFMXiBwHe1TqQEHLtnwQGscZcR1IehoDOgYgBGR3mjOaqfrbhPhF/nCq9e
AM+2E1d2cuUPcMyA0azniHuQp0Sabkalw/2hHHRITqww+aqtjsFtTq7U5yiycwql
09fzQnGnNbVnxisx5mzb6nkgaCtAGfgxtsxfz4EMx1JhesQg7vqo2VBmdnNlNAQL
jf0Qncml6+P1LtOtpcjlCHlsXvtKPIV2AqrBk49oSyhQG6krwVqYsjuJUWkiU//c
tNGX0Qr6yXI/lHTiWAKB2+zcfA5g0h4m29L+Qe9okeU3ljh2j5kboypAAxJ7p/2v
0uUwKIgKyzgUO3KGyJLpc6lnz/m7Y21ibampt7qVMPQ347awHyK5MK7UG1idaG3X
mphjMy/tZ9WvKUiTr70Q5zpFcgGQ0dXG905P+IWL3+rjEPP5OMzU1Q1hkY4PQnKf
OQ0av830UzIUzMAHE8BJUqRCxok/UJF7YYqr4gcZvfSnh4eUoSigLh7a0jYwL+GC
982H86Ye34OtZ6jYMCiskrEi9h0s4cuEMmGfe2Z3GR5BKQxI5iax5oE895vD1w6p
i2J3A4BQNEapw5sPoTfPMHMWZZSj14NVt/9086YVumhYup/wB0jLo2Zn9ccFmwfj
qMx5z2Rhi3+1ukF+/34W6wvmwtJ8h7DwGZ22wh6FYyXjEdFiW7BuCHw7EibRu2IF
jeXVlElGkq3C8ySfcfbsikwLwODJiK2rhaOiqPA5ErVh+ZUN38fKOyiz8MBVbgHk
0jUlAC0zXcM0DyBOC+WawjiCY/bM48JOxs7cgoU7y/Tj/jG1ttG5tjVDASysMAaQ
+IQNfv9uiidJmyUwXcUZRLb3EXgdbVEbnTy2AkmbfHOG2nQSnt608nyYLlDiEBx8
Tpi2eQgKRkt/LSbGSk5O+raPv/CxoWik3DnNjixiGzsmug6TW/EAKqymHHGseKFk
BejZOCRYxGYteAblKJj0oWTY2Jc3ytxvZlUd61gUl7aeylhu1HCxaQo0SapM7u91
TtnMd35MhCQo1R+sBAqVFNWAFAokiqEQkrjErUFExfJkeIM8iWGIFfcr4VTj+Tko
yy6zFL8vXuu/72WqTqO8HVJtCC3zOJjsyUXjaOAuzm0pAZJb/e6mouoLCK27Wv6n
bgERkSEpEJo80p3ZLQdFOqkl3UjJeJ4jtVHYvLlJJwwVPX32FcWA3iPjZZ7WZlgs
l7DdzEXiUipzTwW9xfxzJYaJvmiM80Rl2AR7oPmokXkpVePhN6doD3omPODQbmEw
x5tTfYKzjUdvp5GFTNrPShWdbm52kTZ9cOnCq3g5/E+21AB5/7lsR5bmKg9S+7je
BXpBYGPRsjl5w3KhuBVn8mAr4xYiHAF+ET341iKbgo4ya4g6P20zHsc6mAuMzYv3
o5hswrHEU1gjH5pQHXrKkyP5l7ZkSgYPgmoeNlENkUQiXgpyhdfZIpd+CdvRMfP1
W9sE0gcQUOnNTtrgcM8nDhAu99G56FpbEcOouWPfx2yKCwqwFSSjLWEjzIkcWa7x
EgqSUOyeslvrKHAtArb6Auhb5Dbz/QCgbdWALctVUsXpFuQLS7ynI0my/XO3ED5J
Wj/2gDrhHqnsOqHxEMjujK7r4oCVjuj8Xv14o2vp00/DNL8KP/HhuAK0sCxhArSl
LZc5/OPlSHKN1R7vU1gWgnqiBM/vFIpuXDq7v8tO2l3PPFtqUxVsdQu1Hvz/FqbL
noY44enueDXlY4+FJmzmkc3gZ8MdKvGOvN/ORf7nbMlpymWEasVv1HxGsfqhWbI+
kP9WfORGLBs2Q3pPqU2SQiE3aBfS9BOEs2jQPELowsnNpFHhvIAmz3YyV1BBujGK
L3M1HjWF17gJAQvx23WrsRy/jJCunu4TyjgjRfnvaTWhmv1He4zWxq8vbkQeU3Ct
1JeOje8id9cMTE5Dv/doGJwSXGsMXPjxQmfwBrsWZo/7ZrqlFTpcAxKnY0R6Lgld
UOK8OLChtSQj839xYImtRfLav+BP9saz81G5luz7ir6MWqaynmX5FRmm/3sy7Z/L
os0GpM3ZNu4dxOZSwGb34086aWJ9/lyNF2TEGphVsefM7bzdBWBnow7QXcsiuoPw
GCwCtt8NTOKz9beNPSVcCvYDUEN9hY9uqhITwJzE674T/F72LV2ZYmyJLxY4kpsK
4Mh08BqhGVQe7+ln6SudOJGJxgHjbReWnjtCKtNRQMbK1tmrrotu11zWg7+40iXs
a0fwbL8ZQGATCMEJCFkGfCTohYBxj1BoMy5RE60la7LGUSc852cIrtNsPOgpxkRC
S4+8QAUrvW4G/zGfQitECb9f2Byq9z4uuDOb0pEzaE/AWtWtmuSTY/LjXf43jDQ6
lulgWGu86Hyt4f0vDqqOztkFgm8zs7zOTWl3j7Yvz/j8mk1CPf/Io1U9FWgy6CWe
zITRmdOIXF2bAVdBhYa60JeydLs8af5XMNaYf7C7sue9mjdBxr2poXXv5/5pb8de
9+2iJqsi8poGe1GnGhCCK8qsy2LIyQsG3XcJAK/qwojZuSnqpboe3UW4mMv8vCpQ
re051l+dhS9E4Rk4j9rnHHhOap/Dws5r7lADiTc4X8bTl5AK/opnjlH0UOSa2V73
7g3TW2rm1kuh2R31SPcZwb2wQVUWeTtUdZP7qW2p+EwAB2PSrr0wza4H94cs9j58
uOrsywlgqfa4RNkIYD0iMEtLn9ZvhQqNEh1L2bRPLNNi9bceZlnLzu/9QIcqKUOq
S812/+mTu7aGoFd5fxZ+zOw5XJQeW5vXEmIs/2kVmMAxFCD0kz/CMdMFI0IKY3Ia
whflu9dxOl1YblOEOn5mmI0fXFy4xoLtXNCmQhjJVYBL5MStpkJ59Q8/JiMfc9LM
F/6F6eXuUCKxBXllEJS9QkfbWYy5ItaSu0mZxrA2gjm0788sOk+fDOcZHUZ8fgId
kz9SgrzBPpQQA18eg2vpVCG8D/dXboLqv8ltCp5+CNyHCCN43cAl5DoHmBF0IGF1
fwifCNjsWmA0eTiwHcI+iV4mi3OPMCtrMpj6mgmhc5rG3zbOmy6BVJuXMNZTKJvg
ZJFNyGS+NFNCH9Lie8D5Eyvbm9BqvLYg7SM8Tfvzrjvawo2Y+EIBWNOWASYhubKZ
tueNxohjgxsKEBoB8m5N2ay2QTaVka+/0prt2BssPnCxZykR3kD0Bnn1FAccOkzK
svGe8lZjU3W6puSvXYf2ZswvZBuRU4HeWzha4sAEOh0mEZcdtJk9CMoZAIjsqgEA
O06u9xU44x+aCIxc16tQfWIKcZJyjFfm7M3rEWTJzWQQG5k+7bUbpFOrXgfWEF+0
shqYqv9L36DINJjRDOkCIphmTEluiG3c+POZtfN1YBAhIC9Z9mKBjf1r2PlLqxrT
v6/Z9LgWZdRorcJURvyN8CAov23V9HuWDCj70H5yZEfi9mHrOGRFY3j0T266Bw2A
Q2ycuBd2/RZbJ9YFF1/mLErfnk5D4kMTrEXBvI9rvPDmW7MD+HxBkUOiqmpOHwBW
870/rVex9EC4331D9/4zI/HLBFiI44Oc1ZGSE+LAPVjPrDcEs/gSExKFnO+NRjEb
ziWmrRtNPbujHc3EuX+fF/wi7n2gNTJB2qxAXlVFLbV7eJUfQK67Ea61WA75a4nZ
Hw10PFHhaM3mjcGJoeAd2FEIAUdvo0WCd+Yb7iqYBPfbPXlU2IElbrz5H2fGCrvs
sFSBjMpT+YIbSS2Sll/EpnMESnxKBJj7lybI+1VuXSrl4G2jRoMYNQclmvkXUTKu
zjxpmkPtFQfwzbjvoA8yD7UtUBc65xuQ8/FHbMlu4nTznFJvBxojtMN99QHPVIra
LyryGdF7nf4bVwt30lRvKRxy+xZ3R84MrGDfWiZRvVZh5qjlcRCZT7OlRyNC73YB
8CjeLBdkgur0sJNcdzgblSJUsMekc41aRAIlHLDRp9/06rwSFRgvwqW2ng/iwSy4
ZIkLxlA9umay6s4ni0KnImfPFX+6TAR71hzvAi5sdKUuKf6bLLqxxjyE8lEK6YBR
rYghWM2pYp3ZrqL1UTUfvXxLaW9CXF8KAV7jdy5Yzwwp2WzxKyqwuYJTczLUpgas
2zdgMrRWVY7uIcowHhbkHYvXJxvMY29fyNRLkKre+uq8uVsJqxBiIBGj+RDmpX9j
e3Qpg4BcR5zUohLbu0Lrzlm14bjxTkic9g2l+KcF/lKnhEbSAWffu79Xdp2+PUEj
Dt4C1xi8zNk0Wn9WSd5iNVD0/AJK++cKBNfxmpcU/wBBgEwv/ZV/MGrhBI2B73Cx
Rv6Aocj+eiADLcoc+v/s/GBq6Sh66fkQK+cqcKNwBAjQGAR2ReUJ49WXCr+vwvyV
OBBv4+bV19y+5xrnmmh7cwlXmLHcCxRlVYeSmwAPvdzOio1jmN/ekaxgOB4jupsJ
nJi+stOT9XiJGD4WR0R2Y2bU6+mAAvcpgdNKrts0gTXrg8hXA1y8YtHLiMgV6B45
62kR7vpe5spBmJ7jt/xkUt9P449I1LsmDJrr5eY1MvvP4IkJpIw7HM9TAltLJROE
4n+CR+1Qtw9HdBC6WYrK2zAdEKEa+s2XTiSyj+evl9HSOdWx9kAqZO+WCadEAKyZ
x3zL4p7D6zVVuASa0R2dxBgw7dGOHIYgtcblY9Wt/tobR8a7pPXwmmzNRc7Hx3gw
b0r6w0mzYKE6+wcY4p2jraHxTt/WT/qERHFKJtpyQLGratr9DS4j/dqZkm61iOr2
I28NDqtJ7bM95bcBpviq0ypfbhgRjvXaol25EJCEizADESdB5x84VVDLzB0Gh14U
y39mgoJZ6HtPGcgpH+sJFlDHyoElw2iKZHPsFVccpvH9KqLI03a2wEvWMqC7wtgw
TBghi7BTARd82/J5M3PY5BbswBMMaoHC9u1oYMTdqzcuPZpj6nIL1iOI2ayDpdZG
gVdD0Ox/ERrHBRvtBUZRDWelHwO0MWLnkrOgqPj4AhMmGsyMUW5RLaljCjQFyRXd
4a4JU4pkU25CjFyxSXwWkwTU+9bEiEgKgg+g/u68tNbwc8khsIjhmfrC1MGie11b
Blw8jMoS7Kg9kAYFifRmki7WeeYGder1QVm3MFPjRitH3sT5H8T+3fNnUySv1zGZ
qczKGXo06+O0WBcEECui1g/LGac0SuR5C8ZHevgU2rP0L6/XWLHTAI2/3uG+atEi
dxSj9IJb32Z7K4JgW14w0NmgaJYf18sZ69UDg7vcujNf/DCkwMOXES879zEbCYgR
VDXUvyhm09i9bROtXvw5jOidfT7QeXj1rio6mL0gmsCVAiOec6uVpbudhFdwczVV
T5zluIBBockxBodH6MmKQSG2zvc6icOJ0hIxn+V+u2F+PeJCiRYKuE6OMTJKWTLB
Vd2umxujAiiY3A0i+eB7E468vIvAJWDiLllhyEWBj5QON7UIrW5WdBBgI8/zIN7s
AmtWS73Cf2wqPKhHRGawQRFAuANul7ZM/1aqkgTeEuWV/NtQkAVrA+DWbzWhVhhZ
mx0/xE+P/7+c48mUSFsaJkb9dR0Dfb0YoQSI5QWDu9o2Gpo3BnxwI+gwb/Gi/P5f
lRDgL5JGlto31TqA/fZbP5NcjZopV2vXqk6ikWEdVvBxgPA5/UEMLNJyy9kJjTK1
6nux+efb5YxfeiVTFyV5bFliyLdsm6+2tn1BGeqL5hhd2B22zqm6YJNb+ZE7bUdF
37mBmch7cfkdtHfB5UQMRM+bBHLXPM58rpSWnkE9A+1h0zqC46k1FSFXQ8k60eSQ
QpmTy2Sm/Nd1qxli2snxQsvUAgKM0lIu83eZyoiR1HPvhaHbe/+MakEgaB5U3Uzi
V2nd2DIVD/lSsoWVy1rju08xNXjJ9bvbbL2O/jeSFFSiyu6xznLiowLWCdlOfu4e
/FuwRPKWvXOFe4i1hkf4Wp8TJ5DzRhZxCiRIn2ElEO2Pclt9oFz0XeuoZHO+0dTp
tGPezGKIup1CpOJUe3FPKiv+BEtQBhqYnvLrWfkEH/QjF3DH2iTtR0b6FK6EjymN
prI4qUG5EWr5cuzcn5xHNfIBTZdvpU5RfKVdAwIz5lXAZWxsULy5gJyGKQOoSvCv
2TnKJd/dfv6FXFXlS6oz2XLEa1yo117HdxZ743r7Z974LLffOiJ0cQ1/DQ/CJyLY
Z8U6Mos9CVQqyzoVXgua7nOEPod8KxNT4RqceI0vcR7RSKPHaOHQfDxcLWnwc/Bu
f98lqVK8QQWXO3o7EUh5CYsDCiIHpYNp1iC2zOmPWw/pPdjXi7bd5XkIa0gEj0ZA
qZgLDI/czLFeBbNMWLVRWhx58Z9LqV+PhFT+OzrSgQVF1SjHbgCXWZTuMOIYckcM
grMwFBEVDVdQdhCmYDGvO2x6vsmfgdWBHFOuGEoPFt9bGYGE20FmUFJN2CMOjqAz
bbrZV0hh2I7CHDWFyUlQ1IediPiNyNSSwYA7piTTrW+TOMNHmWS1TTznyHQyJXXw
DsxSg9bMMM14011HogXvya+zRdWQHcXm0FZCDPQkA5lukw8hQcGL37Xld6Yil8AO
EmhbfzmjtCMwIDaTqtlvBhV8fhyHA5tAII4zkG8D9lJJRMRYENd3dI4RfvHIQ7Bb
ucEEjD8m071ByUEm93g0Nw9sofCKZhotA7MmwyhsNaAxZooWj9FguUCi+c69yjg0
23+Rwn/DFWVa7si0fMgGTUvklcLTNkaifzYYxkw8hMA/3FPsc6Ylsw6RA6DGt/4m
6nBGh76EesjiCQjEoVsxmH7vcXxWrqNPUBIgVj5eihGK8Js8DVHdOZDm8xHuPKGT
DM9z2DQv6Yw5lTMoZUyBLZTjZ6QL17qW0105FbxBjIlsumgj5zl8hhJNzykn96HZ
AIQR5w+6O1LhHcQlEhTApFESorm7OXznUTYmdB2sYmua89Gwn9ZjtwdAU08dlaG1
g4vfJVAxXAUPnj5k2lkVwfRIfJ+bDnfJhQG75WAIB0CpDuf9J6jqGgoBZgRT1IyW
8rTAaHtfOF1s/gQbRUjix4KzMztYjiNqTZlIoBkY2L1H76TsuOh1VABqZfijGWuT
MiVEMrJlCHAQnJvcDThlgnbXs4dzydJ/ZWLaX1cenhQvRyEYXNSslR+nmL873+SL
0rIYqk4Zh38dYAwQIA1hWkEZ7ZI6FyzQb7M8Nmf6L02/JDY+2LxPc8Mmd7vgmtG5
mdvytGvAXew/bteS3t2m4J+Xr2CPvJ5dugiILkUbKiPGXO5EQh21BHBpjj+MKFpy
gpgUUs4S7A24XJeyn0UVbBkSezXoPBwYOVsrziohtmS4djybySjl35J89RSAGzMO
2/K0a+L/N79ZuAIOHpyTLB3RQfG1Gj4FObYRiuYW8Ecu78N59YdqOpO++95w8KuF
3IcCJTgXG99VTTa4yXS/TFpFJV+/uO081om0EmiixpNsjTghHh98TlOU1MPe0vXk
X4ZRM0cdQozQGJeLfEt36ZQXy9OVnuHuDnrJClo25LkjFbZY2e1R5eyyszQhYAly
cwd7IHMv39eDZTq6/q++V9Qt8+MmEVolQdDWxVuRwTksy7MIyGoA7gG5KErG2sG0
Z7AnDsnsS8LmdSAUjpaatW3Nb97J5ZP29NFA/r9rkdU2FGnQxrOVLLAJBNWEfczf
1dfWCloRfwz6Z7/7MkHPpLF7W2tUmROH8QDh9c6TU0vDaWn9dqF6PdhdNknkIoii
pKRh3zUrAiKpaOtSnCR9jFSBwZpquntwBU4/6b65J7c8gj+FdMh7zVwO1CTKvsVL
KccXs6Qh8I2y0ln2qv3W8FQshMsw4S191gUspcwDQD+QUWXpCHEyPOTztbJo9DYg
erCtdhH8zuH9T0ppglK1OYj79wXdcovh3gE/iQ2xx5YVLOiX5H36dcEgrX+u5jt2
AzDSvwV9vjhcDEPSVDP70l9vKguqMqreynlmtt76siEIa1ULqq+EAE0jXCB5wcVR
JQ0Ztb7vyJ5sAnCAw1tNTnhRL+GvFJ5MNB4U5EvWoOFLE1JlK9zEEuVWtqQJNDRv
SY2ii+qwrX3ws7sCCMvho2w40XL6TKEvfrqAm0xC/YPIwoe67bqhjYGWjinnZv7e
OuVWy2uhqFcs5J8a0vInyR4EZYhP1/HBLab5mtUwgHYeFpkve0k/MvW5Sc16A23j
Ii1OMxPNTFer5t/hgb5M19MkvVkE4+MJ0693Uik0kUkfZrVRSFeNW06cXXxwudcc
FeKn5xrU2kF6Ur9YZzpGTryuSJzRVNrSx7TI/Io5PHW0+eMcz1MDAD67pD3G6B2k
qhZbtegng+lnDbdf1NclD8mUVV+3UCpNgkhs7g64xjCxTnHKCvmqzFmnpaEMUwxj
tse3pGSPNvNB0OcrIASteXkTXn01MYptGj47EQkd71AXsan+cMzNpFkZFuPG6DHg
CgNLVdIDtjPdYIYFoPKoWot9ZNXWxmaJ3j+sxqzo5Zl/NiIfW6qb0C5+R53rHAXE
RVM0qeDSyxQRKIX2JUosX2cJUWHF9f0toBe8wcKjliCwfAuzhYrwLNcBXxjXPrvp
uEtBI/EYQNZlv48kS9rdU0vByKytAcqCyqGSrScuCvYFIzTjFWEKlnBrIgEjB78a
vw5CBnQo+C1KMdTgMGFq9tFfdmV4n7tzWNay2eFW0ldrbRmfh9OIjenKfHYGaGor
SbEyYHPAJl8CJh0a8L1+rsASuq2Szszq+Mydlcgl6TC2cb3jt2RYR+zX8W55C6Uk
XRi+Pi18QU2czPUUA2z3hZXuVDSmhLDU0s23qAyx2H/JtFZGAEdhSy5c9oLuNrXO
ze0maqhZudcJr/87hn1i64rRLJTuHeQ9VbNhaVCoD/hSbZMRbWMrlO4m1N6EdTU7
mIX2ihJqIbCkSPq6k0FLBVDUzOQ5gVJdnXZQ73CM8jxol/UvfpvC4SkWa/OPH+/I
PL+7+wE2BzOsBpRahPKeQBFNZO9395LVpZdGVe3NRAzueV5VKx5w2ReJSSNvY0Rc
lpRf7BJx1LK1cA6QcvSRQvyKIXG19OAW1VBHsmM814qNtfTl59aBPIRN2iPjHXuu
oOSEOu43r5KIoOLyPGfsWGgXUqur17xOf9YSI5Agp7raW/huRxRGTMMa4ZfA4PUA
r/QSxZKg5q+yQcHz7zKMsMoZgaYthQSHZlETwFAjR9toHfeX/nXxOysWprWIgZub
sQVA0jK+A+LNb+AH/Kg/SxuXYiovdjUdBvqBKQWV5RbBO4ldGUPKWOkyQhi4P2mY
x3C1N1hga7jEwpvwkZos2uZWlVqaeRA6jSqLfGqP2rhzSfwJbDpxI3q0JOQb1551
lbCeJ9mW7a4TvwUBE2Hz0JhC1UST9Xt+84P09uN+J+LUxsyiWwfh2cmt29gl7CVn
KZ9DTil5vo0VOEshRdDEvfW2UDtnaUFlGXW/STjAxVODK5qhQohCSQY7ZqsnLBjJ
q5II1kZtKY4S6EbcSmMF8JqvJv08BwTROfriuYQW8yK4TiedSvtJwcOwRY5C1rCh
We3vCiA0Pc7P2jupjdRxo6mIre2IB/+SiSx5+YMF4V6l7kvkeMW3rPvmpjNdGH4i
GYkC3LeEjX5TKJ4r48xOhpnwix1ho15ToO7680C1PKmudnGE2wyrF89X31s5+b48
rvqMhcb9FH0V0dA5V/uHrqEAjFEsgoTV+ECsKOAZVHwMpQRI9u6lTlpGraaDhW3E
nx5q3fZHd88ZZR9AwBBGX5BXf2RMXcX2mTzCDXVqkqzl9heSYoCsRxVZmgSGg6Rg
H5VRF3D9z3cfELVdSxd1l0/oB4mPo4ntO3889G+c5GZ46eynT9S1lUJooeyGBfAD
cPWkf+UgV6NOILmayVrKC2OwH+UTch6AQ1CgLQzcjI2u5yzc8OZymWODlAbxov05
qD76oloWXNXz6CnLkwaujLap0CEy/Cik5Thik0n2iUwoAWg+dDvpDVKGK34ArjPU
CqXziqWR70EUKGbbWUwGPvUstk2wYDy0/Phh2QAlADiJNCNqQ1D32+1H3CKatXwl
aRlzN5GWqmJVa5zlr30lITYSuU9AucnxH6mD79E8ZsZHCt0yfNq+Pl5fAsmDnlJg
8rd+59+zIru4WrIXSIOOOCsnoq52yoU7Sx8tzemTWLB4nPAUKiMRu/LdbHMZfpm0
EcveuBKbwNDWohsC2js/5EZfcE1s5gXKZzFZA14vvRLLq9g+jIZJrmxiTOjYK5ov
yVsH2Qhhxg82uGMIFCbXT87oHO1a9RNX9G/xXs405tUTwuIGaypTMCgxahQtFwMc
6SeNR8CPZkRlmxanFmCPyxcSI12kxIlgUDTmiZRQcV3k6jT49/xVzzcGZFIpiIK0
C7lUf4dXjvX026kAz8GxPl5zfGNSMPATtsX+zNgtwg1XQ3KpqdgfhX2fSV0EaYTa
3eWHQM5czXpF4VwoYRSxQ1lvb3V+a4vx4WxR31delH53mozGqXJVcyygerENbHf1
PcvDPIugRumqcW5yHdF49G7VNW0hmXtmgc/OTUBbWJkkNj/2UMIUsGwk6cf9t3UP
i1xB5lVA9o7P0Xs5/dx7VD6mSxrEsEGJ9ZtoMDDa8s/txtWeCFqqQAnXgGe5NYlO
o9DPm2bYVYY8UopfeqlY5Uj2p6XJMrpyam6HKDw2QTjz/2c5roReqwKDNfWVU/9A
giW0OeN8chpemeH6+bBOZoj4fUNi0LZQTPD1EcrD2DWWVdDchUuluqs1zhsb8QS2
x2aJrXDMu4roNr71QYai685uN/LHVU08MMZDWgz869KEZ0sRscoXAK9xq+g0vcPZ
R5C2v1YsqJIgpls6APQJFsfITOJo66K0xFn6/rI7eSlxFqzHVoDVpkCUqihEkKoV
fVXEUyuU39t+ErhaWvbnDo0silaWcJnm/X+8n6BDE0VwXrPCG+IigDxtPwO0D60s
EWxP6YHCvaug0KyH82RNRvIJ/T1glujbIXHZIWxlIukKWJldTSOrGx/747bVSgDR
69/wslNXprw5bj2vtk+M0remiQVBi8PwcIsVft9mltoCWSa3K5tO0m4YDGslJvGU
8/3bsZJVNTeEcigo9GFZ+cuxZXx2iAJNnmiJG00F/VKFLSw1x7wmq4zt/5t12wyS
MKrXR4aegCcblwK5fUA2ny+Hk8wG9alfaY8FvoDcRbLCJF/Jl+qtx1ZF6qFwkIRC
IuFPLQhN9od3wL2VdOlzy7WRzDNzmP/tM3nfpO6x2Q8M2yXQNplow7zRYbQZGEUs
/5dGXxpsQG4qMCaMywnb3FK1NrPQCnKVUpOLmlOawdo04VkTAfpnJS1Uwrh1loRn
8j1XIZBiRwt+TEh7NfS+EV4+TogBcuiYje/cWgzyP5ASRcOVxwKIitK434V8iteu
EOOvqD4RgPRoJH5NPVCrTxK7JkLwpXA9inJ4D4nkJZ6oFg6/04eCm8AmIR6HKRFS
4WKi/4Ps0E/3QqvW0P3cqYjlEDTwUfJ8A9g8u6HweKspAeEXJzxkZjTD5xTWl+Fe
fm6PC5Dk0RJelqzQYgyq+0+xkC9O8RyJAAPBT1sV5ARIc+bf4DWU5ytM8m2EqA1M
XXOO54Nk2Tqe2rDn+O4O/nBZdfLFhqNhdThyMW0FLjPdvIQA0f560zsbmSgyg4od
Ks79izyI140WtEzZfAERl54VS2xUGd/StBSsupJG/YYOICA9B0+IzhvXWP5Jnsla
ebaUod0YPSxSep9b8Hpp9+uZ7RDkw9N/W2pDoZ69MKNX3j7GvnDcgCPSI7baAeGt
wfODmKqy3CBuzYihefT2tJ9IU8d5x2QgH2FcEC/yKXJSmTh574Sc7xlTy+48HqHt
weGFjUAuczLCwuPxhBzWfNQLJ6kxlAmU4uWdifi3/rT/xYoe8zPDX16Z1ECjvMM2
gHt+dfq18mXfWB5DTsqQ0c5GWLAz6fE6ciAKhXr4xQsUSovUCHenw77M6M1V/ji8
NONKyBO47WQNXgoyWrZEZ1Y3SofSRVIV8GS+A5fqcOhc/sFRz52jENysH+3WixqU
JEDKhe6zyiObb4TxzlF/IWwtr5bRAYhWwDIV2PoUzRpAeHXHX653yK4XO4+AKOBA
wyu2mfirOMeAsBfXpXnyNSk+UQJ+uo778VXYeeMzCZGf8y3wSGBD9X0s1yFodZrb
rzcwFBPIvO2gDE6ywWDaeC+ZeVMZg+2ya/rS7zz12PGiBXdGdfuWUUEjM+RnCp83
ThHYFDLYx80ZF1hIl5Rn7QSdTXRNQkhnCsR3fgOZOXlTV+n4HtQai/YFZGkABHBP
seIc0W1EsA97PNtDrT/1J7uI1LWamI7cRdPxwxHsm4oMCohHHAVZspExH4BsPr8i
nF3lGcywxVA7zDgtDxXLhrlDCm1/hciAigjMW8eO3l2f7WyFkPaNJhaneWenaGCC
kJKELV2Pf2qV76k993/c4FdFrbH4eDjK/XZ+04TkDtEq/Pv3eWwzfEo1wroj+AP3
JlVlujPqWvWLpZukcOdOtBSDZ7IW6v6R7B61b1j7hjxulhdr/FWtyjk0TxL7Lzjf
bkUiMQTC69mVpfB7EqfSeIu6ljrxVJaG88D8C0In9ck5bfOF01zq6m8VNld4ed0X
pQvSerVM0aAip7pm1WRRL4k2VP6OLGCSsDtG1DpVu5wyZc9Sxj+rmq/qDA18z1HZ
wrF5KrXXoxSeGA0cuNzvFP2+KTGLEGcAEMSvikcLtIHOoLLHc93QB3wWuQqZItbo
gUdqovF9G6Qp1KJ/zmmx6zJxXukfBMb0X8YGPdol7VeNYxjuclgWSBKyzy8fwTH3
mWEFs/RZcHvLLPoVVmwUzIIZmAl7YKcL+A6WBeHrd27ZjcO9As3LdRHqPf+oYm6U
LjpV4erTkkcShYXB9PNJk4/JubMiyLNo9yJeai+8oF8CBBuV+vs4HdmteKlAcwED
3sYnKAGr/ITwvw71ZcddLnIO4lQz2u7Z7Ae9QXNc6wRjXK2Yio+NKHxpgdkuHyUK
ThfD1FYMmDJXeIOBEEOSvNE6wuFfzpdbELjurik/qe4ZaqsmgXzQMXZZuYQxaHBh
EXltfrbJy1DdK88lLS8doDMuPIIhTitrk2ZW31iVd3sYqqOeTM8Sogj+otl6fc9P
k1vLwbBMgpuhzNv6U5J3aIaFhXZIhOriQck7gqs41AdFQoaNMQl6Vqdd3XyVcyae
rYXwdVxqaSzXKguAhpXNiYBDa33Efk5AO4E9pXvdOFtL38GDNtOdlg4bK2Y80kkl
jBCRkyrVZu50gb6EbIIajyafvs0IWFI/2j2NIsX4eZBQ7BGa75/Mk6p03Pjcrdfq
UhcPuH6CfCP9aXfXqfXHDeptM68GEXyKRtyQRAKWqW+0M78vl3GwFqwb1lzzD72f
8KNxSjSgr5skvgFfzFvU0lHd+moWJ2x3aKRsx/EjInW5ENjPvIBNu1oGLd1h5s4f
ecctANe4hUPoIf7aNBzCqJ+PYJfQwh+qZL+yAxGSjqzdA0lVpreJc4h0GAja5RvZ
mkq/ixq3TG44JZy9oKVr//++1l7UzPyVbE4tkN+Lmk3LNq1QkEMxKsPb6VUaruak
XCy1wxsFXatcifss44Y0s5zHziJfXmCqgvZpc55y4WUzUwqfB7y4ZDW3FzUxyqcg
QQv5kIDugR3E26zJrj4+A76+X4ogRy9WYuZxUxOP6loxPoZX5ah8u3tb61se28Wq
la4qk0ir8/NDoSGOKRwWbMJMDb5N1XVnJQ3O8EdRXUTjFFGLCCYO1ZsaPdJwcX7y
bAeojEe+A7cEvrxFLs2xdbDMmUBabFDNno+w4ap+uhptDDBGFphlQYLs24NoG/xX
SBHwPO/zbVw6IjbEf6PX35amdkU+fgdTZAVrextIS9kPH+TAq73c4lGVbpBkz4Bg
AduBNW7Ug+Xi1dQuiCm8barbZqeyebdZCXTdZVbnGzYeTufJcOZmKyt54UtBiicv
ApOqOpBQJIJ3hVMNqYehWNCN6J5BLe3MQ15Er3q+8jp3QeSoCp7SBgDLZLMFxdx/
fcfrco/93m2EIA1T2vtNYTa/klK/Oj50B632ve2R0rkle4rFp91BLhCVyRNDZfKc
dYzm2vcYs+3K4UigsbXKvFgxa2oDpTPINrrHt6tZdRR7Yjrs32Xh+V7LwltmGsdQ
MB1wdrjS4a3HymMk+Wd7wkzfrJqAzkKxv0yxz11U7vXlIOC5Ce+oVe7PuEOcubGS
M+LfYiu1osVSBmjCNwwqp3O+qq/UUJhqyFL1drYmq8WmckDQ5Vwsj/lcVOLF4S0y
a8AMw36SLBTZZg4kcaiuYKk+0Gdmt6c9ZZcPpM/QNP2sxiGvewpchG2q/UBN6Nrc
pwrEsgjiwfPSYPIh8Yk4VqqGKk+3a27fswAfvonp6Rzr/+l1W5qV/lFWIx0J8GKN
Cv0xqbsM49PUEplXWPmJpvPW4n9n5a3qKMlJg5K/WAsghkTzd5RJR1lwlMcQP0n9
OZmqCbJjAlELQ2T/WE/IKF1YWhvbiRgbOlRvM+9Waa8QA/a3AZcyH8dFpHJnRmBu
XiYel3d7OXTga6mCbSXryqa0rFaVYcCML8MJMCQZh7xy83Npxc2Uf8OyQeKt2iXf
KTJEi7sRQ06JiIwzuInQjGEsmgsWh90FbVx0VwHLhJq9zYFyvGA9Asfy/YqxDRHD
hwJTJ7iBu3ueKBVx07W2/FW5cSSZIT1X4GUDRlY8Ei6TDQKMsRW2te9KoRNtnTkO
OmcWDM5QwH7MJrm+S3DEQw==
`pragma protect end_protected
