// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pAesvCR9LHxOI78s9HF7+cE9WOdHi1YsR/3yKqoDu1+CgElGpLZWyT+2ZCwEehvQ
jx4WJTKhZ6g8EE0e6jhrmNhrat3p++vb1edKAYXeQlGQYyCn40n3G1s4RkSZTfZ8
no4f35TcxEEh5pOlx9+yGJmvOsM4W6axMgzFhdOLROw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 88720)
JtPUEvtIM87R6G5egKtHmwEDF6/X32w8XYZI+fwCcbzS5S9hmCRA2Dq0hNe3h8wx
S62E9wdHCpCxvEgIoaHQB59yOZK8N47WaeAjkkLtxwKrsReUpRCOxybhlZpdfp1F
CP+/tJgKk+chLlJSINgf0bL8nDpfUIm+iPoxoGcDLzHsQ0+XcSsZQ2Xb+TZBh1Oo
eeMr6kBMpXjFwYd2h9+mvomU0c9lUbwCDhytuw3MW3rpghTYy1y/1t+ikGj5TIfX
uQSZ8EUlcgZsravCQvvVgjoTQ5apMu1td3WwU+Mrve2NkoLSV+gF0mpTt08tZoeh
x1tv5VPSbGFr11j2sOk/kGz8WCdyAon+SPCy3UEimLWX1h1mZj+Fl5khP2Ss1tY0
i+viLTxCmYNq7UDBwSe6Nhjjv24iGGsuekVpybu3wN2OfWFCfhPWvwmVXqw3lK2n
YfJiXYhhhr9WSFxvGjU+3ssANgA1I7Op8T5DNKRZHaLcT3nee25ChIWodrtPL1GI
DNMeAwyQ1pC3F60437Jl7DuU097aPukBxpjqww2E2SqLvlFSaFHz5o3YLngwujuC
8FTEKFP8D/heSd1EJO+oYMCSpxzGieUNu5NWvqAIepYDrvQ23p/D6CbMM2UzpIic
/LNa7a33ruHPuOkdyjEsjwPvi84sGLjusN063ACtdBI4pIcjjT5inldf0U3QcD3+
8ePMtLb0kqpJf12TXnCUZd7dZ2Rx+l/dYFOv1iBTnh7bB6T34ABaBSQbnWUbopsb
+00PWb13HLgSOq3kXNmDkQJHb69yqLLKMC1a0ACdbKcwTPJmcymOc3F0YHi7Wvvo
M++vtzZtRZDbVkTM/kupJaGdhO2YoOQ+fifNkgad1vQH+04RutxVlFSqNMkiYqmY
GHP4NRWUSgiOApysONjPNcUZfRC0/Vl27MH98JRgnmC2Bf1REbC4hdLBlBXJslY7
c5gZnnyl43VTy47AmbLqXYE3z3YktRGvkxCX54P+kfWrtM48Ud1rzuFvuyKO37Ru
2mYK6V4/2HGWr+i8k6JYrp7bhJsNfQj0dgFeQoXBr1JB4GJ7rf3GWsQNU8NLovHg
G2Vf4kTvXkFGM+S+l5bI4TT9dNk+3+YPz+XhQpyKH50qFUVSoyQ97mAidVyvFxRi
oUQGnSeisTw9D67SoEGxzOIToTPK528OSN99apL7iKPp4K704L7nC5pNKkDQmNkW
BTWXPc0H0K06B3MZc2cYASgMM8SZRklRI9DLqTGjhZxsn59Zie6TwtMWbzDd3juC
vLC275hWHs6FUAbFq0vXX/GNuNlcBzLVdCz9btTJAIHSEGVvk+UYcNlBDH+AQ6T9
WALRF3lJ/9khh5IUhUZZv20V7dxVSZy2VjboLfPeQBrrBTtbbHaQZ6ImIneTFDnQ
vjhcixsm8Wxl3sL1DMBQGclGCTnFon8XmN4qX/ySHxP7jWiakvEXhguZtXbBMQ0U
k2jcLVAjCFghNFoq2cRfn3wjoxlIhHy1hQ95C5ixqhjh2l0/JT6aqUgtkZuxT23x
RGOINGbEnVrtGhPnVK6d7ts5dS9K1noIiE1MZg1KrWoEQcTII2W1Qw4P3h8xLGn9
59mcdWw27h6C19qFB70HlzvLXrYoq6epn283lUvgE0HLNQ7oIHobg3ABW8E9FkYJ
1xCvH70BCscpovUxF8W0nw+x/SGhHAn82T73+4QaXkC68N+7wzuaEmNZlQqmVsbm
BVXMv73jh9qpJowvatzfSZaZM4t+IlsV3nNDVnFI1Sp8gLD/+fDvYBnUGa6g2uZa
84NoAQwEzUtxlyKMfIdGf7J78SGIBgd5SVNwUGCRDO0E6C2eTMsN49IJz78lpayT
z8/44XV4fDytslMBzQtaJBRd56STkFk5iFTWQRD9OQOrNiIAHR7sOHvHdVx3LVE6
z4AfsHPl/o5xXDcZu+Hjo57sHNsMozAWhPeMRXjtj2DPKosgMMWxiLUSeXYo5wnK
I4lIC2NOhGbXckCbGGj1640r90vto4bk6AMm/3eC1BQ++QqMQ/g8Ejtpy7eMfTK0
EnVEobjljj7ll7sCzx30r9cxvgNZGnPi69Is9SC13mRPpTXJna7JHzPnFvn42Uto
Ge2CbTeiGXXBVZq1R5RcBNs7y24Ec3oYkPMYa2em+npXFUnvbciiDmS6cE+IAJl+
+KTK96+O+6u/twbUfEaEn13LSmklcTN0/MlLU0GqzPTrkq9PgrbT7Vgnw16CVwMa
x/hg9F2x+7+llbWVWSv25nnWIaHN26dDrUIzUWdRvUqwQKJWdrpx/UCafx8EShK9
8f9kka2Fcc2qWR6/RdckEadApkdF85d5xwsYySYqrD0Io7lUT7JTLT0A7IZ82GtB
rpJ3xSdk483pK7PWh2YuuWv5qf6B6JCTYAtTS8Rk+rHfEq3L0NLGCoMwGzD2xXCR
+mcFczkcxnRDY/JrkFvIIrOGDwLCpb/WD5IlVqbR6DNKV3gz1idwrwWL/InVRRAV
U4nuNW75268116IrupM4FKtxwxC/tELQQGCzT6HRoQGs4+oz+dcN7KN+fMRSdlCp
5Hd4C/giwQLZqkr3OxycPv/LcXQeHT5fjRpGtNl49KMpvUfI86CSRVCLByZjzVRL
9bBCYHJdZkBWinK0tJXWIs3GgdMQiOZF7SD465khaWDxJfQ73az5pvmwmlGbxnho
wtAnAq2NYetaB4c+N9DBSbOy/luERTnrF7exzZrQD05SPQPqStxy68di4Ve6HYSE
8shFBXk1yJca+o/cNYXAbtoawKtG8DEVhW0OBzJ0ZQqurYCp2sKR5sByYggfdT/I
jhnNJlE4Lq+HJCmzqxNc7P64fgMPEc9i1zAlD6ImrBhUPRyHNbtDvnCbvqvaEgZg
Ck5LcIFj4RkIgle8Kfwen6kN87HYzyHuBN+cX4CNt/9VXV3MAllx5gLCN6wpPos1
GTWgjtUGXu2rAma7/Di3JjPoO11/t/bwIufnqjhi9GP0jaSeu4xViUZHhh+ZcWm+
sqxZIab5OKX6g/yaPAsJS915IDPFlriYzbIxY/Q2eLsYOE0BtLM0xfW5ahWyGcuT
RQw/TA3Abxb5m9za40BDTG094cNMibw1uYsLeiPngOlWDQSgA+5yeLASz6IlNxRi
VGMSRlFFxdmAHWK25A6KmxssCf1Cf+l+FxqBIeQlKV/5mnaYnUVl8+KJLltzD8zD
PzBh1i91FcR4iHkTx8qis93Kc3fOzbeP5CaM+hD4w9Xkoc3fOraSShL/2vpvnmzk
3bMnxXcIeloU+Xk0JNoqDKb/TPZenm2jaXeS6IsLZdw+GfQKSxXkTh4FDYaznVSW
IaL4MKzs6c9UdYPyOPXjGD/wroIrooMimc5X41vmq+wA1xSGHrW1NjVohemzKcyM
YRDihn3y5F1NDCm0enALJiHkfTi9G7Uiw63wrMP0a4NwY4xOLHMee1vP8Ygz05cL
5AItYE3bcp6TQ7lr9SWQbEwQZO5xa+KrHdJDC0rLgCByADId7Fb+fs9e9Q774ZAS
yDQLESqtafYRNbS2e4+lFV3bswLf2Enbw7vLyuYb8G3mAY6zNDnl0ZsouuCLe1YN
VLlxv6nC73rwcsOPihZBRbLsbgJcwoPnLRrKnfVYNHeWRqg1XXKq6MzKR9ViGfx+
QDRGZudxxv7vY0zOBXqGDxSiPQrLqqplututtKdfwqP2Teb8nSMATIeHdUnPYNpW
RQkQnw3MIR+oNpN+tOP4sG/sHAZtyPU+ow+7/lyviuYssXk1I3OqhQnEyaCGHM8B
ZwkVcNAC127c/NE/Xl3LctUM70ZY8UQt4497kpaUYFgei+SKY9giQ096/XZnNipA
+gtTbzK6FExJ9gjjh4IP+1yl1H0vIT9HjKopRovlPFrjRy7FkafSfffboOmA53PG
5VELTs6Dm4yurjWyXLAUD/nCGFG4IS4JfZsQk3u5WGbbzZFrQj1/c7yVN2eIevND
4IE1zJzwNWEs113EdsOLMAUXAWa0yn4nG/6t4lUIViMp7MbC5BeXCPV/Y9mlznwj
Es8UCwM0R6NaKSA7fsrwPCN9Zk35USzoM2a2y3Q+X/F1NjfshMwLW8yaH3bwztww
lxtU0Dt9f/NvVWpVqSDMhpDdtioTyZzEXUp4YETWD3j2vDSoVF6OIKkXWfJLFO3Q
bJXsiDBx3T4POcyuxb4VqnQPE3E6UZcQbJ4l61Z3ktRbKgk+n6YKngV8znCclZ6l
Yaye61YUIwOmeHOGCcccunMcOyzSE0abx/rEzL+vjIYT3PHtflQMUMPPt6w8GN4O
2Z8hFYJhR4JxahcvwHCPWJjhs7Y+n5Jxj9X2c/6hSgGNsn71dN3PeaTX4J4NiG22
Bd73IVZuBS4IRe1+Upl4BPxIxTPeYu6RaPprC7ulU4xEsMcalBZaS3kFpcyBFSgL
8FMd7IalCwRohXW5wdywSKRFIeU1h1S+p02vPKLfaqejpR8Q3KYu0Xr5Le/7531P
8QnUCSje4+Nb1RS8zKy9N1B1F8oXmL18aMUL5iJygCbhjq7DqBIIFz6d1OUDP6Tq
kJktzNHT6dbS3Ogay8/4uzvSqilRXDRIHnzpFSChLUddenGo+u1QnDwlDjn25G/z
UeZUNs67r9LIRwIC3J65P2IAI9LZILHi/kgVhnoC64EeGELC7pMb2vky+mJgEfPV
3U0hn04vTGEDg/k1Q/xtosw2FMYPC8sXmDm7UxN4kM2SCdqCj0V+YQ2aTY9Gn/es
ytnsNAkQI0H6rfMUZN/UaHC7et+HCMczc/via5B/OA8QxcN+DBKAhYf8hIvirztB
VQaPa954aVp4lCmDU8bvXtfaniTmolpT0kpLI4cHQ/61bpPlTXZuT6NdovgYn8Mz
fDlvnlor5rSTN0BrXmrIr+fpc2FG2xZCDm9rt68Dg2Pgorf9DjdoHBPpkLBvRDup
W8DoG3uNAwy3LKQkaEyWwvh86gHqRFm8ietg96celFg3AsNzIDLxkFgshEBMhTP+
MNEieFs8ixhXDDf3ED7kOXwxpqJ6Bx0wudREa1GJylTQC6x0XY489dNA5rig8juM
bLBVshNKKt0j3OFTj89XmG9pH/IKHGStXtAg9oU7SqigL8wi5uC4TDd2PCCJIbYB
peonjwQTYQ8rBy0Uluui2wzZ6LcvIL25er+G3hZLmS/ylvFIFQFyvOkj8OxstspH
/Ww0mr+vPyjCKHhm16wKMlkwfhOmQO3LGR/qcHRxWeifY/Rc1k2TZnHdcVZGJaic
Bvp+qb7DkV5dnqoeXQYboGj+M8nWbIZWjoQeMJ2MC5InBAUsBTO1T82981IQf/Tq
tl41PanFON1o/ihTUiBpXNj0K1EGmRx74BhYZa/WdtdZtfVT9WJLhSmEILVtT2OD
WrLejH60O5t4tukxoRltydhkuALu5jLybIpLPzNBD/xQcHsTK5O7OgHj2zO+mWmN
sIPCCxcHbj6rvtLdf8NIrIeDY1MTfJ8cb9+WcR2nrcR94x5kUDwhqlrC4xrnDb2h
qldKeYzrNX3kHFSIgaOA1ExvFzSnxjZmhFe0V8frgEEjXHFkLu0/BEVOh2K3L5Eh
0lVqqpYu5aRTPh17klSPAT2Oy/IQQF7hcAbQmoG97tWxWk9I6Gmo1sqaJaLmrP9m
NsuZMRdzj0/eAHaLDspAz76FSeZNYvllbDeHLOSyOmB4gQSB2IZJEhIctRXpE/gs
Lj8dceCaCu8xkL7OFfd+2ksE9YDlaMCOmy0YyE3/ed2gezszX/smEi7Wq3C6j0n6
x+3yJ+SmGvccPtMItEkMGqEbbsyad7kBjHYgXnL8sFygvLaB8gxaFFoaAgyEzqYk
6X0xZOPDlJMouLQaXFoXF8uT33dqirnwvo7wR75o9e2lg2Wf2j/QCW332ORfazou
1RH8khjVUUC3CfeS2e2MjDw7hPyQP9kOGAfJ4kJlUhoRHvEPncoojkPjUR4TWg74
h2HOyp27kUJC7DKzYhczxYc8FthnyfRG1k5YXx/bPs8wn6GqmP8mIszZu3v6k/AW
wXP8b/EbShy0hxBLuxxgTwA+fbHtJijP1mqfwJ9lKA7twQdvR++kw8vLFNbODvYQ
GhYOE+9MEUqVWZZaHOWbjUy+6TUa7jTzFE8SsP/pFu9xE2MIiWllZZuyu1RUDyc7
0KRBtS9eWMNpLkmD3RWdPS58XLOf4XoKGWmDiiAeS1sQqIu94Q/4OvpuAAkHpWJT
ujNV2T9MAA6wQPTN3HTDFpi7lqRaNg6O6MXYpOYzdryWVX/JAtze/tp8vvHuvz5p
HMICKLXFICSsdj8HnosgHZI2QX5YA6o5XcLiXMlcBwH2T1XrHUxLRhVdJnAdgpL6
QFRdY0uEi+u5HRJgDLgDWf8Rq1GPYn584aDqTMSk7apn72BjQVgmodEcGVKL2P+h
4i70HVKqd9YThtbF5QqxxqlqJAczC7hlV7FVfBkUMJ7Vsvuq7HDHnzEDZDsVTXny
SvQzwHTxpW8imsta+8Ip/pP+3W+1BFgi9VMJafkw8IRwkRJ3PtU/9aQdEAHtjcWq
aYWWl96vSirEsCEQUgNZn86GCrqksxFi+7FcscIKbiRE7Ji0WG9Zh0Lvwlf9bjag
6L7Il8fW2XQFnzGfZIlVultSkmSwCuyv6ReQnB5X9FbwM++hCvrAKNEH15U8JgGW
ibxg14Xj/Tdnl2woX3ERqI+ORpyRk3+ht+T7eV6pwAp38Vom3DWrg+33YuBubcc/
D0seowd+98IbGjiN/F7MVU0u4HxHsKQXxAbG20cT+DN/WkcNQ82EYmO+zEe+v5UG
xRE1hbjoeMQACXZ6Ceo5CNSlHt6hDQE9f19y8+d88reU8Q6XvQt7gHtCzsWYH7N7
DP0wlm1QfLkAwy+1y4wItbANYfhw2n1uXbQ9Fj1RIJniYe6veGWjAXaWEha5lRMr
VAVLytt9dy4TxMBJdUsDcFV5YXLjk7zBi8Ha/vwPTKLdpq/pyUr8BXeDSjlUNTq9
CKo9teQig1cYXW+xAYyDpUuaiB0rn7/4oB6czClvwtQcYPN7CfTdOjwUR/DOwzP1
Bqsd5N5tobUp9BeKG1djII71R/GyamPH2fk5IkknjH/aTndTYLFzyemTuMEUnn/t
BriDY5f7wpIvwkeWHPmo8Gq7wBl88Fr7GR4dVp4WYSBz3wmIvYSs1hukbakm4s9A
ZjZzrd9UvwQGm0mFmYGp19UsUIHZy+hDYSG4DQiTQtXSjjwzFFkGlkpasnikK9Fj
1Uf3xNHovoOff4yBD8SjjOBzJhuh0mhHp2KH/gJiMRYQOu2OSCDIw/7/iipwwFWd
iXShiXgd9WsnPbb1TBW7byM6eEPqY7ZW9FhtG1paiHjKJCUXHsnhOHmmRfjuzQW9
jRPry0eiSVeKeVRbBgSHqBGTQ3c4E74CkwJYRI4+vLDB/yWd7STcCFc5NTK4tY6i
SbT6LH4F5Yj2kXR2VxjOe9OQkYNMwZK3xd/zTwKgT1ZNaQxwrSJNrSvYzUoSRLGd
WDWFgCN59uQ9oWLdOwqAgdNO7cglnw3DPJb3syFVzUT/oYqkBqid8rTAjmnWP6b4
vKLytTSbGQtS3ohKaHbRR1psDrwh+31Ae8jzJBXtnOc8KkY+xv32ZbnV+pOXFwRv
BvAaH2N7U6XyGo/MBLf+epn1mKVIc9MqRdJki0CD8sozObTfyA2uWwE0ao7Lre4Q
feAzC8+ONjkr39hwmbQ3C6NSlTJPoUOILvIa/BgJ+qux6+jmTgoBTC8gCRjPKskZ
mgFXuytI5e+tJXFMlJcVAFRy33g4c36mYlRz/4nQDsrXToC42c/NpL8kQdmpBZ2E
IPHAJqhgTG/9uK61vIOjKg2AiDUUmorEMtA5gfvyU7WyaF+jjKynE6jnLav6Yy8s
hV76GMkP43IWmcxiODZ5efqiPibNWDj+vLDsDpt4SbNwcBjxmQ9jCYU3tiPwqcu0
vQSWqpou7kWyP9ssxPz3NP57OzN0teTS6xqJvMs7hSVxAs7rqu2neCk9fvJPHxuo
umM3SXeuSjRe726rcSIQnd1gzgTcBt1pFx4ft0rvjj+MUrtGGyZEVW/8LJfndal0
oUW7w/rufaaYNoFZzffrRgTy8Y+pw7A8Apm4GNFFhHnsVgZ3HW0WdbbcyxV6+Jvi
4RsV0YWAHrbO7Ch/9cP3fmQA0GGP6db8UNZGNKQdjj6puuS4lV28RquJZReGxWRk
yNXWiJQrxzfSnuCRJm+T7izzoI6LisCK30bPkIx2igha5eu29Z7T2x1CE+4HOHeH
vyN2KkkyM5usZ7jw4J1pemXiRg6Jspb5n7EJSc6L/BTlyBVQpMy9qIPjNVHej33s
iYJlqVV/Dtq7KXeBtslzOc0WeWAXbAueauxufeh/ieDjTf03VtQWow5mqH9EYnv8
j2OE9QiY3GE2ySeoiZO1LJjvqWto9O2S9PaxSfi0oPInrKaOChp4uIf88h7YSTmu
y/I9SFrU//f7+cf3P2y6fTocFei1+KOdzRVcGOzO0tXYMLIsAZHBXepcpp4VO3rX
IjUqFpq8qhR8LqDbOuM8HEwnhlGrLrfVefp3kprglnxBQFGMgLkxG6t2eOgWAJ7q
dD1xUZeRqv9AnJZdizWFMti9rd+y1o1JbklrW8Q7b2GsXwJqPtGgh7z9AzxsAule
Prq0mHvDX28+fuzayMERvtv5tVR1SwahOPFOHw+EIbJp93vVvhnLRNTZuz5Wb3jS
sDEK1ruFTQVueUogitV4/fOrD75HXDUExYsqud4Ou1m2kRyho5QTJME86qabohMV
itJ1In6TPd5pNsHG1WBRoYQzxUhCBTy14/3CJxFnQdCqsol/Q7Xp6EpwTD2M3PwI
HHxCMaVYT0R+NCavbnwNtYbv/BpQW/PkQPvrjU2m3nAY2C1okZxMstD3sypsDI2S
S/ECVJP2XqvbuM3pBP8ZdroBJwBGW08xvyXCqhYw/UDr2jcc5q5CNQoN5C5b/SkH
V982oBzpl2p8hbEUdi9xT8xnCXRwUUlN9J2KXob9gp63v1w9VrPBqUU656ZR8CWa
VdYVHcCYygRXYyDvCYEaBnlwTuwRk1Y4/vVfqR9vl6uFhSVWTCnS0r+yAo2KBSIN
Omg6mU4bMvbjgDffkbJ2SDpV5e4WFkhgJdOH0ygS+J2m25wKKPUUdhPTV1cx0WXa
j+iEsL7nlPljure+X0hA/Snr4EkH0ZJldIJ4/I/jOhQSEKwwRujrBBYIL1urstMU
1pqDzu3Fcx61ErOFsz3CC/cjHhRRE4E5z2HuerLk0uTMYsnrFTmYjNV/1V76B4/C
lpLNv20fNsUlfMVwH8fOT7Z32cWRzIVdF4SYge/aXwhdYChSTtU3+XE9PSOtjc4T
34BK22q0Z6PqivyEOifGFWcfU+/Hs6yL5UNFvO6Dz2xnNWUD2mMCxrEVjoUrOYDF
2AmNwA6kSJo2XcYT9p30DIRVDVKzf/Y/w0j9L4vGRifvIJrYjAYV09ZrJxlakFwW
qADrdx4nuUY78oifJfzNXWKboge99UzcUfJwJdOvdFKcgtMCCpM6NeJ1r/b9ov2y
BUvWFsSP7KZLiJQUY535asxd4zRK8ATkd1QXWqm0+/KgD4vAYW7TGOFi8c1N3+QI
8C/2TOR1RIP7X2ZfxWjPlq1VGhhbR023lxZxmzDPLsgFfzZtKrCV0Icqm5MSk3jG
PrO4nNUI5KBd2W2Mdq0g+fMt5QgvOzeWbGrmvhc8hJ4MfwqD3bpAlRjrEKV+UylK
IG7LHVwqc5c4Q3sjf/jZaobt9tO++lvr7nKJanWp9YoiVlWIUNON/zHx8i2E9hbQ
qrwSJTzD6TTcBiZF/B1rjmsI/uW85S1dpsvj9nzSqkqWKdEP4l3eD5p8IiVPOxlZ
OCklr8/9JndqJC40mNbZBc1l8YxwWomkME7jrfKDdpuKb6Zu/zF0dYCGT8HHq61x
f/fGIO5FOIm4hu+hMtjuevHc4VVy9Y3xR++4MYyDMS7Tla+r+XlG5bEGnHSxwRI9
lBkmWs0SeYB6IB4VHAgwcVQJfdqhlypcLABgvtO7ViRgskSEgTp+BG6QVIiubj0A
Zia4+kX5pG9BKftZbsXDOjxeHmj307rypaZ7nV/eop4HKz86STGD8ZSuZn/hRLM3
8/n+NKTwt81Gc+x6aUZDdbFWPxg2rAMXB6LH0e6sCrlE3sN537TiI0NMdPbAwaJR
HvWBw/Y7PS1aENTx3LvvF6CRZWtW3cfDq8ydXfKIBCKb4W31LPVNrH2VnZ+bv+H1
qXtwFVKP3AjMIrEXZxAru/woGh+AFNfJcEfoUO78IP9Rj7wlDalwP8vyJ5SKs1Ak
Q+IvbpHU69CsbK7plMN/stBdtshjyNrNOu/UWCEjR2bMPrduwbacLzRZlfex0J34
eh4MqyCazawlMCQY5XkXjsxo2NJTTsoIBC3i3mKltnTNdaO2Vtpr8ZEptuMfjaUN
tyhiFLQr3tAcO7ff5lT72aHmKjz9K1L1mni7YyaUiSPt4kvDn/KG7T62uf7A3JAe
G03oQO9i0qoch19oqyLF5ROW7Ppjx8CRi15p2e8kTrs+Szbc3P7Fv0oOQ6O70PQm
aueN92MOPn85Y9HHpuZwiJLjG+/l6H565fSfK06n59B4KFeCQk+EfEuiSoIWZcR4
hG21K8mNb1iHEwUjZOvRCX0WgYabphzOybN30o4RxuF5rsfPXFPx2jbNHMkGEIFi
qXWYLVHlTQWJDEZYoH1Ivl0+eAua9wfk1Tr9P1ThMOZyGhX/FcQh5RP9VbSCG1Ke
IqeUpBwyC6UIrOLtM9nSeaRxGKYS2jSkrYHSaEjuodO3AQa+8BeI7EIe8rLqB3sa
oL5iNf735IGQZzi+vZDSF8mFbG01DlP8+nj4UEHK/EM1ahiqyENa/1huz6mgeGEc
GzL8lHQpD7Iq35bcMO6ihMkVKukwpSsAv1BnlDYWrIuHYB33pw/ujxG/rCfNfrsK
ZuRgyZhnU2ZPou+lE65moCQLYvX9uwjs8HPnQBIUrkdXhjUzPhkdFJ5DQ1zzgiNW
aX904hvX6dbBrx5leJHlEZmpC+TnKLuTPoq1E28M8UoxoH+KJMMVJWeeHB3qX/bq
NnxoL9lrVg3I+HXCTw8P/NqCkpEuIp75NVq63FryWoCE5rl9dlFNp/2k6852b3jb
S5OB+b6S1+N4u+O1FIXF1FtAiFBleVoIXTuprFb1/KtzLBwToH0ku1LImjuPM7VW
XdaEBtt4+LmnOe+kQYFJS5vxkCE10hBJU20wNqY/yx4lIZmZICDscQMJTo4WfWj+
k21GwITMev3suH7AOQo5csYKODtGzOJsRxl5HKGNZnDqhvDQ75j1PK5Ima3npdQx
VTJ8Fe4UC3FQHJW1ex8VwqNCJqBtvKKjkVrxl5YFTOvdeQ7z0ln8vVSp5WTkuy8V
k9uTgcA+fIR1OVLSkjGOeETE6CFPOciHGor9Mq584hV5Xnvj4Sc7aZqRQ/dvLS3U
s7ahqoCIztd2n7LULNUK4IQvUAGHSJ3R/aCJoxl0XSUOQjEAyX+3iw4/NUA7gQKx
djI9wOsJoIVA2LC7ZS8qt8LERR6DKrSgIx/itXp3K2GUQoxiPW7bsRzOnIUiamis
vTuVexs7JaopA5OHRHFQGMCjue7Yh8o9qGdP5s/QinmA3GySbPOoJ03OXhKEgqH4
8wIhvDcWViGmbI75uLq5ay/EOd+dwPDOW07IZDpdg+xnQ2hJu9recblVMqOr7dgG
Kf8leMpurFIFoo8jIDAhIjMyX0W47h+Z1BH1pZ0MZKbSN9uXyqQP6BkBpbUHPOQv
7/CNbEd7t5mVE0gwtF8EMxfPhXcchQI1qAk7R1wHmGbRbrqrIxfiONpF7pwNhkVc
oHoqrPb5V4vvtWkc0jDneSBTBHntsiskV5k+LtIl5/61Jp092n94T9yFs89dKHx8
IOURfzzPlgif/DWk1Db4JKIeBnsh2V1Rl4adP6MwP2MZUUjoyuWNwWHOV0O2CUKi
6VZeDjH+Si/Yc9Mz3H+mEpsztKvYoq+AptSbiWasQtk2S4jNzuRVqUgHyKKB06YE
KYOWpQOG+CVhj2MMHzVnbYdDDmmgfrWpLAcrs8GDKXhRD2aq+/cxjBcxvkFNiXpJ
gFdxs1Ut20LDE5z+lBW5r+BKBjUGZJK1Xf6nGwFxp5y1FcDInjrEKA0qbGVVfOBM
aatDuT/APTddQPB2MrP4tw6XtSVZXCTSbb6gQrU2GEH6/3ysXQMzxzr5E6C0+lr8
BEHxbHNjb4zDhC1qE16rJep+U2ZO8SjKThSBrtdZvQ7eoD3ur/FeGLeIlcIwwVrA
6+RK8f0oSl9Q3GjTBE4i1e84ek1K2VXGo1wIEdUVzhaHNbDj4yT2HjugclfMu4S7
6NdD7edat7101hNC9FiRuF8Oaw4y6/EMPsLcO2DNYvgmKISXk9l7fG2/CanepJnJ
Sy+TW3WzCtg1d4pMCp29oADlRlugUctY9C7yLcyOEZm1AHVVPJIH49QlbftfBGUA
gvtl7PLu4SpZzrkDFE6n+gX9De4ACM9r5Y4KkQb387M9CZKalLxI1j6tJ6iiyaNY
B8/CgDbxD+x+XoaoZBrD27O3hKJGN/AG3qZje2IrAxkH8A+ynbiuTUQ6jCBIMyep
riUJ0IanL7KaSGPVhEd1DlNdUTJLoX9bF9DKDncN8/s0VzOkQuTh4P2XEjsqn0bJ
errAfGg/M7dg5xmpy/azA8dhQtspJ6XD1+ANLPDcBAoUf2bwgkyhq9FFEYN5NLly
CyTyAAh6nOsVvlZ/x3ixQT0PpoOh35HdWT5BLZcBAxuOTiC865T+YnlrmiiBDkNA
s7CX13/0fktoEdTLnJAb8F9iTmsyoXDpOFXpaqdgWPK+TAWDUku//e5D+8k06IVQ
3DB5wMNlDRKDwNw8lz3UwamcfyXGEln7ltuzUUk6bBVdsH7eZLbO0uyYSZEOz+n4
d6QjrUUxg7qP73FMdU/HQsgCYoLt65VsiCbv1RxCQXTYbKA1r0I8QBqB1yGZOm7r
H9XUApS0Ht47Y2IznLGG8C82s2CC7laV065knQuL7M22TU5no4j3etGlWYzljbp4
s9tS7iSzPflY8mJE7LWyxtQTFJ+UWXhaaWPBSRhi0vsMHQ+uRYnWrZHqbd74KFrp
9z3wDjeqHq0+JTLimdFo/ZKRxE4PG9WHIRC4nd47RdSmlN4ad0B3+WOoVtcQ4dPK
dWnbp5gNJT4/FwPpSlQ0Zin2ThIADOkgo6wJcFmuJxfI3wNvvGfT+dm0cI9LbYex
ZoSTSYTP8LUOAwlJKv6OuzogtGJdLNWgTRy49h8DuFO0A0G8ozEMlMDAKYOVrrtu
D2ELB8wvtYX6MPYlGAdBA4kYRO2sNyXZh9aUjF65lMMjQ/XWhbfORBrZmhkyxXPi
z2HpuiB9yEFQK46oCA6LAKgXNPRpGBvLOKaXujc2OxuyAbYh+7oEzF8bUsZBMdmM
PolZV9rBdFOFkhW8BJLBfPB9ysOpKQvbvhjnFDdZXTs0BF9GByFqRx6oO+nrVFQm
FkjFw0NfKaqanf3cmarVhN49pgZQB3HgqgesNlS8gSLgGRbW3NyLZ43LT9JB1sOd
DeMZOynmPKoJXpPNpVzPv0996w/2lBWLbp9rWENYXVgL3OgS5wX5RzRkqt/3usc5
h3nOakKDVlZpTitYz1b3hVYGQ8cjXi0CmcvGRHi0aibryOfmaO3emLO+SAvEhwSA
pSUycvzUB2dJZyG7d64+4NRc5v90MEybzuhOlxqKdPYeTQXs3vsTYUvew1317LVu
NnLWhxsDnU+i1CHgnhYJuJXXEJETFJ5M5Ok5antIHv9yW5hDPgZ88j1rhc/WVM+V
AlTsa9QD4H5nw1OpUzCmdDSYqGsa1t3R7ks/mtb4sk5Dc6AJXk1AnqxE6Olt/v9Q
eXfrogCFKwW5mozREBoFm1u1MKV+B/QpmF8knH6BR5DzP4YeTsPc4JPUoPvmiXNb
DsnFwQaD514pyNO/hjz87d/ITvrLLGxKG64u1AuYlxenVDor9TR8u0Lqn6oQNVMG
chCbYoO8pHGZ/loVlDKprYjQUnCmYcgbNqHveGrVRMUDDslHpKSuKNNyPPFA6aBM
xT2/hmurc+KhxBc2gK2rcNnu8L0F2lsjxc7+V8qZv/fJJ6EkIqNQ9iSIiOH5JkAI
7kNvHWmHTIYgOFMCs/oOyLGqcUodNmQmRkJCuG+W6dPXdiP3E6+hEAjODlO7Jt6a
VkuBh40lQpftHiL43kRM1hoGQrnULdYfUE9NpvPBrTvSZ3Zgk9+3woyoag5yuOYx
hndw+wbRmr7Jj9nhGkcADcj08Y8Gx7o38cp/18mQqRzRT2ZUMzhFxV/FbPje0EaF
5JmpkcuUfxyUpLHr9m8GE0qWtoXCh+wIadgdOv2MGKXMppYt34MXshqMH38cfAed
/4FBP9tPWuM6N68KFqlG0HfSu3OhdK+9Pi7SX8XZBW+jJvX681+1y00kc735ZoaY
2RzW2F4P+zAlFQBq6UgNc3u6TA03U3jMKpi52jQHa8CGlclmDz8wjPpAV1viFdP5
lMh6nmYyLHKStZIr7vVlE0GFfdC5CU0u2V2JVtp0lpvHaGlx8jUYbzNZaQ6Htbee
Qax3DMKYC0+mEOxoBBeXByDhxuIDWGMM010IN4IIJaqSnKcfpZ0szHLGogjLjsWL
Te4VSLUHDQS8YfcbMaqN9UELReB31P9Mh0VIMbISN1dUqGk/U4wvHYaXccHgkZsX
wqYWmYiRihzGpJ2Co3lpq5kpUV7a/yaon23BNykRX/5i9TSQZB+vCitVaufwuNhj
Hu2yj3uIBafdhM2UtZ+RCZ9UjqqBYN6OVzBQRhgUSMnXYngKwGP/Moprt2EwebjK
U8n1fu5PxGwC+4ucP804LrTtJXc+DHCDSgudl7+spfyrrVD7twY1zU/Nl5Fhp9Xx
7rKaW84ZsHYL8MVzh2fU0NaCK+KnJWnPTFUblsYxIPHcK1uTdOpbvlzS+5xk2JOX
sM+SkbMY7VfV0Rl6D1ij5nsVuaA9nJOwAJR2UWKlrhExqsp0am0m3wSUg+gk+S5V
6S+AKwgUki8UIDi3zxXxfMNis33WcQ+smIR6huHQy++MRSWd0wTSBLP/6zWrII7M
9AKz2zhVzwnVHMUsSIEZzi2MFqK5WJXiUtkcgNSxuzsySzMwacof3BYb0nNtzZhT
wFHn3+pboW5zbBm0GIBCQtC0ouD3c7+X4CteeEY0ecbkuIIKqduJHqUWqS+Jy4fp
ZY9va83xSrxsPlpyArWBe9b4yULxnK/+fu9DUBfwSLKEJwV7YipNn/chs2of0ZYR
uLCYdGKA2GETTCf7Hej+14rRc5VpzZmwvijS/hG+0ZVMaO7coz3Hu/MgQkvgkuJk
mJW47A8G7CPmqC3NcbEkNcAkeft3c+n5cIhvtOi516U1sT5yrfDB+9FFsE260mEs
Ls3u7WHjVotw94e/NwNZ5c1bi+NJmDtrFDeO+XDAyyzPGBWrvZusl8tSg6nIJb7e
h/S+19gpjsoVR/HUPbqzh1NFhzyIXRaCg4jX86UwkdFhfEENp6oT2oix1e5ly1pG
CnNajQbxyxmYB9wqi6OhaHBvW8+sZIzqoz0JLxN4Yzrn3b5v9CxcMZBERkXmH1Nb
HjBLN6Acak6LQdXDOon/daRtDBiaoHAk3k+LcAyu3svJdek86U0ghQ29z4A5DrkW
a+uZmgAMgtDk/bF2gYuSku0m18o+vJ3QH12FCkTF2pbRf7EZWS07qJKnihifh2H6
YBQr3ZIXblbwwpJMs7cuZxNPTGzyHs7H5xSm/q6nVECD2mr2VKRhfI7EeHDJevbn
nLy9lIXf2Sa/2jM7ljaEjJPryaHCimdpdWd+W5QXoSLRe1iKJnBGL9LKUP16xQb7
Nzze4gMJxQbTypvClXZLVSb068aq8PQUG4MWr2/GReFXL7GQw7MVgthvxBepd/4P
dtOfmnKYoEuTrEwEh44Yee3vvpAKcAuUa5lhpcp1Ou5rnZ65vii3gtmflgUMLGyA
quj/of2oUxxezHteG9RTM3AUBqg3z69+Cp3G2n91tXLPMymLo3MqaNLWuJLZT9XA
D5rDb/N20VaNcSy/Tw4qFh2bxXGsOQ3zuOlGqv7B8Qkp8mPyxyUXZaoUWZVcfHM7
kujycxYT9xH7cwZ0PRAIaF9WU1af766rI8VI1ENvgeqGFjT+izDoJdo1SUK0hSLB
ZwNCKy0B3ht7qF2DK2H6Wbt1ri8FJkloN2BnX8I1NMMrE471C3fOGU2UBO0uQTeA
JRuisrk48bUhaWWs/7VDCUr65l8Nuz6G8z+gbcAdsoDzirmulKdfDGBvBCYhayaR
IdKSbSXYz1el2mhO/ES32XFkftWOt1daKvZVFQeT9LGKmmemcI0NIiJGTLSkhXbj
hYT0f4leYyc8aD3Dcm16FVc1HkPuG/vtFGN08t4KJnz5VjPzo2KZqvPPNDc/Cvvp
C4ZW2NfEvNqglZqq/QkLvMD53Q4OozFNww7hg3yh/WcY6s4/pARXxls9/V6dcv4k
tZYpIaoTsnH7+2e1U3K9WPN1HBBcl+VRWiAFRwRd3fJJge80Dr0Q2urEQibL4MU7
5xAxujvexSk9cK4upsLVZtyNSabBs3zImJ8zqYmS6ufcHXwtsomE2LR9zh5h70ht
+ywCdp9BnT+skTMajoVc7iP2sferi3b9xWjtOIAQHpI0lA7o++CoUpigSbuW9rzX
hSS0MJYiGmHe4XTf+4bOH1M3/Rh9qorAQNd0j5Zfy74ZnsbVOFtkEKTGrMsWLpEp
uU9skNbCoGuvhyAl0my9AlXIcEbEqAUkHcPq0acvWWfw70BI4TlmImY6JvyF2NJk
WToVb5ICJ00r3L2DMuHrVHIiu4FQXgXgkaW5rN7FR4uDfsUlUY750SzVdSkKnr/J
tCm9vDZSv+DsCryoQJjQCSPUAAf5S/yxx8lg2WP+5e9ZZAODy7Lhpv/VqZObzGmv
j7voXT4jZ+6abXTrB85ebk51UZx4Iedp4DvbMrTcTrGI9Ynse+JQdCbMDJAEjETs
5B1kDc4rrD99KPETDii1Q5chsZy9F6lve6eNTiSRzu3D3G36sUQzsSQpzSE1Eohl
UqMDnczLr1VmxYo4P9fTyxpJJy1k5QzHusocqmi4l0pmJCXNPM4GZeWEXf9YRMwH
38ttdqd5sDvGz65t4t6hp3PjbLNTzilPxsApbV4Vs4y1mkDBlxJHKaxKQwBT2UKA
CzBqlK8bBHkGoA14S1564egjcLLVnMkHuHwVOuf5lgp6Nk6YTKhVIs60tGlI9XZE
HuTS1Ac0SNH4YedbwksNmXTW9XTqfd/r93ohVX7PVvmsGeFTDY2ubivlI5d5apd4
LGxtuPVsSB2CB4s1pqfXekwG9ArtrgMajYbbK1IlAdpPUB3AALZC+SiluQPCzwwI
ryGvJX7nABAIq0nna1nPYVADMF2e0Zn5CQe9Qe6DQvALW+YgFUJ9RRpzipm7oWAI
kDqbdV4FqeFAZCHByOoymx+AQogxSgZb8ed7UDM4KSsrq1qud2IJe22rq/SQYR1S
BnyXgZwPdf1VrijItmdHN3EP7fGafB6kTlQaLob38GqEqD1B5smNY0gc9SFJpaTg
/j97rpiRUsuRijQ3L5ClUhbUUCCA3/4ogopa0p+oOqoZ9w1qQP+PFelyN0I2rxpS
q5bEL0QHkrm3LukJHYSu8jddSycGMjptMDHF1fa2mNMY1Th25mjUAoM61jpcxT/o
2FPHSY/09wRhSJxOOalRVrRiEv82ClOiiazeqBc55MXTOzG8wCmaguiUL9NNV2db
nSOV4tF7MSDKSz6PLTS4R+DpiGSLfKIF6bbBbKL4IQG0GNq+Fyr5tMtE9D14Y+1H
PIYVxMDvVfz3Xz1jNzXclX7AdtT9RU11sDrQB2PDHSLciZDBHIj3kmMU8s5sxiIt
m9IS0qRMXkgaNVeFa/jeBgko9I5Gv6PyG72SThHrECVDZBdmdgMELKDQtrW7y1Y4
ANLMabdy6bWyIgCCoWwgNnuA53vFKvgSGQ2M17n3HZ0WfRM/h9sDVagQuXHN04YT
ko2++fxFoL9DJLWytOD67PRaI8umfdW7fKLgjdzuyyt4LhD462Y0E6nm50Dyatyn
Poow5vsyfdAHFyYFcYxBneHBDSSy5GoJkwLcsAoDuc/ZfYYCQowszWNevj4pEnpD
oXPSRq9jyOjXzuSQIKHp7NTkBUnwAQbDinLBaC2+Xx453KHogY1fkFn035lTbK9n
33VwzDX9fi5qd5hBAqFX5Q1IfFa+BfpAt0HiHzK9l8m+D/pjTefl+XioMI72zCBn
y5R9KzKiiFda0fP9JVDNvP86+G8Xw9koDoDd4DalKLrhFmZbyLLuvgodjL8JsuE7
ZU0xBbUBoocNWxYpjakVzMGQQhnUkx2/K+utCXef3+ycoKGizsXVp3fq4i4c09q7
e7nv+ynGhncaMMiHohtyXHSI70xKm63Pt7wuh6/J8hWPH2t+IZAZ0eu0eO2z9UQC
iZkxPoh5q0Q/RB5WuGr6lnTiaSWxvptKiYmKZkA7wCZycqgAJG+YB9QNY5SI2DIl
PIriTFkMIivssKK5om5X2S+rjew45126d+IJL3ZqNgV/BO1vRsXeU3ImiIbqtfcb
Ipbn0rNqgLJlkE8Uub/EYvB70GQxP+qXt5+yK0ZHEj5/y/rNW5CEAJGx01U/LCwT
XdFi3zDZj5DkkRDT2EXAU4o3Ac6kSKRegfAK9oSOwmWTo4TeWUzBIcyv+F7N1Sjw
VUKGeQtlewCjC6/KR4FCv+5fd6ttOExXMCT4vXx1WP+3gVxWqqNLqIdmsBY8LGD3
TC8ZWGf4aqPrfdlo1b60RsycVrs/MkWG/7bWdZN9Kzt0ownR6eQd89u3/aNnoyE9
ZDFFUog3yD5OxJX/297a1zH/PUsNiOsglP1QF6Y7a2wU8qB2cozj/yRmA1H1FNOm
zgQskQzlR+skulq5ScGfvQtEhSiCQEWw9YWr7N8JtxMH6MFmrJcBHVBnpABfqT1c
CBOLelj0UcqmbYmUJ6v1FOAhG30EG37yGE75QYGH+UTmzPlwaYT3EyG6X4RiV+6Y
ZAA43M9br0oBgFxJ3LYGmTNE/St6R0PAqB1Xt/AShB7L7y1MHzsR4FAiI9ElZl6+
GR3JrwX3Rdu2ExOKcQwUxKgQZaN7QoxXCt3ZPmTe8h5sXzMfA4lQszzLZkVWQMTO
BhRvxNqRyWODY2B3cG6vmDLR4/EfRF30H0Qiwa5d039sAkxwaGkVbcQrJHg0GplK
sjT9qcwamCcOkUqvuDiKxN+G4Gu0PnQ42Rua1ID42CVuSPTYC+sdUz1O9DfosqWE
I0STUgblBe4UWA2VbtwHRCbzHsFohGzy19M6RxmAmOn3HWhAm4ZtoMMHrTESR8B6
do26fcOolHIxT8zkYzYKQ5SfXAn6ZRYoCMiguWl0lJp2mxhGwkLAyik0AfdPHD0l
FbudqY4ZlUGv2R/viA+/8DyT1hZg3W6GoECD0D54Rmf7Sn3MSQEFCt9MIVSXn9OD
C9wSXkOoLOPfbyshWwVm+LKftpvXs/QGQWobNGw6tuvdtVkVcq5aye/dNQfKeYeY
9ZmPldypkIWO13G41Kdmr/byCgeeQPQoZnWbBG68hyH7V9pBTV3TRvjJMCs0hug6
CxBp5b98O42xFA6p/hUXpHWGFm9VqAii8w4lIyRvIUgUhDJIcMmD74XDHdT+MQTd
cI6Dkt8y6BOLJi3zB/mP+kqSMvWFan2/OK+E2XSylTEAxbWywEd25fO5GZ3orZEY
qnO1Gtq/24hFyJ0cjcnftfUxj55N8rouTLYUaS25jHbTYxtQo1oAMEvVuLysUuTc
83VCwuIQIaLa2MlmC0+gbT7aRAbwJmGjmqFbZnyywT093WBlLjJxuhKu+mLA1uXS
MpOJb/anuV+WDNv/pLm5J1NEOiQW+m+e1YsuX/qpLI2fzYH+YMpAW8B7LKutZ33A
U9/O5LGCA+P73qpk7v2kNi31UG6CsGCWnV36ZdWylIEDS1YzbPr4ZlO3KKEt+RIE
IFA5aGNtlttK82g9OVT6lhOxjI0BSz7CL/VHYFIybBFTI0lt2u1x11/KF6u7UAeP
k8Sz4qBIOiFCrDwbutjV+znzFk8MPr1vxd3JdhZIL21NLGqwfRA8d7GoC6PMmlPB
XRpG8pBnhtNXQ+2llgmejCrJ75jTfOg1SV2JOy5J7hFDvvQteZoWBDYRuGIacvug
2JZDWk8XhMSTKNRJOYyYcwMstyxeWsZ6nx4QWc9Bcyw0cZokv/Ib9nuvWH5egDVK
aZ8PLfL7NJe/js0+E7Nx7eq0BwLmmX9LwpLdj7J1MBN/5D+xQkz6MKbNVQbwvHhN
WReYV5eFzhNZX5Iln59U7rvUn4WE+/BY3mg9lsim/HCP7imCVLEseVGkMSnwmWnW
+PGj7Q2UZFEtCv2UKpJtKc/ahpyhMphUOJsC8RKI4KEe4imaMMsf4rIwf7zJOy8Z
uLDUPoTJbi9Qd0EwlCZiu9Qpuhd0fYmh+oUHgEjZoAcj9pyx27sMH8x26Aq05es7
XtHng+qnGP8+UkUwLrEBwfa3uGHmn/BJ+3NYUvujz76rCdEYx1yjfv6mHFXLggaz
EM18siMW+X2BDbGlTubWwBIOYLZXZBG8aF5wEuoDUUqXvhTyG/kTPuTdVaeyD//o
Jh4GQzx4C1ZYYqQ4ijPxRN5OzvZ95VQq3OqkCgyTwLbCDs0YIgjeVxioVYnEvEJK
bfuZ/SPJi7xeUDWbscx9YALynTntBGRx7zRhjfcCTAY5SjDWg4MWYo+O4SdfcTPM
DfacvUEXX5ormWJclZ8bOQYRX2TKYL35q+ZPsjMICJOS+zrWKAX+HUwMVHbqm/lR
mmUH9MQd+grMmr316E4Ih2FBkGYX4L9SG56O6iqc7sF/4pI3tlYeblmlLKoVZSAo
VAqINL5fpPgElEl3wsu/HHHsCtuq1rZans8wSsxlMk1ujIOwcVQQqzxq4R1gH8oh
ke21JboK08Iz9g3YIGjsyhwpyK75aPSoDTov4r3Usk9Q0lzSIUevxxQ65SC8T0mD
JOmfrClR7aApjDjHSX7EAWHJ5Wcr13naECdJjAuUbNiWMl7cbO1ZeWKOlidLOvh5
cjAvsJDgjERd7Gs+WFC0qPyERhMUbvVMzRwxqTTMN9HUkFPYW4rgwl45DWSyhqfk
k/DFnWyXI/KKOp81nZV3zxp5vv/xyJ1f5kpBC36CwTgDydXXh0Sd456y0LaKLWIC
xBckdLQPQJeKKdAcTskBj4c7Klvb1DQyu6DqaSywnXgXlKGDOaGMLOeG2+VlT+L+
TWC4rkFQ5IAHHf9+blkbT5WTBMXluFQNJiFEsC7IJeLK4rmEgpYzHUvWdfMD1qUT
XJI0qHJCv9Lt6BtiHOuKhiSsCeJyrCp8CPHF0fDm1UEuosHVCsUNQ2dflHtN1Mzi
ae136IiMmIRt++Zq50y6j7qp6I+zi4oT9Q46zGXzuKJemcLgKDDMPxr93V9bPYw5
m0+E01D7z4UsrbByuBjSnffZA/9K8JPT1BP/aXRHNStH/DHPH8FueS2ESIktvovv
B1uH+H67BWqqWcwtJTemImOFq48eZzzQCrfT+LYk6qDI1+HhTCJ48e2iHSjB/mx4
n0ThpZfoOv0QIZemW1zFAPZphU0fjApu3waHgSEwTaWZPwuWd/cb47MZsKCWOTpF
8VKpAeyHCJVYzs1BlUojDaAxtPBh/LueLQTnl1rGsifYAe219iPGgFwL4Yb4WoBd
/MZ41TeRagtwnNJv0/pam1qfT1ki6R2tEj8uT2Ozb2/rK5xTQX58EVzERgBOOERO
ZfpY7BfrbEIq+z6eGNN2IAhxwqVCq7WEvbZWLYJN7x7N1D5KYKIJ7Is4rqBzpkl3
5LGLP8eJfZVbFue9imSHn18JxDh9JIe0MeH01GQQpIjDXcgueUMPphc4jD6MAjgI
MGLp2zX9NzYQ+/Jg++ZJQY2NnfjLXkqzJtmBCwAYbsJMyYGdnIeTmPVj8XD9up6H
Qn5Ca6Alt5KhHXwXsc8eb2R7GI3a0oiZjofeKQgxIN0xf0MLqSHopINJxUkCFbhf
DwcsLil5mkZAOf8U5PtSmwJU/vaYFE9wwJ0KV0bt5OZ8vBqP+MjKXElDY1o9Jt2u
FeDrqRxXfM/7UnG8mRA3P4pew2KylppdI1I1HuYBzPAGYFvkHf/nglnSwWR35pQG
+F4Zyd5d8M4jbYfGfglh2ggXav8B9/imIYiGYBvP8G8fObLPApvjnb2pdeYpw99h
WHeMPnFsi1GN03gM5OPyR6rSFsEt4LYpjn7K4jhTu6CTNLGVIMfEpM/MGpFLPPqc
MbbjqpdwqoB1nUI8Bd2Fklb+K1hdRIjOVzQsMN0iQQJm0+SIGMevXU5REnmgpA/K
5/DC4KEdENoTbFwf3yPijPuHiquhDdR8o1SBXzxXNtmIOx92IUV/VkxmC2UT+NmG
q/OHDV+LQfRy7RvMLVnJVy05Lrq3B+kqmhqHgUps/uxohVrbCH6kA6DuThHOi4Bn
rksWIg0LAgqbuI1bpnWO7uh5QujH0FWGgHRzBw0Ff2fgIrdjSUb0J/w6jI25kpXz
E8/tfx00Fxfh8KszAB4pUUJ8Db03VUnEs7QV3bPcrqsaACGo002vChMuWusL7Yc6
rlrsim5TpgUANzynpufplmKgkmojlaIh0eTHaaA47BKELZ0QXk3Qk7IxRGHkGGCg
btHEblGmED4qGlO63wGxUZ7ZRu5kWrhCS2JbNZgExfw/j25okfFJkuxP+1Nz0xvI
Nt0pFJZ78Yj2510ow3yPigRStaUG2do6LLoSOI8z9/GIvLRdcBwvU+KL/YGYtGlU
sfmgA50kyB9sSz/R6lVjNwxhW6CYo+yuxI7SxoIUyYFcSwioteAfUKdGbUEdrfF3
Oenv1bg2YCfMyQ7M/l070N2IjDZ09PXeX5qv59+D3pIExKm/WKhrC1Hr0CuQ7mhf
siTCpicB7UU4H4rScEiN6drJTlZEbVH8l0ne0sIVsg7eICJU+Rk7SPp7zChAnFwc
sZP+/FHioawH5nhq2BBigI13Ex2yZ+bXX/5LBtxOcucdY5Ns1saB9aqbQyIskael
HWbQ2uwwBrH/SMMELEgF5xPsMz0c+gjTvNATU00LQuFnHnqgLKi9Mk5MoufVfCE2
B7FbOKO/BlTH7gWGP6DU1u+64lp9mi8RGHrfcfR3kED/ANUXBrMDJsvph4tOmqs1
UQRAFCszvxaerVpR8zGHRUkLAWF8ICgJAbTovZfCWDfwYifRkCliQKN9IUmF/+FJ
wP/Ms061wHDBwa6wjLmJCvH9zutRk4yDRk8Vdvi6okKvGnW2SEjVyDfBZnhOuXD/
nEteQH/eLIrllw7dxEfuDCSm4bh0UoC5d3M99iQcLMZ4F65uTWbeSibRiK5PY3Ga
q0QAMSU3HRkQsnlmt+wkmbhAUrzXv1Gtowjfd4ORWe2u4uotaOb7e6PV3528mAB9
7kRNAoxVUiRDIpOg/C9J/1Ml3YseKcIBtG+B4QeaAbsxR3Gk/T6DnAjmZp3R+j2G
YEbS5f5e5WDPR/uY0rWdaSHwkKQlUR+hznOY++NjqdAMUpQJeY5Et8ru7L7GTJwv
tV/DoD2JvEDdtq3vc+EZzlfKUzrmbZXd9thjuJRS0Kaon7Px17M1aRHqR1ImZjey
PRixQSkJa8t1f1H7ypZ4Lq1aNuBlxhs4sgjUPgHFSpkEaSaE0vKGPCEYopE2GO3e
k8U33kh7Cgn4BYkaHofHSC9b6dC1/Efg+KhpN+Jy1pFELRKXxDs7mPTmNemk5/3i
3J/zCV/PJIjyEWRtfoBxOpeYIgochSMRfc11o+XJ4irF7U2rQd3Zl10ccPsaV1lD
ybnvsCZXvRmiw1lCW3UH+1W3BIds/twSzBbeAx5xVzSLoABJvKdIbH6NN1NyUbGL
Ozn9868lXPPrzR9POzFxVvT5dV3/IEqHlW8PI0auVbJu64HwAddftJWoGlp54Hdo
SQjxS3V+1FycROyVY3qKwWSlnrUtVYaa9KZYRuO/TnCFqEPZIEGImm2ngqhNC9Oy
b1W8jO9VF85TrHXUHpodGDs/bVLJCzNstY0K/e2300yr30t/ouMsJuvRsnZiss84
w7dwiSYAPbqVOSAPh+LM/0DV3FcNm8Y+0sm8vpVQxkvsoBKZSzh+Ct531eFPRjyd
v23YaUQ05VbMvExLY3gtLvRJWSmw83/ObCDo3baadOthREVGUAFtBM1tm7D31lcr
+GTUb4U3QA1DoHYxGOCm0ZLHFAhfW2Ouzcyd16nDq327lkT8huupfotoVV9jGHIE
tqQ3Sjl/zr+pW/PKsz9pAOFVmfkOK3qbqx/ElAalrZ318uK3Am2Jaekka8AC2Zal
V7C2G/ukYiTzKcbtPnmGQlyVxR9c2h4qe8ZeYtaR5vWxEn9wL3bihBFbU0S/jJWa
E3FRvtBqmOGF4bTwQIcTPHgiMxzFDo5lnXBxRhjAx6A749rzLZpTgPofs6RGBZhz
7PzxOsOijVPn9h/MGC3HGK/5sCYiC+aL712quWl+Q5dsH+mTLyyZOy1qB2lZrQTC
rMbSvRMpQnN/5sabqEjw+rmwKRr7jDX6LESzsJnr6TXGims/WBVuJb1JehmxGAM/
VMjZgqnkNT2clXQGIVVhJwGZcUlu+Vifn/U4iLo+JUtTbFXrxBfr3sEVHB0NDVRu
/7fmm73EXRnpL+QXS7SfRC/qXc+rldIhMVAXqMQsSYZw6sZl1IMImSTnqOzA6tOG
zIPh8EspBqSWZ7Js7UT9D206+QDxzHgUZt0abgZE9J+1ARJqrV+rN/WmEhLd8rc7
UTjYgZ0XOhsBllmKPO1ff1TW5tPGS2/yqWd9VN8MJiEBGE2QkHvep00C3uorAR9T
LC5pg7TT9Hf/eDBuGZTDnH4BnPbty6MTjfFEfgP5LTdcX1pjjSJdfdzgSlrKuhXp
+TEeJNJoUNWbv1jXuEaZ4YNeHUJWBud0xN9m5GzyTQiMganL3hQ8nAsNGfJ26BIR
XXm+qMRsxTzZzB+vMAMkzX6xZakyGwHKnRMhEd7WGeKvcVOeH+T0FyWLP+3XBWJV
fpk9JYC2jD1Q8+fIs47u+HUWPpYH6zYIRdir185yaBHvsZikfv5k/B2TxKfHZVmt
cLpMhaoj3CqH7jfQrF0JWdJAzoSFcn6MrN1pq9d4R7FbzpVPOQQGqZYj/Tu4Zt/Q
VjiORzvm6pl+tRosJ00VlpHhgHAfJdyjVOjmooF6nVj6+k7Em9lEH/xXxPBymrCT
4A4o2dAPRJbppUGVn8mKzLRSdfJrRaDW7poxMewL9srHC/p4gVyYh3ew3528xEln
gC0flc/BDtleHKaUoDI6Twxoev2C6tG5NE+kcHWomxSjvTlM/7b/rkmRjI+rvGMt
ClhsvAxxSZuLlfF5pFPqLIujJ5d/KdrNYzzsy2t317LDoFKUibf3h5y8KbWWK9Is
HOJ9jtNdtSdnQCoGha7WHzxd/JhMQdEM0MPKZq2CsTvMD6fGY89Ied9bVnpflYrp
VNwTxHumdcAw4JzEOpD2Kcr676kH5HEVCZeaeTvyYOgrA6hOiOkik404aK99I97Q
QUP+RA6pJYMACpFV21XOwc/oIq+/EWKN827Ltyc+Y4OimgxldgA83pqnwkzflwkO
yHXzMng5MRvwJDIWcqVbEV1krVb+FFzq27m2Dl9l2mvfuWqpI9DxNYUskgeVdL1u
OnU5leYZ9/YFDClq2t+smxdUVpzLUXeeRjBrxBWN7/N38F69388fcJKWxNOrCk2R
PqQYG0Q3k1eS9VkYfHjFlxnVPPyHOw+Ww8BRI7tcvJhD26IAEt7ZySweCKnB3s3D
I8Y6TeA83g6KVVftAb/lehD+SVO5yjuteleaaEwEaxVnqyowWUPHBP1TNdNfwLx9
mCskiPNDglpyKvphCrorfcd1npDzzoMv1iXIURMNb7GlQqKhumWKYtI2e65h8cne
a2bFT2mGlRQpQs/ioKdlpDzDQ1MQzWTxgI9F6vyVXSWRGb769t3HrvalJG1VYGK1
C2eaqMKQNZeLa1jb/oOmMCCskvnXQH+pU7Gbi9dwbUB7Docxq+MwADr9H/1WSFDK
4tAFD8X6DtQyffGYmuCocCW+4ni49OlA9inEPKXaX29Bs3eOn/rdOBkiUWOwYKjO
h7LhUh5DXW8ZKuiJJ/xggh363e37NFTQRYhTEK2oospqwu32hldD8fSyoF3YSNUi
D68GqWMeYUN5K91GyxM5VaVT7xDLy81rPCbvuBD0IETNSe5JWUzvhV4s1UvGrObq
XkxFgEiLx7hKIbqU6kQJY1l4qagbcREgw3HUN7fr/yUpj/Ez2a6Sg28JIIZKIB0Y
0qKd/I0iuU5vOEcZuyrYABPgrEKRj9bxJ/i/yjDli7ww9ZGYQ4nT9WyCF9+ZD0C1
/8JExHjb5Zj/8shcNPtEV79z6s824ewrkN0YQOISV/aI6fuN5n4INLUvZLG0M7/C
wjC8sqQYs64Ug+K0lZk7FYDVk5BN/V8O56y4N5nSUBjsP9riczXw6KUggRgrKmf6
iYuhzaZwg6Zy1wHRI2F2x5nBPpL25gli6/Z5rEBTNvmwPtncQ1rcGFMnNTy0aP9T
xpkSA2iBqyFSsi/tl0U/mfsI5bPkrRMcL1PhVq9THMwCYSv58Ys00kW5sF4m9oVb
SMwGWGOdZMk7t9kT+8u+A+7nHn3WdzjQEafvfNK5wAh8V9ch6dRPfNq7EhRNRXzR
amdgchdRN/d/7p+pe6g6CG4OuZ7H6/lNmOb6uCbGj889rGMIgrU4jb+vndQoIaEx
OwDkWcmIm6y2lHhilO1+ttVtZKf75HR8/lBZsHmxc6+0olTQ9NEVXTpZUHfwaBzh
Amf4ygn99s8H++/LHhyHszrmLTnnIiGk0GpObnzIPDyMAOY1jetBYkAlocaigfAk
nASjy+8DdaIvuehaX0Gn7LM0Kf8giddvW4dEybEX6u27Uzn+80184BcbacNJcRrF
/HUUYHgxDOLsejxP1DeHBXle/xp49Bi9koSKrcvpPxxAEIbMteioyZPOQeflRwRs
Bl5FL72WuIXDjdlGNvoXeiY72qx4HP+ulsKrDFsLN+CPArhPDQGhv6A0SmU5eUjK
4ycrL80CWEnQDs8JtFlNTUUnxDy3cnhUfDmH6SdS0HHunMGS306P5QI+4nqNfcCY
YdBSO+JJ1lyToEn0n8T2h92t+0AylC5W9R9m+gd7RybZRkgce7nm98/Xh3op1XGP
hLEs10V48rdxcEtruyP4JP3GNMEHTg5NIaWsG22hrq5ZsQdWZ72VJ9fUWOyNbVLj
9vKd6xfRL93HTo9z5QyS3SLZ/OmsCimg8H0XdNnQCk3GB5UE1giCvuIdp86MC98g
bxKacoSUh4xGDio4O5EC33GhDEBkipVhfF5RVonDX3CKi20jZTUViCcPUnRqDVMX
AZhp0xRsA7I4VgRLIHrD4hsq4GZSTFvgo0oOcdStuRlL1kj8M3kOnA59KJfy/OoM
h3kfXt3mPjHTLHw8YFg/AG6r9RySWSuWtxm46c7A3Jh7/aNKVcfj+0bernmRAxf/
Gzu2F/zneYSWs3HVttJigTmkkOMF7XUqUl9n/lqNHnYQEZ0Mam9le8aoqQYZ0hq6
ZvHXOx3/UtVMPfqQ8wCjmoEgb+m02gZRvpcrPUk1kocSTNR1Au0NIfrSooPknDGT
uGZZ7Ijdl9y0JjZ7yezj9xM1RaAaALjiHQNayp5RIKCpVO8yBfHCLs9CeLgUh5S1
GGOjCTEqsppxlJStDdN6w7AWvNV4U8gHP7O7C+tTvP3v8ZFha4Ui4dEWvFxYi+HK
QqoM6F4Wr2iZjmdNd8A5N1Y5htwrwadBSJgYKJOrXjk6d6lekASYvHoGdqpNEVqi
Cyw18RUx1PI25+gLlJ7lCCxOjSWNus633uwYPv+KNi+C0gPIsfL5Ayqg7On6IReF
aWqjrZA367SxaCvjQpKCInTBFfbAp+l9amQCSNvrUcDuseFEEmZkrq8vN1dw8VHF
987BuceLpztz02gfjyUlHeiBlihEhBPweOUmzuj5P8womrD1BHmK70l0Q5hUR80l
KLylxKR6rrNMWehnOl0kAcMDxdz8oD+/mNAWO2hv5IR6qvKucA7uItgpY+6/4xxm
CKYQ5KrdBTVk/sRglNM3RDdLWdJeFNVoys+EH+8+2Yf2KrraCV1OdYisA9ZmRkk9
vXGjh6Tp6F1VlCO2YjiqSrzKkU36SWT/FXG6lRBDRVkJ9R4ZGelxeoMR3cNkME9S
6S1PBsDA4RDTL/ulm8Dj8iUaGVQ0dU2Ox79yg8EwQuQmKUMTtlq7t/4m5pBEvju9
wWtEJ+z2yoZ2Ew4gelP4Ex6UW5Imq2Ja+U0ApViLWJQHcS90dZrWkRbWkMSWg783
mZ9uAyYLzsmRZ0l081WkFWqNhOe30PS+Z6MSiV/HgUObd74hihPHy9wNx3DK3wPc
jK1CHD5JBL6/ob0a+kfk8h/AOcCbKOEQ2wHoMHVtRzX3oPgeO7afvDdI/gsE1Q+s
ZmsudfsZAOB5x0pyxAjhAUSW4rSlaLh+NHf8CTIJvbQ0vEpFLpH3+JhDFSXEBIAN
fqNkzbcWC2y88eREIVpFdxhO1pCCiK4rlMFIksqnXGVbkXd4aZ3SxSZv3m8IMBSa
+9Y0V6hW3HUAO2p+mGOiXisyj8B+eYM16v4IlR9yCvNFoG8BogWR+9o4XyLPZMId
zqlY5597gF6k0XClv4C3aKB1dnt5V6lLN0fulqKBGmt5OohzuyUcrl1hONvu3YsR
YzTYFHJxQZeanHotZx/nZ1hbFveKTR05r1Ae+SAdF/Xv2DxrgrRR7qev2O3UcQvm
ftmzxs0dKPSQ3nWxbVwR2+cUFe7N/ArqpMT3rRKZwBekyu1ktGVbSce2tK5CwV9l
7hdeY5Dj4Lq1bbv26FaBb8uC6KNadi5pFxPgTPC8UajX97wyVOWprBM1uNX260P+
7S1HKzErwHUQhPaDV5xW2Pl+bds0VJ3Jf5WvvCDa/iTEMPDne83FPRlXY1bx8t42
yiem136f1XAuoY91oenRYIxxK6+/JAEnYztfXG5ioCvRFDZsBZ7BvL+vT+uH4+dz
OtzGC3KdKnijG+UnELUY5fVQ7OxhKHGfp4FXqefw4kbAghjuPz+0LhnjYj44gWNe
3/bFuOpubj1guJS81BP67GT3xE7RJup9+jR9UV0JOh1NRUUA+mah+5Qh/m9Podzt
+/rX99JsozeRHH120CXPghTK9LoUZUaTUuaFpK6vSVrANJMu0UHEaVyaQZJ3ui77
/YB0pYpqkp0NLdpF9EWEMJOSW82NOQs0bi/xbtng8C2et4IriD74uJsmzN6hdJ+b
8cqYuBVwvWx8qAo3A2VuTNV1G9nQ/Y9Wb+0/u83rYpbZroRpojBU9mMA3Q+NflVJ
qbAm7Z9v/wKE8CfwMnyWHOWa38KPlJujKjTa7OuQUb/yDeGrggtOcFl3SK1MRvZW
8n0BBxX3ux55ImnpANipvOzQufk7pZCmRfrjM1rEaBhvBd/seAdhtjz9pnXrDXAw
hQrLwkn/xe+RX1CC72aHqsCvzCP9/Oqivx8HGPxiPSHOq28g7F98WO6m1rjZdcyF
MuTSzxd1JSyYgw4O3+p4BIS/90OnnZ0vaBawX44kqbKDECMSZq8ufJ9iK482KT4l
BXIoeThmHDmGWKVZL/oINhSaXlTvFQDKBYrhMCfvoyPj/OezX8BmbWeq+cAxg1HJ
BJl+UYmK5XdOTzdd2KthNN7VivuGmtctuR2Y2t4nG3QZFPjWxz+NjlHcnXQqEWYF
o+36QvL6ddLe+jFpsICC9gm9jZv5NKn+/YKmN6za0Zin/wLiPs9810Sz7dPLTJpD
RmP4H0JRAeE/WYR9s7UriofQ9hOkh9LFs6yL7yG/qi2NqXm2MhuBw+oRZWrQKSFI
QgL4E5HJj0TYG0g49P+etZTEqUxLzfNEa2YB2PW4glsO3IN9ODMtqByNTi5xO70P
LAafcs61cP9vKMEFxVQ/yYEQsAXsEvzfUZoeTPPkc3iUE3SbbCQ7NDXA7xcLz2Vd
lgb7DXzShKj6vXbw3JkJM58Qg5vbAg6/iOx37HpA5eH3HLw8Z4ZWsK7SAieAbvHs
KwRBPd3o1pGSWvtc+9G2QCRf41CWnNvm9MEGMbOXEquXuCMeVVkIEUiumQmKwpEv
PNI0aFxVte9zt4OzR/q1F6hXoiblBYV+apsCtDrx0RaGWzJ9LBu6rFgJe/MP68NZ
G6sgrAIcCdCrGlRTOWoVnD+aoTdvn/aVdmRvIkgoSAGHvmtBjw6ItnVHkSSXL8QL
TlESJSv9rlfyHOEuTd7nCVNjJ8g3eu7a5S9vWwtDHhKLiTdDcDv0mzCOugFmKPns
6wkHLNtaAQevHwSx6TOxSJstd9KoEV/u7H2qSgOwi9xm+S6Y8m7+tbnwIk8GKAga
hmv6/5jXmusKubO2NMwQ49S67J6pGbEouSJkGVfO7BEy2lNfuTyaBdRaglfM0LWF
jdhUVmgV4D8kJXL+eHn5Y33he/CaWDS92xUNy7fuUkZ5DzPPUoV1xP6sr6KT3WsF
3lDmV0/4M8hFNC+OPvVK2y6jxS4NbtSqZoqp8WlZdYFd+pxHNr2xPavNYwBjoNb+
+psWXNJhgJfbioZg9+7KWfeRzYuaTbRT/JQSw3r3RijKa26ayObhMRcgFlB43B5O
Egl+pCMVUUJ/Cp/7bQuNpCb0yjC9Fz5hC9skEhxg7RkMb8ToG6AkYAnACZzO1uel
ebUejc1oOCnk2qR9bOD/lN6fxehabBIjI4U6COZ2mZzBxf3nENwlt25caOhLu2QZ
quwMMwmkeTURzvgiELldtf9ddf5KWDnwFyI6zb+2Bp8+NluHHs4/WiPezBkynIA3
PdK2B/d9CSOMM6mLfyIgNfVPnVANE0ZAKt2/td3h5K9Cxk+RqNdcSBmoHd6a1Sah
BXIZNIvSuDTsCOmTx44CYfMnsVTCi1JUjksYHMPvxbgMEatQGAJ7HuhEvDCxLKOW
ReB54PrTe8T2rlfAdkKRDys5c0cMTz3bHamZz6U0voBzlQmJhx/X77Pj5Gnpu+A7
1cdxs4x+R86CTL7Tve3PEFv7CO9cWSbMjfg0JPAUt7l1ij2eVrCsY5LHov2lukKb
LX5auG/ALj0t4RJ6k3nDA0nOIQtkjB7AgTu1ML2jU+/dj6Z36CYbcl1F0JZkMN5x
yKG7kWEYoXrfJ7zGmIGp6Z9JKZQUdEBz7WipudVsUkGaF4DtkEOuhp03Brsbg5g9
XlX1GZqeCeHsY4KbMt3X3q5kXOZqH6eAXJgUHAqjKMyLgLUGhfTeiuxhWc7qi2S/
mevP1DHrkueBbR/f+dWmEp/Mci2Fb7aI6HQi7pAep6KZYjHNTPiSSYVBCkYUlk14
N4TPGSV1UHjAqZ0MmmT/i7D02ure878snC7V5pFV97Nwe1IjSuFp7s7XIi4BOB7r
BjyBrD1g2a83L068JN14BKh8FYVg6h9E7o+p2E8OJNc4rY+7XMjgls2AwNqsk0yx
PFNuEw4QHzr72fa5qmVK1TM2BGGz/2szh7XzEHvLfG7o2B4azIDmzzxmUSZq/kiB
xZ5eUNl7OOaOglQygTMvWd8UgZIUirvm4ctMZuGBQjREg4meIUkFtgFn7NZyPe5t
6OUI40P/fQr8e2glYvUpclAy66QmEYlApyttUSl+uJHnS3bMpbqxFXXnrzJ9uF/u
HSYzzPpQvR6qghCkwy/eb/WR61LDRIW3CQisVwMuy7D1SvC9M/t/z96fqV5FR19g
rgcrcGbn9Vs3q8VuNnrZpEqUEgpQlbOFQR5rXXqwSLen+aw/BmybGmNoN8W1zqdx
HsG3ZVLlkZCOuDE/FQd5CwFJnHnlZpq0mbBH3XPo8+LqQ2U6kfrvV9JCSt4vnpex
J5ltvQ0Y/623HfJojHBh9Ybc8hq/gs7Z2BHFTTgXi1gfvs/JhQoEfhT9W7rjVUdS
Wt0iKnsW6LOUWECRSnZfWQEADe9wbL5u+8NkKVSWeIoaGhH1uXkAPCMbcQfInzfu
hCvxZvmhnf0zTqeJzgKA5hgcECpLe1uV4L4A1lgMxxaIxc/5M7mKaV4G7t8t5JIW
HF31glPck7iOC7s5Uis31lW5bioVbWnqDhHeBksurzF7+7P2M24WyDUwMtNMdM96
hKtPx2+LvvQnMYRTEyXrBnGUmt3wcKTN6R+ynlmdCoXRDfH+lhqath6VCyZYw6h1
ssjznvPjFOxPFwTe0WD8YYSvnB5lZIop1t95c9POHL7t8nJ9qQPegpFuGWE66fUc
g3/Dt/9ZOd67suWndP0hXCEURPBwy2GCn9KuxxiN38BHM2qFxr+V4DrOe4smhip6
c1X+oUx3qWtJatLQpAxu1v/Rg7+Y8lomSPERL0lq3Y7B78lKrLCcg2o9o5kAZqby
u+lMnVQruFq5sAlFY269qeLPYrxbdEO3DYe1dXscXtr4nl4BbI7/Z732oCI1V4zZ
masBal4365LkjkD5Erci33+u2uoXUqlNlVFM/CqFkbOss1HtJIX3fMNBcX4TcxqO
w6PhIG+xyh3BNMj8a2oQjJCrD9BJXx2Fbx7FG0QeJ9PN9vzQf1h9SnXC3pf38yma
ghaCCaylN2FAAKv8XYGc0BbrKLu/0x6T92asehfSU+YxNxjAA5KiUMu0MMne586a
8+Fl600eUtnfdJaxNyykgw/a3AAAjeVjoOwBsGGGMiep5Cf7c7ufSnFfkxC5gUdp
nGuVAqeDaw2363YvbcsOQLGzDSY6os30hjnDUc7ZcrEp0lNphIvjk1y26DzOCPyN
3Fa/QFPgN42uesWfmaAH2nJux85dgZkJh5vz+gHtsaV4mcq29O94HMsk1cxDHJwq
QXkb5czgoYgxNbqPsiS76yMwLEe5mFCdO0MDDIxKOA9HO/wB6qMO7dJ4LDfMCplo
xbnk1VtjuhdyuX5RmLP5JjcJcWbMQwlh/N6T/4/POeBPzXp5kfb1Y1JtIU1bUOO4
sVBTnaKI+AzaiLPZrOW//jxndUUHXNGwdi1rkvAkKjMqJJvHbiD1TUabTiFqkdNI
CHqBrrBCH0w5MLiRqu0pztbOMWqnAWmsQlUUNIq2b7cRJl04ZNthsZpl96Nzu29M
oDQWT4gUej2ef6BdhJ5D84TJc1kAf7ZyhaT0t/SeLxHkKlyg/wugHGNxJIiRTVyG
SNwR2eSQZKRVazFp9fKFNg9glVA7dHZdh1XJDiby4AQOT1L4aGhoMIt27PdV8m2r
+AqyRAFE7lmskGJmw9VZ57OqpiCp+AthKOiROVdfmwuxqc8/Si5M8Iq916Vgkbf+
b029dHhQrrhCXJZfQP6B0sozbqGxg1lJQ8sWq9lKZA4wbv8dAddacjMIhnAIWdIV
Hk9XHw/uXa+YR7lx6hW489XkMWg3xQWCwbWRXaqKCmtm7yckg4cGlm57wLjiKeb4
aGtHgjNuj7O6F17tMmSEmBj9wphlUVGjqDFwiHGrpSxnUk6s9iu0yv2e43HTAS9p
hRT7Kf7y7dzyYwo7GocBD8l134PzxbdeWkHdYXQBfcUs2MPkraTEdRQpp2xO7QT1
DMJ1IRxmxLbVB18BMi0YwQ00MQv2N99i2ekFUzFQg2HeoEZRSB/si5ZjZgBrS7pr
gJwUea4Eykmuv6gbmEux8S/lYy38By0Z599gBlKpAmdXK0y2thDBYTqQLfvcJ9Np
Otg56QWwMtD/yT0/vhSjUpkvv7sizRv0OUJv4Hhv76Ki2NfQxCscg4ZU5cTMWq9N
2H1FsorI+8R3q21S1O9Cl4sCLm6eoS3h0/gucC8gxTHxlcmHQ9ZEdK2NlPzbJDgl
HnyG9DhLxQtqtz/+KZM59dxKGEZ/FmXU0oINX7YLg8LeYr0haqt1D8sVbhDxRN1b
RPZdjH4NvFUejZjrpblcuxz7DdDxU45VdBdls2/DT1Cj6msmMCuNDrZDPw3S9Ss0
QJAKMKzkeWdT/D1KHksuxWsbjlk2LtIuJdG3KQiCQS321vtwtpbWlxn3ZjHJ1A9/
XDMpEks+GjcCpRX7oNXjzk0BtwfVOF4SyCxEsxJeEu5aQC4/zMu3oxN3WIujSOqv
4TAnHBzx4ZFxd+Up3Nx+ULdOjpAnBx4UpTve9g/x+dE2gr6a6GeQ+QRIf5dL8xKR
ojvOYTPpdeXkg+OuWUkw3J3kASEed5aT+RxvLmA9ce5OCr4pMnzvfJyr+gsSGNaq
SAc5oGdSBo8ZxN11fY2ybHD7NmrVg/+giFafLfkmCgfKShpXC6GLfPQBSAHwRYLk
ESyI6lXvpgTkzIeMVTMcAWnJBLVMhzk1JSSq3syjA4Noj7uRlnDA3KtWaY8Lqp6u
oiS+qKj/P0Y+0ZxE0JmGUlQCLSR+9PyOW+TU8LPJ0zUtaerns2VyT++GyFVZ3rkN
plSTT2737ku70BFAUNjD9dp88wLb9sbDeWbsSYTFWjn2HIPdjTfSs0JlPf0UXD57
yieXMHWNJa5n5kDRQdZM+0oOw4ihEGH8lueP0w/kC0lhqVHvb6pxdYK5QMe547/G
bMzfgB76epRThTQ26CsoSDFZnk7Io3HneK24Av2ErEHXL8WUBeSctxML2LPm6eJs
fJve87gorC+8rfjifeWrXMUfzvPNfW1KpVzONNmEjNf5g7ITk0Nk8ixZfznVzd5X
4BE791y/5x/h0rWGC4fFc8duUY+7+pSbx3guyFH7NIUe8ocQmI3y/H4epm1VVWdL
V5DFQxb1MQSu4SMwfturdjxqeHhY6XIga9yEF8fXzTp/QsRd9PZ+zN4osy2gKLnE
RSfqy+KuESHcO1a7xKXFXNYQtvolFgK8ltHbu7goxGq3y/QtSLu+qy0W+EWDtlN2
KVUS9fD/sPXj1UgjCQDifAbIXejCq0KWXJm5KQ0Yw9+dMcS3cFDkEVzk51H71CWA
b6xmnfFQXDRWRtIpF1rgUATXl0z4EchLH4DOpiuttOwgcCrv4CIrNWGB5PuMUfZY
tOQLpLgYB407nPRiWgW4Rr0LmMYMpPoDF0ldBqHJHTIWRuTsAWg6+fKUXx5xJ5NO
HNXOeGhhbk6SITgt6kQClzW84/3b39dxwbIysbkFvOxatpYdrcFphOdhYjsyj5DH
PNhNrEDsiQ6wCTa79NzmyiUjGD/uCMGglZS5vMw5g0cUCQlWr44TWncrjIvf1KS6
qi1JahcVeu3DLeG00Oa1aLpFt7ZikGtoS1j84b7FrvH25Um8E+vwbGGLnpfrDy9H
PhVEE5N7yahK2vHwEzHjyYHGGPrpX2IQPsfSCwcarejU/SEBpF5iTtv/FAMob+NC
URquFxNM/eWT596hXOxnMzg2ShcrwmKnE9IvgJfKt0bpxdUwuSMSfVeXybdY0M2e
RD9NqkJNNULHbClG3YFzrDtTeyfTgD5zmLdHaR0NFigXL5UnWvPiEtHGQwYPjOtJ
1N5yu2ksbIw1T1V2beJ0OkD/P+6RyyLNs1m2UpypP72TOgkiADT/cSpycCB5GjYb
CTkMEdl5VJYmYRFl47JU9FxFfsF8xKLKtJg2AEGKP94Q3/OeKJPZPDiUTiWc13tj
9VMfSTAvE+TTvfughyJtgD5Y9FPAGatPmDuWALjfhZ4w4h9+xjqin7TavLnwSV1Y
4xVTAjRH4f52xCFSUHHX1IcsK8HZ41525zUuMXAeJ6Hfda97vVYKUN0KQiCWDdBQ
6og/vF3ORDGw1VkmmoPI8nsxpywDJTecGBRDEDeVz8cLxJwpDGXmGttQ7uJ6Ejmi
QelWYhhyJ/Gz3x9Sk5Zz0CyUp1kCRG3hg3UEdwItKTaIcltOIYFXXL19nJPw/+tC
Ol+wPnkcDIfJurl1y8TUuWj6soDarpf5g+02e0mYHF0xfJsyPWrq4x6i9gs2HIpo
iIiOKr22iWCvmUnUmf+PjfsEol0c3t11Y7SZ4b12teqtC2HAYTQHPfEOmntNtSd3
qzMg5Jo9g7QlGgffLHAFze4fk6N3j4Ttzxzeg2ZKpR/6k0wrzIFCLoMZMnGHHeOp
cqvS0OZXJ4xRQMYwg3xfsmvFX3PQRJeP7saT4BoLGSzLVOomzSSWSzLd8iX5/m7C
gaQihwa7wEbwNHK8c9ZnmKNLLC4bcx3CaimcAHKE26uPW/aFuwjdtdCP/s3Pee3+
uw4ol1dg24hlHUEZ3Hq5Wzbir1D0KdowCulfONvQ15rfQOf1mZS6EK/+ilPLw9cU
NrZRRbMQsLZIofK8r1GNHrWpCON/f1JkMTUZfinD6JkPXuGI3qHOjWk9MrhzPFEg
ueWkJ+WS0M3cxD7WbmnD/SYbkg+eVpeOeZhLLIVUseVNV1Gekyc4pfcFV+II99UP
VKzNYf/nOWexQe+M4QT5qgMsz4zGfd80orR3QMOAF8XDzJW7m1Mx2iWbyzrxgPjY
vTrrniV7qtZMbkiMg44uOWrU1ntaEk+2vvYAcP/ekUUPB1B2r8+n7oArL3mewAg6
V5sW8bJ5M0rJiioUyL5U0lMgAXZKJZZLPj3COHdH1K51yYR/OQvoAPai5u2jMc6J
Si4tz3Ajvosv6NfxxrfWpAlgVZ+MF3N/tHh99LfakVD2gVn53HgeWUxzMB53UqNT
+exg+utYlT8xmu+rNph8ItAowg+l9vNCeE9wM6+qUtqHAmYXXT6UJVXeWh7NZCU7
3vyYo48uIkjH1OApkzk4fcGmuPwvG44FFGPO5nkSpxh228x6+EazK69vR0ap7Fo1
YI8cQdklR1WeFxWrmrR5d5lx6edPnzMKdBiUmZmeeiN+EdmUNY+jQ/35OonuF2XZ
0PUJzjOMdH87qmHNisITln/AGrSqra05s4vlSwaU9hVrUpaGYU1/ZF5jA4HZNxN/
SlcDgRKk6pqzNneTVnTpmA115aqsANdXAF2hgY6mxuqJJrAyXJd70Y6No5rzHXS4
Sf7ftpkberzbAzbW1NNTiOZsfqeDJi2z8r/tE9GAeSzUztcG6kssF1cZN6dUou5r
ldtH/n8mGzsvDA+/VX/8id7C5huaSLvFS5I/POWHmwQv5xaHEJaBn/H6p3sDAvJx
MHWtvCCLnGHRLF/ggLnirqmATnKbdKwu4Pk6UtEIT4rlkGtbcmPqWQBHVmQMYHqx
v+CP2NEI65qS7/rwt05A3YAXZ5ElB9wGyviMxCKxezPILsxEYl5XPzMoR5ZidEJj
0Mp3Ipyo//cMyCVMsfjhRqCGbmuNjUbcwMi1ea5B36P0foHRYJmma/wUU0jVv38T
mkra5Q5zGxxCwpPvShnDKhyTEN8wzmDx7qiUvB7+dBgpsTioX/0KauoNXZBKure7
ABrJpIhUwRX/YXDSrqjywyzYMsH29mZWMNnRT2rGxc/TbW+b2TGSfay1h3vNyzqW
tLhkIJr0d22R5RzIPadVbB9C85iyFLN4QCTxOy37S+Xp9R3w0S78gLNtz93z4eSB
8XhcdC56lOd554W8dOBNoJSTuesTP383wUEE56Xspr24SHmKZBdC98uq54TpVI9c
oe6Z+MN7rOWr/KymoWIzhhOrFWRKL3hOxl/uz7S0NblKTtmKH05bkjvPr99GtcZ3
PBT6ign7dAENFN+Ho0dw0WtGqFV12GJ78m909Ite2sF0Y5JMk5TNptAZo0YB9a/+
5QxgmH8IF+EX5atGC/h5D1QT/FzWCUN2VnTQntwzpopGzoHM8b1i3jDZ8Bdi3HOX
muaEBj9U6qGa3j6avsoGQ50tcu0oJBFGjlLd9JXGudJL3a//dd4z3W7+Ibi6BXhT
rz+9U0ZUf9yVvjT9z5iyvRltJps14rlxXYwMkfCejQ2z1F7meAOqCz+hWR+lGWZm
CzHWzrsanmJ0egOjOhd27ADIKe4PE/a9JGeCaXLga2XHIwagLf4UVys+h/Ifhhy0
U5xcgB1HdTZ/SrUxqLqrGxEUxw0C14VwLU2CLQRvSbj2DCCBBHLObef8Y1ZuriEv
Q2CcJ1G+FWtrhNVtWR+6fbeHmgbaixxJ7bOvThlMBwpNDDv4GIqYT1sxH2nYefWe
3YNplSMgH5P6iKuBAEMsgnZrgnMpbFOjIwA83g7rvh11hJq8a9rstLN8Ha6xZlnD
5V49yy3Uhz7CR1HAbrR4xw3GIoTE5/ItfzijTtkB6dxGFXLx6GsXK4mh+qVewYNL
DAMW1tAuYo2cDgYKDUyGbUc98wJB3R/R1yst1mJlaQNRMleCpwoxowkiW1te5RrU
tjN8Jp6YkI0ChDMr1g7q+rOKqNwc3+pIYvzdpnmzdKX6fDUJYtanuPbzu8AN58TI
wTUW9k35iagHJy5r5hYtcKtQwhF14jJDvm+d0Rgfnt0ZWrEFR6xp6M7pY34bNwfw
Mtlc9p3Kt6OQ4iRXsh3qYt77Xhg/K8EmFMHwPCiPot1snw/dLT9rwK7NTwXPIBg4
Xehpt25qPY0Dlf+4Gm7oJyj5QEmmIvbZEANqffm8GoG4KuzB1To8JvZQwZnXtAgP
g9ltC6bAAq3CLmofDdW3Csnzmah5pfPkThJXuqQQmcS5cpAv0FmpvS2d/cRyeQWs
rkJMiyx1uli8519yu0mTZ3Fw2YK2KDVmOmVfn01/AD8NT8jea3G2+R2oerM5L7uO
9bsxjnYEZA6LDgVOjlQb0FsV8DJzMqxkRmmc6xMzy0BjZSNT+663q9TUjbMN4WHi
QsRZcqlZah5FxKVm1pVejmydyjvjWUOH/qSWX1H/XUSY0Ry4GTRrV+fUe8zjIL8R
jRmgy9z3ENES/zexxRp8ocmMaNUsWRkY79g8n1KA5/3qHSkrzM5pKFDFzQiOmJ4P
rMCGwTIH4EE4DJFo3hzSqXxZWZjYxMNq5QOTlkFVpU8zLPo9W12BZTJMxfl3T3ys
Isd5qHm7niAaOht7HLQ3QEB6kufR2NVM8EeQ4MAtw4+Qq/J5zdegxlchr40tmyWk
Um7VzUNtXX26/CK8iyI2Q3AuructUkJ6OaxANOqyBsa5BsF0uYLFLcsvdVBLimXS
Yg8rPdARkT58WQHUVc8DA1cfB4AAdeeMCfdGGPDNtpYeyLYuGTMzvAfo7asRXBWq
0y2DU+j04GGDew4FIs4Ie+toNn9zN5Wk6Ax+WWAybR5Q2lveoK9kBhTrlvan/Ckk
0PkhfTTULs8wFea0pc+cyrQrKJxU3LUV4xkQDH5bKeB2r7tbGW9jOS584QQ/OMy9
dyfFcnSbG0sbqMmqKsFCOn3j2yseOEND8cRVFa/SCK1JRd9vY2CkMuatJmxE+gA9
sjydBDb6EwhpIu/KmZbnAFOq6apnFQ+dELMlOtCXyrC5XSMczZtDTmTltYKkQmoa
30WunqrDAYvKR0BmqP6i8pXIVUsMxs77dtw0sE32KPLoJ7FLHyB4oR2OqaFzNwLp
o2BL381APK5N0KI7RB8LHA0qDPKb5d4wKTpiNUkDY4QuFHQGsFDf7Palx0QSR3Cf
jloa1vC/qNwG8wKGAqtRaY2ZFbVrG8IBILpmv3fdyHDtl1CrcNBY7XQ7FdpIwY2+
L9rK+CYb8w9TUjY6OV6HX/gQbEGP5Zzm4fyfkU69IBalj+qRYWTo93hOUFgZRY7P
ldOWGKgoxwTygcGu83s3GFXw/KSNGcY9PwDLQRkfbIAZB4V5PQoVBrKiDY1/yBS+
8t0klHBD79AVQ7NBGP+SrTMxyPMAHi9RF4nKQYMvevT/b/E3t3vWszaRypH36dw7
RTxduXSnPnaKinjwseoCejJXuuJQtBoEG5glo+yokUbZiYAPJg5SK4YYxWQomw7H
0mAlhWYM39DbmMgcvE1ZXMnPBcqT9RtpzzTKChmjXOOSPEIX3TtflOnFQl6pNxpo
iX/05g1PtX509bQds0PO9cTuD+aUPDdWAXwQfByAQIyRvkWRYNHm88NYljPmLZsj
A4kuMG19RQvvYS9kPowyPRIoq8EprWiJGzolc/iB6KVPQePtkhOh927mYr3bnLQZ
Jl7itgL4+YztIs8dUILiX/ea6ry9LNwahrIl+hydZ8B5FDlksq6SR+vB505GkciN
8KknpHJ7LUTYXA5MQjolZtfw2Sk+albYc9pIUV4nzOKKeZ6CUtzwhZlU9N7RMPNx
X6lo6aHhux4DyO/dhp3WXK1fzcpYYeTo6s3lv4G6XME2+4AOhI3v5yfjznsUW2RK
ScjbY0r3PDizv5f+fdBF0+RggvUKnPJPZffvMd5nrMBnKqRKcMC6LZU9CilB0Ypf
Jmv2+h4/wXVfjJ1m1Ba0Gj9O2/7Y+AHoyqFrIYfqcALGk+BRz0fieClWXOKMEiec
gphVnue0xf62ot/oeASsgytd4Hfu7WDlNy6vnOH4jLnvnF4K6OF3ggVUYx4J1iLh
eEBRImNioBsSIDK03hqJAQPdrZrMjTNKRcXgihDXAwgeOssR/7tL3EiB4Sg/B3fN
lPYIx9aMls1bxPaoFbOd9/qnBwxD+DOSj//aPMjr7BjONR58lWaS204JK+0X8pFV
xs0xOSLRlwh3cRpqBbUNuQKZW9vi/BJOHJ//2iU6kuewxXhgzfW3VrbllZg4gsS+
67iQmErMeJyZNiF9F4NSTeEYzpI8YX38WqsMje/cXjkRmWft6fnZHakEApTB1UsS
2YL465K5rhW5/wX+sWF7Or/ph6Fm/b8aFSsgESOyxNL9Jn9rRVHhOUgAGJr9M+5U
R2TqYakufsjEL1Ty8vXwe5iybZVKCnUKKy2MgIPXvUcyYEKCaSyrAb3mT+DAwqID
TixRSjj6/KthzOJmTr0fjfZshl+nZlb5+4UtbwZ1sbqdArWEKPMk3pcGO8BEkLrm
WREiSV1WkaM0O6l7aGG1wokkdHmdKq8VZwVmyqzs6TG8/xUI1cXOI+wkWCKvsLgc
5otJKzeoEL7hhN2tY6zdNQUpcWMnPPZF5sL6GZ+vXPUcWaPBHk8QyMDMf0mxgO+v
ueHNNONWdcKH3BItxmbafww4PkqMg+XL2r95uG1RvQecfQnroS3Q0YJTIxBHiJig
YDktJQOq9fFzC7C6qSdKh//CXRr6DCg3tpONzJUsJmPTNvR02MjbgYuu2WoOZF6P
T0+OEhcusFbtBX55nkI/7a/gzA3kdlYdxFdqxj/DuJxRf1pMfcYXEL4p5FkcB8mp
QuUPR/KebCmHshqRlA64vB81JUj4TGr1llGC2PwIBngnSPri0qwGjy9j2qjlzAyZ
WWTT2SU7plckasfvCY1J5RIBTQpNj/Jw937cNkUbHhxuMieXh/Hb9QwET1M7/3QN
MSzqBCgTZlg2OyBHVtuFWXOv+zri9QsNwxXYN8YH4Pub8WBiJPUs3lIza1zWn5ku
oE3uznf93G4XqXkKMDWrQ02u7bQ7nt2mneub1zbH+w8PFUlqMeO7R+kFjZGy8l6C
44fI+eX7vegV/7KhfVZ0CDOvBMjrYrct1gDjJeMMrNvy4/VTqXc1guYWTn/TTAvC
chiv/W9ZOHATu2RSONKUB3uJAJHFC+jtvLdPbPMttYRIWvif55AfiVHXhFNRlAUw
EEDb+WlWkJddponxuFkCSn+r0+uGmKz5bAlvMS8Pa9WYjATLCh9s88Tpm80BnYsN
1+RuSgW5X3c3CuFW5IuWxpG86HauOf9ALkSmr13KjIW8wrcLOu55VWLgbEK1k0f2
5dQFKa/12lcvN+g6wUicOD0PD1/5xmt75sMiClWKQEpxFejPk7pPgZ5mIMmsq1mJ
aK3ER/E5lyphAGH0hEQ2wFJQ52GOamcsN4E5lr1W3B3meOHEp0FF+y8JmsDsoSc0
veWiY+By/scHwBWVyL1Tr3FPSQutyHxV4dYBydvzgwZrTa7jjTsq3304JqkrWzsV
PGSYAAuv5RZBsDuvRUvc7AZc22BI7ObSH34TV+wedBJ1A+qDwj2tbVXkvDOgNyht
uDA/H543PxgLx6g9gMUhOpi3GGwrnniTRuKeXnmGMch2s86uxjEwHl7fubQLms9H
1AT6+MLOZf2BqFTTsaubxHuIZFSDSwVD2UZZtyYbWgdB32pglRYmv3cj66AzRT1o
ob4jNBFbYPZFmrxvotZ3VgTkmcahsRe6yWv08O7YUpJwMrjK+/Ql24f9NGCYo0ZU
rCRBRZ0CoY7fWDQCPpX1+ZDNxzDJZDpOFlduJ98BwJbYADlx8AN9n4VCgMFrPjG5
NOshBVrIcbhfPlC0t8n2GmPikAsmOUhOgdQQCQHDQiM1m4p8MPo8poPTmGG3AxqM
iqAeN0mc6kmDlWdJp0XLAeFrqgUxTzEaOCSc7jDsys6qvWP63IlE8oA4+B9DeWHD
zTpvtaohdo9yj+vZoWZ/6dyuYzpBoNR32sIOZ4nUXoitbG0WdRt/yZWFqBSRVYNA
FGhvP263PFQijkJ5UHuckBgj7eWdQJxIcoxIJM8vyvcMxFDeZUihUjMciW9y2bRV
Y9dVVayz95zHYs9E3Ep8Ao8fSIRmWZZ17sZ8wUjdpd4nsDw6FkrQsa8H1rv9Ieg3
RZE9Np3vU6cfENdxKAN3Td5CyvZCOEh/1XIhBvp/FzbUgFJCIEv8CPz+KJn+wKuK
ndjVM26lHym3wUEHz7uyFPUPhQuK0biNXs8RJIt88nN77UoYPguXry4s+AJhE+sg
zsxhnm0xSe6JHhhcJoLw1TsKS5hFEMsQAD1NfD35483Mu5x/tICWB0rm4XS/B7JO
SevKapu7TNt3echk/cP+WxPz85jXwRiiAgzslYiXvphTyPOX3zrDxnEzg+soIYA6
9bPBLYbtO2D1ldwEWAdZU84FFN+2EJkyiA16KxTqo5PlgPZb5QMiHaw0FUs0WGaD
rHKrRIXf+xuz4lhlPnLZF5W8LMwLwQjJHygLUY3wmZlrATCQt2pGsawYHBk9pqxJ
AF+JGK1IuVFvSBQ5i8Wv6EToQ/AgC80r/WgDoLEu4m5G56LjNhN01mDd+rlBo13S
TpAbFkdrutsSUihW1fmxxqC0OofMmqOHppCbesoIasdX7fI1L2QRiSP7hybvNDBq
wJ+e/QOFWxrXIY3TsY3IR1jSlg2Y2XtLDJsO8QvBXt0xJOHfeEMJUtsVjFmGU81o
i6IbSS4B6NuYP/ID6AQux7+vtU0bPpY2ySCuKdYZzowrx5neM4a5z0psgBA+Pkrn
t5B5CVbkQSGt5RK3Use7Pj+HXlgiPnfEIczobVw6skAxbZEMtx00a1CWxH24LlmT
toXibVHnZMgETcoA3hw3sOIjHf8MbFSx5uDeFWeFbVVO23Jg3k2hZs2Ch1EnBiiu
Jlr6nGG22YEUyTTUlNW6gcP2tqpjiW7ExIfBznPoVkTsDYLuPLHGAnqYbF9u6wk7
RyWcK+seu62drvK3ITgnNw+JMObOCI0FOiXYzK+fpE0ViRwWq1LUT35y+5+ZxzSM
ScFtJfCig5lLZOQxMNvT94D4p6ioEmqpXGqZkbXUzRDnLKnXequovY5LXlkTweSW
BagXZEvQQzizaM5O/OeV+JV/hXvwa8s8fRsFyA8JeEqiZhzCe1mSra74nNvXc81Y
EVpWUH8mkTK79XlulcgQ6LEP/AzZvAiGq9nF34ZsOiuJH50o3M5CqTBkNbyv4ZCu
czbkiUeqgLDOp2yrAjl3N0StL+/B8mtdS75FjI2jCCb+8m/m0tT+sZMohtAT7F+u
6XpkcA+w5phFLH7Xord2TOu/Vka3a4H8kjAeDrsXXg2vcqlbBjEpDB0HI9QEQBNj
9c6V8G55zwkxlg6/7vkgowx56cO/JmtERdX2uExTdR1eqgbJg405hmgl9RkHcCWb
VylhJpsDzR+NvjxPKtDvfKlZLvs1XWpwIm6CIancF0KOp+RUH/j+/jHC8+/DdUUe
60aiRuEiZ/vQHB4Yah+OMzazBkFzCNNWfyFKWFPjBtpZ0+WimLDMBJUD6Ymi6Vm7
QOmYCUhIjWc2mRxHVUJdojJ+FnfVmz1lWFcttllEY9qXAy3OoDRuk95ftln1j224
IVFNLIKH5D8/3XjlOcFPYKvNXnMYtw3YRV/bFiryUAyeDl31bXbdIg4PGzFySUiJ
7uAl8M0vcr507o+7GB+CiFr19sxSLVlHwkFOUtlLetAAABQ1y261iu7U4aJh7o9N
RQdWBxhrpxL1tINDSRm0klYNlpKKq0dE4nHFMLQ5mCNBqS0w8Y3x8apUE709GLPN
Yfhptyu5oenZ/O0+YJrn6ldrTr8XbPBKjMO6SV6QyKl/u4N8YIvg+4dzqASggfyI
Xwc/vRxeBDK7w2g1nHYPZ6I5Uq4epqAtmNN18X+Vd7Xc+dOThxel9CQZ7QAmwHtu
PpSnQsUqnNuNDhRkt+uNF6XpUD3x1senCM+2PglXXYXAKjzQfmDeoWgbEkvDyUEg
O7qjS6SyxjnQFaY+8yb3dW/8eEQ+SolecNcp+2g/lVwyRw8s1RERrkF6f7kgitcB
1gMFa8DBLILUCGa+T37057zDDosABmMuk6WbLgGY5a8mBJ4lKGy742g3f1qtUSiE
s3Nmnfzp2mLEgdXDVXoxR0ZdSy+zRoSsMIlFVaW25sKuXrNXlkoAnaeY7Q6DJR/B
M+B5lI/b/WGA1gJp9rYwJs/WxSrx+gkd1w3+7Cf6C03ZVbE40VigQHb1Wp6uDRz+
3NCLQQjiGPJh+df0QdviC4jFnkfp2marHWXUSMMzhaeSczhF3CMfyMFkWasw2m9m
4VrIoJPI+I4L35AG7hwiLTHwhxWL/Jt61jJuXxZNxMDtAnEZz9xE8avo5NzE+ylA
TRcyUY070GEj2aoRaxjdi3CTk5FMFlDL9KJD7679VOSUva6TUV4fFSKJ5mQSGfrt
HZbO0Rfuk5+my3J/y2YF80gaYz8TSUUv0+aHxJHqlL/47FPLCW4Hsi9EH9yXw+FR
rlTJKW5X/W3X1+pa1aTNzzYclIIGFKZupOc6176I7uQfUH5/fRZHBMQIaXq1khmD
3OqFMXOcK3Q8iOV3QouoCjIX4k3Bo5kuw5EGUrC/h8KZoqd8djA3lQSZr2tca5MU
9udbWLFxiO0P1lCs9nl6H7ZBhAeuZtWzRS4211/pFADzkZIqdV2xcEozrkG9hyGv
RlP0s9h4YLf34ZGjy110bOYbekmxb+HtnaN0nW25Zv8k0su74WCJyU9gLvimlU4z
UpDKGuqYP1q26rPj4I1uOtLtHTZRZF184qZt4FTb1dypEZjHddRrXDavvu7sJ4Ev
qVFF1+qLjMREjsK7zr7vbeC6PKFtBZ3o7BVETzWiwoIMclvq8dn6Q3xfFM7gNkb1
K6zaJKA680C6mHPE4Dp4QtJPdVAN64JodwUGTEkUV7ZIasmqm96fYr7sqSuN9VY4
60937CT8x626qYBjHSNVhgWKrmcewQvOaPwdTKuCOsmEa0Hs6vALqqtOu8aWf4RF
AGe5BfhOLITbtznkqiMtl+9pB0j1vuWn8dsF1YM6bu7yz8sH4PzNJZxS1IRlpHEq
CesTQq6EA/G57JXB4eIiGUDzgV2wXHm0C9fTh5XzHfxDCnuFS6+J8loJJZKVbvmy
SGD/ON6YjVdOpONV1GAppkMIESAFAlRWEFBQBN/VHI4OzvNI+NMKXBPrB15VyTmK
tEp7uV4L36B7imeL/SysJQqXRxKAN4Qc94YQ7gMedP5mBZvlfnDPJHigB4pQVV8Z
P4cqCZcUPk3yWeg2aOx/KbvH3MV+hJQxlQeWRJ4teAfopwEdSLiDLdvmXdD6CC7d
rC7GX+rGVl5+wgeRXPDPID9zycQG3R5MoNOhxbL9ozyhFgk7rpGd8ArKKeyLuHOh
RsMiarGFSLZOBjfz8/Zt9gAnYm49/DmiYxXXGQxpWU6cM1Pn6yGjbXQdMm8xBD9F
PizFAxv1LMLqGmZOq2aO4k5BmXEtIN5TEEcnntg1vsXJGxUeolVT/mvyNtj3wLgN
kT3DSf+XCm5wdwxI8BzKXYgCnlIyVl/cKx+khL7T0ysfe7+jLsDzXOsl7jM+8Wto
fsoqZyJnBwmZ+PDzwPAwkjMCZ1l9gLEmP1AcnoTMuEd7eIvuzKeTqlBFBxmx2vO1
G9tfV9xoGlqihNHiiyFZyl7L7iGyvINTk6HV8Gt6eOBTlr/KPPcez32I6zE+vP3E
aP2as2q2WeoioERpGEJYrWPD3Y/UTyRXQn3dhK9fBEEFqPXSCNkkEIgF/k25Aed8
zM7MlXk541EuuwB1pX14gjhA1aYF8weJwAdT6roOUK3ivzKeL1EXfrI7Ix530kQ0
4IQfjitIDe2SzNc1RV55i1P2Gm3a2ofxV9xSkuMBKVlA6EQKLp3NIMztu3JPWDso
46c4AcRx6N9MAiD/3kVFOp4ZCrxu2Mw+nSfWc1KrgKOckBMst8T1KkG8rXbsaxGB
rcarTVETtrITozsc5N4ocQqCBP9Rga9irE8ID8XJxa73qr0vDzAXFu/T8HI2W6+H
CDSlBMIVo+WpGWT3R4REE3TlmEAqR1IekE7DeqhHjpWRHez6MPRiJe7t0B1947S8
Wx+dks0UlmTpWhZo4/2u/LIkSfcWWQxxBTphhl0CdL1s2y9p9aQO9Z8Yg74X5DV4
/TlruTW9bw40uCDHxPMZjAxpsWlAdJc9eSBemEnEh1CFTmWBPvbE6f68tlqYr0OQ
YAOKCWHYlIdt6N9u1btS8wC9Pq3CfuZHlZ4zkGBKY3pOybVCenwBuphsBFCwK8dA
h0HYrMgKrABkOh8JvhhRE9TfR1Wc22EdZrDCz3SSe+PqXjr12y9XfYn4t71PNzT/
iERmWZw/LAYDU2i4qxDDjuMREtImUrNCzlaXnzazGP3TKo8F2dGLY6DqhnQIwt1a
qBWbiFJ7HgD84BQ2usKa7Uz3IkOykCMlLMAoYqbt8D+bUOrf/tr1n6Qml5BK8ZdK
RWr43i5wUeUSu0uHDnURWQixfFHgv7qHLRPJwnKJ+7P0UuOSjsQIV316cCUlL0IH
LGTI1DDbPPzTg5wfOPa0QcoDN8+kuJa8gHFQdQOiP9hOOJTPW05/K6W7DLOb7T32
l9bUU2iFsVOEhHsf0ghlUQkvWTwsl4GBSo6jxYk6t7huHIFaBJQJTVdEjidNTTxN
7YpCD7Ze65IlSd0n+Oq4Xcg5/qVWZeIK4stPAn917HDratvgHBjp0NR4bfVYWsY0
qarm9qfyfBJouTaxc33xYFZ1gIV1OhimTbDfmSHCWh4xe28VQxCvIlqU/0hxh8ul
587gmtmboUouDqEgBWTY9RgApzyDOr3ulXoPYHNOyXhJNZcOIz1w9VVq2/KXHcp1
miFQ8WQcY3lRbQFlZLv6tfoYky9HFcgk038nuV6SdoTMiKPIUvKBm/P3+lvRkWGl
ZOP8mBxQJZnq1nwSdRWDdaTAkfhg2uGwoImJXLdwAURlXfr3n03XVE/juMFy99SA
V9HXo56g945VvMj8N7I//7HsIpAZIM3qxpS99BWQPdLN6ByE0pHcoHgdcUjpiTjG
PyvIb4NQ8ECawVAd3S9EPPc8Mh3FYT0s/QgwmMFVdHON2bQsxpEUHBYKWgsnYvFl
Trp3VDcPCtnD5MTWV7bxXq6xr43hzsMF/gjY4PcT/1kXJJcc65c8Tadv73+MxYyO
taGg6sLzndfyL2mcma/owmeLrWqGbi0iln2iag+uqVwMyRTF/IaK5BFE6aLqIY4n
0CXEMT7RYCzhBZbcv2fvGnqxmCZkZYuD8wwyshav/jb3sRzHdT/pQHBc6g8MiP9Q
MWpXdVDsnKweGuJml7OZpj/PT5NFouZ5UThEmj0KmEZv5opDrCKg2X48MZDQAksj
TLjq3PUI54CNlh+NtR5sX0nRvsYecNguLej52RNjzm+iNMnnUb1j79Xun3XmaMcg
eAO4rhR9Y4zPcuQpqbMDXEsygEPeVi9JPWBEnbh9lmA8NGV3kCbylc0EsnKZ2qZ4
/zylmetuy99Ij4ByUZukrYR2XAer81C5A3ZONoXSqwz9Rlzw12qUSsbbphO+pnRa
CKKtosj1lWJMp0ek7cuhMyRuBoMXS8JYuAikG57aMYjzZgJJ1Fw1RyYgLa0D7Mvs
XoqcQKZRcdFdlZ+ShsCihObzGHy19omxB3cK67BP3Dj84kAgZ3zFRMOl1ngtyHCL
P+fBnHvA1vgd7BOcrppeoYo8M1u/AGuc/UBBwFYM42it6xaT28F2NqEdbm4XOyjc
DU4BTwkwjHokxm6sNhmw8ZLfnmI37Ppqnxc2Gr/K3Sw3Df3TE4tMXFfpkmHHNqul
Vqo5xNeP6gGZEK9uJR8+6hdcI7O3jd065gwnYaxsnJ4XRfXwN6WCaKG4m01BlQMc
c6KYtuL7uGiDpA+cIGeHXt5MpBK30hKY6+bCBqsvB/ehro7NYcanjbZ9DRYw4u1p
9auFsvXd2/bxMvoDrd99K/uEZgQRSyIt/ikWfMpBHq+tUtU6wgDmiGRZZuKRdWuL
G/d9pjlmWFdc6Xqz5XoscWi+EzjyRGpdxApZMeSng0tsvWhd41elpR+2EMbU/wGE
u8x0VEHT2Ut+M0WbozKw2ylLcnvcZdqOPQM9jOLxX8kIUwChjME83onxjHNWS5za
cGAJLU6/mn8O8vhMfxrLGgJYQnX8NxP6IttDnQ8JhkBEg9rkc9kt1WzOhVhTsWWc
/c/EZzz0P0ls8fM70vPInrujE6hSas9zdpUFGcpRYZuYqC1cj4xPshHZ7m/tIn+K
OI889IknfUJ7cm7OWTS87oG1g7sZSWJfSoDP1aIsxMqA2j/Rb+wLs4XvVLvNvIBA
zSFRB5bqOjP4ZdZNY8WHJGWsvoUCHBaFKY9WVvQQrFz07QoOUucbC8d7KayB3nTv
/nu01PFnBjNdhvqntNTw0hPYj9XbfXpW10t0I9l4rj5FszIN/KwuUtONDhXGusQ+
dG++RaHxxqqr+eycuUqOv8AP2Kn278kdoeKW61iDxGbmeVM+3YZiA7/lRQ2DKTwl
th3TqI4IUM59E/pdVxUOayswOl4iDjv+ZgIS1MMlFFxJ3SU8bgEuGyTLY3B7Bsyn
gtOTeymdxt0xq/TF1yAc7AbQ6sXiLmiMRK7Bi7bcHUp5+Q3DFUOwrAKi/vqd4xM1
9wIQmO/o+V3ST5j66OwDdhmHUutXMLLRdotuA85bB+KPNZsaPmJkqaJpHictRTog
4CFVfBgygFEpvU9Q3g8YPE2grhXS9CeKsIkXNsqs9pZ9GCx0xLCfgkXT9p108h+4
t7bkYxM2F/eCGABuEtv/XWcVX072+QbhaFE+zqAO1GqL8yalOWObYfSqYdMVQlKq
z/Hv0DfzVV7SzZ/jOnRCczsVqHHjtBjwUF3RYli+LxhpLit6cVoCbG9JxBQcJsv9
x7rAbKYV6i04JC9EuA7pjR99ECo+dqM79HT8Aza5jPNfzobZ/Qoz18QMbzSdDyCT
RC2ldmw6CEvLi/kchg6BgSdwkzB8kmaRa4cvum3iS3/DkOVDUA8Didc0Kkws05Y6
NFu1krE0CgckzDJ3sQTTAbetPbEMfK2t1LbEGz0wo999Nidadpbqjr582tTIEzTw
PCh+q/7CZXtjeTIcs8Qt6U5eGrNZ6zCut+oIH2beVrRhOp4EaImIijTJAGik3wQI
Vp4pyvA1VoR78kmTpSPfQ9D2UbF/e60TgOz1H6ewdOapZmJd1v2X0hhw0XT3uzHU
F9j/c6eo3pfRcMO4scYKTC/kiK00+Z5U+oV82l/Zf2yWx+ubqqz2l9dLMoDwHFnZ
Jwz7DDsBC68zX3oWbWIc5uTLbNyHbwGGdfIKDJAKnirGe8Md0Socp3jKeOYbumu/
B3KoqShwdQ/ow/xnTOpH5Oz/tV0SdJbFx1U/4SXxETCqEWiM2JRKhkf74asJ/HUa
qpkxYoN44nauoYI1OsdIwK9mzczFEVPL6840HRWW+6rwwWvRAH/zCFxEpCdVTHfm
IfM+xlNS+4yjuoDho6fPKU7KeNZMWMiOxREXRiQSeJNrhSpSoWnZuXXBekS8HKw1
OiZoe374d7HSqjOaEqjS4F5bTcutg0saFf2r/obaysR7/3XJTEgy33GYI6xlUvvF
cz/+EC2SysaRn/fGtix+8OtjT7tFQwuE3RrCRWamZ3LzlCe/5x96mfFolofZQkce
LkBcNH/InFH94oCY67cIMKxr8/ULcIn1Y5uIzdc//mpZdUUITO0MshG6iqqxTvt4
mzl9FjVr6Wp30vuOlzv1rpaGEYhhY3viFY1JPBZy5otpQoT/C5bCfPP9kO4N26YQ
yZNd88FF78delLlsTvyhG+JjIsbuPrulf81N7aRjhpK9Unye7kxOYLLVOBIebW6D
u2GGuCDdJ2IJBvt8Xmfn+jWGZLcKMexwe33srSduLZ+zVyMHmMxkflo3fg8inLUb
MdjBnJSdNKNFlyRrQD+tpfhA2Cwpi7HJUKaQmHYP6ETmj4PBtTh8Ff4gwfvpSzkI
jm7YUiP7t5zmP9maylebGCn8m8ur4wjfqZ4sTVeqSwKkH630HVxZQ4N7EUhGT3hX
REmMLk0wSlh/ywrBrAkJIw77icE4Wdxxe/PvBoQFVl+ZADV7Kx71dM7XJGglenBC
3O5GH8p8WkVRsj1NZCrVbQ8mGCl1U3/SjUbMsF60fvfzso2B/oWAqJ2/CcVutlcd
9T2EzWrnbZlTqX02HE8ijoAyulFnbFVe6YSNu+bKp4IPt9scswbjep5XIGIofnIi
4hwkY8rotB+iV4IzHq2v+UiUAwnHCjionYgOOyInx8R2mNPpRT+Hgc9fh/iY+rU8
Zeay9+hFqZ40/7c81oDP3nky44OGlsqWzv0/8oFftt7Rn+L8paO767sM+oyVv2nT
Vks2MMnd2HfD9WD3Ah0xJBLVYbc9wNtO5O6HekWSUBsh+qWF8BBFCsUB2W7bXedQ
gjPMVERB3rO5CXZUL554A7d9010INwSz0jTAXjTzwoEHZ6aE+CYMv80J0znVwbli
oEWeQ2isRyFXYz6/LRQF6DD3W4jEyZKAlxP2YBrXsD7grKUcUV0+RbfwpUCvT3VE
OgqXqUMsIoNdH3R69SYaHZzXPPLm2xj8hGgjfTnBsIrVvpkJiCcSUlcDa/MZArzF
js7M2vvxBv18nf2mEmUQkPtif4IbyVpOp+2vhqvM/9JyFBiUJgrv7BK8yeFuWBL1
8LRfxOp/Z4/+G187HRMxFmENaRDbZB9B80KKLS8uSCjHTjJLVaefiivIfR9S5eqb
j1zYYyelGAWJUrdJGLdbqAFwH2836kuueUeLMaLSimYPZAxWSA41zZ7QHyGh7w5v
V3vzoXxduK865Vp2daJSfb8Wiuga96FSpfLNFPNHyA2DeXBZjddtJoMJOjDU2Taw
OL4U+llKziUwWnmGqur25UIVG7CJ4ZySmNt3hUU3uspaCkt9u0qWBnuuVPDm/VaL
e18Q/ONYxh3A7YtRVm/ZPvuiov/Ch6TZOwQIFZVpd8sdGhhAVwqXI3Rkiur1BD8r
0GBNWUn7qN6MjXS9HEzWZfUF1svw6rirHxYoZrPDLIaPLt5o0yACnVQtCHyjA2kP
KSiRGrkLD2Z+rS0PtHlynrvZjxC6YxPxWJoTXZUhm81BCixuS0hwZKoRSA8UAIZH
9rnHiD5XRdkCu8jDOC1Z4UBW+gsJefa/o84IzGz+61EefFYdLgvrizNeFuhClOzA
VvcpHfG82Ph5HdIwtU5sP/WB/K2suLrN77IPHolQ2syn4FPWrxPyAdDdPoBRrfBl
OHmw0S5T1ZsBU6OcMZhc1+CcRcpIqY9YnVDwDduxag4sgWvcoaGqhm4lLOvvOteL
nvQHeX4BuHo94o6bkIag6/4b65Cpz0RBKfyByfjalYccYjt9Bm/0Zu6VWK6wNyb+
4uoSDFYhbL1FrM4Z2kEaS+J5oVhx8izcu+omrbyB4KRmjG5ixP4/iRByuU/rMqqb
iynGzDh0/J9ikE8gaasiTEMi5JC6MuQqHX5UxrVJDddzhTDdYlv1NO2440rToZyO
4L6N6PbwwgllSO/3ZpYq55a4UUrBZhFIaJYdWSwptw2OlvMW55ZiNGOOV1TT0CI5
8iqqQrfAd98rlDlWf/uUbB2uRl4ie4bcwifUb1q44pFf1GNZ0iQSEFKHK/d+dAMp
R8bSsEyz9PFtCtvyqXDAMucpqwh4vSzAGFrLva1GkvCyfx4eRohYsUZWm1g1MZU4
ligdmBkef2yUylgcMzn7YziMHobu9ge5ItX/oKWe/0GStPjzxNVmlruXPLQjTOvz
58PVTrYpp2yN+F+QjpTUbhKDEAScqSOJup8DtrSqCstbDWQHnNLA4eK+3Ah8RMgW
Y0PI5cqgi7F97x5nAL8qICd0yrzH+WoHilM7ewExbuNbhiHf9LdWVBEA7ydO9v1m
T8HvIBQqBCDVyACOSosHJD0KE53H3uMqJEwlbeLSUlOCLsj3Dkln4dzFQ0qJakDc
lD4fRzwdn8BTo8/uGQwzPM7CIKT8hr8VG1YgtyYrbx0p38oaWxtDmw8+qL2xFfRS
h+uAmi/gx8Wl926Uj8L1SiKOxx0WqGFZmIOQsIuY1eQJgplT/Ie0b7xI4ygJ2p/J
NPAbFidu8EwEO7DwSlgKs/P5QbGAqOFHAD3sin2H58Aeia9sFACHPIPvr3UcbiCI
d2MerwMFqLZXSV1ZkwViFopKhOpC09Wk15S0cr7IQbvsJ/eS6J0pkyHuziIHYG/Y
87L8poH7VM93Hh/bIYG6ekxsulM3naoX/O0ZmE2Qn9lutS/grsv1LWAHb1Qhhv2J
sePyL3iAm9dBxrOZ80M7WfKLwhwPjg7S83phygS0HJkjqtlD7k8av4iA8MTcLf+D
uGr+btiFIB1Nr56UcD8MIvHDTbgxg5z6maOGF9n97fMKUMWjuGcMgSA/QCmvj3MN
aCEkXqhKN3itRJdjHD7z6gEPlcLG+COaap/8yOvXQLf5SY/6PCrdZoS4ge0YnHOZ
9jQrCeDIvpG5uxY88WQA8+X49n8B6Xdx2l7ldFnGs1x6hDvlXxs+EBs00F6Edl0m
vYjGss7T2VN/i/ofo4B2xbgtt8nbNRRpGVpn3nc015MJAeZI8pQGp/stiadjGtOP
nh3gMw2UAHb4f14H9Hwwt62eWRjk0cT7XiqmYHm+7q3DAWr/f8089VkQT/o9+7iK
fK7JiFkTj/aDmUEQ3ZFWdW3Map54gBRZ+EYIgVJxDJuFgi9lo7fvVUfl/i58V1D+
iBvMUAUQhCtAuQPqVhiZKuOxPoRvUH9fAm+f8w506IL1fxZsEQQql2eMZJIAMzSt
1OZTkvE60ZCm/Gm1p5h8vxCYEdujgzKj/KCFdHXZLhvxQYe/MZ/7CaMymas1Ehc2
9vlViwNrTm6RoBEeOFWoDR5h4TO1oXVpkJ6n9wzanWQBv5pLfrcv2ItqIMgRqFUa
D+cAdPHsAQEsylGdpyoU/wRRdxUiF8uuezf2cj1mWXSaGb5YBYI3otY65/cegdYT
iLxoFoevFtimft/iGRaz4FvZZIYbX7MfJTceTO3jtP0ERX6o8dFPhx3pebL2YwhO
M2noTNbxY/8jO4tsHCgHLt7yUnGGJClZUTmj4m8mC0XhJx9XAxFoFHfu6J8PbFXG
o6NI+B+tt48w4VHiZdY4T+mXjirZz9Fb7yMSCYGCbD9epDKnToIWBXNCyLtTpZA0
v6UrOjaDdB4TB04qHbuiWOEweAYmeb7mEo8BNbViugHsjixX0bj7lzoYnF3Qdc6o
Pbu/qqBG67JKtGahjqaDR1iy1HHz1rXRkjqD9tXGqTSE1BUe3aTQN6TFdT3EsCgF
5CW4G/Hm00uNWrVGTeSNxNrc8wdw/0WqPfKIyl8RucyiLQfXbudBny6jdSM8G40Z
8A5PuK7nQeWg488SpW5JJoAomPrwNDxCUR/SfVMjasRMVaVP6ijNZyjMJ9wUWK73
XrUx8nbrLhGvS1urZfWyVlxcJoqnRQvdJ5/8UjQjrOA7/wpOJsLRsyt/A/mMtgEo
tb48G7xbXMwfY8ULtTe577UBti+3AGWfCSMGNqEVXxYdLfkBqOzVo2ZTnaZzVCIw
aeWWemLYGQi8JlsaFYJUp92zlnUoLZRHTovPSH38LB+aH1y9a5hFSYX8oQj350q3
h1AYCnYxVQxjLcqaH7abpSnrwNBQQPxDFI31QtaDjD6iNybKncY4N9qAyXxkFouQ
2uptbmx4zc3ShJxzEWJeQV3hQvzyjO8/1i1kGYVHYghd1ShYFdOYy83N6yKIImfj
DQtCquSbj58Oh0RxjgwuSPd9lY/btvDB+1xYu380Y70dHOTwbAg+s6H1II3IkV1B
XkSsJ900n/8/LDACFe1jZYQj9yUT9eRepcvIsuwQocAK6mh+ySGxw1Qx7vMwB1lo
jwYmomBjhPFtId88vMDrY+Cfh3FCocgCRbp2/WKgD5h0Ke70rFl2qs1/D7sPGvyR
/dLaJXdiwuZJmddPqd911IjAw6oZ58oiZQv3bBV3CQZy5Qfvv3/8dqNqTT5Tqc2I
DqProzyHT92cTRYwx5uf9N7lN0ZhcgTlseH76UuVNjrkKOOkZBmn70U4A6NPxSkX
qmOmbhLohZNVkR+NTnhK8E6I47VCcO3Oy6K+qeTUMJfbJPAoWNFYGqyNIUmA9sKr
JCtUSubNF62MmEkfynI2i3mTDpre/Zy3GPjzKL4EbLdTxA21dyelk67JvjgvqmB/
+hw414UVk4gvna6Sh33ojPQcNetmw5/19v/UL+L77oqvTlX8J2kl8u1q4zV+AR2s
2khJQygILKDq2j27pCorXpbThJJxZ8Ohd9y4AQb491sm7C0Ll958I5U1mPydWPBr
7+YHUIYwuQgBWjDRsyyhBo4PauHXmSI6ZU6TtM+HJFs/T6XzUQuElCujLNEBqn6X
gVay/tFaV4xA6A9dfwUAuvsdymRR6DabUr/wjL7xuj8ku6eUC0Vul3gvn6qND3BX
hwy4FvjBkrGunw36WMsHbkafeCUHng3j207yH1oU01cALXlKWwD0q4FdSypPZZSh
f5aaKoMErPaP0dgS8O8MR9X+8fFA9m2RG8rsLN3By/TB4lplzYhqlVbfftdRa2Le
aEHiMEWUG1htftTcpXRPluaezfUUc+sMFcWj19dXrxxT9TvNYqqvV31zcWxdxoPv
oDR6XrotkyWCUukFwe3nCl22R8itl6mpMeJbTHWTUY88JA0EXqvJFENtx7klPfhM
urJj830riyA8vOKdmvT5S+qrDequ67z5UGYvitveTX65F8Pzbiwys80YA15ayIxH
kLmi9C1aUJ7jn+npTUgXmbYG8YGARZHaeDJeJdEDy+fIlWLKD/hDnnWef3/4HO/F
yaohPMNqkfv+KYXwix7JV/OLtamIjS3CgzbzZy3YmRIEQnnb7YYh/o5vcfB1Scwo
c3SfAZv3BygaEuQWzFBmowc+nDcFBUW0EaYPtP+rzBE6fJGUfDMYPHYGsJXOjrzv
pC1o6YnZ0C8c/g1+U6iIJsNY87SH2my8jN2QY2uiIrdqC+rzsIVYNyuCwZxBl8n1
A8+YbuSn86I4awD/rsJigO5nbXZPvC1XoVicaSKm7DnCXCgdKPg4D5/WQ7FaRb+3
JSKwELqS7PdN11wPqYsUyRS2FNu2mAOH4zgjfSHvmPxOxeUGcEYsJOfyNQMUQPkz
udMSITk6UQrRku4MqGnCiX3CNIFITdcqf3R8YnCT6ukf4AnQ9AoDd01derjLwX3o
tCuWuMab9lkb2r8HfyRTM+Xd/H39eNje1J3mggpa6jtznbnuKnUoSrcs7Au8FH1+
e8uwR1ob8wZOd2zXlh5zqV9Ixb5dlqDSx/m5Ltp+nu3Du20ph9MSG+zVXqDwAhoj
xfm0UD87emim7Cdu1w+RfDFhSbQgkS2FNNVopbgOH22pNKyVtvRHIaIYItLFXvvm
++cyQo3qa3jaZMUkMdpQiD3N8C7eMZV3jXOuJCUQFEAimdk7qb3LcLiveP7vejP9
bsav7g/8TUwYOZMP9l3NaxSpiGmdxSdQSOG2V1DErf5wHTwGwdaP2WqmFUlfn9A1
E08vJgDPpH5Xjx2Qx1xZhAkcJ3kL8Vb47i1OVT6Kqf7vFFr2XjjObPP0+xyNoNIg
eim8s8uxs0NKbdP5p5I6RK8hGfInogR83Hv5xa3D+zAF4QhT1HuFthmZoZQRTdLJ
qQJBYGuWxD9ATYLTi+23t2PqwNGcmBw53ldSkanyqH6rd2Vg4k1q5/FLfyh90pMh
xODmcdc6pSYToY7QVL7qjTA7kd0Vk/QKoF4ksvWWSH5GmwLp9kkRFroxUSJ8JZ6A
zoAhVIfDVjue8R4x4NS4Zz75xkHKE4tYu1RtViVvmTNuhFE0qH5y8QBUWWKx7n6q
IHpqwu+aYtjG0+URq06L9GiWO4yQ4oOSlH2IMxjqSHG7nQUd19S70sid+76pMmfn
z5bXuOMup/owczGcD0sNjQyHjEcSqWAvjXU0Xgp49Km6g6/l64MJGA/ilzSgmio5
U28fXDw3MR1ns/e/JbpJUpdkDJW2DpUkAgNF1WT/8ISlMfe5eQ2Mn+sypeJHMzmk
DPg2ZCdCbMdH4ApBtzysOnVeidcSsHp0tQTPGr0hVFo3hfVr5o3grmh/7KtZB1z3
kL0b4GomwowCUcC6QXMKDOtRoiH+610Ohu9Oxhp9Vm/t/B/7BMnCq7gXNqU7NkJH
Kwt+J/6JxqK4yndYtl/pJMP/stLeLzJpi3y91inNv6zSJz+tl5YT/b8Wgv5WtVrD
F0U8tswwQuNT0n7I07PHc8DbwNtlgNT5iGw5zgTMGYRJmGiAyGbSrBVnh/hj9W/l
ERkUloGB6jpjZqHJNX1tSwwsEwxGNNUxIPAwHKmxegJS4/ucDWSQ/Chvhgmr6hZk
Eymqs8N1weu6UwofIJ3zQtMr7QZJeqeeLQUCdRJ5feXbMiCgEpkXBEt3pJ/F42SP
kO1oG+ql5kAMqLPboeAoFdBE84CZ7cXflgNsOcX9+DwLeEmbtBmI3DvSLxmznNdU
WDUbtaCuzfD8tbNA4hEU3lS1oXzcliVIvm+AwZfSHeLhFi1VTNrx/4LFTGcaMjRu
imoSmnneuKvThl53PF2DsjQG9vbyW8hEVpewYqpAker+gTWzvuPkS6SV8Y8m8twM
bJzynE/NC+amuyDoLfIHzJcr0PYrxZaLMCF56uo+eSrlcT4K1ebfLpurpGiiaHaC
YcRAp8j70rX8ZU9Nz/1IBuB9Oqv7ycZp0RvYGGOWcGcTyO8TWlWoYLaTwd8y1PFB
1rwkpVmvKZrw6F3BdMAeT+TpOOF/TFedqQfh8v36SWqeqcWv67ANa0TsgMjHp+M8
NdAkeSfCu6GcUvpJePQtb354PlTx42StOiPREjE7C+2e7rKUZsZvOAO63W7Rc4lJ
/ifJK5Kx0DROW0wC/85y1dX8SnSWAoL/DzZ7MTa8I3ZkqJEHxNbhk6noQoyRjI1r
iAe0IvpBe2ezc7KUHQRNtRWtrzNSAhVMZ0/7nz1y7iUiLxoEHVi7YEICYOt/MpNR
ubaLW/2Y1FdWRVE/o411jlRPHxZvhXdhEfByU4dE3MdV50spLmBFmeOOe5DHeSm1
EXsVB5V1JaRbblDjaiCcEqXwWMwOp6oF+hgZFm936Kh7zxbab8goqXQgLtSVgEKM
qe2U/hnWav+xMCKu3dCJDdJ12aVuWF2MUFkyDYHsU/nSyd7BJEriwnK1IutzGpvv
hRnlep+fLrL7rXvWrW6qFDUmpocdG6O2KimuGxSlz52WryJc1qJm7JsYptx6PxDb
wBvrw/TxYdN7ohSc1gWLrvgbqhHH8vQsOluQiieByXOGndFotX06Cv/iTH8m9Fx4
+HIt17n1GoJ3UvCsy45/phcj2pziWD1+OMPIR/iPpUUjkSv+qynEVR7a/zwUEX/+
/S23UuPa+HNBudL9sNJeB1uAqVAeBMfPqvEgLC06BrGHfOXWdUlPGM6aykxvMWVU
y1jo4e6lBSnsdct+KnHNIQSbxWB8M6hlKXFTlZ2OYaz5G+SRqpF1PVflMuaNQga7
C5fA7ZNp7UvQ/polcuX5zpwDW4w4dnEbRWYVEz7EjNgPHEFIzTxhPE4aZYYE7wJ1
/DfUaBze27qhs9CMM/v/zqSeerIEvYIOH+FwN9wOLFUJkrHBpt6vpAGGSPXlmGM3
tZyxWiMgrHzj01qJfg+63/c5Q/kDowLdzcUDJC6kJPbQHqti7s4+tOcAdWMQ3Yv3
5WY4v93JplnhCgp4jPjiy9sPa6XQtvDPdNI1MY4qkelZicJEZ/abXfqiKHT/OHTJ
sR+arJHzaLhd/GzYAjXtCiSlsQghjt7ggyRiMy+gjrTi9HS3r0TiIpMb4IeTLjIs
WIHz3snUrJsjINGxLxA68EO9MxBV3g0jcVgrYe5ZYuHhkKDqXdJ4JZKBbXNdtGu2
/CwfCGdqHlLQ5nN8mkXVatwlG+znNaonYWgO+WTcyziFXjwAsPKEK7n09PWA/uJj
Kt/pgjDtIjEr2CwVX908EbOR1rjTZzdLeqpYcRw0EhD69RP425cMbWIMj49wDjDv
RTGm8Hs9ARNZIcxxeRsEWeQKZBugT3KqzcfOYCF3LjIuVLMI4J1yOt9KSdGDt4QG
c2b2xNqmN5UbCxRtYC+SKWwYeDAM66/nHGhSlQsqcpF6W0ZSt5fbPpOINsL0wSr2
CI77VZyRQyXglKx4ToyeWJgayMflsfZbRuj4Fsw2bm7eGATnfEj15n1hJcjNsc7C
lKYVf0Gd0lpj6gqAPZ+GFsVRW6FERuqgE0QsDsceXw5kWbm/cl6quU8w5NeFtOpZ
ecmc6gxzjt/wLjlf5M25gip7QLCSiM/xG6MIDus5b5YxoSxKof1Y0jZTYNEXKwEb
+HDIwWleEQjmUgBOn0iuWqU9fMZ0YTWZFy0Sv3cCLh2VV8Qvi7HRHQS4+jbGHeQi
6+7lKGKmNxNtlaqeJlzDmwCXqVbf+B5SOMJO8NAsSGZA1TxN1S5BPe/oP7ILjLoz
4au+L6GWtKP9upGAN5+P91xLvgLv11ZZaYOPjoO8TMOVbkovpcPq574/6eX56SgQ
VqF6tZdCM8SM3h8PvCmnxGPeVgwc9ho8sCQ0bV8nOxh97YXH7LBk9IG6IABFPC60
2MvmCkjRTFSeEUBnmSHdZhMPaxIhk9Bu/W/Po5FadQ96uzmwn9Bf1YxgyBuhWLBT
JdCEzFTCd/hhrArcu6ODXlB4TYZ9oJw6Inbc+7AUq/6XEPFB5kN492ArjgomUSWp
fSfx3MJ38hp+8Q3CpyhfqxmBB4G3Xr0GWYjy/RZgD6KtqzWh3WUsj7pdQXcqDSL0
+e2GBHlw0kQ1C4BWB7yt6fUW+Iay4mNUEHjmKZcLt0xLiPQm0hIjuE8sViZ0+O2m
P+Kg3jWwV7q8X/YM28KRhWjiNU3N7B1i2LTy+N1/ixLENge4d+vGKRb7mtm6G0Li
iBAyUBxgFtIOQiMKKLXe3g7aTwaOtbSoxT4OVsgN+X3dhBMIcrKuOkv/X3WGw5U/
Uk+7h083fxNKk2+Uk91PnDw0PN4n3U85YwHYClg6mzjkvD5WgZyx1KiRr8hRCGyw
HcX7kAvhuKRYG7A0YB1G5g3xD/42r/M7Of+iwz4vZIGhXefuh6E3butYVwU5vot0
isun0bjQzQtAAbPuQlcREtwIWaCn8ic041EQuGR51KL75cTwzHhF0R3ydV0IC7OI
XLp8HCwEPXYVR79x5s/AHDL/cR8cQgTwmpOB4cOFI/LJ/tsOdSiDNTCw68h4Jrha
I0GwXhAoua5qROavDxKcMvOOh9cM467iPFifNXXDmKtpaDB6GsjXV6VJ+cprVgDm
CK1AQShwGtvq2xDSqWKLpBcEMGE1XpaO8IyYzVniitkc03AnxoZzayHc3aBA/qRy
jAQbJFfX8iHn/Fq9zZg6TYL8umLNVClVKCTY6zLCpvaeo7XPD1Rm2DPlgoCsSai4
y9qdzQLThS0E5HKW4PihXbhZAcfjBcvr96vvOX7KT4N5YvEs3yH3HfyMnu+mewL7
LMWXUVNneeSXEMj9nI2iI6queaOKRmIDK+TpzDGXSUcMhLYADrExzG/+IwEgREqq
bSCYGDFhK4WxoAXZwoirBXBT9tE9DJi4CTRkbZQUc0xU7XQiUQHDQ7qOtIHpb3al
P9vaqzkKJ+MG6PVTomTiD6mplovYYl9QcBj3i40u4bybtFW+nnN5kla7EIVDQmWz
p2UwcCQD77MZrrLVrpyF2l+fueuiLdSu0dVhBH2TfsELtQj1cCfaPvdJaOp2Ge5G
duojpGSIGZF4MVZTUsCwu3Y0NVO3pmn1m0hHz4IUJfFWPYtpFArEvxqhOQGKCKej
fW4IjI6NykAHxirM0UOKd86EeUsVWS93TillK+1ZJe8FSOe4DeQDwVIFGoaG7DIl
zRCuS8wMFpSXAO9xy3ndq+GkO70W2f8KCmVclZR0svTdRbyo4fDRd7ZG0oYzIpVZ
dx8DMORrqt2ygLEFBDdcmvUxQAUhTB6OTEXpq/KMeEnWagCJyZ89lHlAWKBOMFXR
W86KwGGkQ6eflxg5Lfy1cwupUDX5KDn/HSMqzFb5wEJx5Q4+jUqDNmHoHyCOzoGu
40x/UOghslfFjHFdBRKI0kqrmqEsIhE1rNnWODJkTcIiCO4+MNOdhcSu/0hUqKer
zx3HURNP2+mLKbr+o1tXkXdcjr1iNX9CmEpdkwRQQNqU/W3/O9k2BvyDvUxUWrRY
x21FrzUMA0ttRk0C0vbsFS2Akkf6jqKbdBPXx7oUrgVxNOQoXRIffnlgekpRG1/c
qpKpMyyBMhLdE304tvYQwCkBzTmqEeZnKCCeGIeM5VxhWx2qpCV7557VwA6cW1Qz
zov/GukCp3yX4MgKeImIhNV3K/DCwduxVvZuNY34Q7HIFU0Ng91JTRWkiLkl+Jxm
Y/yIj+xGYpy9YDwyatKfrUXHitT7NpHRmT39ehyW5mI7q3EvUIoPkxy28bCQcbLD
+7OpcWRLFxzmVeNZEfarE/sM/Di+8hEG4EdNn9cRX2yEYgXlpP8K2r+0pWnfqNr/
Xj371Q+YSGVbir76RQIJhDsh4jr4DaYQLV1DtqQkNFvCG8y7eAb8apIeSSgfnySD
EHHYHlEfbOs6GSiniq4h1AGnVc1TSjrzfKN+6CugpJOsss6QPQA6uCoMBXj26sHW
mnX6hhldrvancOwjsV1qN9PS1xVJnnzDUlyWMqcffKEEjOeEHRgAQ3cMUEb+mms2
3AgNhuUM/MiwX3KOUGa8H/GCaUT/S1qe/xTeQcjL5eeXirNCOoRqQJUO94bpz9jv
R5OmYCf1CTuUMparWj3xvzguPxlaQqAtacaWj0EN+d0QlOXEAqBC8qzFxsdbsdr8
vj1pyeSa0xe1SfIPu5i1D7Kw+JCL8M5/5qwuifXkidxhAlIrg7XxGobDRjRRfNaU
hRahq/92jL7JjGxP+FeEt7C2F5JprLQa9KiTj4lP1i4h5jKwP5XDNpL/rhOtQqpl
/uEEvQ3xDDYe+07fzVwI7CAH+C5BXJZoGkqYErmxmaP5bgPNzL9+5xXVGTIydRRZ
PdM25RAXN2ztBdh9B8aMiqVMDHFcJcdDfEUzJSVRZl6fEnAmxUqcasJmwi46SPqk
HawO4xTmY7Q1LBnLW1axcSAViT+iWnXafrrM3YZhRmDNs5PyaezZIYVQNoFlSbty
Gac6dr7Mz6Nald3DKH7P9MBrqkyhZG0neQMuxGuRscbTIzlAa9r60dwFo8vFZzI1
0fi528suN8bhMxIZZL4yACdOKlnnGkUImgmt78a/afGeIsdWKOV5EQmJb8vVrvf8
ulVfP8M+kZckHMwhqL4bLB8AZPOq9S32sCT2DBoXDk5u+h10bIuDpysDua4MS/9M
AWWaGGuU2Verk1M/sv1Y4hTZSjwZ+kKmk//QdmKixVqw76xLYOnG/gEzqlWAQd+h
vzhtO+uOPGYYpT4tcSruwAvOSJq+OzKaMSSvmDeeXSYDm4yzABLyl8MtDYAas7ms
fWt6iRwVgigeFRC97UtUTSLj5XLp2KFLUT/rpwjAzDxiUBuYTd3FfKFNsWMel7Uj
7sp+MQ/mw938B0NsxC03h09f01+iHuU0X/X54rNSrqFY+yK1H43mXGL6W1YK6KwO
wL4bpPmu9ZNVPQ5OhS1LBPH5iv91HRsyaYKKa/SGa6gak9US3B+1ws6BXDINRK9+
wj3vTxnxzZqQ9m98rW85gHhthfhiGriIeQOX5KByfiiaut0vJ9b+PMkza8RJEyRA
sc+c2n/RyMXNuQr4PcqmGjULNhgzv7K+FlTe9/hs7wRM+7jlb+DTahUNtpGVXwDZ
bBkOrlQU6OzH2XZvq9B521YqoYaeHJxmgaxCRVD7BYc8xGkbIr5MPfOBuFSnn21j
ANVFM+qhQNZ6QgXTOuEbAMorzK5E1OypFgPTJMOGmmqtpI6oKjm3juTwyqEzZe8X
l9XfOYn5naOFFkj3oP7yEmltYt/3JbTtnrLjh6xdqK8o8dSWc02D2DMAlE2DfrSi
tiWlZhv7Tbnls6sCh8K4Nj6eCmYCSYhyRLcIsrRjnkveavkDpD8c75Wgp9oZwoIV
f9N1KWInUaFu7L8tUqxdQlmINSH5g/NYJlqEPQ2S3RtHnV2UXj98axjKB7BdYDQE
oEouVBq+RvOwHTOXCWOkCgKd02ehDi1fR8Zt6LwZiWInQzqL6tISB7KVAlbps3a6
+5PTA6eu7oSSXb2EFRCMk69KsqnL5+cirLv1qlk69N57hH4d1hBZERw9da0l7Ih+
FTvNIR1BvuE2DIPoCq8yltDABLby6QwW8US8Nr0Eixvzfdu2Xuw1PMIGrlUlnGDx
N4istektCXd+4TBzv61XaEO2NC10vyhxwFnizEfpNZs7xVZdZfl8keDSHoN32PTV
ERl1fqY3qN+PIivEI/MjTwo2KkbzdkD7E99Hf57uj/h0XztaIShTu3Qp+Er0JBrb
35dBf/4EKgtqvkTRZ8MP954SBJGTaEYGpbb3U/mZriAnWXDhdIHG1O7gcPag9yyJ
KOWWaX7fv0cvI6xbYMKgwLvElgoHzZJhbjz8nOb8ZGq5t1RYPl6Q4jVl90f3jlT/
b3Wrsjq2A/77gYpXBRui9porckpLyyesYIbNiZ/mccCSQw5ujYHbxddRFE2stjzd
jLVJ8pvUyoGeVwE6r0Ntbv/63f2Huk6rndDVJd8BfmCsS8linnIyLF5SN/WsJmG8
0blkp9g51sX0HA5++2Zeao9fLZt+t32/kiIe62v57pX06h5dGQQBXLt7+QXEBUoq
uBCtfbt2NaCd/YM+7+jcGHCyKFYCulUQVAbF4mqxCRKUA9hFSvV5rKWTB+oe96h+
0maCVjcmEJOJyKWCoDBSw/aJi3Jl4ORIJpadaoSb+8j189Lxtz1TghAiE68vHRht
+DBURee3sAGq5zZOy557pmfBpR4XLt5P4TCvM0IcmJ0Ux58j+nIGiuNjsKLqmfO/
wVC3awAjykMddqM22IibPq/BGg277Fd18Qd0CQEJJiufGLM0eAXM0fI1tYcnNWYq
vtpChuHXb0YG4xvsGkkNzSVPYqNAC40B2sKz5qaA0wZOWzkUHVo3AHA1jtFzlRkV
rBw0UCj4W2ruHIIhIjqwR3CHh+QTaClciyeHZt6MHdXXcObHSyOWzqwH4MwvTNNu
vsVnKmYdddbgtBc9cEzU+7TLz9gghXnUOGHBZmuLWj7twsO9tNXFpemV+nr0Z9ud
7Z43KXUkZCdqsjhEib6xYeW5aCTGscanqsu7h32JscxbLTo6e7YOf3EQjMYf0zmw
53FRf6BMbvRSg8exQJitWjE+gf92UwnqTWwfnE/+XdtwCKdTvyEY3JyJx72477cl
Jhg6hPMwGY07TtSH9dd7Eb5XyroV2h4rt0NN5UlZnK04ydWJ1RyICjYTVYA/AO+y
U+tX79DjVkv1tWXNZuyJui4MfsMHDCvO0e9H2licOOhWe68x6rw+0p36hxMuWnW7
c+JcqO4iEugJJMAZZuZZwBBp3h/8sAggTwRCjYAHggIQHqb8ADzQsLJ4BcnjVI8D
jhofaHIzjoqWBgjYpuql8TF+LoFtm6O7tT+f5haeQMPWdVzigvk9lMBu35LnskBS
4IStER1eiFRg2c9A5XXfZ6IwUEbwiMZv1TSzVc4M6mlnGe1TOdQ4xcEWVqVaAN93
k2lztydE1A8N40oQAz0021eFHCKYZ7ROXAa23Pe/Q/eTG5gQHyVzbyNtEtc6Oa1O
cy73qMs0IcIkFgGHHeY7q6GI9/scveqTEqI0yqEEBUyVMgpGI8oyUBQDJP5B5RkS
2FJaFk3PSxf4gQFH1AlznEpL26763I/faDDOevlfUr65xtZQz1JbGikl+yP3+0Fo
PQnWuXKWIIdRyxltNiEXO7oJefldPZhcNk6TesCeJ7jiloIvu1Oiu/oN990Irs1I
cStQrd2L7ReXan9QeCZumJyZ0tyLE5dadY7P+lk0jX2YsCoyPgeiiUH3PkF2xK/A
EypfgozWIK1XJL7FM78ZeGpxW+IF10L+3V8c6AASDruYoX8Lqc1wqAtvDnwxgk0F
KehEXdlL0i915hphGo9JfWt57wcihsOM2So4sS+CH5RIFHosfQB612UqNes5nJp5
QbyU6QT2PqDOzSh0DaWlufqZiDlUKLmXbJ0JKThaeDbgppNciA/FHUZxHeSF3Azg
Rl5b7utX9ibDg3KPVD2AQBRDl3FFPRKCS7lBUvq/QacfzFTE/x4Jn/QT3qKfwIl3
yx7VgxrKn6UysDLyge4h3/JJTj0uB735l9uSeDlchPcISQcpzX77T2UMJVLGSVHH
ZjhHohaDoLIksGYn6Z6OhKDD9vL4YBXdZGv1ktadipcYBEUcFuMAIsqw5188EF7D
wTNFMM2Uq0BSofh/Jv8jlg+26niLdGrrG2U6F1K0tWcXSzmkcnJp2rMzuY5mfwgL
bxQrgqAsHNCG9Fh/dHTOIes/Ge3/vD8IuQMUXUiuJNXVohS6OJxbAgW6uodjQdT3
CLIWxZfb1PXFFgrpcRaxmLujE868rJE1cqAIoTOGsxU0smRj4N3Pu5AZpCpe3ccJ
FIxYJiRNzjX4fwEjZuxywoWsYjp49WVwjy3N+k3UZxZXNN41VdlyjUplW/23s9ws
zah1Gm3aTMnwCWGt0Ly1PUuGgaAbzPR1PtpiCLIczCX9PWImjVkaT3d5A5XQFDvW
soVhwRIbs42CChudGxzgRfy8z/UjGtHZwu8HVfIM3DkCslT17i5MPj2/exbqJcvM
q7KdVOe/XHYCCC1tBU4lNBZv5PCA8EyzV+NtvjHtsV81qkDexksGoT5kFUs/TPwF
+bxKt+vcSHRrg9pothxUg216rqCXU1zPDu/ywu8dhAriNTmCcAvgeKdM5FvP/TmV
hWKN5HwlLQYeuxHt3WckXTKj/swFjEqFRquGUlCqRZM7MWfcuOHSkrAl5SpnZZo8
te5i1JwYXMzS8XBsM3Ol7bQaAD34IcOIj9nSaAFE/F4/02vtzYFC1FElxxf5DHMs
6TQe1VOTmtEd9gSZzzsNGpTDYSCKlK8yFHeBQb6uybA8MT/MLjFBFsknZY4JPeds
UCZX+x2Yz65HqaQksPxNwZI1ffZNuOdAtlt9AInBQ05kER4SmRNfHgiHtO03DFz6
ji63GDntHE4CSn2egQa0oPL1mJMNvemmiJKTRy7YsoS5ZcbUucXz5ixhIE04yhjK
1O8Qum2PSsNT1oBcaDVGTA1HSLDWs5r/kxCw/t2h5Knw3U4+ri+na9942JWKJIV0
u3DaIBgpzTW+u1hsTqKHhNRCMl/uWHuKGN0srPPD8wf4THbQf65IwA9n1FNCQU10
hgKpfX3tLt+OckFXHUKjWKbMOaAAsFUdhbX6LCtfPy1/UYQJ77uBkaGGRVKaSsry
D1rcQIjKnG8LzSWiR8s/RHS/Z84BE77G17ari952xSMncCZdyW8Xo/V6Nx5BRDF7
NRxim6EsD38lRJclNtr2ySPOFD9ZFLOr/9X1m58QuvRR1Jxgl6TdvbU8dsWJ6uGw
pNKE7zXej9zVzq2A4XpOn9q9WLwG7TtIQIo9U6lw5C0oyQDpfE6HOebF2zx4SC2p
jYMNGKy8jXDrKZy0ldLB3EJOdZeZRdFXRvjNfWUhH2cMdDnXX+2AqLWL2dt0wqVy
VE41BfqAMHi2JALUDKvey9XkjON/dcdFnjvbTGktgsD41uMyIIpQXAIFvhtxPVca
cnIW7wc/rep9E9RwDWXQebzYHpfehxdRxtz/ODWYHYKIlMDQMY072Qwz/YRxk39d
JXHnpRvCew5mexd9j5nRAn7YKzZ24WlvBokupg2QhSiO3EdlOhPHvdJ6ktGRkYHG
chlhQro4XlMUxze0wGxBUrAHOiscHKvxzGW++KN/HvKgc+YnVwYO1+1GxrfQpa2S
ztsmhK3t0IsE7GRfm/aUe7mPGRnImAdwuhXLmxjNljyR4A+VAdIg1mGPG7Im8Mkq
YYgRZmdPhdXXZ0Byo4vlGEP/21Kh1RS2xE7aI5yb/hKYTjYTUAa/2Ry/x5ZvEfJF
WPZ1Qsk//fcsDjMW/7zouOdJ1iVOYFloy022K4iV4P2Xa+nWR2eyHd2GobxR3hku
HdG4bTSjgZSCxK1G7rCgojEvchjs7PPy8SJcICBC8SM6U1T53jOxQbJJsSRAPQ3F
IJbZ2JzETWzvZCLhQMT34m67symtefLejrUOTMhFaj8RVUikNP6Yvo8+KpNPrAe6
Kf3TzTt3BewlyElIiKcmdlTUAYQ9131qe1n5ghSaWn8f1MzYRo/xqak6UauZaU3q
r22CHClIPTfKxup5izlIsdxi9ZTgvjyQEXoQPU08GfX9CZYMTxN/aPkzN1qCGmwB
fO9sHINQNr1ebRBIWM1aGRWuM60dlnZ+NZJIwqZGbXCFnldau7eRopdKjCi7Gqbt
bq9sZRO/wvPSuE9tMyEIJ/u7+E9shJE/yeGH81sJWCn628Ap/JnSK1/fBUsckLg9
JgB7BFfiZkQJopTrl16WEdBuPwDEkxh3WVWWREKmGwU6HyjpdOxeGKaQlRKgTkDc
Dx9Tli2ZrAy8a/wLcXvxLuo3Y5uDNTcK2QntR2qKZxGAdn02LWsXPL/0If8XXeeq
XLf/5h94OaVxoEf0+DcBTLEueYZVWRRav2Nrqv43W12aAMi0z2UsNJFpYnrQIkIl
Rh+bWoI55g4xHgis3bJQl/32NbA6JAa+GZzgI2RMt3Cwnv+ES8ZEDxtqSgHM1dGD
Z2IZwYBsefJCWrHf/JWEpmm/3mLrwdvfbvuezL6oXa0vCBTaCklS1ijZ+05rpbms
YUD4RYuuFskWDtvGgIyJhZK9CST78k/FgXlCqL3w2+XIyhGTKHMRHwCuHRVCnox2
4BD9dzf9RFmljRb/4KRkHNbsXwfy3fCtQWt6ZVR6a61og4XsZhMUr57y036kBOSA
VSfv70JvGNzGux3Wed3qmbn/uedu/ipHQtGQJs5c0b8OdmLDBk122wWpHtMlZYPi
k2Zm1MHpXbWGaBB82WXo9r3GQ/P0fW1zC5VJKSF4oZOJWk6nkjTLhp3aYotKeOm3
yaAuTQzXJyEEzAv0kYFZ/hYKebzCL42cmS7ZZ5Z97VHmWxNR02gLKjMd3slGCITZ
AvvFPi7EAXn2mMZpSz6ZkrDTsyvMcF54bDUN0/S5Fd4zSwZLJWvX6s64PErSNqVk
5IcetXVZEnKlb2NTPSQ1e5FgTky5Bair0flCXyCiLBqAYVLINlR+E38Zb3Q9OqBn
+Y9aVOgOJEdSkP3OGaEoz9Oqt4epnUmSemYYa7g9iTo/lBZziwM4IBrHHZaE3kUE
6svv6sIglWEdDFCQoNrP80EqAvAhRhgOZdhFhkTU8AzeYxK4hrPbxuzv/JQJ73hz
vNaOSN0Eox9U1YBgy17vnu7dodj2sMpDgn0rTVLkrkXRWG+gfokWwc3xrbN8WDec
s8/RoJohHMi/RqPq0ZcOTGs7ATY78yW+6FflZluoRX5FnvmK+MdGNdY6sAp2DgAV
Tf56ShXn4ZuvcTLJ4Brx1jWy81FRc6veH33oxKjoZLPA7INkNmTDJtBVyFRBhdtG
oCcyGC89dWF/wDTimsOEGZncqGJH7gf1314WtbVTzsXxCziGIeSvaT1AUofubdoa
k49J8d7+PIk1LpAHIW6mXV6PDUNXEUUgl2x4drvRX/OrnMKENFewW3ffBpGGnN38
h91uc5zRGpDd4Md9i0qIK7qOTZrGtn8xaLzZFnz/8DTBJ9jGKkDc37zeU0Sw7jqQ
dy+FuDqTV8Jaf3LMT39chEvQYD5tzJKyywJmMdMu9brp7wv9T7/FKAoudVIUTtxW
9SI8YUL31CcI2c/WanD+Na5kitZGHFsZkCME6ERt9/j96013Xv6X/I6AX6SjUv8K
4sWakjtjm3fD4CF8pehvHlPAJe7mq4gudOFlOAlZGFj9zo38fklzljxXDMg/M2ZL
rarNimlxr4l6Jlv/CABQvXMqEYeyWXXbA5XAm3AxFyOrAVMVIqLu3fvct+rM00bN
GqM5PGVgyKLrwpjTGYUVsbhdHsLyjj4NFqL3KUl1UxRzMSQfhGDlzpL14DilzjGX
73JZ8261Wcj2MJiJRNuRPyU4zTcMQBbDttRExe1oTHvgkbxz990Z2ixVkBrraj0g
d0Icby93moIzZZ/3Jcaj68Jj6F6ZOSYyZ/GRluPCCCRwQ2R109RWqbG3Sxhxz84H
9wEp98KHGdxvCc9rnUcq9eXjsdQpD1AOpDiaq47S4lHfUzby2Z88egZ87v8B76pC
fJh6P6+2LEDd2bG8kQVbWH0EIj9xYl/jbGz1HOwTeqR7TUpbvwR9InFUkHjFzJsd
y6jBjMKlyKJUIWljbrraEtCtrai7dGCs8FvYn9aP09zI+Cq1dT4NoiiDqzCrPFKR
+tOoGeslSPMLf4fJ/zi5bOj03hZ2csiTrVOiFUrLFtb3/FLIjjOsV7AIqgPphni7
maXBK+0Ub2lZFcn2MFTpe5a9Gfl8j7r5NIHujuDU8ry94twcUYF9X/G7aEWIon1s
lTBwOhuGhMYZgbHfxut6R6FGm4ZqjnKklqhPyiZ3SSekoFc4Fw1jEw7NpFhLxJ3L
98YIco6kwa2ZehXYsHlX4P0OSPixljmDm6vSxADHnj9ACcEXvNqmDpnvLHOd7Bvy
dRFcbsXtYnhLrhCP6+kfG4yIlV9DUmgTotTJJsyGTjqrDMeae+5kSeVC/niJz1Zm
nmmksyiYswCB3pTDnEmMaCK1CaLdqQEZihOrHkoo3JpcngRltEuSqvMuz20WQ34k
0sQFnbkKTWbzmaKsNnuIZO/IfJ3CObkrPRjUMuH+xRs/LAMHBRkK2V/AFuJRVVza
xb13tbo27XtNkFEdWRjaRBWzyHBSgQPKH8G3H1dTyWkUgp2L1jglhimvB/TCxiT5
P6WLVRQgbtYczwaLzydp2qu81LQPDLFddlMJZo4f1P6DI6qcLjMKAxCh1xoinblx
2fdvY9vVwHKUcOt3OM4R8IA1BLCVi9NH9xB83LQIbdXl7vmtyBVjN7TDsEooXTUc
pLvhElMk5XKY5HNdDnBt3oOfkSM9yrDcM7a4JeeTWg7buoFHYoKDS8EwcjbcaSD2
f2ZdWY5QeW+M3z9yVprXmf/JOQRhTdoq/YJpIq7kHDt/AquCBLAJ+poD/PPnbMPC
1ad0II1PlYEyGvUqEy9UI8VUZzf0Nc1j9UUc6szysOyiGI2pM6RegtPgImahQZBP
lXJhni/p0TajECwwToL7tH33hdvxgp6DkTvMr+TQlsckfJnZY8lfJFvmSJFHTddQ
QCNOmT0i7/Jl4CoqO2rXTXgzyvxH5lezCnGNMUA2ZaUoW+cgWVnGqKIBfAEPo2h6
sGnHnBpKQPi8arHoByjG21cAhWwDIX8U8vahE62IVSnRySW/Z29Cs5Jdc02stJJi
/8BKWhtIkwYy1aOTVZ9aPS6bewZgy4l1jjlGuNM6JXm1VHUmzg4PsGPv0cBCvDTu
oGxWwYxpJYxqSrEEL0NQvvubVWA1P+C7yk0EPxLndbvcaL/eRzmpbDVIvXeys8T6
Aa18uDtAnKMSyFTdplvq8qHgU39JTKJ82/ZKQeK/J5zXwHSWcKMZ6dlB6+d1tH7L
PF7MPvJ+RGOnT6+yuyEjj/Sq0AVKcKDFHaVIOhGy1VAcnMoX2HiSIoemHVNvhu4j
JOyu8wsLxNawPW95Ux/+e698490W0NX2W+LqP2ahQpWpeCWneLBjkBc3DKA8XHIF
4GvJeJwTiismgQ2UM5emEbZkgxmLYFJcPMk4nK5enG0ui4LCf6SPu0+7us7Yjnsq
kTAVMgvcoW4z/++ZfHN5fXoJ8FOgeDH79eZtMKmh1kE9SM2U5d3ZbgIxYun3d5Fl
HRsqn/0BdKY8ujF6GvLRxSUG249SLBIaqDSF8+ex2UkT2HSApTlQKaifASGGT9yj
/6XYOl8+juVTTY/Sz7I29d2elT83leSLwk6lsacNVDIuAzs2D89wl57UxcWh8ffM
aeOwZADHYx6UmAoZ+4cr9uiqzKwQ3mjJyYXfNBsy9AVm1JJhX8FvpolZQpYdb3vb
QsaxNWd9hS/1E8Ao+6i3+VA0+xn9U3/Rypvwt1SEYc03Qcjz26u7qJG1aKrLK4Oa
6QiAEjWCpsXFaGvjpaGbkWOmAxYFVfFGVR7XVmguyglwW5nVuKErFT0qNMOECBnS
kDnNR/wMPa0GfijiCq/KTj1QPle2tuh97pdXkV2uXJJ+R/jSuuQ4wBlDbwlcmmX6
yP5fFg33vH7/KhzpMjVVGz56mvq1rOk5AEm2aSwDRreg4oDALS/iLpVtcOM4fyLB
z/+1RWkvCx76ON0/mMu4ShXdkHG+69N42VzOFXObhhpE4CahDkJxBmSHb7CvZfLH
rRB4maDs5tG9l+r5K+uiiqD1hYVrbF+UT/4NNCcctb8GCTTi0mqtE2X2XMA9bLnU
FXzy+EjE8oIrQIFKIWWUj7QdzJWrneqdwkS2V5We05Ac2Tg4LYQAe7X6fN8oiQ/A
TM4P7Oc/eROyBlDyC8hXmqrTet9zkmIkd4lTIp9njuH7Wvo1AEto/CgJbAuIM+i8
ZuK/OjWWyG+12ZsHZRr6PGiDbN200s0plarUYOrHT7uR8XHOtXRHgtn2zvyQmI+3
XNuQVfEoRP1WPIrjQoJ90dG+ITv/SN6V+9/LyoblOwMaoJWERerD55wLJ7wuv0F0
mjh56+vTRnxzwkgQRtTfa8f/dSpljtIDgZ/9qQFV1Z/s6xSLYBCOx+IK8ZU8cPfl
gNkchNsOivMUpwhxE65pDxEWQvFm+aEFWovTHp/wiXoEHFEt4zeZxliGahCBOrNN
98I/yi4s+QMDvT9zGO9nLU3WXV0Gudc5wrAsLDJBb5q4gWww4/UmOBeuRIAJChEA
yUxlGGI3FpShZnn4qFgSQCrPfXApj7itagf5FcZ6ExllU8QCUZCWwKyh9nVUGFLB
pD8W9JPNPHcJPNOmeYyZ6a+BljaNNa0iuw1/bzcPC8Eri2pIzAZXzPOtNp9rZUC7
YVB7ufsA9RVzm3smmoB3B5nWL50VAmJlAEmWooQAfwLJEzF5NJ5J4dL61brZW6FE
KEINAylMVnb1vaVvvx30L0ZOjNHEkp2/AixnCelwrRqe1DeaxgC55t1Nd3Jf00EK
GRJXR/xwemMOIBXaQNzirJQhdTdDsTE6gSLmYgHAa/tS/0g9Mi2Gh5wApFzBjuiA
fep6Zkpbw9iNxDg7wnWWNtH6tAxJKD7cIFPOCzbaefLNO5EpsKCFSajzQpeORZlZ
MpBqq0jrJBGfV2ZtIIZn7IFgLYwLktM1d1Tyil+ZJ+UwYFR5SU/7WZfh4uthmXDI
tLTrEnenVVOh0x+LUhSltk1EfHCCah7HZbmfRe9BbvfGcE81X1krG3s9InXq4UTW
qBu3lPqik9jPzKuO8/Gs94OD0tIHcqjBC4wMd/7Wrvpupd7T2oYX+I75DG1THrda
HHF91uUuykTG6qJcf8U9ll8u3TFr9Ne9Ykp7xpXCB4XwxbO1RmD3k5ycYJdsXYqD
hJxy+ESTfoVmxAzZjQmB/SyuS9C6v0MNDLvq1ramj93ubie0rCZj5Pr9bIw158w2
GuxYpqlvn63xSYTfGqRGFPpCTrZHvg3u8wY1wyOLXqJlUC2IjdbCOeCK27HgqMR5
5OSInx6hevGaNQmDWRsWWBmr93NLjBY0RxOuk2ZD2wJKrpgpoJD6G68kDW+PQAh4
53NJF1XC68/58WA7pQuZMz0Xw4NWBqvE8qLNiBLyWSjcnypc3XZO7FAmBB8URJIy
4/0xxeZg1jWG9ecntBOJTJ/9pGFZhzZKITGBHKccmfmfwm+4nESob1iQOr4ZUARG
ZbbIBOfKo0U88o/hY9ya1mLLJDgUHeN3MLpU4VPEwrBfGPq73c4V/zHNffp+p1g2
0EP2xvhmlA7Id6mQ/OP2XydQ7vewrbd7QjLL4I/K0lOSv0EYkpWeRxKBaBiwqkp1
FOcvAtStxNzsXiY6QjlG5U1UbRXaw4Ik5Oj9Qq2LSk8tlkr8S4TC8THg63QNwn4t
aLdM0GYS9UnnzpiFPcxeft61aYzcsrRKxvvfw/dDhzdBjP/39xn8yekBy6uzrgh1
GOu0r5yXpg92/g3C3Iny+ehGKrx8OYkcPSk+bBJ+ukTQyLUIbm2/MO2IykjZuhhQ
yyOaiytnmrG5Aww+ByuuVCDYDeBqUNDGM61qJ3F31/31Ls+2kqt4eiXc7ssSNw8x
+UC2ebw7EDcEGGiXzA9bw5nBGz9ic6ddOCzjJBXvnjCpJtZWMRgiJYPBtcdhO08e
X3CNlT+tPl7fZoUbDiNI0Xjs8q6CcQp57vXXDmOnLX1/N5R7HzqRSEpbdfxBX0JN
gKsaR/tfcJq/F6HsLnxC1Rrq0o6+PAJDoL0BHnGmVQO4taQYnp/NhdEZNaxS4PRm
KbIyeTqcAw8jRO1UP8aw9qqot6okC5alAbeRSIBapu1ISb7kj5Y04TqLDh6eA+v1
kj+cMSD2HD0L6iqTKbDIMJb6pBTiHkPNWOJZ0jXjSCIHtroQfW5oRb4FQm2xP8Bp
esDnDh/iAXDPTTRiy8Kz02g+VKlKf+IFp98+ppXP6+NFX7HwMN7K9TgF6766yaCr
PCgWeZGhArGvUntIMztqmachDr43mnOHNbP57ZfJZb+1sZaxcmNhIkkovS+Nnb0u
6ayYEYKzlcEGP7fsZLt2cXLSeI4+H3KgXGN53zvsDMH4U68DmMrS4exRJ8xzCJ6d
FxSP8hwziEpy4WbNbdrf+wuJRvHh7107xOMF6goPVFtLZM+v/99VXT6z8wKssygO
p3UWmO5Csike055aWvUPaJfLrzlH19gU3LD7WwGQVt+/QrARDae1XQZgbPU+eQV5
e7jE2O8SeDIwWhJFWRWubf/hNbjjV2Zn9l4Bzvjvb29wdUm6rjXueF969LJOwMer
Tq5EGYGiLC/b61grKhMxdbrUMVaa7o8cTleUZYZOlxKpIKHOnmSmby3V6F5p2Q8t
X3MgcMl7FUO+B4DDLjY5AFgoHsVr/+KS39kG2tTHDJiiQ+GONcIxdk+Fg5Djom+K
p5sZEwpgGCul4+0BXQFpkXdeufg2bi+jiUIwKywwCe9uA5R9AqhBZYtwmmqs15AM
68up55ew8z04Uovui3X+k7M+YqnfJxtXg3aKTkMsrGARom5HYEpdBVuzzkF8wFj1
wECoZcj8pTx6W1X3HmwLOs9wHG8w/kv/XYUaHArqwzVR1Gu9bTmwbuF9GbdytcXM
uqIYxTPRrnIj1o+WM03EcBp+X+/Vft3VR7jZZ+kONhN2Rffm//2eq78EAa0hxglW
tKRPCkxNw6/GHiKzeL3FANfdM+SYMzf6wGff4HOQm7r1jYDCdFB9tM4ngV0FVgC2
+A18dpDainooXnjT71eMFJtYWkNIFGDxdcklSH76mnPvmQXEQVdkPSBcIcdbz0qY
5SDaQvwhM0IePwsedBBCxqksY1PGZiC2j9eGk5dKxxUOdiZcCZZqGdiXrwrQ7nfb
q91IEbHOitxBkXDS2hTk4orVGAOshAOrQfDqKuauG3WKdR8qbJSxzIEfSvPen/c8
ZLogIumpwwRdHHhw5WVocO/G7svASR7qAk42pYh0+8w41XQKNNdOujLkJPSdPTcD
RCD1dFs8VJ1fQpSpgsGk4BXX3UObE7aNbuSANdAzerP1bSXQjeVvdMek6mP4aiuT
ae5iObuayHS5uh4Vk9fdlDxg3JNIrPyuXDWiZcvJP/BqfLRxOTlDt82eMC+wwvmG
LJIl2ANkpklH+2Hlp2twr5U14kyL3bbdQmRSDpkSHd3SiqIilkkaYJ0POwd8Dwdq
1kaaYxNVooUsZlyKpsenBVln1aqVPTboicTD86b8ycOSQLlx8FD9ltySV1k4NizM
sFKY1VLcZq0LA69CPzCXH8ZYUVajhq6RQOWPr5HhnIcjumI8mPM5PYxF5/td6C8c
tlY5Uc5qKGzK/kE4anWTO6qoSS1pfiXRJfKOMgwVCsPZhBJSlVDQBualPe4o1/99
YUviSZWnCThoY5VSriNnmon4n2Omk8mVelRijmukGV9wOpSsCghuankInhSvjoBC
M7xaaLFqdYoyt61jksChS59V5rp2ykR5XskH2N9XyoBWimyr5ubHJDl2KFYCtiBB
k23mlxvUqkKW021AEeSj6oqYPOyhBKytjkwmp/C8pHZDw13kXZ99AETO8OZ/qpYw
dN9MGbgClNYvmqvgFkJQVHn43bxmZr1q9q3/5YnSX0EhncQXkLZJZGhkeSDWpwsI
hcTYCPtg7xFa2m3KsL4rO6x05dArDztqO7NFdbCi/2HcT0lPp56AMsljM0YUJOv4
WvmBvR64uYdp86b+O7ZZ+Qp0QQPRQdForvWZWbEMmAzVG+anZoO/zLdC0CgesLZJ
h4Afn7pKZfppJyTiZxLvo0xRjy8Uhwqk6Xqs3maOynKpWBtEFoMtmaXoA0BFYLbq
Lbv1ZiLkZhMiSc7T1vdjB2wW4n0jqHiyuf5MAG0zNDtVxintp+6DVJTxrAvrzRig
p7loddcPvAdpA+ikh0S8k3cMwVwgJsNwSEve1JQr+579e1ePlteJF7hH+3lhItce
yK7UOqi7yvmecYxZOMH1U+9aBD79aQ0CIOZ1W+I7oiLKclAvxgOzQjVsxTFEJstC
PwJ4keIT7Zb5M2K6CVRiyIQugyR/oxowPF+cNNt/Ad+YFtPgF0834zOScUGZmhLd
YUIsTg8ZiZXc1a+YWIsFGVFRaPwfHLJ4BMc1iCOAZ2zOgJiyMXUS+ObhzvHp+S0I
CcwouTalT+W/SWECjWxCXMhxZRpY3v07NWs6DMV+wobq3eZ/yG3iOh2OUsZVk9G9
UiZAKxR4LlXzQx2/rDebwHn8CoyVJ9goy6o850zkUpEOI5Q4Gw6gAtoKMn/6DR+i
ZyN+BTV9KcH3e5xaclFSo+UlFUep8+/9CQS0aqX+Fn90Zw+FT8haUv6rwAg9Xm8l
Ehx//5J1DOj7mCxn49GWw5v/gB9UxFLE6fOAtzsJUNHt+0LkAdoBfYEbkBjxlpC9
YU25Wsif8gC0oHmRKWKcvlQ/XHc3L07C/YKxZ+brZbYTb8d82T4ddapg0COs0rRk
/R8xD4Rq2+waN/ury4dkMWIFhxTwKmH2hyjEa6RPtH5O50RB39A+OaI0+h/SXjQv
cTFKyUfe9fsw12Z8TFEVKHOWILHj4ThGqaoF+pQjXqw+0iOfZzbEoDsjpiRaGmm4
phfJo5EMOilLfezPLtmizX5fpMPJEFprbXkc+gyMC1XDKD7yxlXMFjd2tAx1rzDQ
nooUTj49BO/BVtOE9TIEklwZ1//pAbaAlaJLKt6EMbUECnvcurJauwbuB83/kZZu
PvOtpvs7Uq8M009mWbuf1sjKtmRlnl7ydm9H/sK+n18Hz9qAumnXoznV+iAxLdn4
c5ymZcoe/qIfojHTpDcYCzBXR29QR0cl7KzAYv86jC/rNjfnFZrCwsW3FwZUlRAA
BwgKSuk+iUTC23GfOQ8QwnMZLsFVRXrZkTunDAXvaWzoOD5DFnaOoH03UlwvUGQq
R9N0ZLHr9NXk9Qku2AfBfdel1+AnL7bwTh4gwNo8FNj1kM2ZSI3HaE2gEzD8LkqA
6QsmM/wxziYNBbevMs7aWj4iJnCoQlg04HPMOwaIYh62EeBDC6p4L7u6orIoBJa4
iAqnXLqNxJi/ZbtyKzpL3S52rbvi7AEyCLZziLnJ/mXapzWuJ+SdMOdODiOPq/Sl
qMcBnFovdZZ296TPgTu1drWu4W9XCT3OwqZMfUrdJCyUXOLBs65aeuyixdhmisUZ
l95GK2MlTC122WB6+gF4Guiup08nfYMUSULOk1Psi6Mp3ha6Mean0CoTxPntSW6x
8zrzqq7b5Ow9XiRhvBFju5UNFKT3xYe01N3+EjPGDoTO1Qm1oKEVuECLtINGSA5j
6Bf4DCpSrmkjk/uLz6+/FxJmcPLETOSG8+pUZvwoNhS1zVLxipuwnAXXKpm2DN9J
ZaQB+Djkeby+Ui3b/8I2CixbBLfKndzikVJxAjEgjLQPFAxuhD7L9wxam8lB2Y6l
cRr2Dh1s1b9IPC6UYbZmvHrT6Qk6EQd305BjxEF13BpKuBvAjeTCLYwaCcsD24hV
k/i880M1gn8bVSfKK5pXDedoJnfFtkt7Kwjb+Ye8dX9UIhxhqjD4pIdnkzy2YWiJ
a0Gc6s54kbL6kzoJZTZSa6I6KiSaJ2BXjdNPM4uICZwCrexO5Tz/Pgc/+8s5lgDy
S8YoaFJEdjYA+7MCDAGPJXNa5saHCPRRO4+zyY89oYXaS8ej9e3/t3NymMdLN4SO
GMRy/pUaZPY/CTKHefL/g0iLyCTc2XmzolasY9MRjLO/ZoNdeCCS7sDw1metMoxy
Wnlt4cUDtXF04arH/MfEKPrUbm/MBby+XVZxD/mDh7eA2Tj7oceMZYKh1bRHgoCP
zqE+WTN+bKhDX/6gjdRzpENAh3tZTFexoX/bUR6jPgdw/eHZAGX++yEUw29sOfc1
k6RMW0/pSzhUdHhIG62LPzVnG4apW1aWG24kwQbAzSPyCOf0jp4NVxqZ3jzvbpNN
CEWUcfkqruu4YPxu6pR8HTCf5DiJeJUJcZymFmg0mUYgFyDxCeErNeevjdr8si85
jTEAR6S04tgywDjYBAkB/lIPR+YGNjXkgfak25fJDJZRnyd69z3lFvqVqhr0NSpz
fJzy9qmtdDQEGS/SccsQeDifFNLF5qjgi4sOn5cRNEeClDk6RlEmUw/GuXwSE+3P
sU2lKNrB5Du2g5P8AqvgMk5P0RE3ZnzCJdXTwIMTojAFtTDbq18lF6MXmbcL3bRt
2lKbV9u23eUWwSPvWUha/IrCYMi2rf1pY5vx8q5vK/UKs4tHN75R7zAzPfcINgQe
SiduBJZMtbTJ1IeP0aBZjqKOQGW/w+Ew1h8V0FLi5smGW/PlyT3iDEiFMCP3+kqU
wyeXlYl2Z+EoxFkJXVC7rpSomC2UViriIhbeYXzHhIBUHJGaRN/5GlMGGT25T6UO
ExdXOgNSZvMmSjL/k2bc2N974+567Lpmm3Bbbwgd1NmsGVt5MlrtKDLkugsy3ZZA
/VIlzn/OUEEUnubd05jlsrUeNTHUh5QM5Qf5xzGEuU2hRO8KMJMkLh24TV1fBOjz
iztiBpQM73DiRvv5nlTqzWOVeV0a3qArYpn1clSwPUGtwxQKurjaFPTooHxUGize
mE6ku0Rsto0Y1AIfU2/zl3rUymmQi0DgV2pCdoXw5fsDNTscAdkcpdHClXe4NOVb
HsQVDUvscHKU3DDV1OQQvFUtnnjF0M6X/8a3yTRGEXSYhSZNred5iKEOgG1KUZcE
aD74wKfU+7n6Vx9i0hKT46jqsf7GUnDKJOizASaJ/S2R4vkvcpOeDPHeuN3Svx/D
/luMDxuGGcfTkLFqcLlKQOdVnAwxeyGqIuIBC/G7EWfajLEjzFGpe5ik/QAbjVe1
dT4iTh723Pnc5gutpVNWgWB58ldwRtmqmFyKd1BEQTchZP9ehay6tzE7fiJgR7HN
dQo5uCxVyrkgHJ6r6MnIRbbjXC6/swdIdZxHk/ZN1wF/b8aNE5KOEN6ooc+Kzj9m
sqSERdzdWMDNC+hbt1EtvHLYJOX9PXhYjr98YSkOfG89PKPs18dictU77Ef75vTl
uxBTm61MgzZW3ZxQZUVZo3kefH3ekOTEnSADx27Fb8yV9mJRn1QTk3aFYa4XWbsa
ERRc70AnJq1dlgYZwVAtgd6NU0sr+kCpuz4755jMaB2M8clOQxDUmqgrsXv0Qe/w
5fk+8unur+8CIuipzyXh7KL30umLz7gP8Gfy8GBfdEkBBn3KpfFbwWKTsMOIqic1
qF6U5fbhP0/1oC0O57A4jyv/weyHUJJ0B44n+IUORGZpDUOnrMvOwNQxJFjCr7wN
8Rueb+x0UBPB/zH/nRk0vskkMHyKZ8tjUNCO1B/IJSd/ayGMuZT3a1g0dSlYRFxt
PhXEr1FMJtPcDpDdgsKIl0BsofxEz47fMfkawCTX2Jw0hMLEqr12DbX+K55Fy+YL
XyAm9v6oX0CcrE4R/zc6EE69p6ABG1bQKEVXWGbJfvdNlbTDFEtOkY/q3bTWxrPX
JaHqCrmdQfZQjKBqC2oXSan7v7r1juwkmWO58t7AD9r62BgX+txSND9XM0ZC6FTO
O2OoS04AfaB7+2JrzRYSH/HrjGowTFqliUsXggmXsUz7b+Xv9RN8tevSxUkmnlm3
iDw/Mfy54OnXpwYTfaQMjnX3AFsGxGQ25QThYWyi/Vwog24LtwxH01JfBXCbt+SM
bkfF3zo0xfuLJVy8YJKLFIO4YJ6tDODaHhdouWDzUb8k8QIOLbJkeZBzTdbDiU9F
AGpOCH6GU16MSZ/MysrRc5sFK1YW1KLfXdHf2Otzp8k0yq3j+koQfHSrhOmMurZF
EZ9o82Z8HP4TWcQxD9LUXEq27sQWHAAgtZNPvD3IyQV04e2pqOnUOj932kQ/aMUc
T8ifTkjevEPGyTdCyK6/I8/dbY86cP9ZATkAgyBFXgB2xkhd1GlAZf3niYTAxzzj
8AbIzrARFIQbdmNeCjIevoFAfjXHZAV0JWqv/YfqM2i98oL8FtOTllQv90g0gBW2
y8cYiaxKCEdGDoxcAd2km6mjiTrffB2ASxnHrcMikVjBIVwIrDsyeWCUvDNMQoQX
s72d+x395jD4Ek02bTdovgIF7mefbT6isOMEdTr01XOFLj0GqE6A5oEIEIM+Wsb6
iNKf3i4aK+6a8LJsLYhLkuIUj1PTHTXpE00ViyIvQmWL0XHb4EIuYQmzHIYKIzKU
fJnB+zQnxIiSZrTmfu462P9dXo+Iu+Jrf1JVGBTQZsNEsQyIbYm52jBBlfdf/y78
ylRKgbP6qBqCYML2HQfuPR0Mx12dZYwGoCj8ExZttWAQ4dv76nVp7+Ci3siLpIXt
v1vEv4l/orULT/uJDF7qZ2XzLiCOrX5eevewRJu9JzWIhJFzol4h8wyntW5ifeyo
AtvYbgUnLWz7P07C/X4UmMtOHIL2ZDStgICwqEOfoo2vPTmogw+oLyxEEezzzuPZ
nhJqKtdkvhN4tytV+ZLOaiapIfN5hju8tLjAtDmkyM0iXq1hO00+K0gc2WrPHBC5
8Cw9C0yCAgZp6o7dg2FfXragLMSVAX4wi7MUuj+0LCvrg2LOfU+t65ajWMUGYWwV
BSvxT5FhCOg19WEhRZ+429IfAHLI9Rxw58MVXIuNaAqXQh4qbYPmeKgltmwxrjG+
NQNVuyMc3eBtiZZQBH3ExvGjIOHbm++xBYJP5QgISBgav3L0PytGRaIsx5rxqa6x
fhaLk/APRduPJw6OcMF4pbbvPY+yHbMDRVc0por5H1sUX1ZfrK9c4s/X/bZNbbzz
iCHA4oEQCAl2JmgbtxdoIdE1W8gODBX/GWk22sWyARyStATq6UJSeVmgguJzW7dh
6OiWKEyBDRhessyR2PlAVpwoRSmFiiYoenh0FhG3rLWkp33F0AnOhcBReejkvO/o
wE2umYf9ZQEngFfuEw0CM7MmsrZ4XmGheQ9oPr9OpIcmejTrMPxwJkzE8P4dqYyw
/anvmOmcydnEh3g9UaaUoNVa8V9k789BNydxZ4G/ZBJg4clsxYTxi3bAd7dpmC+n
GPGilcOvPRVMY6AdJf+9hsZHEGadyBE2q0pE2Deg1ixSFwY0GE0ULLSbnRqcxnt9
VBsrHx3eyvTxY2FiYLBQi9Z0cx8FTmH2tDz/7rm+sGQCb/noCtaMqR4QwonmzbVI
AnlsEeGFH8LJ1T1dy+gqWMc54S4hHXr/ajhsFAnVY88F/R1qJcZ++a44Al4ep2n4
7oFCb5ciw7Gr8PkbgPxthoT+68iGriqsiwhogy4dr5OdZu0fWJViJJX3DWIUI8Sq
WwH+MQnB/aPskYV8q/FwZJLJTZ3ft151jNDRhqqmFEeE1gjvdJFE9shdOFBiK0Qr
bPowpDch/3yrjmS82XToLoCjJ6c+pGnW3d1IVtdzbOtQ+sQqkr27oPhgmQtY2T+S
PMCN39H5ObudBsoCLrgTa0EZR+rB5RpTpdYorzf/StYkrLorhRg3CjAY1u75/CUY
sOB3YdwkEHfQq+j5aWN085uyGsr6nfEQ8D5pPNXZSaqDb0Dz3hK/xrRLSQE+lWJl
tXfzBAhRdRqitB23vjTlHaiwsPsuCuxcCliCRY7fy0mHQcPyNWMt3l7c8ctyREMG
bketFRTc5lA4bn44oa2nxtK+dUCJF6lGzX6dnjrgzfukOUT6Yvxf+6ZQAT2grShy
NqxdDtOCppMOTdhAYOQOIy7c8B1Dr99mI/qha5pIkGSE1oKi8RasYF3JvtRqfWPl
YA3GZ7QenCxAdjCBUUulbjXm73pimaAaq1RLxn0nAkORaXw9YXnl+HaSi+vuzTdR
RehBz2bPuPV/SpEAhg1R0O5EI5XYB1xFnZS4cZRh/d64HEkxVuW0EtHbgIsdkrus
MNT/bIXuQ+otogXWiS1TEaXmrlbdacBl/s+FN6mfixGP8ECYoIyzbEOmhZXpyQ4Q
kxyBiweXIUbCG1CVg/C/bZBokBTWylSiMn9SCx7ryfTqyf+hyfp00rpLZZLcyfHF
p1ZqwE7TT/T9S36JHQD8q0mirJ9+iD+1Ytg4iPp7uSCihzuhoaiAASDdPB+r3keB
sMIyBkLZNBLizyXJsZh0zFOWhZlwIoZtKZy6w/1nSJ4y8X7/0XpTxFzqo1eDWGYr
rCIOAPYsQjbvxtydMDNH3uOCJPJSpMdRnpBfoqYL7y/TAcj+uKIBp+3ZGAMYIv2+
8ZYfRC64X9qeyQpjq+iV6it/p3fd5EqZIZ1yTwe9UZjuBWw+mz9XRp8HU8CBF/vF
Zx0ldiNGfiSwrapOT1xSXWK1psX8SE25BNC7rtqdMs30jx9fE8QdfPCxy5N6LPen
b/gtMAmBDAtMyTIZWEGoZ1yklolZWkrMwKNSG5bXENgAHj87ywVtQhuZvtI9MXai
FalX/3mLPEO3CH6dYv58LdYRXtVp00hbwdkC3gCnJ5k0tmREn9rmcPpugEqFG5ok
m5mfr8jBDkMgWPOmH/+m8ZQmvHNIy4e9PYZC+GyPmZOPlA0YnqLcWO5kBl71l/Gs
TWUVPtqJWHmPMRiumbcRwr+s7MQVIspgWEFehUUm33wZtrtS9UgO8T+6C/oh4SZZ
9+8V0/Z8tJw49WnYgkuh9w1nYD3VZB1zrokTVcSJV8YK4+YwylfKPKw50c7xs6iZ
1DvP9M44vpgQc9IIOQyaRAPZxC2wbAKxR36CLl13amOAa0BxEqGOGhUp1Yga3ODv
x5iPAD1czv8qmpvNg8H+fvbX0heNZFHZZFI5oVCxzKaRYwqVoWEV+wl4MPFym/SR
JozlXTk9mZX0vFMEHL8YWvHpdkAJQl3OIh7gs0qv9xQe4ld4ArX1xMJ0Q7yPBQ8b
pK8aXXD8mAQFR7PL3lfYfuIJ6Zl3mpITwyKaVqf6UkWmNimuDcXV8kPFwnupRw6M
KpPo8GmIB9XyDzQFT0QyFDBPjIf8xZblC0bQyu2jxoytAif2k8goDbZrsPVyl7ua
c5XVDhLIffhZgsnUx5sLJHp4BsSWbcHd0T01FQUkzfwuA4vW/5cruOxgd1TyBgX0
feW13mmZnMw4oMAhXBeDUy0/Y8qUDhQpVR2Pj+MUIR/wrK8Enws33LAU+wQESuVZ
EupgltbqWMjfbLTP7fYSxkVYHqlhuU4KebzKdgxcH2fq7FJbddrOjSlwYMFyzZpJ
n4OTgu8VLQ1nHYsesvSM9iglATxiSsrQL9Iuu0i8ebW77eS3sEAKO1+0fspWpieF
r2rRQn6JUklTg5FzcA1fPVM/teDQgdgVNmvzJZEkjDehdMd9Y1QUU6g4TSdwRaY2
cR4wauj9+PqprNh5lcMUr/DUvv1bL5oBKm31PuowxcIxdSmvtsv9imuD4QjcjD5E
NAKJve6w8cJaaxHMXp4d7IwQ6qSrOpQH65jzbPerq2Hd1pvIUCfb9jlDl8eK2maf
YOd+I2yLyKDJMl6Q+eNLZw6MOSdfnI2Sp+srknU9le7WNOcu/u3uLa1H0CBiO6qH
w3XJM/tR3tEz7L5vFm+ngc29SGNJZa6BFMtkrQ1dv2oUQdvYynZZOcikZscIpUqh
9qyMHfRUDj+o89kDAq3gjHeaaDnS3mvWXhILLV/d0fQaUmCefagP4dZztospFMVb
G1wyiQ4yT15ESsMwNr8VeajLH76vA3uajvaCvZHGTAgmic66ePN8rXTVfcGIcyMA
RebKTwX8dS/7azEz+OlqiDLgVCAtI+M8vNxXao86hxt3fVFKst9xbep9o8fZg8Mq
uM3M7MFVXd1nujRCxvGZRRqbTPH3Na2xrVySKbVwcrbzcl8uHhuHnkL7Gk//EY+C
6qYi8WyJWpE726VBAwAEg8YRSLH4dPbxjEmEYtZBx1X4WkJNw9scGwlUYg6BDtdu
+mTL7ItWKLSExhSnp6yN67Pe2+H/5JIkU3FEAuSl5ieOxmdeWHJ4xa1pIypEvfrg
ptyCVDrs284xJtFJm5327eq3sgRu8a6dPkzRGjPveVwynxHlaYmSQ2v/lRQw+D2U
B8S1nGbIVIwEp5IgCMgxpRDUlw5jdjsnF4pz7D5Yphjhggu1JZaYtupkcH0RzMhG
yvWSJMgmOYz0Mt/FEQEZrYpuEC3hDbUzcBZjxvY2/oUmNToM4ojndYP6kfd1TKOr
TqmhJucTwYLgwLOCmOwe9yds80/BFnBn403XPy8V1ukx3bRtsW+eMcS7T42fkDj7
LhOamJ2jWvQZ6wIFctp2WQ1/9SBvafpaz2mDqZAeE0z1nA28UPJG6CWkIQC+2I/p
Tb8IM+EE5OJ+4dpJJ4AnfFtDyY1JprStS1OKV34+XGu6QN1qA6ENlcLGfFtvMnEN
mAWJ20VWvPxO/MFgvX7+3QiN/PB3M+pbIFoZ/F/jnQa8eBWbrzmGdXvqBd/1LXI+
LPz0mBbkjofOV7UJvVjcCIphQdMtsinRVjJCcn23BuQ+Z6miEX0hZQLvvm/0n4Wh
xN8ksf326ZTAiM3soq0S3XEkc5FzIZuyMYFBNswFLzGhcjoBbmT8mbNnBHggpf0V
Q03MiFNniHCtV+qj4j+/gZSPDRvmS9uZ2cRmJfGtkurnXqYEcv7y0lJtJJPINcvB
UVKRinwk78odqT/2xhcadQIQ5YuOGcfV7jimAaQSlQmu7F/c8yxSEyklgf2XJ16W
9rvdfZXDCZAr/iUWK6Yb5uM/yjyuXNgq8A/vKvSeE3nMtmwLUeTp/tunsGVr+PXA
MHpM9C6UfCgA5PCF6NJbFaAuwFQntTj1EWezyIbZlp/JF9ObZm2QvLpWWaP+ltpK
FhUPCoHQxjSusW3fWAM097YcaIh9Rp3VQZoSEBlMR03ZrupZjaq7wO/YtI7stdid
Akhe0XScz2gXDdjP2GTwwje7OgMV0Uv4bXxlJp3vkjDD5jD4ocaQxhp+GO91TJ1q
bZ7I+khNJEkeHZP3m0XocIWOZg6+MZko1WvWhI5e0RVB5ptv4iMsMcKt84BYpDsg
lACg6dk7y9wQhdpUCkaP040UmHLBzxWmUSYDeAcclZSQjos8/VBG7VdwhtaIuD80
CcalgP9ppD1MB292ETK1c6jlKOs+pjYncrVh7ydN9vSvc0ELe8jNWx1amJVUrkOS
qqrVd7dld+23yM2JoFTm0943hg+OZwOzc8pibLpD1rSnmMvvRPpsuWXWOsHxILuL
oBiuzBXTiMy4gA1y09BMpoLA0dbVtUAjAGVbpxuY0DCW3aU2C1hZTrcU3vK3YweC
sAqH0tIrmlv11Kodpxd/Iz1LHbeU3vAfAqp9AlzNY2qO7J5pPdCYihS03BQTaXtD
zeDYfG2JQ59ObUEfK/uAlto89BYBnnlDaqCBnXyNMi4X5K38aAfrP9L1Mcw+wPJ4
K687bGgoODoD4k9c+LJb/bq2kJxYHuunacSkY5wCvbYMwtie67q2qdo3HZirnQzc
1kX9zAVbFI58hpikNELE5MVr9nZT8dGcdzUwJvywqUVTc/pvVPn4Ez0OYImGOBCR
kGX4Mt/VyPZvq5/Y7xlug3hP3MwSLUWc+44P2wmIi1DOINSzhHisPrxDm0LCrsZU
kSKBCi95/XtTF/5VujVaOnHLOgtzv4NvSMQS1MCeQp4Zzzastdzp9on3xdH2R41E
58VPOOJntYT57E1INPEry6c7nQlo1ZC00zgaP+/UkKDzVLlMism4XXOgD+nr5MXl
pZNqd67DbDKYWAPz7PzkbTbLTyKCprQ8cYZ8oH2ZwBxf8XpEuwn1R+TMHpdAex5i
pQljtjZz312qlp23OyB7OXxxDN9nXOhn2BQwAeKZTrhqc47LaHmbGFtaL38E6Gag
gwE/dygXNZ1rjG2VCWGYoH/rmX53ptvDjrG+m8GfNdfLFF4nIcJ+sCFFKf6uiCas
grC0tH9m8oQIMdpot9W+C0kb/4TnIQmrF4sS5YW8UZPHlgMi5ruBilcU7L+qBIOC
xEwbWaQwDUgkfDl7FYrnRukECrv3n216VzVIQWjMeRJIYdquRSdPRmsWkdvBvh2r
c+BemQY5W0L2QY7iVd+qt73FmlpJwtyTQFw03BqJOl8IoDXrW2vAwISBk/6oys2y
VHwjGBe6Lwoods+IZBE16gWExPWTWJ16IZASgBghirxyONK6C4KAOGNwFs3Azk3z
+Eh/W1w8XhwPdAclLIgXfl14Yreos+1KR4RITO8SF5B6ixSWHmtcFaABU4JXYHlp
rtWKb19l381a/tdOTTfJym5BSjWSp2zxfNysMAzXLltISzKveD0ff6FTqbpz5+CZ
XXi3sVTjoFpqa7OTNBZzDqWk1nMckXGI+UGOY75iRJn5zs7wScbQ5mSO3KE3xXnK
4oMfJjmzOZQ3l8rlAK5XsI1ehf/gjDK1kz/CttFmU2HUA3u6JzHxsWljq/uCsIU+
hxlM2OWTmo3u5qv2mzwZDpsUsehoA6h40HlY9jvuH0WTR7UDjeYR702aefSR3Slk
eLG19NoSzmqjw4ZSIbZ6vHf5CZCLfm76bDq+H3UoxyJhRV5ojZwLKV85V2ZqPEQ7
wleMF/spco3IBQD2Y1rC/nbzyxCUcu5FGBKYMQ5FGEZJYFrCAjgqQyVvxoRsAS3B
dBPNEy2YOpjB5H2UVdDS9fS1fqv0GWW79ETUkaF6jxX2tXNKM3upwO36quYwEs60
Z+Pr4DSFs+aBgePk3+n+2KLrAYZ14F3ovLoVU9etu1x4AVFdWlb1gaSpuA8470VO
UA/MEwKpRhjMARkW3gVgP6PASU1eL7B6RrJDV7wQHiSKGe9n+6JjXuq6KraKYjAK
x9+9j/MU1DoTpIFi0m/iloAWUISQyQ+/aN5B2fewRsmJjf9LGCLeMpoOo7VL3fLR
LOifElqGoCy9RJc+xUyraBV9ZgCcbVKHYndZSexyQq7P9cwp5dc1MjNpiQ2kZP39
qIbF9eBZH/PCQqQkvwip9Vf2r/wEg2ZBwQy0VhehTOBf8oonYSUiP1koHD0s6hwO
dRzadsgA6MoA1VaWKpWEo5dOIbNbSWUdlrIjiu9XPMIt/zOJM/ZHNVsl1bQMIU1M
pT2Cq7h1e7FrOVFLrlYdP+ddfVNec1ajSeuuI4fX6gKz2okH81SLMs1Oesp0eCon
OuAvAXBgARwFL6uuGeQ73oUKV4bHQtEs7LNLFNklnYEnyRYz8TpeK6J1elXKL8WB
kt4mYjtzLK+/7EDCxISfvuLyW5DMfxOkYM020sT8z0NSTN35RaNEbhlg6+qw9b6Q
qRmzhROzmP53EUSV+5/IW8nep352Dbi6AOlXsLSi3boG42AQGTvHyu4o20Koycp3
X3pinccU3oj4KFp22G8OBb0SQvIMMCMgr+8Ao+Wei0g6HWIUjo3ECrAOlsqbmWUu
NQAoETndiC2Z1Ze2hNbVs9jrc50hL74zDh1k6XsaraHPwPyvifmrP9LtNif/SnnY
Nyv8b+JSb9oGINSFq1Qi+9a/ykCnQy/Req7ZXVWgMFJrVRnfde2Tg6w6o6olbX8A
xNZ/6L1s4R4Y+UoqMpKy3wJdT/rVTBx043gMoUOCXiaofNPT07mAHEQHrOluJJZZ
WN3dbW8WDl2MyWV3GanbvTCX/cG53bNNK3cZocry/RZ6FxbCfB+ud5TAPziBBkZX
Kn0C6ShW7LfvrnoBFHbYjBy6r5bSZ9/nzmuJGl0PhUWukwDwYae1f3CGYqnGrggk
bBF+FqwmPc52V+BSPhwpkG5E+yPEaxqsmE/rzoBRq4xJRht1SIZCQrkyNH+yaSBF
T9BpfVgXFGSQ8ErweOH2hbrwehQqQSl/dvOUT7QiCl5qHL6oHGQtqabNYuftqDOS
gFy/6+Z5x/lRjImwAno2SzTGP5IAQFJfyouVxm+Gqfsm9pe7yZeVyGIQ3lj9Mjxx
mQNcqg5xNkfW2gDDkMgQ4BK1w1N2WlU9CELwRDxdw6yQH6q3ZUr8H7A5FeyIKsz5
cwBdSvCQY04ZNWm9n4y+k3HPjtx6Xg4OJv0OYxoTTHFX1vrVrsPOlN7ZRzH8AKgf
5y9Cxp7E53Dmxq/6VX614eSqupc7GeI1pJKN5akBXRotxhpmEIWyF3bctXzrk4XI
QCMS2NtdzJZG2Wj80xR9ZtgmLzR8vm5T5d3Wd3e053wSr2LrfSqk3+PTkvRUisHE
geDkBccAJ3ZSO65Yh1zbhrB9rKNDToP6+78Vq9XaKt41zCk5uLeiRtuFeXzksub/
MkgwMnh0t8cL0mt+Vg2tkCCJPj9OTcAKpI5cjf3NSi7df0VfnB40dL9I+1fxKm/w
+l3wqijipAbRxK469BQv8DXqUYMpkkP0U9k1d523wEq8Z/MciK8orVH0lXGmdvYN
Syp5pUGu6QrGGrsOKIWWcQFyc2Gpbg1yOk9pZgUA9vxhyDx520gLlKddTYmfidWp
KXUeQbWjm3utO3tyfcWLpPEy5EsVY7bimiuV1fKfLnZ66kU5k9G+aF/5lnB8Shs8
J5JmuTb9wBSFMnJiL7MQa+nfKRHYJv+ZO6mhby3jf6/KY/dW4uCprtmOgfxtjvWL
2V/9IlWp8rxgjd8bzq3FhhFsiZAXphHWuVdEN+5Nu60pmfLeLw8L6rm+fr6uVKBt
Ucvs3wq+dgvOWMBj6jzza9F4h3hmxrhINmm3YZIFtlFQiTtgddtvin2UFelYBW3j
aXKzK3KxbLwqigOP6KRboUahR8HwxVVWBwsFQ52zbfHSOROBRrj4XB4MxLkMQ2yR
YHyCw0/D8mhaVUjWYRdM+GZiawHGk/ZQXxV1BOGqrInbnHpB6lz9CGlO0//E7QbZ
7JgU8qMzKdBWJTj7WocNKK26TESf4iTBtRJVcKqGaJzoVWncZwGa/A4Fc+zZawen
v7WOCTnQ+I66jmYT59vHp4XKbQVuj5J8u+nKxcO76AIgFHhrNt4UQZjeie1wlDQC
mJ4vuSu/C/7xPgLgqHoL/aCF3j3+dPczO6RtXbp9xACKumSpSW3Rx1SoRqht5Nw8
MKkECs8lcOArIO9lkZCShUMZqNNAD2rMfdFw72apH1jGMglXQSCiugJOOtgzf/sc
x1hAbvskTWAxaqFBTyTMWvmW+NMo7nAvHhhCkzkUKxQPPV7Mkml95PafrLQFjoFU
2ogbhRgNeDPRFiv8l5QruoJHWWAJOyKfgxklXNsIVrLOwkM2ahdOrWQ7JhHl0Ril
q0UsWaVV81zuwR7s+CNzzjHQDmrn/FKm+y0upX0znBfGRLPNlZGt12G+B3njZpPp
6zZdE0CEuWkrPXPvZxncUaoKuv6lreh3hAWIc8xeCQtLp2GJZZ60e97o64SdGU5i
nd2RqraTgLghecYVW0B1+jXAFTbYtfL0hm8UutPsKz5+YFdsTzSDOjq/ie4FIRdu
fulSr7xckYhV84sMipamab/pZl4w4lO+6WpVz+omc4BaA1gxjNa8kr2JTCjsCBm6
U5jXLARp6tHP2CfVkhSonaPlTGB5iCZBvoZGaYOftO6AhCJb1IYDCnpVahiHlRiI
e7gSizVzEy3F2A0w/fB+/bNR0A5iqwde7tbAXJoEYLJj/GCWDVSEqj7UeHKMV5mp
6diRk7397iPb2NGNPtUScg2lbbZLVHRv73v6x4cPAsroEfdIlQ1Vs/h1FURq82b7
YO2nD4eLoo9epK3BRzeYRPR3GgAkU7b4CHkADtqtyD5xmrhiS1QhKjEHAyh5yyEU
KJTN/XvYtQgvPa5r4wykxny96DFhoLa+G6ovLFV2epyQ/pbY+hgiXJ0L76xsysn5
FVvb9igrCwl+VP/Y1JgNFE/VukJpo1eqhJwqI4RiTA3FmI+MP5khsEYB201pRYEB
/jPGA/MxUskt7Z4v/LbI0VJlNhiuSBgD8yG+XFtqsVFl9fUaoQajFUvHIaHZG9NX
TJPvctr5DbxAHeZjJohpZQlVLhRmC7eLCtpjhQ5e666B4Mf09ZCWwnvjYuMUPdbg
0K7F3m4mLYwqphZExZsw5dS9MZqqckb7O5dZobh914crFx7QQkLKqkFssgahwYKM
KHVhIu/grGAHNaQCu8MLiqBfqfwYmBQZhRaO4gr7lR9ysULlPGFpiI31DxnjqfMK
sLL5ZafQ3EypZtdwe6o4aM9SwqwtneoiF4Mb1yo7u67jXB1EpW4KAuome4m0Q5u2
qtetd+wPqBljxUACr7GFRIZco9LFUCs/DT9cIVqkMReFF9CoI7YOyUlSxgBZZw/W
MMGZeSfaekackJDo33CwplLbjuBk2dRMKhM52y+O8I9WquJiwqjPkdRS8B2TrUFY
+PbKrUhusPPkwZpWeZMUV7rWfed9dfNb8IqGpAqiDK6wyAtgIaKLnCT26OQOKyUO
hMZj3W3VlqyVFrwKRcO3QEzIPVPPf6+SYapAMa1BehliJgZ3zqsotqMOUidkFs9D
AqZoAi3BhTuQ9G4jiMwgZTW4DvWoXKV2MOze9VfnWmEKzO/JvQy1T/KMS9NAHG9J
2vUe66jweD5svAfUa8lZs3qYJFigVqTqXnIERb9GMkCewlxo9jNh6gFgp/xj+O/w
28mmlg48DpcWy3RFaDm7hy8/WpBJlhTYY568s9KL3TT1L0bKKQY+r8ND6HH5mjLc
TV13uSlAWAwOBuJdhmoPWGyfVDn+vNBH0KzL3eh1fbfgnrTPbrWiy3xaTo6cBaFH
EEya3TOFYeZ3b0DcDiwIfYRuGvLgck/6zjH2PLBiasphA9W8OpkS0YP1rIlqyCtp
3UpI8gJc75nROjkKTmFId6fhFqdnM8T9geSUepFzuP3WC5TFhzrVsi6pt51pq5R+
ZrcMJmvAwudpTnm4Mqc9vbGxPi6EBMxwrhLv5+MlZPFkqGl1WIDZ5MboUnPwBtkN
05Pnsyi+JUVVme2uCndndc54qsqCJgn2fhz2gnWI5BfeuT41YibZ9ccG5BT47APD
aUHB1URUwAx16wUiK5obukIUu8wUV72iPrBMmUbkh2sdKNFgbIQxQldKngVQxQRH
Xp8nJbplfFhQUJ5M+jZJajwZx95U4KaaQS4qd/26owM9moMSJlevTFOAB3mmICoe
bo0GDOWMwrO5xq8e0P/lC451NudBKIHwoGH/RKiDWKmuXjMruu73zTjzN+k6WTEW
akbLD3CHQhGpIDuconWl38AWQOnRqlx6mphrI/MAif5p01juPZN2tC18wostAItL
Lld2A4dXm4oATbXUImoMfDCdlonVif6Kjl+hcJqQ2iwGLAD7yJEUVeqEC2bSxpDw
Hcpx+x43c73EN8RKIuIs6siy91xDssPL3ZnzcegbvoJEYQdqwui5HsKb4p0TLahW
XjWKtFElsHAjWfqsKOITApwfAQeFRxXwskMvHzrHUwnQpUp1QsWeYS1FDieRzhMJ
oqjFJUsilZPzMqqsaji5CflGTEB7nktfW+fx1u7K4gh3qSAI6Pm91QDQL9j8rjQE
vN/r/4xOFoj5ZADzUKf06z7ff/p8QimlIrliwZDfx+nHo05ALqiGu9ScmUMlcxot
Q2Scmsy89oZVJzMOWAdmgMl4mVWt7B7EZz/Siw5xCTQfyhgZ0H2KpRXSlJEOUITN
S2Oe7vtGbNnsUUaJVfvmg5h5gDpZ7+eC/KW3jU0RjSwOQVStVhLykkjLrnWKqscI
G07guWhXdEJtcwINXVFuD8KoARWrMcLx1/O/Pk+ayt/nI0h5sCFXu4sEPua8k1yj
YBnqZXfgz7Q3JYYyYI1PDSi+tNY/mkBGcOKWOM0bFicoIhy8H5RUPb2DXMDx52aM
gkp0zH5SHQZifBL7ckVeebvDOpG65DRIO5xJVU9KwyFNwgpaZT70lFeFzFmku4X5
1zd2XuoxPi0w7ZG1M4GHDQ50ASGh3d2fZoU/189EfAoP/4t7Tfb8oOM/YNM05oad
oz6CzRqa7yrbxEFd/2qtt/GR4wluRN8lvi2Fs71ynyDPUydP4ZI1jMG8H9Z3ViVQ
PHIJciLOyXJX0vQ+PrA4UzyKeL+g1juS9Y5y1VwxPem5vzrmXX9p2j7yYV44muBa
Vq2OvU9AiztpwRUYFdmwmlLcWmSw/h5j3RHYnZhXyNKMWIYQl4w6m7j30bx40xMU
ylTt9bL2Q/gqyekP/lsA0hNqxGkFgipqCRXXOhkVSUO+P0fligEx6Mc3e1Ox5Juv
5fc3cYneDSAk/L/F0ni9snEIkndkkL/Rb/tptibiEkkGBgvgjltw2TlYa4ewv5/C
9PS3vCzKiyDNkoCQVeNT6qU16tbMPJRZi+p08joANfZtn3nQwAzjcA8y4mmRiqzB
bXUsjru4Aj8sv8J5p776y9fXroZp7Efo0Xfb9TOSHBCK6SiIupkcMQ0OFLptNtkk
WeHy40KxCIPcKS3ZiaXwz0GVq97yPrUcSYETnUK//PKcOQf1koatYCMckmmUQpAh
gK75B0wbED25Bv/s8zYBSONBTk/MhMRUM0dgHYyIZR0CEZGrDj5NblnaHyRxU3il
R4Z15likuc9e3a4rEi53Z996K5ZpW/ASFTy9mvmFD55Zk6wkQOATofjd0ph5ZSRf
A4iOom508gjwcJP3HUhvuMwdI8tQYLItGLhuXHGiTCi5d5lfs1ORUzZ/s/1VsaCe
buLcnrmD/SoCQsKVygPwDd58j3RG3N2vjhgmo0hilEpG2iU8SqizPpZRTVQRyvTC
Mz54Itkt1FC7gXWXm4ZLhgHUo4QpBi7n/ax9ouLQM9m43r3gdYIIctWCzfagUw0/
ffS7Vi7kITI9R8i+7PZByEgvO3x7gYfOtXXbQfXwBmLX3waqFP5R2S/bsd8K5RnB
7vyHiAXeoXb7yRyRkcSMHkoVYwGxy8sCExzHwHg+qyGHmFZblOC8+JcZvy5GYt4X
0Yp7MAOFvPc3Eoq1AswBoWAlzoOxlYC6C/1NV4TLaGYLCdhltOi2qA6VFcfon1Rk
vD/rOBgVH0hregcteY74l1GWP7ACpElv2TFeqGc6xMnGjUcWcCGZck+Q/+LU4Eyp
+pYuDla0Miu0Rg8PfjMhrQp5METrtfVvwroWbh92H8tP5d+Cr5VRiccqZoSAu3YO
leOJZjRMP2Ws/6cqMaALzTXAS9549OKaDrtaBm9QpSjjpCn8maQAz3vKWIzex5t8
Mr51CQz34zPGxTA6VCGhHzeDVmlvAixxzFc+/Rmf6aPZQTTtJ5dBuMgoiJzFkkHl
Ed0olRBexfZKvKse156JalwdljTLWiqxZrt8YLPI2l6iUQ7nyYkaQytuKyui3hi+
rWRSWLqHmiS/MJXFe5ofsprHFwcWfWNgLDu25HlXOzCMMVDQiP3+pMe2eVqMjA1n
XkVqqDfppcqNkZ6AbO2dV2VXwxx5smhS9JeDaZEkvE65mJGOjXCYXLulaKNLaMiV
KGWkSvdzZ54PnxNV7LjSvpqow0q8PytJXPgxCpluRZ/nAUdfsLH67Zb4AAG4/iE3
9yFln+r+XipehSPl8vI/vuAdtcmqsC1IhV0TfruP/hG2w8ePLH1FP/HE5u/zwj+7
fVSlf1+N6gd+B+Zy3uwzWAhT4mR7qsM1N4VS5tzfyaOdPkKPTVLT7HtgOnJCl2ey
YESBr+IAsu+Q9X+Yy8sJlOmZWKJQGq1my01hGw9eZIdE2aDpgB4SermF9CCHGUow
kXa4ni/lNCFADmyVOZMWMPtdhSwvGkLklKWIdqa5RtqwnnX78v4i5+OTxtZo4/KZ
iWhHW6+OGYLxUDhaTpZHDAoKGRjCf4gS/9/rK3LMMlRjlq0Sq21RjCXZ2zGSd5he
KJhViPeJoahIoE1VVcJAC+IaT6/6hEKTlQFFQ6BomL4xpjtYS5X5b+IecpOMFOV+
vAB5FvnqtM7NGSm1YceVmJAjTu7v9DZFv4ibvEgSh2wxWnvCY5aFqOzEVypGv0oh
W00QVJJ1vRhjs8aO9r7LaVCYIbZzBnDLyROyXBx+U33xvOKmTvFU+UDLXAhGiU9B
7NFUYnJnhmFcgfS8pk352TzvFUczmNEJlwMLQu31E45E8EQ56/ODgBodk2hR/kKF
4RoceXKUMrgTN1TSohiC1Snfj1A0t4BL2gynpOctT33MTvziBG3ZVBYrLtYxS9zA
uaTDKF8LXQybg2ZXzD493vecf4ryak0UI2uTHyy62xyx0nBrCImsdJkCsBHrP8eU
xqF5vEoxz1a7dnnNzzjGIxY42wpbLvcCr9KhtaWS0gvOAH6yyibA3jiPkHkt/2q8
O63mtPZoRwRWsDt/7i9DMGf0wiAMgOqxKpK24WWmpOK9pHofL19YP60nvl3WYu57
8iADf7aknEDATC26NigjiUEt+MkbdO/nKP7QtTZ3+ID9xs8D9KC/bIgxubM7/p6M
32xnbnq+4vSNprCVOecy/Fqm61nRZVOlej8Qn2dTa1ODzbJawGuh8C8m1WhHl4S0
94zc079vlAcVytOIVeUchrewNt1n0jmC4dWqHxxHXjjyxoPSMFRplSpsKOoSNiu5
v18IUyQ7FNw+creFyyDpY2oArjbHqgf5ilXykCyt67GUi+hxa/Dv56nFesEg2lWP
MGb7ooKDRdqHHpKFnJB5GmskL6TYTVY8pvcfQ3Dy6BCmgs3tdQiNAhwu6M9J8vB5
H32Wlb27jV5feyuA6zEMPGPTD/Rqum+NU4pOpSuSrwAmbTZgx0fd3ESOgHkKKiEV
sfy2U5nUsgeT/scL1ttI6V0sFZQxc1ZZyhN6UN7vYpgdDtnZWoDgv8TZxcMNBZqy
cXqaO7Ta0coKodEepSwFy9G9RClN08tJYJzgqk47oKK2n2DZi/df1qFf4FtS3LGi
ZotiPxLKzfJr/mPFHCLs7Dqv9AQTZmns23kF43bHbFgXy8OzSlxTQPohBmWaDjq/
WEO+L5n2lPI7pFhVEuCTJZ0+SQLpiCal02jn4vt0DB0tfrYpcjrMpmCHAY5Py32P
ATnCSNpD5zrSpYkGI6+GLZZOB3PZCNlNKnQweBHszzSjxst/INGCG4nHJ807H/62
YOFSfF0taExeFdMowR5/wkE+haZvdTmMfZcmAyuj1DPMylEHoSmfAQoW/AtNWXRy
0OTg3CSZFBubFBIwwWiPTBlPoAG218IGyRU/RSJrWhpaOF+nBTVxIfWOlHyTkd16
cIrrSW6oUNWyOY7JqoJM8H1bJ53KHFd6pFDr10i6mjr5Zx4bmUF5L7hOIRU6qml9
TK7hwUXfprQ0CLmuvx8Ulq5e3Ma8xnsuw82YYSFbXHqjY93G/oFELD4jK0PdCciA
8nm3oj2B+YEILYdtpKdJhk5792PK9bFpfEf0DY0h7B52dBePu2LF9KCE0USBOFv0
NMVPE/6hQyZQGJOq903OkrNPjurYpchUY35i8faWRQusIw/OYZBXA0Gza1SYz01f
BjwML490yJhKzygVYV9fEPEC3L/3tvGG2hkqx5/Gj9dBdZ80RkGo79upX1Z/3vBJ
tPIanuUtPxD+uJ/I4UNZRcWjt3nu7IZ4d78VXSeegtomRx+3jnJkkElKyEB75p/B
8wyY3tRGjdLZBXdUeEAwCq6n0zAGSIHf8YytruWYy+jcSmgpLEeYJN6TlzJqEkTn
RByi4BHKWaOW1R6mjBtXOZYcR7CJsD7OfFIqT8g4pUFaKyPyYEx9JN0szZq4lH+F
39lXJsCqgmAIgejjYMgojYRP0YykJVb3q4r8bCLnFenLnZXKKYPJIx8cQPGNbK2W
vvZQuPl0pdhKqvLZCOc0kXyVmF74kr4b8utIhwuq55kJUJBpeHt4ofuLzuRqtMM7
wDzbpkl7jiPQNS5rqhRYVyXgWQ1ejr3MvC28fuJ16uhGk3idx+ziz695MbSn14o1
IQHbujlMHRdoP2WVzhMHRWLJ78S6DTGairPoU2Dorh/NwKdGA+LHjrMRyBRciWly
Omc2LTsh9g0nzHdMI1G8FChcPfFkBGjLBQOxqozCQIOyHEFmXYucjoHPRpZNak4r
1nIEK2M4rNtzVxnBvB1pnz4CytJm0qeyPEk+cg3bxYApPANe0osbsmLbzea8O+6u
Jhi8QxC/huPQRsXRjILzlVnaHIyOFfslmZgFCZ1vXlWmp6xsFuVDsJlgiylJMcgj
XeOe8GiJzBYrwLgnTHcOuPumkkGKZmCqu9+iXS7CWTXC8ZjJxvMZJTUqmf5JzrOs
pf71qZE3IoFlna1tBV7ljkEIzl/IpuKontrge6PTK8mKbAhTCf/tVFZE3Ud+RGXU
BtQUPK/wtDCchyUnEXXIy4nmW8FASCDEq3HIxb6jGuSVgqcsbK6W1MQb14YGvYQe
BEF6OtTY7tuXVKiZc7Pv3uR3Q7drj7BJndVmLOKtmlhnFmWmbbIp+adfYFfdFSVG
CPTddSdRQRujF8VvtJL28l+e8vNQWgu/eQdP7YsA1yTqgXAwIz/eK3d2uymF8cW4
jbgaMHvZzwL0NWlkdIPl1lQfA2jB07w54nQP4Pb0PfcunRCc5n3r4iFOhLOlCRGC
adZ2usxxnGwgI7kQePGme9hUOCLKmYB02GX7btvGFYoIRj72/uO+u672Xh43+EBz
IJ5JF/klzM3WRnrOoV/2lj8hSgFNejguznJ+hgJDePjaNNrA/mEeP5qOAyNTiMSQ
1GIVYWORaL6NXd60qxP1MKyNzAMibRM8cSu8yDW/e6eTXW4TUj/Pf4yaAnNTTnnv
sLYDj4pMYtLb6Z4l8yIP5OuLzjboSMtMK1bx+Geu5ZfgHNO8TpqCWst5rdt1uM5T
eRo+n4qjM8muCxMvzonSb2zNuGhYBNN0ztFKdU6wSZOP1wuc43/a92XdKXncY5rX
3eMCeOsFogoRHSSKWraZFcFNLSnF6IaZJWjjpeuWeDS/uICSXHxFRloM3wW42pvt
/NvnWVBZOCyCJbZOYuJTGwHGJ2ecvCxpRQSfk7uQLW1Oo/9VtXjSWuyPIMur6Amb
Mjs00Y5q28cqWkqPcBgsLks0dnhr3TCDcNdk9/3IDWkuOiTyeqy+7rs3fhA6ef05
FTpYtXF+BDSVu6WJWAjmCYvJU4ykdrrP6RUNvWJjk090ygsmpOczhI03SsKSiFge
RDDJBEtGkINAgY3OeFsTBacN2NQqyp+SgcDT3QWG+NK/Nacwii0AIkk0qDEoJJYQ
t5W+T7CNma9SOupMaQZLZ/r6ldysi51RDBjbGf77PXF9gFvmJkaaP+RoberEz2wr
4wkrSDnsiKctBucAQBaLN6H76n94RsRNkvL9q7xQY/qTbM80tI+atHmaXwBcRgRq
OiTvg6zD//sK7/IbIl0r5t6YB/ZRwLrqpTm4gmhtdQlZwl8Tu2lAu4aJfbBC7OwS
Ge58BhREPIGUMB4xr0Zkpp4+Sw/wy+p1PKOlTtN5L4cPerhSc0DbatCuOm1xBWxd
CP/272B9h6kZgRsF1T8/t2tF0AhOtc93ZG1kXQWIGWZ7evhrWYLYSlMHz0/YaFgj
6/uVx+QiveEqLTXPSMx61wbrl18BEqumAcZPFM8t2w5cPYkyl2if7Jru5RYP3cah
ui8/Se22nJoExJ6FZuElmPYRz035z5uNDC3RBy1YBbL+i5u4lDoQuVtKq7RxspOw
ZEkFBaQ1tiBCeMPbHMMeRB7IO+gTXenYYWMzxHohKk3YetWTjQtoN92wpiByaKEk
fkCTvZ1R4EyvBK8GQHDu3/08xa2zbXsyQg6p1R5AR2YZph7yiE7KvpcB410/fNas
WjVuLVSv3mDz0PWI+wVLw2mPAdlPqQTfuvtEzAFrXkjgd4dNqGSZ1jzpuDhSpKyI
PfbYZwF1ayAXVKv10x5ITUbriRecNj+DMtzSl3GRzeHY1fjJqz3/qkMMCagVRL6q
sDYRNS6SMxEUBdH6165SaG/5bcC2pFMlicWj1k+EqeTHibakvXiUyetLYSBIyon5
183Amm7SVnUyDwBYC6YfLLkk/B1MysvQ0TJ/bqIZ4VescPOk7UMhtoD0Ff2PeMSn
dZsCKryvC3RaB8hIGNMFvEeeuPCtNhkJ1G14yjW8CVF9C65rxSgQbsPMMl0Rd04A
sJIAHTcLT6gnICeQFleJptaLRuZ6bZ6PrejKB5yESOubLve3Ette7Q9Vk75gNFOS
133TZJlHD54L25Pk6AqsyE0uRgweEh1G/XeLrtv+9zuw/B+AJAg+/B6+OCqfmH4M
DK8u/izCG6nzzdUYwuYzGBlRN0nC9Kv5SF1lu/mQ70J/Pe9TfDhw6Ym7DnYYiFZG
JJAYLsXUwrr4BaHa4Q//yvgGUdrABZDMAwFvlu102s0byh+BILjfvk+v02b63KF0
TmLwtP6nm9RfoSWI1guRHuu0IxYemnx0DCzDhBNyaKRzN3iv5NZQ/3KZIWrt/sYV
8bLI1iGZYQ/m9nOXk2sf5DOLhA7CI9L9EDxTdn2MRJHZ2wdF4jKFfWUr+dYrmVtc
pm0YFwOCxFM5xpj2IY1qI3QbKke2nUC0qm/JdOLBokuG1Y8WBFFOKBYYpTQOnK5o
C32KEzjSkwSQw+nvM0Ejicc7U0FfSZxBueBfmFPhHhLMmODOfl2x9LzdUsVSbLAx
AW3LCFWN+2hXbM87cw+EY2zsFJZZDQMMdh3qtUAkCR5JSTunxFela+tNp1LfGHtU
EWCvCsH1VjdH3crlE1erEXUZ9wEl0Y/K3KOjAXx+NOonGdsEVPt1xpMZfHnoJY6B
MTpJ1uh0VeV1goC3I0xQM7QyQ2bGdLbHbaO0K6QGrabhgHM77AqENvHXEno4ey0K
tkrAErbf0r4xEBRnhMOnNacxE2Gw8YBLqhC57eIYIhdYmiMSOjgfq0nA7b6hJ+PF
HAv68B+QddOcCQMhyi7wJ2qG+BB4WL5td1oQ5Vnsz/4zWtCyFIJVGN56YVsJf4yt
NvGLp0KAk6+DPVk9mfI0Nsj/CZFnN5U38SBCIzwIZYJujHPxQRcEl6L3XpEMBHhC
QISdI56N512bma33yrgaj5lU7VsZi60p18J8380rHz4B7vfbscklzLdJA5J8zTXw
8a7IWIHjEekIxrNMQEDF7HABFQnTdL1J2Lv4Cf+2QUIWc+YcSbnn3tuF0gf9+ccA
zYSJX9ePVvmkIWPZpChZzixkfQB4vsnvW3J6NwMsB5DcNId66ZK4pNsJxeCPEzWn
XM2TD822B1jlxeqRgnAcUa4yS1XPHCzELEIYV/j0MG7oIoh846XgDgHAFEGsh57s
KeuVkUemVaJXtatJ9AyfGm6qK2LP2eSepBEE8ChAxHI/xXuE88LMS5+cYZYohp06
myjtvUds5Q2gX/ur3FIcX3tNdXWgjB2zh188mKdHzkQEgW+gnobbjQWGjt9sBW6E
dnScr5YdvcAWfMik2W1ugbs2MDzAW3ZBpZZ/UROPNZTJahPK9aXCxtZTPAjsp0Rw
ygTLhl4ufQkdhFWdqwRP/j2XcW7j2FiASOzN62fPfgWR7HOl49fKjbjDqBEYtCAv
iE6Y0Y0R2XbvJcrlWMQNz3u70QPN/wHC1pcbpqAVHtYbOeHZS1xoV49b40gPWdZC
Rv+s7Fil5Kc02JN5xpQMGeRwfiXAIXhBlRja0GTE8p9nEXcJB7cw0TjDMV9QR5mS
6XoceHHZBqPIZrpXX4OZU2bBmHD9qfcoWD1V6QEq78qeVYtjJXvotB5qA+7ExY1D
+UxBi3vbSl4gDWR1kEcYu/zfEJ4yfbzaZGx42wAiydxVRIKWyjZA9eddB+tjulON
HEvBuOkQIEwueKGlKQUYdwtmRtvmub3oUH8H8hiH4yCukFTarp7jNOYg2xevTYF9
VL0gatNLVzmmsj7u4AEsQDg+CG1KbLqznGiN/lAbyFqg0YwaGbbIKH5fflryHx9m
gWHiCHdqhcOygq94EB9pAk6QU7v6MCUrT7QMXY6C5FNJCqiMdWDgy+FGFW0w3sNX
V/8YZBSIubls51CZSjxeUbg+FUR3aqeCkzQxjW+FR5dWlMmzu5Bu/ieORnP2j5wx
kvD2Xobike+w/9dc6OyunapzIHcOWJ8RPEVlPJchET6/TNdKUHxjcfvmyi8rRL5R
+px0SKjoflX/lHE9rXEGjgJI0+2Gx6mr1z8ar2MkhZjN6RniwjkWJjsN4CYU9RXA
0PPaWLb0NUG0GSLsLPUTwbVIJ2IlklB8d0658Hyt7Kvj8kP5nL36Rhzfj1vWLC9d
PBrW8THqq/NruZY32bNSe+hmFgHVcXh6+mJ49O47GjVgJ5YiF9jQj9q3SlgFB8yQ
uZ0DRAdn5tRXTe85rWSbxtt127ldDI6sGO1fa9yjbwIap22AhPqD5C4nSGwMEsqv
yKpeXG/BBRxYQRjLn0Igkl4uXOR9gFd0bGthEjCY6nTvJR4xXNYLXcVNuvyLS9SS
m6Bzrb0oFZ7XvMwekWiUoc+/QgexK7PFT0M3AUlr4BCbyk2RY02tZwkV7seklahu
0xnmOQTmEtOHrm1kSsnDBK9treOAnehUDeIEU2l35wdYjvCFP0tyvPlyrHb31gTv
68j+/Pp2cqWUEPnJSyoQ6H9yxA7SwB97adL20myILdCWui35VERmwrc8rVgMyVH8
Iox6UFHd7GVMqARes9FmlbkUcKdsl0towtrZ7Y4Zagy/Ao0MIL0vdRMJk4WdEEY6
W9tcTEqnTt049ZCpZUhZ1U6i6W2aLvU0JNUGtq9ZfW0xJcSRYkjN4I+aCXJ9Hose
KL+b34i+6BEm/hgowMx1U+0aQXPm2xaTQYOaSa44srlL43/2oEaENGKuh/2BPeh3
FExRmJtbALiR9pMd/pk6irvQ7ZpgNoudl+RXVleCp59GWAnJ0DsEs56W8uvV80DE
KhqFWW1LqgissPIi/iCpnmJ4aFVtqXddJBZG0m9FhowIgxb9FYkE/0oF98YuYw10
xWpThbq9F3CiLMNK3M1lbC/xf9IkH9+k+YnGdf/4X9SuyJIKmG2WHo00Asjhx24u
yf90p5mU/NoG8YEv8nOqOWZD7EMFmCZq/H02/nOvGf2IBZY3z/nHQnW5MD7/TnTN
RmbcA5IXYYgks6KDE1MaPGCciV43nk7jh9sMuTXuJ5aNUNhmovGqxtlL5yQT6T8h
OnoWWIesNNyYf014JZmT9Q1Gqh5rUPa+hnLqipcvMVhb9kcQogcfwJn6KYpQyhu3
5Iul1BQ6rx5GYANpuzEfnbAdY3kWh6dCG8pyVMkZZ65C0gGF7x1eHPfRhWjCx/8X
DYc26lfi71l7bioHf6DaWhrVzjTsQ6AzpdC43ilK+ImnzFQjMoOkJ8SwJVQmXY31
b+H8b7WTA3KS1K8fYvu/krol7qrjIDBPbg0nuv0m2/sVjeJIJvMB+6Kf1fh/XAZX
3ffKzobs8+LWzJXLcC3z95Q6OjW23TZTBjB9POPKIoaRFu2dPIscbNuLXqPw+5CB
bFmTsJkrKNtwgEcdzldElpZmjLJmRuN86ZG+Asmt2mBCjGCxC/FCr9LPnxYpu/ua
At0x7H41Nnzh7wdNkan3jMdsgn+ShCA9Jdf25WMVum04V6x3JdfBYcSrnXgzuGZ6
ROiq4uQjpoyp+VEG8i8QxTc0MvmFIa5MlYRBfEqMdXva5g++awFdHY2tNGZC8OyW
1i/xWEatEZtSl6/GpamODWo7n7fXs4abl0erwHz0eEn/FajXmjEvowkpUvUbH0/j
s3+Mjj0z5399BwhwTaxeFqSu04FETPt8xxz5ZB5zCPSieucFCubXMmhlvouuKCt0
lgW/LTa8sw8AaA+RKM0n1VpkMCYE9Y3E+95xQFhwnefG6AlU1kc1b9p2UTaG4H8m
f3PRijUdmQxE5ORxvl8EdzB97J7QI2UVv/3GxmQSLen2kyn90PhkXD9t9oT3/cEa
GhCp8gZniRpCkY4kTE87a+EKbA4WsJBHpj0A6QV0WBENILuRdfj+4eAE4NY6MoWe
Y+NdCIvV6Mv+6HJw42SaqDXnBCjPMalTKGhMRo1gtzkwIQKqp6zAZzGLYVQL7Izz
OFWbxiH+RFKWAtywiQ3rmngM4RN407sBWiaLJEdZnIwPpExVsDV6hhBLfUOKufxG
Pxq/MxkuXDxQyVK9aeKr/Ee0tFyEboXsHIEEqQwiYBoqdSGhSUYXW/xPtQy6jlXm
bJGrYzsm+uEEKLrJVTXcbO7naEj1W/SRCNIMOUstyoJG+sN6AGyaVD8S0yQynjcs
RejLU814cSwgSvtPb93QVPic0hrCsY/oYOjZTe+KV1h01SL6FA73uL4T1tE9Bzgg
ojtkrC/LwHZ45X7e0zK3gxL2cxlubpdiSFglngQKWhJIu3sZtoeeJydUaoSDfWeO
mKvpRKmUMNLECPK+FWTOmDrILuvJkeZ/ScWA4wolGbd+ReZMXufOtFHuHU3nk2Ro
PmO8gTEQm/2OJGUR7PZCzDYW6icPLSyiF0F3XJmvnVpdjRjC15kYl9xDdMUjmGRz
1Rq4+3GlC1ySm4t4QzaIHQg5TC6dhz+nUMq4jeVYxlvlaKz9ZUW7x+ui+3W1tm1Y
C7/Is94yqiKN1MMDzUF9+Nv0mCareo1+SwCekW4lYSdfYGULwLgA0FT9YuquO8ac
zoUfVwP2EC19swa+c147T323eVVlPM5XYTXNRf5bkPczuayY0g4TDb1HIkxOw4QI
BMymoruBf+hqvDWK+XG6Yi42LH1m2X38GdHOGLoHHWy8ssem+sZrLRqQ1II3dVXI
Rzb4RzfC3TRIcC49i7gbOHnwQaYT/0ODP+pGNFtY2k9E0Gpm26hKDxzo2Mlso7sw
GyleG3/2w2GtEzlkNcfdYnaR61Amt/ItYapBg5UlnHUtNa4gkb/F/nC8qDWg+zxb
uN9hBanqm6bwn7L5HbIXegGQWF1h3msKylLKteOvJXOzU5vArg8K758OGnPKkQJ8
KK68rfTJBUVoGfCJiYmTEQZHXnQ5XUGyplEVM9t8kgO2GXSpky/V2dIgrB24TaEF
1FAcQ4lGph+fkzXV7ewH0AB9VPwfj0oZ/iacc86tRmYlwppAZrEPr11MBuRb+NI4
sTQXjDDxOXP44Uuf/4LTCA6Z2I3tOfHlSbYQBJxvZL6QyLMwDJcGIKm7cLusIlJ2
r3IvA4kUBo5K0GUpDIYIgrCirAbXynd+Vz2Qc1LDEpW3SUhKUC/7H0j66x7UHW9S
5n9kgDYe3uDQBeNFDz2FwupZRXT9omzt55XZVQ6jWB5Kb7uud8XkzsWM7yEfD3Hr
iN/Qdlo9qPWLXoPwZkGNvIce1t3jeS08s/JZkZrL5XrA3Ig7fUUqcJNEYd9cRDCj
Fc8akp7hhA3C4dTfO6OeV3WFcXF6Ixjb4y0+v/HeG5JaDnyBr1jR6SSH9j+6YW/A
cdH5xff8aM/+PYwwiW1/XTwusuePRcS6hTMWIp4umP49h8Al2Uec3E8QUfPsMdaL
e0XqVHDEsHyzS3hIkDnJH9lhJ0hnLbP9Qe1TizYJSekWj6sgtfmpqoSsPasl6ur0
+UQwYHLaMIP8ynH6YdWxH4mDfcB3V/qBi877ukBGX5Xm8UgUrZvdwQQtP5EySPgk
TW+sd+5omElSOs9xqS7GlMKqMeMb+Y/mOkQhcA4mRJx/dTlShcUqZNPE1Q+lga2X
c7gnkBC5ikrEr28ZZUkgm/uJl+JT1W2z9Gv8wo70srRcowTzRPzx6/KXdCEn69Xt
Jb1TnZkHl6zsUwrrrb8ihWAwa8GriFTz/B3YgvhLqQrMih8Mqfdwa4FAHmQbM41Z
fe9rYk67VvFPoNY5qEidi3VhYDdvaF9hcZHQjdEIDNAvkRQz67rM0xNXXUkCyD2Q
ADMAuwlSpIuQN1xOzNd8Gd21XccbqxNPtxB75WToHM8foa+nfv5SYKIsDv8LwFv/
wwuWmkloeoSgbPu89iUBzAo81ij+96GTs/NWJTF6YbVSbtdmV+1S4JZSo2SYObXj
0LnGCljRBxlOaYubJHaoYlwpDVFH64fj61pGZ+cB0OGu5SLw2E7kMHxptNvdOjDl
CpsZMT7bu2KGw0gAQOsEm1/uKngw2Nbj9KuG4MkLIDJASXFvzKIpmlZeNGe6P2ZK
448OFE6qaW2SYbLt12l4KAhB4vttd4WIaKoxOeV2N74flf0YYJOkTiGnaXKLYegi
/dWi/q4y0ieWCeUo2oZpb0RKU+HENceNhwa79MiZ7BhPZblE6EG5BOMyHvyznrNI
oBkDVyHd9m67ij2nNoaO62FCja1TP4U6PfSWoVadljXDD38l+QGds8n4NxrEcisP
qr2RflvKSCLfeFaaA8yF5pdf4SsODfNrdOP2ORMX84v324+T86aNPGnhszgFdC6E
05w11dq4yqO0GEUL+iM5zkLN0eYcvMnB9hUfW0hSijp8aVcavYGBhLLL+TdljI4h
6xGSUrRYSWw1fEcyRMbWuglB8E8gzTpyxyrM7ZPAu/3dV8frCO1gLaDtek01Jegf
J2zP0LELOMjz+wCrIyzJQ+sY1oFTOudr4h6drugJGAr/+3690hEEvUEfgVsQ8NXs
atl1/tE/RSGhi3kLyTkkSojuleseBEClZMo+hjiWPxFXRX0felofavAsSP0EjywM
ZDOrAAln4kWWkmEhtY8mARHFNdZyezb7owVd6uMTVxPWJ0rCvyTomrAag78DAQI5
ecHf/9ZOBd1E7xnhVOu7t+cJIO9elI1NTfP6OqQZMIzwRQp5WegxFwXcUc2l3O7h
T+ZVcXa6Y9RwIvNC/g7jlNwXCwivxJhges10FasyRBVqj4bJNC1/rO7+nqytDak3
wGVFO+fUdoSCQB6xr0cIqumT4rYaGbq538ggZ6tSpzNEvomjlMTOxxKsD247o8WT
xOx0oq1tW7D19mHswRaooLd9NQkPSFYWDmX2vt0oWMScBcObO/ys8Iqw5ONqQxuS
zDkbL6LAKcFD0vodTyNsYWMY5XusP7oeOMzWOIcFQwtRGS7QD0BRNpw8WywSaUhl
eecLkBZ0zbwMVM+6kae6l5XEFpkkc271FgT0xyYMpvJedwQIBeea4HasHnGy+Vco
D1/91gBRAZF++XkCtQTXhQccU/AgmayjrOtdnQHG1guO72dG80pYq45sBdC8JfAB
EheNA7rP1wRokBptOWgfH9qb+53QaBEfRotcWw9FOV20Y5mInymQ7kkDsAfzK9w0
6vg/9PclE685fbxwMsSngmBb7KGrdErpFgRQNJvuPuHwmxl/RViz94zGDTfX8zpW
Q0fKEZBJ1mt0t/siAVGwxvGSHDeontrqOh1oAAlJ3w9sDkYYnUuNDKN5j3atUqrS
vFDdHeC2fK4y1M/dmTdJ0ipKsQyo/zVyqiLUBtjmBKYcuKGb58ABoy9mPsegQDNP
ABm/6BZalZbQU15iCN03xYsk1xhvOTG8wdoKqbOcNdBil3E+eAKb+bhSCZ7blvG6
JQzzXpyZcOuFyZscxau9ezWS8WIBsvEK0VeITU/IiGThgLfq0zw7znA4vAeVtXbV
dP8UwlqSHZAQMwEDRKOmU/Y5d0eriuB6skZjN9PgUgIG52fUxGsqtzDphK3z3vTC
tjlLrnooGRymiOTcFScJ3i+UxTn/rSk/zxcxxfdsyH/w32VcekIXFnDJyKYcqfUI
waObKS+jz1mYlgy6KrKIlmtxggJ7Lap38l5xUj707V2eTSImYCDi+BwwoRB499jx
EmZIeQ+9s/OB4kipwvFHSsf3emTFgUWxHW5W75OWa0CUVOl2jYL9b1lFikGmUtpn
ubKUxHEZ0qi5bU6f3+bK7I4rMggbzwY5DEpqFj0AKQ7QFv6Ilm8tLbkYMSLFvBbO
icSks6TjT6wM1sY/c1B0EGShUSAgpMZZHHYVooPl4iSJGJZG65v/RPyjcEhZzqj0
tmEQjFIeSLrAhEDa2CqpHB3Pg5rKraliAokgkfmiaBJZ5t+lZvqZWOAoumI1AWq4
7EennrrCn/hrDqGdiW0jeyaPPHEbuow5jZH7PGwQtW5mujrZ5RD07jG0AVvQNNty
d2ZaZMfBcDcJ2U7hUUJuL1tb1/2d8E1cSnbTDYDFEWhFKaKXMa/RMsF7llAlYccq
CgnNgpa2S+TTAgLoACuD+0eLlOfigjeq6TWKKdiAa0i4LhjSNUsbwXANYfUpE2LT
efZaqAZODBmKoY80wvEKd4in5FwAfhsfvLQsdgh6CgwfJD6Y5bQvsSAmTB7W3N4d
82zGD3AaJos/TdFkiaUYEHreCAVIb9niJpJFel4RGmNQuC/nWg7VrJGNyPqphndo
k8g5GV5oz1MGp8MIT0lStmz+Xg8q7wWTULtAWqHkuuqOMt1Je/LM4yCIrZRWzWVg
Iim3P6MBPTn4xSbzdVid7bVHauk7pLdsZTafRg6gXNe6hAml6McuuYNKobSGj9cD
P94jEUqz+pN7wT8C+uopvrRmRo8P7iflUgy+o/nC+sDWs85bKMfKFlcnuySmMCkL
b6YcYjfGWmsqRIX2dk4/vi5vX1rWoyOdido1rZDvqls/PfchGR+IHmODURo0X6+U
yUiHCRAJ55tmBjOmaHhMYuMWv81sbluwqqR7rm/3slHkDwhNdn28nvo6jDRNRC9d
KEeyb/cewXxDKz8JzQqnwvElgF4WUdZiy8a+qFBKtvU3jN4vi9eAkBz7MUO/S4G/
SNKGCK7DaJ0OII+QoSx0eyUftcwKpo7+RWzuQINfIj3Xs6T2jEPFZ7LA6O1eqyGv
IoMGq4lkvwoTaI4VM5kbB+G4ZgeJRFWajyKoOGFHymUYUAg2bGaAHdqMpv8Oh4AV
fQGWk41OGZrYV1bhlDVrAecgy9TXW+VOhK2/hZpNX8B76asef6qG7mmlySdiYpO1
rmFW5ew7vTfPCvlwwegdFStBa3AiTJx5DCrkhZyJQCOBHVNgVYxQsdq+Y+i6yc6W
k/vc3Ky2of5YTw9YiXihB+l/LDhVnPRpVuwCRmcgHQs5VleqKFAHvIGdW8PsC4tu
e103q2IGQ3jJA+D9+OHO6mmQCtqmhTLkNSxH36DaUxCAdmyAGo1WPg8uuXGQ8WdI
UUdEeJDeNpmVrnCyhjtQbOaEDwsmNb+MXnsYFqySOBj7KBvu7OGfJkJLiN1rJhLW
XgvUIOvpbwDuyE64myleO5pHV8JsalTAJvzHf1G5AFEWx2+NZuoyHSwZ06Auf7SC
Br5mkJ8mg2+uF4xODnV59sTg9M7Ud2A1mG/46GphW3VT5Mqn4h1jntvnK0D7Uob8
G9+YY2d0T2CrDRkVnbC26gwGtJewmkNBzWZb4aM6XVHdYLlN0yx6NN7OUuUJ+Xxi
dj/ByBvPcVNLUOd4ZiztEjJquWsIZ2+IsqbMsUlX7P5O0sLnwcmfshZkTJFbXiAD
zIh3j5RWR0k2l9K7Om9KzXLIgpSqDRSMadUlrCAy7JQKY2F5M/CcqtQDjErnovvE
MJaiKzdG1tgBoMDyRMfxn1odEYgmPyaX0LLzxNZp4TRLb4qhybWsz3b/aRkU9T21
9gWQPje4IfOyZJBY+zbyi6z/ZBS+P4jIB+rDHPO+qWOpCvGnbko9QojSk7JZ3LV+
fgYpx2Or7m4uGqV5EdHQwHEP9kuolZqAlE7Z68fWRYpRMbzUbGQq9r0Kg+e5SdD2
P3kIH80QdPE0fglyvzg263ydFB9wlw3SMCL6V71WS+Z6IxSSPXlk5AHUCtHnD9bc
QYt55cMBdtRnvTOWYyUtFbKhG+DCOKYzBlImpcj1vHP8IsX4U5MR/ASzChEcmdkF
tZqOOrn1IlBPYlVKBqo2johiIuVcr2B/xVpBjlqliGkUGGNIyljjMfEXOaYrP3gT
3VbgMJNFuk0uXjH0CyKVTN7S/BNjYN4n7frAvlScH/6fbFtJBd+PHa8CxoghE2Fs
Yb1/APCgBMGnadoDhayHHHYcBt5Cv0hFpJ3Nr/6LgZ+5rHaMCNSehNbNJiadh2n1
sZI4wOn60qSq2nimhWUAdgclmyk0TUZb+vDWHwl96SINYqB8++DxsGtTUA5ajXqv
8XyoyyAY6nSZNHNuxpTDDCs84VlkO107BQt2BfAWFFrN58aqVD7RPnVr2QEdFMGq
omwbvcv3FzijmtxapQ3WgmUlKrYuhdTjHbyv+RWqM7eAxntmTyTBu5edcMqb/pki
1hpd/n2r0HWH6MeaQeEuXOL9+rkGXxJiZTza6+MbJ3CBUPiV5vsQi1ERqNLBhbyf
j/XYQAXXcS5OJ5gZhkQcowEOJxXrAyHcpvjgr2FUCwP1Ec3BOC4pBUb8FPfgsPZb
XtdncYVEVVfkRSEiddh8XuiSPvFgiqmAmd6ml1+ImUAzCyUs44ss9PXbcgTUA6Zy
kra895Vx8IvkiXUn1W2NN28QKeBiDR8vbzBIQQKKiMovlqBlJdRAPFPh795aKRHJ
0e0MY31j6Cw67Gr3FUkQ6NhhWoiXitsRfRyYGSNOZbBWBAaomnTkw9HusFgnYYRd
4PZiJVvoRZWJVlXM33HMGYw+JiwVJKVRrFeRgJfkTmXy0XlfWpHmh3nnDOYoTx92
uxwMLkE9wxCEFP4opxjsVFEUDHwvVoYj+RYqIvTJpZujUVT56nIXzVk9+MR+TINg
obm+Fo0dZogVnEz4XHDEa/FnttaE7eF+fjQavBh75xEDSKhEeoV39hvBH3s2LRdn
D4tR7+n1xZwlIQ37KvDtWXs3tKS72zZy1mP3zI+Zc43QG18KNBSf6Cq0g8/3DAYY
bEHii19hosOp3dVkRvxPhpxdTB1dfDBLs14bFF4xroDlGMW0UPan45H8xVFvxOBR
8WWLxXev34uA4Kr/dgukpN/N3Xx8NDxrC3pZ9ivUP7Xlp0My3/5UDh3ypGhJbPCD
Rg/qO2/dtep2d6IGNKAQRcKmJFogi3HbrF2GC3dwzfXBpYYVkJkJMaDo8IZRqxBU
tEWmVVYgoE5Af60coBJ38CXyYh82rWZyu7Hw9bgDxGToC94gO3YlB8ZTXVchyLtK
Jtq3zUrmSejw6dLNlqsVbvHvBGAXmN8Xl81W3x+k2hujZHNyaIlvJC/GPrw+lo7d
W5yQzGHX21e9cUuJkgXYnkwmiwTM9oEkp7gkJoWfGepUQM+Bw/9Oem6u/GuLjCKl
4N7qID3qdi3HavjRGros2p/FpeLKfe/Tu7MlsAPtJBRCvD5LNNt6gH24aP+s83AK
+CuaGcYVYi3aF4t9ILgd10DX06PwV3t0L63IO9dHWnk6XG6W3CiTofrRos7c3m88
s1PLKRTxXBqBBtJ0odw/lGG6In5RrxiJZ3SWAyMfxfh6ASaNHYo8+f4O5OhQtQUl
2TpFWtYqCMzp4Eu73f2rb/MWS+YfMRsdjg6Co3QoqI9pA3bNkuokUuE0KzcpkOP0
5SQu8SGs2NQLeuxpQnL/C3NgtNp/xGBOIf4rFHPfIWDE2u3+isi9XU4M7J0WJWPp
s8H/LJZgVyU+a7u1ahun7Pjq7JfvzWDyeDALKnCe17LJmd8EiOhmS+TEy6fFFoJu
gNRM6OOMWSLx131V1eAsv+Vj17DdgjTtBHH6eyfKVo9QgKN1EN2SlgAKvROPvTHI
GhZ2NvKp6b5+bRUHVgyhF+SLSZ1hMtZBoR9w2Rmy1eZpAk1GfvkkTsJ7+vCLNyW8
xk+ESwhsA1w8+C+ZpUczykka7uxdb1/u94NHvSdqVtLGLeWNAB7PmrZ+3XYx8FpD
wcVbodABAxKlSL+dK3cN0pbA30AWBlPbrstbfb1JRYi7fP2IaDE+G9JNT2CLkxVU
3nVxIKbD1JmhG09uQ9MNI/y6CHX9pDN0crkHpL1P/a9qCGdlIYKhO5mQ8d30Y3nh
fX2UGMgQOXLhD49B6UwLEpuhfqXAFuviVyg3OTV3Nfls6Ed9KPUGeKnj/ibsgU3Z
B+n32vNOpjQF41GS6dl3EkBh18oPYO4hVktyq6AYMXIJ1fdh6vaSWhRjLA7phSIV
5XPml30OS5YiFVfc5Ul7kD5sfP/y1sTFFcdnuu1ETENHOF8kzH0iTRZJWPuVptCB
GP/J3A3aOQsHINyctEiVbyOUQ7D3i7M7kj62pLtOu6JdTVOJ6JQbJ/a64/OyeXoW
L6IgNC6H8YV4WEj0AI2P1P/X7n/JhzjZJsH0z3Xdn+7LB/N38E/7aUznuznMcHKC
FhQ5wH9E0YHIkmmaKL85/DeLen74eLWdKyxA/vSPev0w6Z8kdI+Sd/eQ3m2PAlos
UsEFk9e/4fB+lvs5GLTrc4qQRSGfZH5YdXusZ6OwII1srphpp7VkqFq5bn0REEFX
GNk88nocTAHR2pF2XXO05FEyMAjvFD7LEyotjxjUlgs7ZxgRwT36kyeBS9fG6ew7
hu96fhuIfeKrO3BYg/HicxdgKO34ilTfggSB5DQP1+6+UamVQBrW6wRpGTXehAIo
Pt2MptnI9cV4VwvdD6frqZm6jMRkQhZ63m6LXdBR9uOpIGYe/ofwMnxjmk53CXE3
pOm+bZ7afQPq6S+ttg3zgI0DjoYwSPQrmH1/ahY31OvOb/U8MI1mh6WAu4DWYLpK
b7PXUxZBqRD108cHEH5orppqboZjfDOQ5GuhP9Oeyzge4839weqjYqTfJ0YvPThv
bAGSLQDav7iBbmjSxNxZxBEMxdurX+rlVgJW9vKaX3u962dXuDQVKQmu3mAWnoHP
nuTHK+SfgVygF9i4oGRw7tQ6PTHpu/I/5xp8fn3auGsgJ0r9CnidK0MSlKqgYBYJ
2l5u3VlEhL5jDhHvzRnW5JsqToYJ9+Tzdqs1HKgJSu4yCCF/YUQ19e2FZjp/awsv
4qmt/b5dZBxHszQ4JXTmpEiTpunsiBZTLE2pZZOK7og7E8rKsrJWVS+jyS45Ruet
sNmObIuji1r02D6nDJvgRCRtytgs4WwVrszdeC2H+FGkTr/2TltkqiEW0ayy+H+/
XopS2p2te9/Xsy4FvwfjeLIsD6+O/Lu52ahtlPtzOJG10LGqAATY67mxX2ibQZEp
vBXp+eG+pPIBVrz19OkWmsTGPHiIl4sihAx15+fM+HDdPvBtzL1oKOF3JauYgA/w
LsSM1l9FKCallOdDwOqdiDNXyy4iyyI/OtZvSz37+NmaPCzu+ek7Alsp1RiBjL8P
Fz56697a4bb7kLfzurUgMOxQxqywRyiVfL/p6ls0694yOCs+2w2csDvSEujIpHcj
ULFftqxnVreDanOyWv8jgLHUiftRbnJJKeVOjviBGGiFOgm0Z6NjV445LSFkTtjT
Igrud+BXSz0FpzyDJNR7zmIXx44PyJU99jlt7NEBt607xBZ37xao4Iat7biI4dZX
VW90yV0Csi8hvJEMmxsmp3qjIawHK6eN/jKl9kR/S48zovO5b3kKJYyna8RETxyr
gp92nKcjJYxzy93X816byIK5PeQmOW/svCwJbmApcnlr1FOSuRwikhNXYOtMcyv0
eGkJl5sbVkeyYxHCUGLP8TypkfKTmD8WD03dXmlcIyYbgvSpbS6lV3hyCtMZuBmT
9K5EbQC0wZe0vwCD+8/JiXHffSMm7A34oh/mV/+bNzuFAmZ+p7e9OR5xNs2+rih5
VbZ7SQ2roofYTvTAYkt1PPIkwZyWpIFiYchy+lfp25cFPTGwjot1T1BHp/+UTvW6
XZuTJddEaYKjY+RDRrlwzBCnlOn/0UbTRAqFTuApMSnB+tdJB3fmBxlbFQNk/6YX
XPFEvn2QqdR5CFfZa/Hq0wCgJOwRwMnKTHQ/KD2XUE3f+FW3w6ny7ERckjTXO6C0
wGdi7xrJGrc8io+50FUTUHWfiVfzluMYiSd6U8tHBFn3261CF7XF09KwDTeShsoj
81Z0Y57bNmThdqQRWPu3J06d05ROsX7RBYbrUCWeJaSE00tCZNxR6pOry+jJJr9f
jOro/+khbXsh1k7y6DbyTjWgKAZ7xdPoGPTOuzs7E1WS0JaUD80uPf730oGHmxC7
HHaAfHz+GxY5MU9IiXfy0CAw6/PgBxfJ6ApCfo/fPWI+byNLWM9akIn95WPCmxmy
8vufMR1d86ok79aRAxIFCvReYD5RYiTexucrXcluC3k7c8WJ36FzRIK2IrtKdYFi
0msYUlJCJFRAnuIh+thELE5Pg29c9JtcewbYOzOplkSIql6kT88UKDgXqIsG8rMK
q8jnRXhYLG4jz7fd0JG/lO+KsjKeVpc41cID6Lg5YmSUuw9eiJ/BD5zyDDZ1LSK8
Txs+liq60z7eF0BdEkpGuj/ZQN9nJdgqJL86IZfL0xLq5/piMYwS1gr/e0A+Aq1F
gmlPaaSlRS03BbbXEsSLvp+wI3pkVj1enkbUr0BHP7zd4bYzwG0nr/zTgC9wlUhh
rmCPPCZIw/glLBOqKJH4q5YK7E6M5XLv7S27nQ+hMZS5allg7bv/0bEXR0nVKCgT
eF8/xFMr9zeeNNrYbXjn9uAJoHufAtPSfvGbs8EWMGbx2znQQXDAOMh+XCCXp6dk
d7gP+fWpP499z15nIueLHMDhUtxx4+YsvkbCQp9UDZAttepKMc2Orb47SNXO5hip
wzFLwqBf+pCCJw06wqXVuPEXgLK/LIucFBh/4skf/9fFt7CLDSAnuWnaOR/K0XVi
CmAVljD2rhO/MeinYx1jfWD5isMZslXn1lF6ySK56rh6hVWgNmoqBrsDeFKhKqP0
QN0zY6abrM68g32yygoFe7SqVKnGaFDWth+LTEdsrp5JRJcArlmWMToKF8FfMNMw
lkXihGsyn4kyDCscPlveHG6vmnTezNcwDAUPj+sz3j8DVWN6UaS28eUaiSgi9p7e
YiaAdFPkBC3qb96J2kWTfq1M/xdDkUoTqGxps8VFVdfKSYtU1dmmJmpWnTDVNlCE
+MyF+082D82fFZOP6kIL3cGhRJfPbE+Bz1TN2KJc5eXDrAL4qBeJiUFJg9PAfdHf
jwz6Mml0ctH8e3a4fviv7VOVr7PSn7r88aJ7qmZ5ynxfAwcZWLykHVCheLKm6YWO
T5nfwMCKaYfOedgg53GlX/sXp3gsPKEQSCWX1fZIN/wY+HtrAV/AOchQuKY+ZMX0
CAR2LH4ghyhqUk4jTW2OleqWL6cw7JCeRA8/l41NX0XOREcQmFAn1EvT66PcqiJq
5CvVWCJI71uQ/Himc4GpqWxWNpk2RDqPdBPTfDCnhFnpFY8vxjjXvONOrN1IBMGY
zxwoNqzSE+jXlc7egDifxtaa2o7kkCsRHduZFZjfcSb5NuZ6MLBfNIfL/XXP2eQ9
atYIF2NyWOlQgxAnl5bUJkdcMBfeFqF9N6E4i9s/fyGaEff/xL2quEHfgClnWdDC
b84SzpyTpFdSul4MJbhVYFCJJqpeBA6WBWwXRrV86xsum2y8tbw77td+z8p1ZbJi
ljhklKFXskLoKu0AJnqJNmhFYSdv08cN8ozRB4XCCA75E396lLm7aUPLiLFqdgak
TmVTBl/qYOU3QuKmAho9iqcCyJaf1s22Y8sRiOzYKuascKzvrMxXlxbzE074Ahbw
ElzruvZL4YU8/7eCTTj0JnSnqZ/9NgYiVwuyzYNWtc0QchSMAUTqcHPxtTPnq1UB
vLrttZemcjaqKfVWVWK8VWYTRh+RE/oYhVT/NTZJRc4qYZOMwCWxwm160MHOUpcz
SL4h9uf3onIt1Uw/r1zdYuef5pxCCP7GWYYblDI59cLFP6rtGCMKu0GQzXxvNahB
clsEDhOR5hYv1X7j+yvD+aqJpxW17W9gQtPJ3cNLfQd6FznetnpnRvNn3Ws4evOw
NAqSpVg7VRwSZ5Pc4T81ygroLYSU0tHaNTGAWzNZxqqT+RUN4s6toM/bENZ2MH9u
GWCzkSIL3VRUDvSynEmFWDPtsUYnms4KWppUw1nc6nyherar+ofDF15uNID+OEmR
znfAl9kUtMLrFP2FJMJuZ7dnyrKgn/YU0NzlYPkknvBser4fx5np7kAiTQAlgUXS
QPSFXkGrC/miBPD4Iv5qgRmSclx/UYpagiHj6E0UGKTJFtDJq6Bu99cxmPatM1nb
fl+dqQdXsQpcGZL1+UpA6yCwUSysyyMK2yvd7mn40ZXYEixv6TwUsViNjo2E3gqv
odI02ppIVenoaw5h1RY9g4tHH4TKsEiOISExX4Om11JiE3ZTmaTYZW6JnrT6mnRr
gwKGyJu4FUHJU5q9w1HoicnVHl/Phg0tJNRuoA4UliIQ/LbL9qKurWsMxgZBKvhg
2kRA7bx/C+wiWfVclmVy3lPAWBjkomlg7HNkZPQIiWRtBTLim0L+qqSkvSiqYAOk
HdD/n9w8uXUCbwmqXeCvCCDfDxUk3ppgthBpt8OvAAEzNN6A4BhzwCt7tBMgkIp2
rklIk/QhclqclpPIN5QYu9QQ50qcVsyH5AR0EmoVJ7aXUO1rASNB4haMeB7pJ88R
RXhYpZpL8XzoTPfIMPGNYS4RGQ5Avb/OojKJ14SD8pvrqykbtjfRmU4xGv1fYGsK
3/yDdSu2iEL27Pqy0OxCjwZo2mGY3AVmXN2vWP9ttSKq34eYWIntm0TCC2eFaCiH
9BF2IvFO2UaoK/oU0PB8gKi90+ue6/qVkulVCdsDNparwnvThCAY6BRPEDvtbZHH
n9IIbLaJDH0B0OK9UEWVtATq5mVne+zYQ5Dzjj5Y5VCuvapvBUzNcIHnfZmcu4Zm
sM+NySGZKElmXAY3KMni466cUwVnXn7Umqary4+FUM6NadjRWFB5stWAMXmnBChB
wM3kEqlWFeaAE81arfgIXdMlxbc3/xBz6GjPaRZZubewDPnsKCxDGgmPpfBDsjnR
psNDMs1kwY/R1bPPMiSv2Phc6FnBpbJLRuZkkwfTgMHnUsxY6eY69e0wqn5gsN/O
goKzqt/3f6LsvqsYl/k8DAbwz1Yfriohilcy6M9HzGRCPRAbrTD6WyKML4OSvGAx
JSu5f2xzby+MKD9uFRX2JB8iFQ84EsMqEzFZQTWMaQhaF3OH62Y0Gsa7B3TvaRLn
Nv5QWl2z+Q6Sqh1pZjKDa9RFmK6nJArGup++nVqAFdEb9lzoT5SIRFKE+XZZTbQv
HWVI8+G1BtNohPP9QFjg/GTRsehZ8HHTkdaEfgwCdeYxEAm7hmsjCrjuWR8TzKls
K8vgLm97vtbXUtMb+yxHJqt1l/3euWQhWR/aMyfwLzbr+b4WITlwRF0JoClHj+jv
GzKvEL8eERyca4WSBAdoDItZnAQEWx5mUPCwemx9hP/uf7VPyCu0milBmA5XSwPV
Y6r3rzkcFnWqYEiK/iAP3MQcdg4tJ9H1Sv2xvvtDyhMR0uIeDcIIWz+AtZkKyoVE
kbOm86U5IxC6IJ7rsgyZjLXQPVWleyRO7j0SpvFHBpJ5QnG/jIffSvq0Evcq6VXX
X45elKyM+cWnhLQabRyRFk8GehMOwNjcTvJt1Zkp4OGzJYm+A5Am0WA8VZ1XtQf9
mzu1uTKuSmrO4CQSitAimZ0SIquQ+Ot3rsmTCl0e7wksNuswqQX7kUUYHeBuT0F3
6lG3+Ptubq9X2Sw2r8bsz4PmzeBG1VKayZa8SrTiGtBvlV+JY5fnPLrFbV1Qg8W7
FKGFBC72VFCBD/dm50tN21Ww+8qCAHpDNSYF6FW9eHXn9m0U9fVDHKPtnH+mTSaH
QPQ8WuTj/ved26VEAjf1+T0yYZcsaXsv6dtCnZ6HU/TBk/9SykOCSdpMPH/vKcV+
s0ZrAAKofvpmddtXuO7fEGfHYv6R4W+4KJa4bKFC016Bl3nDxVMTvzQ5vNt104k0
XieVkbcfAl5M06FSmeGKElrHX4Jrh64tzcjJg01EsbeHojJv5MxoZkH3i5FOLXZE
yeeQjgEVmJObN2qxJClkEl4glKEqu5NoxPS8Slmchykyg+xVCki2gOdhwIaB9ZVg
rj8QVOWifEKGxEbKy1FwueajpHF3KrQje4XQAmfditiBazm26UrkCXYow6Fzhsay
0COHuRbxFv8fZLhI7Ll/hr854zrsF/UIYZfKctKRqqGsjONE6fybLUSSJSqm8K+O
1OmXGsHYEuHlaNgeTKbjXBaXYjUi+BaGkfNF7P1b+oq6cr/Am+s6pneotgrjxqdL
el6GU/fLasMRFsYq2+j4B2T2U0uyfud/sISwWs5/CQCJNvePOqq+xFOXtsuVVn1K
pTGCAc/vzbzFchAo/qjQ3Od7Cm59eKWH1RkkCt5rfa/I+MxW/n484fRJ4E+iAOdR
aGM16zkC/c6XBWGs9E5BuobaNB8THFAyVxDYJ8/7g8fdDJw0Lf1e5DSauM7NcqNB
+31XSgKzXLz1Hv2oiEkF8e3YJTJz9DmJwwxRd4i1pSptXgKPtoVd7BsPzL1K0ch5
YA41BM5jXWZz5ZDDl7Fxre9PH7bgpJW473EXtVEZCa89BL7LKGTSxYsdIOdY9RpE
mzoEJ5MqJk0eQ8L/EpkiO9MMJNg7zDUa7RkFX/VVG53U+CdMJX2TD+6ITahnNUHn
YqONZ02sHYeuc496TUIEjQcLp6E/MTE0qI0Xq0pbhHbXAafOCin7OffPnYAVNcsd
JvvMdzfZw4uEi8+TnxfUcb8hlSLtIoe3KmGzrzYcsf0uUeZJSVUw8g9lk6l+YLLU
K5eOQ4Rmy0b5oKxWn1aQJfWdbMWoABHbOfDeEFBUHW9cXGOAgPv0C9bJZouVWuP8
O/JlaDeP+JsiOoqrniGuN2ho5o3ZvOQ/ib0RtUy9AmWejrfgHP6lno7H3nurpcnz
EhKuL+DWXHfZSZVlVyJAAE8QON0TlqewoLmGENXpdOykvxeokJcFT7fC601oEDh9
x5POvo4QXL46k4btMQ5C6lw6ouC4HrVpwGvlGz/S9xO/BdPkdzhW4oBdRsMW+YsI
KhMoghdTpV1RnLJIaZbm3Y3Zln9meVTLxvK8lOyGsUEFQmDq0nWWoi3FLc6ieGDW
d0zUKt7fqVGhWfoHBOfpSrL5mm9TuQV8iJAUBcX2H+LXTKrlUACn04iltwtXLPEW
zVXvCXATg9vED0wTFNC54ocWj1thJLOUw1YHEe7VtGX5lguPpADobdhfmvILh/fe
RlU2Xu1VrwJRZPj5edyrfotYzgGkNFUle3tHDXFBgyMbsh1NHZifLEh39blPeuBm
HTvKA7LNwdXzOrisMXqHrgP3nNgxzuKRbeBa7XCGzrgQnjBq4z6ZnOKHlaVAWFwq
7G4k8ZUw1NpO14wKzsvA7i03cB8tm2EnqjlgpDgNisoRMAREnRcGGd+DoNFXMr+V
BOoQn9QUgjYfpPD3SLC10tFdj+pANI5YJazD02rKt0RSxYnDKurGf7cCYLKb5Rdd
xuLrKR9+z1J5GKOtnGqbTFWv1Mb+Y8sVlJjC9Od9Bqw2O6a1ibzQdzoIYRshqNan
90wMb0pVBGpf0uL339DZaeszjTshMbelsBEN/3+Yx0sZmkjVewndY06xGASwB292
qrlR5ScsNmBtddTeAxSh8T37al3fKljSVLIVx58glo+sU/yi5v8bkJBOxlzX8cB5
MFF4ZvY7HkXbxh+Uxgvpt2+4vKiNL5qR0R75XqiR9g5bOcKbPSxrgis7W/FbXaoF
h04bJusI9PJ9lhb9+UZUkYdSitrgCAIpFm2mrCXfOqfM6vcdRPxM6inVKXtBXsX8
ncdBco9UbAIJDVMUrZ/CcFeEdOy/OwsLngwHgon0k8le/IObBZcJNAgemicCzHTu
sH59CQT9mA9t9x+9/P0dbsOXhPF+MMRZROvBRIdFF7W1C9bMYx9BdM6H8r5LFnES
nPEVOZK5flHj7ymx4BGaqKKuf2Y2F142Kj/y2BUfVjwDei1BnXQLqvSU0ejTIFFr
k/VOpF4JxjTBsUiVOTXm29/dLKuWQ0+FkVQHXzzs6w7Z0jhG2kLYk3K3dM9PFE39
eBH09AonYhq1gbHtUNak3pDY7HoiO8yCFTFLMoh49zW+IAw/DccsvYE68TYdaEHD
s8rB4zfcA8eckZe8lm5981earZ6sYsflYUz54el377uyhIr/JtL0ex9ZFDFdhWG5
SsPuGO7DP4NTUedXHQsZMOga97DtMyZEO+snNHy2go8zGPQTqKWJD3jnFkYh6I8T
K7YZxE2ywhXmQ5ve89r3WZbm5i/1QBoSkLFrD7K3zFOU3MCtSxi9fnucwjRRdu62
0KDp2tuSU5IIICeQhXUZnB2oCWi1et4kUv01cvvi+b9O/r1MDi7GBwGDsI2anO6B
QXox8SxgDdneJg05Awzi+UND8h7lz+MdVfCHPdFI2SH0zkfELlm19eiOtvtaAMId
thTjJNhlZn8/1QmP9XzebDaPmcegZBxTv8ZdAmirwAFqfNMZaQCZZ1srXXS9KtJZ
n3MzlIhlAdJtJggtZhIk186uiDEeY+BNJ4xyKwaoX3p/tG4WxlJiwHuMRLjfhub1
u9ZhaX5los/3IPW+HHyoM5pgK8OZ8KDMLKWYi20M1UMERRkDelIIJOd/7y3GtfTn
Zed50el9+iV+vkd6QtwHPWSGxOs6UY23R2Jjo9yLWPPPpKooLBYhJMLUprCfHsef
/G32aQdUWG3d8sExMW772LPRTacgFg4x46TlrZSDbmYfAoc7dgiErPmT8npbyvA3
6LTvKegHJ7pyozriz2yVvU/AXvA3S4BtV6UInsLFfFN5bMQUDnSPrAd72g7Dq0W4
PrsIf+mTlgrEOAslJq+wCQkc9lePyM7fQTs7D4c9hVt8yYiqZAP+juuX4ucywROe
z8O28nmmFsN7DoWvuWzLOrz5RepN3GYmQUxnd/R+GKk2gbpMpjdWTFPdD05YxCkm
DKm6LXaFC7W34i8y18h/oaHAitM0mks1gNA+f8pdYaflXzDcyFFiRLZRtlVsqpS+
uXK5aANdJM51Z3uTpvaqOm1VvyjT7SwgWqV+lcp6Dc++v0dRmCk9OQnTqjgsRRQH
Lu5wxXsjUcEtcRpOCqb56fcRKBl0mtG1/wLaSuZMJxjGM1S2j6NalMPKTGETxmbh
jD23d80hU7mtZoAU2fg0gXOuu2euH3REUDmnqZdhHRG10MWR90YbZvaauP07zcDW
WhdPpWV3sFqDScRGiHUnaQ1feiUWp0WdLhqLZ/pOdLDpa8wrHkWRoCifAyoUZEzZ
jx06rCuzBdR2qcB/TmLA/vY65elyOjRTH2k5b28fSTFaqYncfu9QcARiP+Bi7qjQ
6qJYiALmbEVAF0QCLlfxRcTKQFDfzx7txCfz6Ygb13wSlte3dO2SypYkg/2aGdiS
Ej/N+bGOtlFHHd4h7aUHq9+584c8vR38jXTrqNghLVk8iZRzPVNo+n5usfROmVW/
TJs2xNm57VeKtvdTL/2t0m6EqbAj3igph/M2y9mxG09LJp0D0UIuU/xylnEejm4v
eGt7nXHjJplisBhJR5+4FsK6TNwnbdrfzzsQ1Mnysqnh0J2JZp426N1chUDtNDRV
sZ2ky+s2HThBAST6OvJGQ93limot3Rte9id5VN+Hbvk+PuGLAN24mcJ+Gbs8P1Z6
miuidi1RfAt54qLjXzgNyTfVTlIrhQTm2+p2MCkxj0OuV0fzMWGvUQn5NTy8kW3R
XB7eKS22Bxlwws5++VYjvszdqDneOZSpvqldT8ZZOG32fW9k32KYEIhahSrB75+/
VNwnIP8GeMEE9/dR4Ewf+/tAiQT28XzLIDB3Cv0diNqYDeCLNFu+JBIkNeFyQV2n
O/zqr59nYfe7eg0FN64PeA==
`pragma protect end_protected
