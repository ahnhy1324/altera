// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WLfX58ZNm20ujJPqltCdChYixxMR0MbzORVeLA20fvnMr2n61KBPw3MbTGlILImb
RRJ5So6rxZPVr4r2f6BMJM/c9NQ7roQV7RKznGdxwPSps8OIwwEfVQkWPRcOwjui
J9ZMB0Sl7guly1B1m0at92GybxW0qpSXaxUTL+dHRRY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 62912)
LI0KjEDAePLRC3BHtDrtrMX7+rxt826OYGhKzc5Zobl9qK8XlWR56Px/HBXbZJT3
Td9MqVzAxPo++b+xBgWSrruGNiqFko89cGhRCCdSrs2GmIdc/hnqaKo6Mz656oQ7
Z07yUwzmCQHkR7fB2PBmyBr/SfseNSidgEOILvUqc2i1ly8SjBoBXF1amGor8YMY
unAEf9TL9CM1rJgJcL46neHncwJ4CL81Vl4wLC9Sq+y1WrBTx2TX/izMRbGrtn/E
twJOtZBQX/z3svIT4vZD5/6Biu0Laucv/niI8aiblodhRtksy8SB1UqSDXLHNKjQ
WcHQ0DKOLjpRjssCDpqJk7gDwmOGQypNZ9uRhcbJk2mokIQqiTA0p87+oRM3OGlb
sydZInGv+Nth3wXU7oV9lm8bRnQGotIlI7Gb0Hx7DJlDRGBGMLv3Kb3FLHSy7fxY
a5kx50ONHOlWd3X0pJtGmcejj3LfgyDii+2rxkmyBhnsSxCCSF4vhNwcYu4U9G0g
e+YGYf6DpSb6McldgK2UFP4VLB81mzkx0ybjc6pxxvpeYQV5DoJrTZ9w1m1xm6Kc
rDpZTYEokvo+3FJW0eFmfpx0VYFbgGEW8Y+jo62Ze2VyVRZ/6i3KO4hNCJXdj53J
7ESCYa+4vcdBENlbgUaC92jqO+zZKzxI3tRfL8CmaNitlXuPEj8SZHnwMKnyK7qc
n1/5PjaRH1zkVtKzdCx5LA9SsPz22+XdA9PgX0XyS8ok62YAUKffb9V8tWP0P2yS
ZJiK92Q0k/hCzLO69eZXtNRrxElj0jWTQ3IbpdJN5PskVNj6zHF+T2fNYx4gYFQj
xwovgwsdB1gfjzRvI20Wl/H14fv2WuwIlkmrzprIUb+36cthOCFxlUcWyI88otHs
q8ixrW+2MeRlPIzHAOLnQo0MW/16vXkMGQ6i0WtXnERjOt+KSyWjZD+zBpeRvbti
5Fyjnf2AlkMcCukPAaxC3HHZDH43ghaIjIGdZNpXxslkgUb0vAt+1W/R9wx1UDXx
BJ/gVZiircdAwDxhL/HPTKk6BkMf3xnY8245RRtbylnUqtToSrtazTRocEeqHUEE
yCf3HJlVdqUXlXM7h3w8sV0EQx6As9n4/4nDKf1GEVnMmGRRPLPDqdaFkj+jTGIo
KswAb8hPkxvw+UOSEQLdwhLp7TK1Et4m3INSSXYddujPqqnoreJacQykmYjJ4j23
HdkL4xZUq6vQnoQDI9dGYIMk0lmRH2eOGL/xI8T7N2zNIMysYpXTK3TLGFsAH9a0
mV+F5BcyQhrzvh/stP/p31T7FGphC60sJMtUubnV3JJauD7t/QR23b7oGxkvhueD
/YFplNG3w9mEOCoF6n6bLex2BP2EQVY9m/+Hc8TmfSE8TxCSfCA+aBRsf9OKDsQm
N9Iv40i3S9qVMWo6RM+gZ3IpHGlxsZIRG6tGyqORGywKtc+8DMwkrlYqAdAamSnF
awSMH94ZhrDTmTcoTi9Yk+WbaFwXFa8iJsrFJXj1WVbrUIAHnJW0zntDah5O6UqK
AjmCJkJvTuK8op9psD3EV/MXvtFUF3d09fnJ96CO/ixAovnqFLPeuVY/XuDf6LKU
TJIHQu/0ymRm3RY7jDQ/ioAF7EKC/2XDLfb8Rovzipc5fo0sXu+7SXF9WXR0cHD3
y3DEIc80cSJYAWySO1irDJx/suMmVPOfUDZn2VfjcCAh+3RExtMkr4OGQeK8Phav
dXBDPHs441tICZaWDQH1BuJiDmp/CEZorj0f92BAV1oNuyel1bXGXa5MtCC7Cx+A
axKAsv3xO0in4yGX1TD1WnLsOvSs/YJmmDhPM9npZggGrWrNJgldulnYeaBfCiEb
820dKiuzvXb/6ogNey0gjcbFQcTCZrbdHqhU6aSdBvJkOQqxGdVEh1PNqkmGajUS
bTcsP7yEAWnsevgjcLVvTSdyUUhvmgBHSVcJim4Lqh/zFGmyLwcyc9REQBgXhTmb
XFGrREoRzEps0AxY3IDeFrZaFDZHr7TzOAUaSdWIcqJai4Dl5hyQXiKFdPfPgR7h
fiRQdla2ZSOYCNTJVpZfdkuHLWIagzdH74yk4jO+T7iCbTcCsMBYCU/3GO+3r7vZ
0R3DXpUGueNtakdpXRx1xhTwI3u6iZqZr549hAeW8iORsHNHZNFv8vOsT6feNK+c
sYjJXpHf6Fx/sFHqMWtTpJg70wXT7pNVgYkUfOoDOWx/PG6od1a449j87NnxaeZk
//uc+u4J+4BJ0JqlzJk9ecF0FGvlBU3yYtgWYZJKe3nfxWcxZBn6ABpBO57XvXC4
/pmUfbgiLyc2EmoFkaeL8kxUXkqXLt+6sTRddYZ85mm3rhhKGfxhBL1wp+A4JelK
eDzs7G0od5hyLGfPWZoL1SGP3KupSLtdQ1oJJGI6a2Vzw//VfwYZjorPx2lsj5wZ
q/RhkP/AHvshEkgCxc5hM9tTVdA6TD9CG0aMTWQuVcSw+O+I+/IUCUBRlgXJjG3g
wskQ3KZ6wuMTweGKN6nniwKsUJeQEge1TKo+qU4kFg4VtLqtm2sF898giDEG7C0u
kMe+klABHVvxRb2QnGnVHDwiFLwtiNKo69Zagg1LxTIhFXK1Xf0MgrLxTHgasAIU
0tb64/Gzhzas/F60wg9d50convqOGO6TfVZxhefLcTcih8jkQ8LH+9PqYOtns5wc
9adkqyUp3INidRxGvIT7UXJMxWbDEcyUHanRAg+gZ5HVFAajg3DDdfFfofVgLPo6
0hx2lPmVMp/PPpBAFhSVpXVxiFwFCWEUrmdYEEgKK1FI63pR2UK/sjtAHTU914Lb
ZMtYo/2ffMguHqtvtCP3rMb7jBGs3119rt+rweki7UnJlhXVwKQS8iRMo7c75BHd
Cmc6QsU6NyiXezpCaR8gxZ0slQP8sj7J86BJp2NlHJVsJPqaqvwtNZTVVQa/b9fZ
2HLFgZZVMymHYf4IGuLHmTSB+GaJjC98XH95/sVYGtrPrk3qyg4SCkTRrqhFk0nw
lzpmt3TPUAx6MeMeG7aLbRovGhIcTP4SVj6aCJAAylBZoIPE/78BoGvTQUIuTcA0
8FD9bxBIu+g2C1CzXbTTp66G6BcHqsbMEo6vuvWDQkd61HHOKyyqTfeqFljkWI9j
aGa3FVt8MH37wZ4WFMYr2hJL/NAzt0P1v3aXvf1F/OUxRiQDkOm7ByuKzDpNbJHB
ZHmTGG+fGuHzjjk7k2gHid/asOY6yB2FxkNTqu+U8QUQ6oKPCPIk+ZkDBiZZQZ3Q
Ltrjz+SPSP5PQ6fWjHWbkw+8ALs+XuVvlZclawh9TlfQqQugyWHjr6tyVJgjl29c
C47CL+Hx51KEPl3FOugfMP7FbeUKjdJUB75cRJx8om5PvNPfT3ttkEnnIgtLBNw3
mULCHika3mFXvc3dnSnghiGA8/n1VdAiKR3rKIDBkgfWtcLw3ThtgQsVLgjHLz54
xod2splRwcH9wxa6HxzAGAHgEBKuhOw90Fh1TS4MsynL5wP55wFxts65W74URVTe
zbT6RN4x4Vw77JxM2g/AQY9p0AxUykUxyghUpw3QdlEZh76fISfUdtJrWtS2sOuY
gde+Wm9ZyYgQ+VsVRVSFc3T42TBT2yki/6ZEnJNwiseqZcIZS3oL6HsnlPLHKlLh
bYNsDYbwLbFOVhGrpg7WsanZNDLRQtDXVdS0GsDzM7wTzWuBmCbDNvv8vB/Wa8vw
P7OQXT0Mx8AsUAbMsx69AQC3LsL+6S8lpIVI+OyQcER6SsdW0E82tMneNRoEBPnO
iUx7BbK15FldkdXyRAlGraL1DbZxy9ZMGZIViAaT7FKWcu7/fn2vlgXGcW+q2p8L
HdAuuiCh+8UtyeiljcjVFuRWeZWLbDTJ32lCyyvIpJBmb5PiONDQHPg9jT7oFMjm
HTPjUaBcud+c2Oy3gUso0wJQO8A3uY8cmCQ9pN7jQ8PanP8F/s1GdJiUY3geV03h
9d0H4k+QO3zr/a8SF0aj8P77ZUGnyrX9e7w5h6ABC4aeE0eIIHD5OXTkx2wZpX6U
pSiquee784DhntoYjpS0MO/YGPKaPqH0dvfki6ooPplB8WSfQpkovnC/16+dBcND
MpUlQ78uFePgESRpqeu4WfAnDrG9VupLFxgk1WHiH2cVISuWEaMXatbdQGM6jgjS
aqsJxN5l7hHhL8iZ0+h/ybfUps4Vxpdj5ZSbm/STg9JcBlpk3JSJhwoHmyUJoaSk
sYyLzaXPRkQB1Q8fNiTNvbq9X5hIJLtIwqdiu6KnoEnjnsiYXLevHoyFreuN1brW
McbuI3PXsCuPLkcEmur4YeDZWD3ZHQx3yDNULu3Ul2FcSaHQaJ49vJgPUo0VNFfh
WUuoOOeI1ZDLW2nofpwAAMabXQ4nkJJuLljkNzVDpTsdypNgtevWQo/Wq8DgruAn
ehISqZXbPfnH5QuXxXOeXV9VZJ+djACs0vEbLgrT7y/NhDYkNfg+kt3S9Pcp0CaX
xpEncHRdcWThC5EYisb0YgLvx7698s5NcNsLzx0G54VZU6VQhEh7E1r8KfDDtkYH
hMotQ2ew8+h6K7kEccUoTgNk9MPrH4Za9Z8LaUIsHzoBV7TdFTLy5H8f8qlY72fW
LMUc0R8KG7kM9xUqfNPVwtygfbY2a1aYdOQCjXXqvW4OwYylIg/+Ke8ZmVEczfKh
YT5AGJk0KkgtKzNKzSBNh/viAez+sOEA9fXne+8oa1W4BDNaF6D7ELrlr+qenv5r
IZnbVYHeriXFWxVWlgX67kHDEBEjEZaqp/JjRsFfH3ETy7jFci9rSF1DZhi3EivQ
oI8Lm2kzjTHkhD0rzeJD00PCAyMbNiRA0OUpVFOnF95vWtPpYwDyyObwoyLrsO+m
SiZDot4EPvNRilo+QlRD24xWap5le47XjuzuY4bVznTVvi3YmJuJU/Oh5gav2rUG
R8gmTWh641gFK+uZIRt4PmBwSFnD3ljnqSrgjZwqpjbrIRNemE87NukdcyrIFsYv
lQ9qlOzqCVNuuTlwlJY7PpgrRQobLdcW/n8Pb6qWU9XzplQ8fw9+soKaJSuS1hwc
Zkslyz1Ux7mrQHHQ7r56PiLw68QpaZP29qXspaLxhjUgd47XATGg2vXqG5+ldWGb
aGZ5tATZiZq4uh1yHcxYxwwBOIsBkqNdSV3cEX/BVgzlm+LbyJvRljznsqUIfZgZ
kZtX0dum40jC5SfDzaVzBrc6e6ZYNvfweGLWTsgfNn8zd3m71puVmGWUHAGHpwIW
lJQoD2WxLleLh181+SMQkHMZA4J1b2SdQnaMVZK7x5pd0wYrWO/taZM2vh+MCodl
AhUYrAkDX/qFUMkVLmUqAPjykPZIs3tITHEylO9q20rOdr2g+ESQwOogZFYYexqP
7alCh8GCVjTA24sw4IPINNKAkBAU5tJiMjnZ7+As/oIR9B8tdeqHW1P++4AsIXCp
KUgZUMD8yU8ESRvcV2mb60WV2Xwg0xfDtTmzNHgVha5m5v/49N+H0yj9+I8tvpxy
yzBXk7/OB1A/oesuZODXfHrM5EMZpT4Dmja7HWgQhP8yJ2sl3VYFr9a1auT7r7SU
tpiAAi1CXgtglUf39WQIksg+GQcQLQy4lyAucQL1PiugpbYVRzDDVbHkTPK+Fmiu
2GWVk3QqRaNaeSkhnBCKAXE7B3QKe2o8pp6crT+Hf0Kyq3HNzcGbx38Cn27YGY4d
NvObTx5afSrmvPvQCEMugOyPyNWq6OyQN7P7rlm6hWIOwM2lP0ugOSt0ObKbUM7e
PRz9o1Q/AmZQIsLl3Ei6sXp89M5pFog2z+9oSCuYURPHXXoakuz5Foc95h/32USM
/wrxymaQR3+9O/lD6GBSEtMsbXmXbS4EEFX0DaB2YxV+yV6yy4pppnhskisih/XK
1C3sHEFCnHbJOs04Kvlsuw3TNfZZe5u3ANOBJtP7sNkMNBY5LBxkeFvk1l7h97Iy
Gzw0yLnuC5rJ/MjBHChiXP1A9+Q6z9dP/ZlosSBYDjlabtpKXm1i2bwzgyg3frKH
HCYVUubHlBPRhrdmc57bj0sOz3YCfZjqNq0CfgAWs6BlM2EuAnD/oh6BhDUDbFR4
QUo8yGW+F2LCKE1pIRc7g7kbdxqSwCtb58f+xAYfQ2bBzjz29jW81ZtxF9kDIbZc
+sxOOP4e9kPn4jD8AhXVr0L90NP55FfeoL3yOG+YHhJKOkpgRN8MOwDCUVM0xrns
g0DS9jllGaXfi8FST8doF8Fgjtkz2qSHUVZgrMZaynXRj0dgwx5KMIW7aDbRssBA
jLvM0J90QYmdRrGEhHC/P6xoCmjNX6D2UIxTZkIiZeMetp4NMx3aWCPVjnaXSoG0
S776LsIEnJwUJorVP/yNvovLrKgfuLFO41/2wLG7C5OVOpEnfE/W0TgNk81KuYia
0mvv90gZTeO2Jvf01iRipYbEWzCZOOlN9HQSn6N3gsSSGajpReMu3m9xAtpZP86V
Tkg70aj75ezH2DIIfdDi4u9X3B+oXW3oW0FqqdSTBj+/etfqXkJTXHMeq4v4P8wb
VtLJj1hofEQOP4HAfLEwgtZybaORx15BwWeyGli8BQp/jseRhuu2O4ohJIF9fO9J
iKBbDBBN/NahEYZAIJNaEGXvP4fDX3ktVKB/wKa/SfCdCZDNsqimvcBsL8kKh4qK
T4IJefjToPIvQQBDaynBu5qa2kXFoZwkCnjogWRaofzjivekIiujTpEhk69RChlX
RFbe4DjI9DdW9n8A4mjjFqbePmWGismN7L5ZJKR4UStQMLl1WaKguIBOmlHPlUqo
ymsWrrt+04qx33Oja6lwVLl3zj3ZYB+HKnTBzXSiQIJbfkc3qLw6Tl1hqTCodq7+
ftpKoMzXnXJMPE5+48AT091YYtGSt9OezWzgRoJzhladA8BeSaohgJXFqVdsxD8C
7UGu89fu5zdoBaNEXx2+txwUKW1prnFVNZz7Ras+ztf9MlxAoDLfmFwc/htQ0yuW
+0Nq1/tCnEb9J6ej//lrLkLdkPMNYPPv9ho41qw2G3rM1FRM19tjjKxPtlBqUEtH
tV/ZybCegz2BH8U+ds1rtZ9aFO8eebAtDiqyJvOkZ62FlGUF3vx968ZYhcfyOws9
5wqxUfFcHuRxUG+9AlmJchhGd/+Zb0b6zL8apwdQ7IZQrh9vrz4XPz5cxWvSKKD5
l/dbn0bj4BfIx3CPN61AKJoP0dYhRMcop8x/W1YXg5nksWVYiLY+fTGHfJ0LfZ0i
oS93J6bPpdAf4m90+6MmwXqAnXFdniXG7yPGoBxeSHN4zJzWBKG3nPoWla24XL3Y
XNHAHd/E81vVgsu51tjtpVegFGqzTTWIFQ1gT969Jx1ZJNSA1w7AtUQcGYMEaKwt
Lzr2mOGf/dGflLAYqGqWfpY7EP/1EEoLKCNE0NxeqCdLflZuP9lILcknufpTXwTC
g2Uk1G4NLWEGnnkvh5RNTd4KvwIegLEZ05LTSV/fXhJe4De1Z6RQGfT2904NgW0p
MvEwnOmNWB1gZvhzxMJLsM4rSnQL0EWwKxNaH9eq+2iwWh6t7h9rk6hoWuQplKWQ
CG2l+8DtGDKR2IhtqUUzAd0Ww89EtgSkWVryYkHtOsbz6473OqNO7jsNjqqCgZ9B
CL586hEP/B0zrmISkqF2Jd2iGaZwsjJGOzwMnlUlMqUiSXDzcld8p8dwB6NTGw3K
hHfQHAh7Bm8pn/JVSVIewWkG5J9ovyv1tbK3UjjhUcKkD5NBj2dLOKL/Bag8+pWZ
5RRRk7O/7MNO8hQg+lK2IY/xaTenkbBY2vOEv32IhrF+kFSiiqy9tjgFcxk2Duuc
SuVVJabxgAmmG0oy4EcTo6tJ7V6qEpOn2kg7fJOnaigaANyI5kdF5MKHh2Pqit05
OaDoTmFPd/CUF6sd90hHePTkJb+RzokZb0e64G1iUtvvn1c2+0epfEpt9WcXzdnX
qL7XcPSFKT572CS+G9p+/K6oIojXe/mu2U8rf5zEy7wfpdEUvNo5qWVTeVY8ZYDL
DUiRym/GbaC1rsL1lj7JtuYFZlw8t3GwFLSZovMyzIFSbB/pRM1bOKQ+WzsRfAjC
6zkI+NNw50qjdB7z6ZwbRkIWOExCoSEtse/xShT+//PPWD3vJzOHIDxm7HBFotwf
I/7EOJ6GJgex7AfXiJC+Q8pylzq7J0l8vNkbLvEmrqID7tNwcXxz8+2PBXh3SeOM
qxTFZBcImbQw7sNV1I65w4e1Qbv6cqt/5fJMo7QJY4NDyUbgfPVSqd3cpaSs/5vp
SCCvzVpZzn2gW9n2R2BqVrKkfRieHZy5JxBU99TWOFO/596laX9DeeS5dySe2VtU
pbXt9nEjVm7r6BmpDtimI9GbSwpX9qFUItP6WahHQkR//WjE75rpM0w8UCjKBizn
8iKY2es4lWpdkT5Bm2l/HNtkYD3HCDo0wBBsRv/gO54PG1WdAXVGP5ySAm05F8EQ
zfUDm1uLncVrTEj0pV8YryCnvL3993SqG2+/Bk7oMm6L/MIAISdOoZsc1Of9mtrt
shasDammpUcrHeyqnJ7QWQYF4q1joMCP//DtsACGWKlKbx234BEzPSFClx3jkjVJ
MARSATIuVRaCYx6il1x2zTtMSEXMBHtZNO67ZSRMKLdiFGe3QmrVvv0XyOK2mEGI
EtnZM1XURFz7ALMO286dKHPvgTdddlQ+2xBxlkTCL0k52vzpPMxAja6Z0wycQof3
vuw7SZakzLFlT3uk6VRIYwUoHJPmE7X6dQyx4NVXz33TRn6lsMgcuPNMy10P/csC
kjghuA7L8Be0W1WjqY9sSkQx+Gs6zQ2fdQe6maU4e/r1R+exLhHUUJZ5CAexnImU
H9Di6wmqpVKAO0J+HwQYn3sFbxY7J1VbIRbS5CcEoFI+bfAvjn8xrCmGJ1S1u+3Z
VifiSIhKt916esiDbtoLSvI+/GKL/NPgQFP7MUiWtyCgaL5WS+DRam1SYlIFZgEx
y12V+9BGxWZmxE51QkFEC9mX3xqgu21+w8/+cEAYVdkbkYuP+xl2PEw9uvr6sjQs
Ick8qGAGD9V3OPQH18SW33wTZdBGdg614RO36qz1jlpcRGXkNKKS+3cBvU/Qaedr
EjJgRuPKrwrgM34mjW9L4ilozaZ8cAxM7jTbCTvbiAkIEz3k46CTuDmLcdUzG9K7
DHerX9cXq2r59FuNMstP41swCikrxA+hFrxJyKm6A1m8+WTI9TOIfHCMYuvHMzLW
IoHAAfoWkR54h+BoZTc5Q5LCPjaUNxYDc/fnyIv4EOXD1gJ25LCGHTFz4cewEqHq
zGbYUezqbpeNeyyCBFCTBCYklAff9kVtL5iATj8ucxlOKq7lIgjEl67s6ieTLFTP
YmPyB0y1b0Vv9BFMS4N6+eNB86Bb7Yz3nuv5FggfRJh2CnHzHZpVH46wZ8/J5EXl
qDAuZstqMdbKkuL3qbZJ6JGpuM25j/4uD79UDdiZotsTBJV7Vf0o4yIycyZot/tv
rgLQGBwZK7SkGiC2bOa/3TtuMKwy0mb1jkkMPdasv0++Eh//jpQgq/vOdzlVH+WE
WLkFw3F4VMcIeES1TBZKduj3VojgVflzz33Xd4mfi5obS2MSIv2gfdawbcXdHH44
86aQaKLpZXOv4jD2rlemOeB8mW0bLVAKV01uxjk094Bb9QXEH2nuTS16HI5ASEtm
8Rjn6YyxHsQX5uC0j2X6PLtt3D7cd0M8MoHq/R8kdgXIVc6cb+HKZFAz1eLdzLd+
BhX/LHcN0o7ObPtD+Ay/AZ28HCWhBdGbUKKR0aptuhCIcGfKLCQ64oNWvs/llArX
XnhxW2vrah+zp+0Q8VE8pgmreu3EybOkPJnq5nMg7bLwDvRjowsctBk/60UhfbA5
9ekog1hYH4TV75S4ixozTnqtUD4Z9f64cmisxZr9hLPTRxeC+TCo16dTfwXXX1z0
wFYgmzrb4OBd+I5PnyDC+fk8xomi48VyC0vsceWU6RECvuyMt7BmoUkVGViIUpo6
b+JKr4xfJ5TQ74TGARf+IK497r+jIr2cvFUAkJEvz9IWmTdlkUOOgrlnBXF1BNzF
h4YOBtswYbgGFaJ99UP1acwqWqBjqHdtCsrZj6ZQ+Yyl4F+bgO4KLCAzj6vkpPr+
zRTTxHepIq7Vam5OTBBAO4wgyI71uib7e51jaMLoZdb6SCXubhLgVCrHXaxGREMp
8lsA0v3D/1xRCLk2s5qTbGMLkDCy62UHeeT08AuF3K7RpKBN7wQPCJscJj4y1nI7
UUCQN/Ugto3HoFFEZaq0szkms4axLfcndA24EgWNKWZtPFOgVRB055IfhVs+oF1l
9d/vzBKdycNKeUmHk2M3fbaTG1rReRikf3FCoC/I2qQh7eYIqdAbyPusRT73Atm8
mo8ezjRQ9A/xlowGpUFV03YW+xdI9FxTQuMxkw8Zu/bbj64bRe18UC72+xVO57SE
Hm2REXC5nDr2l/OV+SxrIySfvd23vh8QYPyp7llE3kYCTYF1yn63Fr4U2AaILs/s
siUgQ2FZuhx4Urknvb+emoJtYKDfJcPoAM6N2FPbKElPmRv0hcwTCntVIhMvLsTe
uDYihY6jpHm7A0y0CvtTIFCnBOukaJfVosSMF50ar+P5iZMQ2TOJwEgCb1DoUSSn
pm8efSfK2JEhDOPMm2z0JvviWKYbk8OmGCnDUaUdv/2KppN4JjZ5uX/oevyyYYsb
bOnbPar9doiTybQQIfcFEmpLAq5xEYGFRsMEA5XsixkkFwJgaU+RnYGeQ4oWe1Vi
zFHdKztgyYP20jEI8VVKTZrLYlfwhOQnT4CbqGjkLXmh45SZC2SPaO1uT2nclcYb
gF6vKOzyt8dkpSGBEL5IK4dPgNxMCSwZfnr1AGTb5+iv4X/cMdbucce63t2j2UhH
QxI7wE5qQ0Pt3lKKAV6AEBGY7pyLeMWN11bght/qo+DnCEztYMvFPZwIRX1KNmW9
kQQBf2TzTamB5yt5XPd7eLQCE9k3OBeguoEgEnpbyw0PdkWtAPs6YU7Drt/cQ6+C
mn85HJDhQMFVfRdtwOdvJ7TDZT2snSfvQeZu/mmJsxFezhTcwf4i81RJV5YzXOPh
JqXBmyPzZcF/xI8SW6jklwiHJwq3HCPHYLbHcrj7U/oOSiatNJF0Hl+VwxYP1GaC
clmn/qF47fEzqI/V/CuQbpHTvaId1s2pWZaJiE9J8ueXVRzn0SSJwEOy1R8tsku5
uOokmOUDXrZQu/INVs1eqC25MOiGc4K8jdYNALcSMNXiDi1F9+kTTwgTj9+wdcaW
sbPZRFCa1eZsowYazT71/1Bi5Os8vhh/suF2gmjUY8F/un/+1eYypT/dAuKLH883
yVxYw8o6Y1Ufus520ztz3kf2lVXOGSUxWbwCespxstO1T2IuHrthD/NXsYU1R4iv
MaGvb482V+lE98lO2ddI0w861K4BRCviuq9YPM9HuTjw5tL2M9vovinXlbMcab5f
YfnoqO2+w/qDsoQTHhgfctCkWyAmoLcP1CqKyYmqdDLILBiU2j34THOZzvPKIlSP
tNSmE58/pCAxz+V7H+Jy3cQVv7dUWW45OEWXqVxRL9QXLtXEWjmq7G2soO8ZEgt8
6L+uq/pC5lfUH8CaQ6rWMkZdEgpgeuJH8ZyPChSuzn/dIa47PuRJUUP4bE/p5ndy
zvqKy2WoAG4shfRmJMGypmDD2b3VoCNIM3D1CxGX4+akAzztx6Nvj5gOUT/yBdLg
5y2wRqQ6Pu2o2t4of/i5M2cbeTQbV5iY6X9izcgfQMuaKVaS5FTMU57kaZH96ffQ
9Aa/s5K1qBr7hxMrCd35xC2m+dBrtSXqMhEu+B0ozdQzYVbjTGH853ZJ8hgGU+ws
+cQ1R8cBWgDQsfBozgc6eMq6E1HDmQlsaJqlOyLAPUm3Y8iGul/dQF218oKW3JBq
7fDi3PWCj2iz6dWBiYhW4V2RcJJUwgZi4FqrnfXGxaj/27gKgXrai8HXz23HE5OB
av7ZoSjcNq5L7+YF+M1McGt4yPC7SvKu86wXOgiJ01ePftWQiJZlCap3LE7H7den
A4PlEmlpYgiBceX1ikkSen9+qla7su8rin1WEUyEmxKV/MVkplk1Y7kP4gb+uXkv
fWcAMMV+FZpc06vIDWhfX8arPBcbrBoEBPV/3D0gpbmRoUrLOD5eY3B9Np+xn5r2
9A7H6DWYXka0i/22ne1Z0WSikWsg74LAwMMphc1o5Q6oqqV0hi+E7VXdJ4T04qOv
AEVhAhDFZZLXWLUX5DX5qH/O+1Hc+JkG0iHQJCFTKBDeAQWWy41684zZGhqfrxGE
8XNy7ZrMrjpwj/uTbbqtZp/pmpKOIAlAsvYUac6s0KzMY79nDyQC2oXWN7wROP9H
zO1hr6P85q4NQfVTkzLkTU0tIgSqh89T8GCxQjr7Gl5A9qWdnuNGMsKT/MoV+nuT
0sma/fQHT70qVJGcyq+qZfGTgrtcVTCWUIlcxhgvs4BolEF5JOZhlIGEIC2S0C1Y
O/8W1rnRaWRvA1I4zME+zrkk0N/KMKnHHoTUZSC/3aYmJTVqp7dAbsPCX3khRfAE
JrfEvpJHY9dRfJj433qR1pVC9VxABgr9oyVPWwiA964W/jyH/Ex5RnI9q5beGHST
VFefDrd7qd1hNroK3szhtsU2OtKLL9boto8jT/PjM+1yMP/fORTZui0/TwWNe3i+
DRdvLGcx5S2MYzood628CmgBbXEF7IgTHtFL9JSaKXCI+hNwmkaD9L4A0Bn5u+kh
Ef/8fzcVyYA917MzwG5Vsx11rPJchkgMiUtd/YkUxTu5WnVA9b3O9IieDPgEJ0aK
q6lrWtkpJAnIb3h8tSSO9VQ5P3yG2TT2u3ccm7L+tA4vE8Mm8JGLysftEiF2Twk/
p6LHQX5/h4Nb6OCtkTphLlJERr1t66JPvpMnlQRNjbguXeL9APdEj/jMGDv7Kvxp
aEQ1gJ99bYr3YgqwxNyicUEGqFF2t0efmfwnAGA0922T7erfbrEclL4VQgdPucFS
dOuaRTrgnaua/fvt2CgB8TkckNySKDFl6hHJNFVsHy8kB0epCOj0cd6ZcbhHhXnI
l/UaMU0SyZwcoKVu3h4zsCc8fiCk/5YEzbBkUAzAM1mfIRB8Mzw0Em3KRHlwr1DB
XwzU/YXt2kOMkZy4uglfQW/fnatCOm/qpck6qBQv+ZyB7ZLkrjDs71zz+sTwgzcS
nr0OUpp40JsdZAkDq2jLDnwcKzvo7BK3TVDDqrr7dXc3v6+x9yjznalz21a225bA
frq8gyvdNo4nNVcitNWOQIWCxmebhhcWcBnX2wHs4Rzce6FGUm3aTYXHtBy5YLtQ
YoHBQl1TFpICTfCIGQNm6UDbrorqM2tg2x2o+kRDgrDUwcXo3fiGze1dgwL+VCiP
4vjYha0yP/CPQafyLI+/TbZV7YWGseyMu6I2HyoA/utMhx+sFOMjc54o2/ImhI5d
ClTReOqYd5cHCepK4ZRvGtNivdV2IA7cQidw4SP/hegdjJ1LQeLwIo3H1Ltyvh3r
D2eknG1msSUlhjuyXxz8wps2nJlCWsiJ8b3FbVTKaHGXA8ILCPYOuDCn4EpYp7i7
IJWjrRJGdUssjKLph9K+TV9YYft5xtC8OMnoj7WjNjof/b9DX/CSD3k3KywNX9eB
HIOP4WHl6pQNs0ioVPjYed2UFKPf4s4hKQwB75mf4xt5Kp+9J1GAYGtbE053+HVz
ID0+mFWzddD43tjbxuFOat/Em2Rk8q2GpFHppmpjbAjyehC2wFFjfeaO0vaFUauP
J1omMvGHgoPAy0TM/ZlT7NM94Ix8q/nDn9drthtatF79xTuzQ4HeGm1F/h6GeuYM
jcmTx+lSKlecQ1sr0Ma41WZgRRC71NJPOzcpDUPWACA/Dmxw5/AsNDsWWmDmaA4g
FvBEVTwWHta61vXIQSjqr6idi7GJB2poAxqAyor2mSYp7S/S5zKJHPFrUvSdFUYb
I+jAhA1nlG6Q0sO6F2A5wyyJ+nJjPRiV3tPkE3pYnwtue+1BG09ysBi42mw06i16
cB8iuIeiQJkcay6qJdn//EFfJXDi7o4bC4fDglSHb9LlP7tH1FcXE4VVffuegI5A
Np+DOPXdqnJlQ6bY4pksDU1l+G2f0ckPYyYVjHpRuh649eiMjiFLbOjqtd5oNXL7
IhY733tuFMc0g4YixIWZ+apnmCbstquSOgDWBvOTw5MKQHHNVoNK0EURAAmNpotT
RHry8hRIsZNjsVhyImggsqj+wWO/lLtBWQvpECGGRHWsPNivYR9axRQcWKIT7VWC
QcT6iGw5vDLVRk+E6gkvoW6UWzXnwDYD4HFYzEvYiwYsZsU9xEXmcupJSQ9Wlg/5
Ba00mFsOqV5i9RGT44DsFLIFlid/Ox+alPDUQniRReXbO2s51ShT9evMd9rAWmdT
RYvnm5Z5O3Xg6pMWw7MHiX2PKIuYZDZSL3U5UlD+JJKUISMgDhSB+ahxE4FjyhWz
qDazFn0MT8IcGbRqIyq5bkwuXjs8nlW3CprdzLbMSuQg8S7ffrRllID+V1RWBxKd
NUhhyuv9GfzoeTndR4xTbSHhxJTDawC3Nr7qSIRTlQiMWwLitHypyx0MoEc+sooc
uVQwkkLFko3YpLgGvEX9Hbk3538+Wq8imMDoAHPvP4fUHyIJNA5kdahh6BfW+VIC
adkY7jZ/nZNG/gyEcV+vrrll6s7es+NDTexVgYDlbhSqdwttrzkrKcYZSR4/uz97
FpqkLbbY2192X5nNa6HLiTtdjLjN7569dyxn46FViYR0ZYEqX1YQe7ZejyXYopVm
xoRjOL3nzOZj/PQb0DIXwQsurM+cESjCjnBJcib45brHko62rYkYojHpS9aGjFhu
Z52B1dDLbi5umF6mEz9m74SpR0Sg6gWNVo2a6yrzwdrEjoGdDZ01rjdmTx4aKu7U
Lf52hG+4T1/LUA92ppqYmQqmsbvYxm0q1ArlitxruX0dJxYOfxReJWV58c8P9fry
PRoSELgZNVTYNrhhbL8UQkuGKjy3I0/Mx639P3iHfwMst/m49ArduP81KZyipx9O
Liykp84Bbk/H0f01oq388NgF1DYJ12+Q3WH+zIptHtUXiKoRAJUWRz0Ml79oB/gH
79OKAAuCRsvYXAMcBwRBX/oip30ATr/zZMpJBN1eL5LHo6l2Lf2Hy1L9r0T93VLN
v9Gmtr2dnTOkGbI5rTMcYNKKYutcNKF+4NegtcqjccGGmlEXZVsGp3im1bCTtAdG
FBqSmplE4h+XA3o19gwdglFY0e4QusW0IgVJvpJ/mjSP6Ku3rFLcX22CsLfdnu62
c0Ws6msLmPDUATRtkrKXVhwJsaShpgip5BDLOu/lliWZiXRgcnotg6GFTISoG0LA
WXW+BD2/eyZXyU6r6o+VlA7Av3ELJwfxx2PQKHX9XA1uDHgZNYi6u3WRcZNInr41
sOFgLpbjpUuYYC2xkUUeIJLVfBuj0wcmBp5Xd5v8PIjNTenNb86vq1YpQNMhSe9j
q8MlUyaivDtNzcROailJjLjcQhTSEgD/GVR6spLvFJzjHl7mhv+iKGLZHg04RbPJ
glmR8fHIB2O81G1ZwzRZDlKz90J2j9JQDK6JtAX9Ol3446/cD9WFZY8cYtftJntU
q5UhZdkcEmlNA1hWR87Zt2AttrV3VyHg0mTMRR7dntfx+BMB+9X4e/GgrmQ6dVCd
ZXxV0Bh1QahqNyM8gpWGcggLmdYA5cQCp9gJ2d7kvVyFlpn2P1N8xhJW36pb2lQq
3wUyqua1GDL57BPhep00LUBXWXKsP6yEFYQPl6PKTYmrWvwz8oE7I16gtQ6MAI1b
GIbyfPQeelrTwL8KxSvEDfu3kC5ZpTCRZ+t6BCMANPs/Dj2UER69NYi2e7xXJ0e6
HZErQoOc8PeGb/1FdNW2VMbdlVbFTeBKVKsrx9y3jyJ4LG0vuOD4gl0+sfszHKnJ
xISOl94psDlp+FWwaixSrzYh2Se39UABJ9dLP8soLbaXWczhY6n6ktHtvPyrjvng
VS4RgyC0lteV0DsCaD4tH0YmLWunmdgt0ODYKx69jlpyBYb1MH/8N7TUkGI9AwjA
xIqxgiqlPdJUbyI5jCWy0LZ+GP9MCT5vmsTrvZbY2iZurTNJQGyyiOwBzjnXJFiZ
kg2Gq4PUqM/zxsVsclgB91/bArWkKfYb8KTM5o3Kd7nFCoi0MmT4UUjHD46Ueiuu
OWb152paKZPE2n9PpGm0oS2Ux1YDXsadyx/8ZLrl/ine9TDkyE1P40Oy1wBA+NjD
l2P2e8bY1iUWAMcPUn7TA6dkFHhW0Aqpu8WFzHsUKUFCGc5WAwvOAnwGIDrqbxvI
53YF/P40IX6iMk6rURB2ZjQdI7BeNYF6+2PQCIKZPVF8tceIXIyBrlTuZELdbNea
cwRSGbuTexPO8UL+nQmX07bCE/vY7CmPdr2VJOUWmTBZrExPXgKHFqKEBQ0yKMVu
yEpwe32yf3TAlLwaWnN5dE+r7CIUZbjS4rswP1ZW3TT7CQkFi03S+dVcilfxlWiB
B8RXbaOF10bLPLMPUwngOzKQlRvl3n2bAFD/3hl3ScLABAnfP5ZTWKWlygCSuzQA
hpVrXGzZ5+32KdwhzT3hhHbsmfakYE4WdIns9n7DcECOG5+nNyks1j5hntL7BrV4
0wvYZE376yHWZEvQo1Gc2Lqb+uavAn5IMPneCfPP9tt/yVXEWFmnlOwmaAJtzf6k
4cqup4+0R9DeiNQXYQchVr2B9/CL4c5+cAFUuVUU9hzyUO22bpA4wm1H1IPDkdKz
2vCyRRW2xXdc0bH79QBrQR9V02iygsIGLxnKd9c0UEM10ZF0tOHhmWfW8+qQ1fhn
afshG0oLVf4q6IcCMDHvoeCMyYR758edGBswTux+DdbinGBtsct5TJ2CXbVFOHPn
SqYFpHCSIm2mq+CtF9ZYHIw/ga9FtFTPzGuZjqP6sgAyyZ8aSQqeL1Sav0FBEOj7
klI1PrGLewOhOFcud/atlC7b/alQ4hTO5vG3qaN50xQX7XuEN5vJGR5yXrLQukqa
1WVYwKQHRp478NF1FiFcFyAWKCETG3HifjqkSsUe7VGHpLC+lzbMfhTsEVPFT/pk
LgFz2/A6vSpADMAVjKiSJSpqMseTR7YW+EKK4trsQQQ6ew94MzGNs2cWckbDW8iJ
5dsa+Ng3dZpYPES5oyA88kZih50R2qd/Fyw4tE6o6qz5QLIJuLZRM7o/SQcQQCsD
37E3xRyGTTcs++0sB2NcZ9K3/XCXUoMcxmm4ltAt9kvl4vKP1i03gfI8eGnHIgf0
dE8bLJxeIPssRqJ0BGmt1cD9ISXr36BLnyPrB1b7kLUzTs2VcBBpQQ604zbD1+/f
s6Y8MCi+5CUTOJHxAdLVYg93g6N7NmWuWL1jK3azKdrjrDJkvvhcNXcymaqQVUkN
cXuBrVnyaLindxWmpPBThIpra4+3nwhD3ITFgw2ikLpuuJ3eS5uOwkt8wbHFw5sr
MCiQupXNb8W9VDKTIfT2VT205jCabthOEZS5J6X1NOTEhEOXIQjO73jbUyiAhiyf
0wzXnkEn9K8YrDAqKn1L50SFFlSK4DNlmZ7frFWxRg9C7paOU6+sc0OXazmFdXRW
GNdx2JrsDQcVRRFtbbP+5Ud82nhI7uLFEM8AKvIUxSBnDrztbes29MNkUDXxss1X
RVAxO8QmgcoLoDiv35Y2dQh+rFO7mgm0Z6Xgn0pWrtAvGLBUFZQjHUMvhWFfJU+e
xV6v8a61ZpEh1sHDrG0PZ7ajfK4RdMSproFfaRFWovA9qlqs5W0fzxhnJ4gOf/q/
AZknWloe0O1QyVwej3+RHU+zV9J60wNxV3jJnhrIhHVYkcONw2zy0w7MAmElAMoQ
aXIDByXvmhdOzBfF1qcRZJ7okcQtl16IDgmfLfdeK9Xrivb86pcfZMT8QmXvql3w
pgA3RR1GDiKrRiXIsRUKG1KNx7BMC3SCZD1itiaT/VmMJmYMhKiXO1VjOqpwY8x+
AY007ToMsTQZPiVyILR/uKh+P9yt4Q3mymViF2WZFxWgina6z+xPBvRufyaFYU11
2bvyojBvqOXkGFjvezUODfZIuJtAA2mops6N0cMY3uxh16RvbofoLBhzR8zRVWc4
ibOBxjLM+jkabZoCthw97Jb+7lzyZkfEVqN/hQyHGx5LuPtCATIZKQ8Plen4rYAv
THkPZ4IPyJPGW6lHd6dpQhUwqHA4OLo42J6HdTtwgmijH9KwrTUtHG2MTThsKOGc
5dHt462D3TL+qtwUEWJ6f9qGm7ONxdpZm4/2ulxuQS2DVxnGBI9nBbFqrdl7wzsI
8eNwioUzsTaoLt58B1pNwO3eT3PNCo1YtkcERrqZEv8on+Oj4W2LHd8XSOdxncLJ
0fyAL1eqxEO+4M/svNxum0+XgnecdIg/8yaqiMhE72pCl7qqRNmhLq1PdveXtZAw
p3LB3I7pcH6qIbv5QMpAtNo3ve1IAF6YYSgoKLqGNatOC4v2aBLMtsPYlQI7uPRZ
2x4OYg65nKE1xQ4U/PMFJ1uD9s5Sjc/RbLwlXWA4MpjC7H4s5cbS80D9FzNMAm3O
WODA/GZULfaHOCoreMLo9IGesrPZTObMs2TWaJv8KtxfGTXZZ6laTeGavFLgWl7P
EoChY8LvZ3+QcpuBOChTLkd7E105n++KtUhtVCW571grijVUzGGXRZRXayFiYqXM
RSxtzd1mbb+LZ4t4Joqxxe5iw9+pF/0Js8Vt9oZKhZw4mlHGjeMLagVhuMmH+hx3
c78Ec9l1uW1VmcHwt2DffxkjEAI2IDRmwacEzj7i/V8kX4EtaUP6Ym2w5uGdbnTx
wQRVL5oo6/ZEqFgseCksrWPW4SmmrJuk8EPpnEri+z5LzbUs06GsYHi3UOt6qxfE
HSSK+m3GuUCwiNBDoHUQ6eUyRAD/tM1VHHxecNu/2ai2b6kR+3jLDf9/Y3OsDed9
b4w9mpvm9mXFEWqJt7PhA+ni77tVTDNohTTbpeT76glwr+D3tb9NviWWkTm8ONfu
9OxxSb44QxPfBqVFTGvZKcUSdVS62fO5pZBYhFB9uIBARsnuZZu7kcndI9CQW5EE
KkueokCpiPSb6UstAihs3586a3xVMh0i+pezeRNSSlxi99Zf2JVlo4s+6pqdITZr
9Sa8l/YQahygieLRglZOibEIFiWSVDIFM5xFM15qQQgWiXQCgUSys3VNT4Lh7K7w
voaX6CtuQ0B8lDZmARUHiZeN2nByJzLEg2PrS4tSMpYzopxMl445oC148GJO70Uc
G7VZ/90nYPwv2KcaCxuIflPy5cO9pAAwsWINbIhrCDWwvwWVX51H07Cen8HFTNwO
yCbHQejKjFk5USlJ4hUFkAlvwKz+PJhj4USFqgJnRqOqouIN3qeI8SuhjZAruFXo
nKQFBriKeaxOVIzv+J6SgzMlEGMsz84uBuTV8aCX7dDyBOxJr/6YXyQOzP7gKwb0
9EfOSwN8m/nkg0eoQx9txcLN9VjgAuQ8bYl+phmj9o4hUHQYouqPJVipXiO6Uj8M
OSjE2atmtveZ3+i5OqjxkG+pE/714SYRO9zADVWnRXOqpJnFsaEl/xLsXd96+y6a
gUjO+YJnf5hCTXkGKwGbTn3yZgO2zIU0M0otuuxCqxFv0T+AEWiIMJqLdDKV/+MX
vgYmBk5FUjUigcvoCowIlW/YAodie5VsedaSdvYp4pTX/DJt36vAjHZn0I8o25is
42l3a9BB97bw41kprnXdTX+ZxWvYe3/P/lyrog30csGWng1NFoQaQ6eE6EPbTBnb
1K5aJWG2w9qCsr2LjPVOcFIyJWLjEaXl22jYDxAlDTNcEBTda+6HLgmeOFJ3hpmK
aJBskKlJTmvJeNmP2pEC8B9K2/MydfKga+1MhoPuYD309oG9McGkn+AfGeOO/t4q
4vcBgC4qti5jTaxTjWGMUJQ2h52W5v0kfHEKTT4qNJ5rtO0FLj5U24FWFB5pXg9/
5i3vwqWksiLj4JQndB4bsm2U6NHDGmEsDLPXwxEiSLuniAkPMne8RlfzYB36bTBD
AnOuw7s0abJ2PQusTKi1Vpsl2z2Y5Fc595VBHa8uttHdjGfh6zs8k6E5TEAGyBaZ
3viMCVFQObEyKj94fiWCR+47Gq0CMEKKVU9+/QPcBakGyBTX9Yq9HJ632/2W1w/U
FxJ4U5y3UnysCS7qzXLrhGJEGCI3nQ9UbJuULOkQc4tNYXaGdeBXRKFWUNkoFFGd
M41uxgCh4tXECHjuhNKwN5mUISAMSMQe6iqvupUKMp/O+yyBStRKzKViJO3kpj04
9zc578KhzsclFGf9wly6oeUfA/7Pt5zxeAb8ulHyF25Ht3Rl98/hAA4HMf6EGIRX
PQMOoHz7ykT7ekDMsagZjt/XE921KzhVE7VL36XEE/DTW88+FGTM65v4U55m6kjy
AuJaxxRP35YwFfhBcmnxFmSy5xyvJIf0kFGT9/R5uNIjbxJny4qk3VnYPar1bWdL
ez2EmlsVShwUCrMhbP0Vun3IRJLzB0j+NTAOX333dujmPvaoXRDOBu3AC5/HPkO3
jeCDUZ6fDiIS8V2hBMlpouV5xHRPva9PVANuA4L2OlwU7weC6U0x95ezqk157LOi
zplMB1wfBezGLqG7dj92ZarAPSbwaev2Z0gfObJiLXO20gMmBf4LOPim0eTvh4D6
Yagx+YwKBQQwXgEHOJo1hWEvhRunDxJLvuwu+OHwJKCmxBqoarMEe7EMdDh+q53a
QoXeXgG3wdt8iOxLmfky3ZxbfWs9DwEKaYtCeZPMUghwrD24UQK1Kbtv4KK9X2GE
q8j8Ue2gQh/5wYk7YQa6xiDtSczwxpDJqxSemZCh2zVjn8ldBODhAijMEU9Hlx9X
Nz8PKtticzNFkEHZZVrpAU7Co/2SX99Drj2LFs1AtDsrFtqV066QgyeCnSFx3GnD
4i82arPIZBeEyeCniGBXi0QY3gs4QUG/0yr3DC5SqkvE+cAH3Y9feL0ZkB2tB+ok
jLkBpuhmPszSTvwaGcizjhNrnzNinqeI1XyXMkZZ1ilumopcWpbNOoGfg93u4mg9
98Aow5b7LrXOTYcCq5hHxUW0C+ZsEnvvTCh5wxUt3/DuDWMzOKpAqtyGvibMLmq6
WNpj9rz83Nzv6NXC5bTOCv/DIbeoOmyihkL4I97A6xF/4hzd1638RIx6g+jIJ6TA
cZGbcMa+jY6WU6d5wOTaIfUwIjHo7YeprLpMQf6MGyFeXRuzy4hkl9SCTPsQsXO9
zZxq9cwDgFW/4nAg3PAfgoMQqQyPfWbrbE6zXSNbTqPHxvQvExxQVr9qBYDRIsga
ZbDRreV9LhDxoT/YoMaU/k3lOVXzI1Xth2m4wm1ZLEUwDD5MLloZHRdGX5lvIA3O
L9W0tIKQEdzvmNibBrIYuCXGHPVfxvV0ApNLqUIE/Ep+EiTpisvUriBaz5Pc9luQ
JHviOtxgOe8BIgyioQ7KlhJ/8dzgLTY1wvZu3rxBOdN3Ugo7hcxGS+Hrjg2i+Yi5
p8nix362LIBTc9sND0vcv/o0opUrkyKlliz+geTKEAyEvDuoTHbxd1Mm6GZQd39q
4OcrBIgbwyhj29Cr+1hUWGXJpV00I6gVjCtrYn2OCcWXfNqhPHMp+xv92+3/Xadx
sfl80NfaSEawleuKgA/QTvAoUzWYEC5lpQaz6yvvvmNKcmoiDVBiBkBMBGJ6FF25
3mzizktBsDctEK3K1uw2br7UIaQlFecwW/HdJtRbUZcBfNEgpWXoyVWyln0I8ayt
Kxg+5cNz0lWcHpbnKoCqiVLFWeevFQmO1cSA6RtzakzSg40oOnsK5zCGQEdLxUvR
d01sNVII554pGJiyQOtSjdpMEjo9NMmBpGbKq82ra8LBi3KZAv/Iy10rfh4jKTe6
tNnJBxpC7tYQuT3LtVNxl1iEVws4Z3ie+ylsfbCv9wEWatBS3XBA9KfDo7Htd095
uSa6iEAgb44Hqm3sgQLsaUkq3ZfAXl2cZbQsHfVCmzZNoB904/C1k4f7+VrsBFPV
guJ+Hcfb+te+6EOamfsszf588vrgQWDkK6cdNeYaB+woR84JzpFDQXPR1Y7oZ1yD
lxaRcfjbWi1y20NWPEgbw19zSjryOnutkJK0dxnzHw8rpwzNN2+muxtBhyikB1vZ
jEs9X02UvLxmgMAEJlWs7Wl95Tg08NHmlAjy6fLLrrx7Mz4r6+1oNpAjp/plvf/q
uHBMv/ZHUi6yQ6TUBibR0jcpRllDHr7fy26uuyZQabrIeQ177eJN5DGltmE5bFjc
pYGKjigBrrzXN3jvtn7ap9B9lDkiLFf6BdQaHdrcPHcn1yfwim16RsArBjYC3ol7
FT/0tc5sfUS7I8O6MPPuRxXcPLA0gYlXxjuoacGaDllJM3zDS3V4+y6sn5OqoGHR
jURhJkfn+mHs5SpsBMTvfsG5gk9Ul5I9wBrW71R2GaGjVMZ5D4aw13e2kzyN1ZCp
Be+7lPt1uUXiXT41QWG/M+VNc1N2fCriE/fSzFaArYXHXn6ELaMsiS0iahgOPBtD
+mbGFo6ArC2kel3KH355SwQ588Jp9MkOiuhs9OoE94h7Jjp5TIZCRX5O7Ulepw9T
XnrM1K9pofByfNbJOASOMikio9wIJTF9hvusa0hoa2a1Ajj6ETnZL5Gm20bZvK35
obX4Ni3N6Dwoi0+79o3zEYsmACJ/MC1xZFyIghuheEYgRYAHYuUIBD3v2tgofjo4
cNK/5ZcxEbOAIyCcG3n/wEYKysLRpYSDAlreBzMbeveGzHExr09bMzCHhm2qJX/E
0eG9f983herrvoWpleVHcxxYWZt4lhJGUIw5WwC8yRLVlen67TRFVj7FhbGCvdxA
sbsRhS3/mceP7Bvx2ifmmVnGngF5EdZ/5EUY/5BTyaLkpKL13e6wf+wIMOz4UH+V
GnOWqBAtVH+2Bd3CDtxat8lsvLBBvoisV4CYWKhbDKJVKRBLPSvGW3qlAyjQLBsL
ppoO2b/snFDHqSn+YfnZ1iRhN+PoycxTPuw7irQY1N+P8tDSxqq1bYw7UjFWnkDg
sC5EWx4hnzL6QlIYR5ObRgVmm99JyljPaYGiinFftWDMH2kP9pVtP0x5olpxMkfI
jdAOrqaCmJUkhaVmbn7rFqRA0YoLEVZgfpqurLJ/7hIvwsQGcMpp040Q1mP2RhbY
u8cbokeFqtnOAn67tEQFy/qF3CDqMQf4rKtUQ0Olc1G4xPQyNKs3aK19Oqd0jWxz
H71HMwsMo5py4YHjTnIs3f6CZ/41tfxRJqxrnAMFsloqtMmQRMb/DslkERqgnNeJ
Oq801h/RDrNj+Yv8pzUN/yLEQ4+Zc2TegGCl1Z4kycb8L+p5NgU5NVByhENBwsZs
TYkg7TQE+JqGOr9k8K5dh91dGAtb8cNRkBwNdG1LtJ0BF7J9gJAxGCGht3naJlwH
b3QHXLZ2c/7h61m8xf5xH0R4Nm30a9ilLOmb7/tdzNfjpGP7Ef12RuUKJLa95TjA
fE4SJb1g/stLSejeEqpSy/ZzaKxerHlU/juakmZI8ihgW8cTyyt+xNZeV5gfZuyQ
s7cj/AehGwPmc/sKLyibitTxV4ZN45if9+jSQkFhSLipcPHLWNo2oOtLmsEKKfIm
ARlM/Cke+5ZBIXARoXHca5pdKI3pvBexGMJldzvh26g27W+vntPEc+fet081NK+G
IOyZZ/Xs7jvKl+IHOjI6sc/NFmwDlgraUUb7QewOPw3kJauhJt+zqk3OgORGjMET
WuVtKmK0tKoJ+0wEFSJ3W7FHbr9aG5bNZBIA5vm+MmBdkRJ4dfpSPLcvYECAASH9
vCaDHEFlkHwB0ht1/obZpPOvF6E+0Lx+f10aCpS5M4v2Mkgz2FRBZk0BWwmQ85uq
DLAHA7QD9G7CrR65F5DHYXFDVTVEqTRBDKXtgjGkZQ1asRiZwPkpTcEIEAD50HBw
oFr227HHfQ8KirLt+mq6ofHjcz1eVbhUMOkeBtfzAJJjUR6OhYf1bhrL+b/Hhito
otg2bOfM8GpC5yRqbJgqIrv6GioXFAUN7pkl2l3iObCJPz9cVasnn5O7EMkvt1CV
2sb1AwSisEQ2hCqZJ0R6EIwiQD6LEPf1wGc/ioXYHRDi8NnDyDvo2oEmFDuGKMyX
U8AA0OVO65UYMkGi5+WX4EAxvVOcBSp921la50bBoHZDsBPW5Cuv3YODLQ/GjGrS
tUNajzE2crDFh4LXStXArXIhMzhPmY0CZslNQiJFbSGRKfKTKXkMnz86zIO2xURI
B+vZ7KXEl5VzMhiVPEMSfMka+fqsdZ4BMpvL6iHyJnBsXnKyhbfaMJH3oOe9Ymrx
wiHiqGZ1x51O9nyqToX1/5cHoLzRd7y4Hm5rKJxcUGMaALS5BVXPtOg8Nr18RHeT
RJPJxHLlZJpp87cRnHgSyXToVGj6aeUlul3zl4kfmxaEff1BxAVp2UgX0A25azCz
sUQABPiFOXSab52oiuifwgyNnz4VnclE3+6PL/C4xzvlafMmkGgRHRlUGdGVhYZn
X8qegqo4Ea00tpZWok183wHLuhm3C4tJTWGD2o7EqpLWKcU2m9wCeFUvy8EqTP1k
RQsOISzke39/Mj0JErHPjX5BgpejH2XIObkeBTqPCDwWX9mgbznOH1FVkbXE7y0H
h4PFLLT7CyK6cT6PRH+At+V/UJLYoSJorgduFcv0M2V/p2iCKvi+VGKfSXNzJqmi
1ZLnAmvhm60jXHhSMZpw1ySGbM5TvQUdsjj6b7JvQzsTOR7j2xzVpldQp+4YERlI
k7oy9Ntq3+CS+jDxKkaUXU2P1XT01WjNU98atTi8L5/6AJ4gPbnXyUeTB9Cav/8f
26CUZniKuH57e4NvBEVLfQ/Z3arv7/HagBgsFYVO/UeS+1B7Y2FJLTFI8uTwHbCG
z1W214VQBYXpT9y0sYAlyAQ128d4t+sNIeaIKkcnhqTIbm/+b6CGzC7a+NeCtCSh
gsMFzE69Davmk01apOFkOYNF49/Vs9BocHotQWRTcOuMwYflcQaC87cjkqAfI5wv
CbFX1nXPY5wCsUWT4CpiJlNY3/MlSxotYOQLD4KbSU3S2DqpnxM1NkEwu5EhSrLv
ge0tM0XyFcEUsIKXqLnl+TCp8pc5kOe4SDysZnVWVvO9OvM/OUmZ1L25xoQ+nDKH
xYKJ4gQAlIoLwaVUeMnT+54zJOUFzJ8McCxaxvBHTPXeSBZQmadhv9z5Nt//LkQV
SWaDm7sjt0TUarFvRnhIGvDpDQx0rgR6kGf4xjcowca6ddh0R2uTBrKzAd8KED/1
GzP0TjUoPSxHCv2/uosCOZNSNn7UpF+KazBQHJbIgb0quZSKIWc3MnhpfxupBi71
d64pDtARBsEHsD9FRb8iQJCyg277jxp3khDUrtu9u6Eji/oE/La55NnY1aXtWwve
S58y3L4k4SGPF3s0B+7hrsqz1pVVYy5oF5kKrxg6Q3SUT9AT5HpDSQrhCxKXIkBM
b3XV1jVnAjtSU2Zhj+jgYqw7T8Tfnr41SPPt4o3rDZ69Ah+ssLYLE2RsTaicOpii
LfZEi90CBLzj214AgzSnvd6qAOvq7dfnHuIEyNYZMUuYvalwBeY7JKgyfWhttxiW
2qaIDSuqA1xAWN6m/kT9svcM86Kg9KvboDImEn6Shp2wSbc9kweBAgi0Tq54sRLN
jChLUejQM65AINwU/8YZzlJK8uXDmPZR828jcrT2UbLSN+UDPUuk3/OmwQq+MIw0
Zc/3YPbrT/hueHtWostxqmOMYTofpGM4ZsF7MRTmr5TuSVhbgZvLUohdzni+Kqr8
0RvvcI7drPFsKYOhtVye/zWBtFNTj25Bpjn7umZmk2JX5roB+hSjgKK5At4iL7RT
93OgyV/KudPa8QofVxi+SOEZraPvYRsb0GQJD0D5VsHkvWHWe5PaWJywEU4zMD8w
zULbCkHSoDaZSSFpIUDKXKguP8sIBed4R5afROM2Fg4GXvDvhHHAmt1ffS5+eTzW
sGzJxEiMm5k2x0jqfZNvsXrIdO2fohobvqAK6lSsc9/gAILijOzzRtbb5/ps1NMV
LlsEd0xVQTOaFRl2EiJDgo2YwhbhPamV9z71ATF5tJZUUlWCI1l/Gtl3s/intkRr
Bnbx+dPFhpWg7DNUqcAH7TautJ2s3tbrkDft0itDVCvM3l5u0k0MoRnjvNjBjNza
p2N9/WOyeYueMzHDHBm/DvmF4GbAaQQ8D6NVAZxBbJqjZS1bywz+3AHUcr8sTofe
22359DR7ocs1YNiUoHnfD/2YfQ66vcUn++3VS5A3PpfqcZFyQ0EPyPhVgZlJMtrG
+IpZ+kiNGu9mK3MpSJjQxomOmfkHlvU93KcjygecXGjig4iAwR4Lwhucnj5572IN
GYwLUmwNa8uyTFOucuFhWTwH4nvWWu3dkbRaKfwvmyRPs/tOPcu2sdY/7IHMoZvT
dy02jvLZSk320UJG9dnbvhZtiXvn2JXZ3JNsgQ4+kTLP9qcJ+c2oflyjDQ+HEOtc
y87tpr7CStmZpi2qAWJgWhi2tPiWsxCVow2uTj163d6Wb/gtTQuHdRfbjei5NgCl
zgqClGOfDJ4H7/eeCwkM9ZE9A7uHmc+a8W4d2ycI4MgqZTNfa6EOzHc3h+LMLis/
MvkQGrb1s9yoK5FQvHhEnXj6eLYS8vgQXcxLSru/wvoL0ojtqo/mntLAygmKTss1
C2vQOSrp0RW9Y5Z+0F9ZsMFEA78i7jvO/hczhPhqrrrRRUjkowqJm2EPZ//qNg40
E491uh2Lksn5yYdvp51o7hMUUyhrSDCRunbbm73DIwE8ioIQskcgMQnbNtxD6RiQ
141/gUff5c7Ff3hjRwhIbdZ61s4qp0zDTOj4CY/XOW2mkh2ClBnAPn4a58pvSil3
QgB7RrkhLFCrniRY+d0RgxeGgU93RW33zSnn1ZDMb8tIFRLQ0OTUaG0jXg4uHVJD
ItlvpGbBx7PNgc21a/+HlJ+R5GUJQ/39h8b6w+qWNGTB9KwtP0GeGvHMHR1Iszpb
l2xUQebAy2clM9WqyH0PH71YihzQGj7Ujm3vtB/cbY2eRzaGd8SN4Akjmzv80mEE
UCI0pqDu7T1Yp9mQocqLBCKOLfUcsa09SpgBQtz2n97H52NN4Lzp6UIDWmN6+fqP
WVnf3M4DFN/T9rfv2+JzHS1asWKllVTrV6ndnzA66AJD4+UK7jOREI/WPS5le1uo
eQ3+6b+lqyp5WSn6QHwanziqtbwVo8G+8tveZalHPERS5ZGAQKSUwMzaRzrEptrW
DvEspk4cR5eaTE5QhTpiTlo3ZNNn5QTZxrdY2Kcqhxuljl8hJNgN0m0rHgIBaVOw
jyq2WkS67EJygzGTVNilSJQv55udcxcvPC9WOeeLKTaA0PpC6V6cKLRTaBVTK+Mg
DA4HdScRyqmgTR3iQedliEQcAaYQBFKblraqR8yCY/ZDee95O4F2fO6jmamOn2Vj
RUYYGr6D5mV6wuxSZQ68Ojf31ePgJTSrwtD5YuZH9h1Qe98WfpkCQQbxtpIY0PSK
CsOj4+I7Lhncnx3cJEl9qXQJyYxhQ3i78WPBKH7xtmXHUV+bvEERjcwPPByS6Rn9
+HljU/22xTzrrRMaphI5c53kF0u5sUhkvgRuEzA41IZgIsE5KdGN8IW24S25KYNE
0U1DRazQeusI3uvRBBDoDgbsDafgsH63wvSqD9HZaPagAmdv/iKnAePWfJBAD8HY
sb9SnY8720QyZM2pdkF+O60JuB1kji2lrt2ta/0XLX2D3NExUYSCdrjfeW7fQRZe
1x1mZB7STiWkgRbUY+U9uW3BQMH52lDdHR406n4BzknZ8adnu5f61MKD7JrH/diu
EPtwhZzPt4rXTgZkeQBUygNxxOzWkrWnu2N8j16hH0Lt9Ei8s70ty4mt2NiZcHDs
9VMx5mUTQXdkPAv7SNlKeZmA20jO1LMUq3wEpitmszshR+3RpYZROo+vmk6kdw94
Ao2P1ygJSgYcC4QNf9d/3Uzf+yHvjnYm64vKr7ZuFmWvSRdebESmzgcWZQ0pR8F8
g8waWUkw+bPpQM6xGIuTFQ4aB1BZQ2nAnWsI8XO0tSDcYjUZl7UKCmI6WLOJsZ54
RROWNqJ7MOIwF/FH1g6lsTkUFf87XOL5ZufX85D74nmWV0uKGPb72MWReurf1kBz
kvtEhtqOZ9zI+R7IOq7h9w3YZXM7O9HLxlqlLNP8xaSsPX1cFq9MwEdf+V7EBKg3
F9Bb2phsed6DHlGy50h+YBjGP8JapRSWjshwqNZQQ+1xmbdmSZ7sF+WYCRNDAq+P
NYje++/rcRWveX+AdON3mzD2DmizPMqWUwJ2OnGm7rmWPG3sti59TuQY9ku0RlJo
QRR03xsy4g+At+rPx010Q0I0fviuPU2VCoNLKj1aNNPh3VAOHC+D+xmeWgIdcQBZ
j8FsiWXH8brgbqEQaLuqGW3DGCTc9k+YJzGF8WQFbMAFq8zvTaYI2Xmw1BAkXTEj
Rp1qm8YiUSwqIj0IQXV0cSCspnqfd/4OAQQlfKaV04v04PFJ1yGgcfmbuFFCL9uf
FkT1GSjAA1RlBPS8VM4fwmm5MeU6+YiZyISMeiUF564ErDib4+PjuAFb9pyDvr2D
fIKHBBx+XQJvEXKfykZgriT9tYECKebY/7N2gOTjgpc5xD9ULEgYiDCSGrqJE9pJ
7eYrrI8gLBYjY6T4UpmFm2tTKnGuvlbJT1Q5JYeyFwYXgLsAMc9mav2WH8BmcKN2
yS53vDPKSjQlVVWlI2tzfIs5L8PaGXJojZPFQdI/AEL1VTb6IVP3uueIdHzdJKao
ZgJ3ikonl4aLsOnWarDqTtckhUoPOKLK3AdpZcoHZZotNsbwoUEAYyU3mbAKeJKp
BujVWbBHlz/zwkYQJvEFbuj0V7hC4HTLMhTz44cK7x84yv+nEINJiKYKQAtTF7aq
62/ecettU1pUSU1RzhAVsLPoIek424RIR5rw3JbvSUlhtYqTSnDcbmQ5BcX9dAT0
2cPJLIliK7V+YLbxOtYJKsiyZBFVMI5PrsUKatcjNZdAxS0fL6i/TcIVv5u59t5y
d5o5B9klvkzoo3ipq02BteubPYQxX8KTYBmeClPZPYM6fRbv5t8EHxpEmsoIicpi
9FpsCxnwXJG1z6c45ghbLB1drd9FI1yt+fIbvhtjlpWXHonppnVRlDGmuM0t28Pa
FIbT/V7H0UQnol7wCdCe+FayCqUsun/bQa+jaEso6DAUiXZ3oeAL21YJ2GbiYVRA
do1JtQywgCG5MYbZY3/7maG6UOkuqgyso56ScLZ9iu6HLPy00WoMjxp8wtpip3W/
cD2M+/6AC9twC+sZIVYUSVGeAWEBKWcrzkfWoiErJ0MZ0Ki3kAq9Ip0jzbFmCxWt
tttjzOApZIDpO263HqjbHknX+f+CbnUfT4JayxomOQjmabqyd63+ZdU5C8BHk9j4
qfcY+3pG7pnIyXNAUqT7H6JfGaVcrnpcKcG+JfveeNOeRjgz5xwLkQdFAcXFPDg5
1ypFWCuIhYrW4oSO2c3cTFccROv9OMhMzwgsVMyEuX1lpfmUVJqnO/FUTV6G7fvd
4TwiMGVao8dHrUclFVCOrmJ+9ItW44DGkrqEdzxtow4fUz2GxXRrDFofXPTLuGih
hYTRDtvkgZecp3HpBWHUeks7xKmFkgKao/lLWSG/5LVVj20lL/7QOEFs+8k8ztbp
gB2d1YdoIAq423zwj9T/aC/pBtekBCOQv85a2cZyICwoKrkLwKfnw1lfPBrHHgDs
XDLxCjHj8XmTVLIGSVoQsws2mnlecI4B74X9GSzSfmPgtas6ZaSN68TrKQ8jm3RM
+RBoYIU3R5xcvHXwjmVzWoK8xuRp+idzlsAIUGHwtRdmDCRmv40FBg8XZ7B6AUJb
wozr1X6jH5StRjrRQlVvMZWOUeR/M94Teu2yJrSVQmM3hKJN+SN2//2hGpVyfDdA
0sCvfC1eqx6f2M+3cBADbh9AihRY0BI70eI3GxV/MClOVjCIbMljo3Tn2GZNQz8k
FL71MMIsi70WK21AoUkOCe8I+NDNmob9oz9R1SFZLpjGahU4IfBX3l81yxAoSzFY
oljF9jLdzZaPudqlWmRwFk6U6NqvRRICI6j7cNkD+Mm/P7OxnpUKApxwaoZB014a
k/pRdeZ80Flf2FbgJ1TzFbDMsF6+I1EEayzSgAlQG/iekCN2UqK/u+XQIBgIb9vR
ozfb0xlELa4VLlmBWwZpIU2ftk5ezROTYyQyhOMMydNdwckfvptFURR29wMUDiqx
p5AR7SHhaiPqQosbWYpYvTNBdUdMWyKAO0Glu9gB6FRI1G6Y5jRl+MZwgiryOcFo
6P5xALIqhvxOOfco3fuAZ76xzhEQ13H/SuQx7iK0cr7DCzqFctE/a0rfuWDhZ+E3
K9EA8iyOm4MQub4J3FJYdC6AQXAetlulbk7GtV2R/0eU7tO2wV/GdCk37USPE4yG
CKV7Esbnp7cUvRzmFSvl6evui4yUSNK6C02ELgGj9hoXLAW/Avualw7mo0LK/cUz
d2LB4Idqipp6UNHJISemTGSag28SwXqtBRxZFIaPA4EYlkMUN/tpO0M0DiNrAEX1
QF02F7AWtU0XDC8h+iLkbSfRUq6H6m/ebJHZBKsgZVKsy2q0scqkKRZXNMsDyOb5
hpt6I3nvaJ+u99DqeuFDbfHUXowVAwdI9vKSK5iQAtXAlSFX6423UOa0T/GcXC4s
Tth/Uj6vLbd0gCqDPHQ07/C+mQa/QZGV0zpD6ufaARI6EL2xKF3TTYKEmxQNPKh/
AJ8z7d1DnUMhFa1r8AMwQa5Z0g1867uc2f/hcItBKxGw8RLr4wGc/DHq5NINNUB3
DpuKIp/IszDY4vtLsfjLoR4/kdWKUYwXrvrw5u3xdD10mSX+2EzPe/fJqWVgUUCn
b+ewQUsDQN+clbOaWNR2aF2p1tSlhCHgi6bjvGWICdT16aCn0bvHKNWR0WNsayzD
EL6UJuQd/2lT/MSlcSPuvQIMTtxIHSIqCBpEPyEC9SHOMxMCHDilnFwFPflIkPe1
5XFOP9gAvCRgwEiXGfaJhN2NRg8Y4aKB6HT6l7j24RfgNLlTcPZ9vQOVsVb9QpOd
rPFFlfMTwl/t64jUDZTLMkWHNiZCtBTMQnBt4RjOSuiInRapfBOtJjpJFwsYmvQH
Yj8R1fkwN3Wne/JIOHpqbqGxFlX14ujaSVvmhAXWWntAUNVlacF9YZvNOAwFVPMN
25XfzHvqQAAVDzddy4nwTL/7ecslqJO9CcmcH/NINv0yJ9e4Y4yA9T7QsxZaNGzp
ojz6IqBM6btX8kQ+x8j4ZjSCa19WhT8pqXfAx7hFKthx0+J5wnw111GsJRx+Jiiz
0Pmtpn+Sn+iw0GK1TjOYJRNzFzQgf3dmHXv1CcjjRsPLnmswUHBHvgLW6ijPlegg
kOqQI0ef/rneCV2kPk9FN7NRww+H+kvmoK/TLrooyxTD8KwvS65oXG5gj6Fir0/F
QHZxZvt8t1j90GTcga7GDNK9qwJztpuBWhxyA+oN6zQN2lmxqi10/AWkIzPHKViQ
xzjrYIrui6YrQ92IGkAlJpznCf0X4lEcQQBfeEiXdccBk/3VIkOynGb1iEnSsehm
38Zu17kNDCbnklGzcyv5yqsLnzXN/8VWi0lozOmN84e8HxUdmYPf01dNTluL74Qn
MG3Ncjg27sEybJlvMZqnqbptE6vdv9xh24ao6+CWsTO7ehYhDOXPP6Cm37OM36xP
omuw5i3r1XKoB4L1CxjspVxIr4Gigrf6cmcAEG2UidSIdMBotiLg7XvsRoNg791l
r31COECqxJ+CJr+dDkrprC3qVdTzMHFcZd6qdU7Cc+Hyl5HL6ZCJyOCrWIHxAwD1
K3EquHXpSopDEJ3RXWaYBjUT26a9tZOKsPJBnux3gG2fl/MumjnF9z4VBh64Jvd2
gfP5Sl8dYRnEa8yXGtS+JIXlPEqDpAHwNsf3lk4nuqpUXm73rNiRPv9vgg+BuPO7
nZ31NNbzKvN0CnumP/2cIhZ2eR22OMm/qmpX7755R6qF0AyPd3ap7ZsCJftGqZxF
evIMoFO8Gr3AqDq9lBp+TrAiFCsk9a3jGAb0+xhjr2+fyfPUl4XS+3u8Q4UQ9rQM
n2s8rJGtbsqPTQgPf8jqdXku7me+FQsZuz4uzfPZEu5m+X8C2ofgWSYRUWIaBJz/
X5/rzD8VsJ8KuWB6tB29DmjctSt5X/afhze54Y3m7IRpk3uIylGKG96Vk/QznYuC
dIgqW3sDpNKCwR8R37SVMysg61nJmhYrH3ZqWZi/BAlzdmlH0UnChA0wJTFMUmin
MGi5HNSMdfEcMWZlSYJ5lsm/b7Oo9o/xFTOH2As3HJxKN7etCtJ74by5kbvxULWZ
reDu6iPS6iET7l4U/egIrf9dlxr19npslYNGCwU09ei35ALCr16dP3abUgxn109c
1LnNzVDeWnUsEpZoTN9PqSFH4o/+FQ4iza5Is23UnQjAblSrTjZQKsosjNcSPqQB
plPE0vo6VoFk2X7MQ/TbwrDSsk3RGP3icpsp8de9JLwA8B7+NJNszyyxULJIBu8X
VFcoGy18yhjviTf8k+Rs3dekrBe/kSyaocwGECMJVKgU5JXS5r8q7DF+FyyxOeQh
8T4FYnkAT0mCROycEL573NV/f0YYByKJvbOT/ShHjmTJKKnWrTVoB/5V7yaUdiM9
fG6CLJtNvPLRjVRyFlIeajlgzzrTt5Tgh3za6gyNizQBp/f+73jxSxi+2NyIY/qR
G21+NT1BJYfZD7ma1pBzeJ60CjlGiUIvDOitRZa9lamrFswiX72uJO3GcJSAfoTH
qUH6PMWxuzO0zjYhijaRf8dUdcjLvLTdu9yRza5spbVdVmTbSzErMVZrgdFfILsG
R1mE7HM8hBUIxXFlfFDA0OckS8jv88nCRZLCzzPVlah+ft7yRCQyt71zeIWiFz/Z
F9itGx6sZyCjML2fuCbygXemKCIGoSWSLisVg0N6AZaWsl7bnI3S4ogX4ZcWqLRx
anBlTxi5mbqMuaDLXQCF4hgkke3LVborT9kxHaDEUXBK92+mNn9IDsahUEqjarQ0
hhewSg2Lvr8sYNKD1AqFX2P7zz4OBKCDmwyUjKL1TD8oJUvO21pp4nU3bkbIrCFv
GsFdLvU64b6j3iad43MeLPYh9uK8haddA/eew4CRvPlTQ5tkFgbCz0pkVTeHTUb1
PkVCALivGEuS5BX8x4hvO1vA9kd6gxTQBH38Cxh9XYzKSWGFY3uiKr03E6w1sxxZ
R9bexigLU/Dhq/Z0FyJZjRZqGGoAYjBlDs7SKLvt8h3IzFNblBfXpLx7JasUN5xP
4040LQMvnlF3VQVxcSFU084Yvfhrdfu0TG40S2hcr5o+pGpdrXwiXzsjew8bPu+T
lvxxjnsK7G1blq9xBAnvMnmxemNE96S7vuiLlvlio90kmho1Oawfx9BztUVb+0hQ
2oV9x2iU5B5ZO28SkBGujOYL8eadXOM797uVO51jhuuWrb/YNoBCmdGh3Db7S7Sm
iUkSjOpHOjwbn2enpiKJ6czLboHMRTRr+VlA7HwZlNUbXgD4cPAnCpFe1yIKP44q
H1BPn8F2ZnaWid1jSwS9GBRNMVNpdkc+64tivrc6cltMbEOesReyuC63Ho6PHZ8H
vESGFDKotQBQjHf03kbfg9SWI4MGRdNZ7m8joHN5mccLVe7S17YX+PkBA9W6v8V6
Dqwgv/FmA/cnI8ptaSXSTc9cZ8wLb9U7AL6q/yLndlWc0tBZbKoSkrOXdIFDJi1L
tv57IWgOGkRSuq4J68gBfJC3uhty0SUQWYv5tR62HJHxHEnXpAqyR6PqzTj2Yiip
3rQal+k02I6+/8BhXncEGHUu95sghv33ClsOiqJ5tbbm4dSPuH2ItCQ7YlWMoHzD
qHOGoNYfd5Jt+MMWsbHTuyWiwOs8pjT5isOGx0cp2W90lqUaEVzqaQ0QhRCLPJIB
8SRZJzXo/tNu0+vVuhIkN/duCL66EUklxL3N1hthpuljL0IjrI0m3ehtLul3eBAU
kiQidGhQ7QnOJcI5aqLEJblD6VxEjOJ8tLELLACdKcUd33VfB8j7l3lwBXtX49Bt
gsf+8aBLVjd66HCYJGl4SI1ZeokTFdK9zSdM3QqQDtOBEbumsgsUk28J/IG/2AsU
+XRiQ2c5D1xEfeO6QuJh+JkS3ahUybNLvDjXughLpz4jMdfkOyyKEjLsUmgeyn2r
Odx35VGdk4mJ2cimxHUMw11vwKaAcRgczNRtYRwBwF7jmZtC9igb9CiL3b7uCk6d
6Lz7fyxP6BeUD//QRqYaU9LW3DAOumvfRuNl3aSo4aZB322uI2gg9oEvyGwPwT5p
6vjfCxcM9jnu7FWpxguL322n9QFvzcTTYJIdy6MpfyMElGi7Yknw6wVtQNh2oZ15
Pb/PH3fTXJX8x74a9sfNZLdeo7Z+dT8RUGPD+KtEWyV3fYBjhiAcn4v8Xeka5DQk
qbwxVERZpBp2yTMmwDLB9y5nM+U+F8/Nm4yYLj53QlGKHVkj+VOxEK3dPKGVoJNG
Yt6EH/WLZ8X8KU/3RjHrga0Flft4U93bK+HiXnNuSp5tjfCmwuKR3lJods7rEx4k
4ohwbm8mVhkiI6qnx1GDo8FmqPZ/E3cQ8tVQsqcTvyX6BlsjbG+1GVXam2HpkFKk
ld7IO399k6gljwWwudFzawcw1/qlZpzFsFiIqrwYfSW29LRtii10FCwKZdsO1ZEh
JtnsxY3qe+AUBP0xgjwSEqZ5H041ryDk02kFAXZpYGvyrDw+P/gA7DUxhrLhgkg5
ZtkN0kCTXe7bwsLkBYHSHz26cjzt90Suc32C+M3APgEUw9uTl3KniKP+JTkCmj8V
z580aJrbp7etBw0lbJVXqJWRmJXHzxqADRDJG7JipybmAtkP5BVKglFqYN3hHLx9
W2pYwYDNhtggj3UvnxowlWwxZQVw5QhCChDliN+J7eh0VmlvQk4poARvMhXlxYNK
ywnHnK6bHI0LtTbmY48ZZNg7brHeni6SXlSZxbVCSp/+RtQGuUVfv6yixI4KMo/L
MTRoONu3BJp3NS7aLgACzQ3njey3RpRYyUjC5MWq06fhOt2+mI59UKO6QW4AU6oM
OQhFU+o8rfmbVmj9yh8LTa1XVmlj5jE56HdzbY2YWH+Wpl4tqU4r/541Mz9oap4o
FE5dW8izOBiPRrDQNmMy7N5NR42bWsxBWe0ajUabgXFL3ztvf+n5bLig9Vlgb2Lf
Y/8yalTGimYkCMpo5jHmpTBje1/K6EGrqRLchioRL2OgPxwlKnUakucFkC/qZty+
JaqbQhGxL5hdu7LwFjgMG6Gp37AP6h4i6WGWPvx+Hv8M/jdkzhFciQL13BfYGDs/
GF6k3qDLb3jmEAKyADMDASx/up5FwRPr51wDNRq1vZVLKKfYj21KeuVNlZbM/Tcg
d2zwKBc4ztDR4aEV/Hq3c0JY8oJb3fHbqJlZgls1URj+kpCbghbopgAq0bXujAFs
GBx2eYlxvNeCc1dcnvj3ntGtFGQJagkhdX2Iex84zDpfH++qAW+93Z5D3q6eZDxQ
d4aR/5lbBwLK8xRsjA/CiyyFVtUeyF9GXzy7w42GtxtO0fov+XMucwPqXEQVmXG2
ExmQUk+04qQNQKchQueneHllgt/bBlGt3YI78Us8cXdAKl1ywcwETgdteu89wSAY
015T37p2mLQ7yCsJMnLINVy0KvGDgld8Xqc3QB4n3I0qhsMkUVpdG63nmeVr7dKv
/na7pKZaZ8EbInvcyoDQn6ouNE+20v8P9Tw6gJI1M5pi+9RBVhnSj2kEBzsUoMQ7
mT6SWHWtJVGsv/4MRfzUKv6Eu1dEKdmXiN3F1Jzescov6LSOcYBxTilWEWeZklcJ
H+Uj4mzltYgByljDs6PNxbZBPYRvUCLT6xQNY8IArO3nCMJPMxgIlb32E16n3bkP
mFZIPsJRgSVKj9yazAF5ccJSWyVc00QHVAaYzaDQJIxvgQpNY0mzgL+685bys4IM
NYBYH2esp6xnSOiypLnZoMGihrDfXtX8OPlrZM2DptTY1qVMDGlfTuXEk9ql51XK
TAAaQwRsaCI7K+ayT1ezRo9JBFvnZkE/JrJnH8vVz/ZsGxKA66p+wt4i4HODmFm/
3ToysyuXK817deI+fLDT3XGCU5C2AjAwv5D8ASLsSVV4/8FA2rQwNpjRb3Xm0etZ
ipc1LFdlPoj6byksgRdGRmweUqt+TP/8JsI0S+tXqCiRZ7zGpk73vR6OpytVmktM
naTtgkxa9P4reM3pC4UrKwDZN32vBSKFzzqYgDx9tyfTD4oXMWeGC9ELc/zTDmBi
g82EaEI7cYq/VTdXl9HWM/hG3HSY/cwSkVzy29GH2DfMm/Z1X8jrqCYNRQgpEI0K
tPqvGTTchAuEUOaWwggVUQG1gbO8dsDnaFf4iEPtrJMc/JsnND1K/yf5whkmKS4o
h9Axxj1aMKeuIj/WP2X1AEdWYfxzgJseuk/xtM+miG0jhsLdlppPlkppvdZsAHOM
NhXavefkO+Pkz90fVR22TgtUuLMVJBis1d1xZ9oi4HAsQPk8z4w7Gtubj6EuRklJ
pXBDAdGnIb1mLUGMjKJVyxvIQbSmK7Sad4yJ3ve3OHqJzkIBKTThWo2Cu+V4rtvn
4Xbgrjd128pZZMG9ZatiueGl8c5aQQcooRkzJCkgyV40MhSOgnomXxON264vt0U7
uxS+y63EBhLhpz+QXrijdsNLA6+rvW1Xj7Udm495SB11yDIALMEqqkb6UsElRgaC
ZBdgQ3dfVDqrdFs8/ux3fsCiwFN7MtSHYUMLOVR54ab84svJ6Sv9hpWJB5k5ALb7
zOLOWx5KLNbos/MO8qMG2EN2tQ9rRj6M/RQe5MFWYoTTGbKCmJX48pnibo8wO4cJ
LgGXWO6fP7Ahh3zuotVd3jgizhRaAGp3bI7jW5yItehKOfUUFjKuCWOodVwB2IBy
c51x3noZjj2rjTnHG8W5dLRrV750vOD27yZl2giNLPIvyteOnDUvcMJUoOqmEKDb
7wNtHxSliDs6VU5qPLBLH7kdw/Yz8W2dpFhb6jLiyhg/5y/JcdSaWm0wjDGqEMOL
Gao4+c48YJgbZhVjJTyN+OQUTwpuPoohR0HKsLwQBhJKwZcVIMLeOrt3h7+Gj5NM
vZkVrdVv4TjcHJrG3iNeAv2sq0u45KMTMCyPUAQkuMAuFP3R0RxXl/zIFnyuu2np
g6reP0q+1V0djaSrj3ilgybeClDFv8V1OGRjtHso/UlTVd+4aZ1frxNp7Xp5g6Yi
cMK41Ac01mSdXPbmrYo1BrUtnOFoSnEnuvxUihwyqbmMSRcnxHHh3ZCnxcTaipmq
qiVN5gxbAoIC0eeDvVcWrFHfnVMggDigbNTKHv3BHtQdFYJP5YCtPkx9ObNFo8zZ
5uqBQ5e4MHF71MHGx8hrcf4uTJbCkCkLxNUhji/hk5+BJOZu+ud2BOsxl1CAvfSg
meSn97rDd7Kahx4HGa/0TNB2XQF3dt46mRJGepv6E59sl9Q8K3nsvNgFvlA5M4Rn
d2pCRIuLjMSFHN+/t58Ok/EED22BomTp/A5Nv+WWaJ5uWy1DWLCs4oao+bvhgymi
WnC0XVIAz91t4CTRROvRF/ddU5J1C5+Ii9sOnW1J7IhVUuk15UIAiOM6moMWPX8f
JlqV53NEsOTxJbhMUOvQXVcbpmnnLug4v5WcVIS50I7GKcFIuuvDXkqoiXEcK7La
lV4xlqwiKxu//5oqKXiiGQY647UClNUDZgoV3Ym6enTuPKwlo559fAxADp1lUKpL
TOAKR0x1OsBK+bGjTVr0UUa7h3LDhQLaLQt2XGjfaE6Gd/2zolI9ezv8FAn7SvRT
eHbz2XzIHUGM9p1bTw6oS5tqwnnJd5a9+RCqJikSA+WAQ2hlFBuCkwRkpvEnDhHt
iK3V2lzkS73QivMx1uRSoNsDxby1kYOTlAfbNdwrarGhG0aLuwPm50QAnempllpm
by2Xvmv0HUkVOCM4VhUUeprBPQQ9hBtuNpY3t2XhbrMSPfyVtydQ6bJG2yjJdcXn
yYw7hB8R4KxWM/v0pPjbvL1YfPZV4ot1LuUooF++u9jvTJeoP8ZHr42ZlvmIV1Q6
ar+k7ojKSPGAFwWZ5dGmhodWebKYjb/xR8kv9kENLbbP+Fr1sMp/P11kuNu/DwbQ
GO5zi06HXWrIfhGzXTcxFVax43Ojz+wRTp2KWy61g9aeoz7xPGqnaO43Th5qnwWZ
+4xWcbw1eNQZCXxe5qZeulEIyGDk/Rv+S6byXujBcfxuyf3/Ud9yHl7CxkVkPUKo
fWSq2eQ7qYlTl3h8dXRPqUecy7xVi3sPK+WeVaMD11TUZIBOMlWNrcSBdhLHzlsr
2OX/PbWt+h+QALEjLp+fjOl9fBxIZQCDImWs1rRawZs/d5S37WN1RTdS24RGXrKL
92jqP2zHG67J4j/egSDTuQOA9eSKa2lx95xGulSifOeiaUTWv4gD76AAbxyWp89V
WgiGfM6Pz/dhEn2C8SiMjOkMKCsz+Vci3CZ/ZYhnpCNoAHv6iLVpf38+/Kcv8UOh
47gp30SeQ9xxR4wcZUPV4IOFPrlbh5ekY1ZdC1NO5fZAhQ2VVNToyYmBOaWxbnX+
YuWQyo4U6BqyzkUqHaV0q0JUfXap81MpfBnDo+IXbWYFrCDPaJvaqlcQUVUANYa2
3xrjCu/Kxx0HYbi5R8k4yBx6b9qTgHWtV2lFm9PkKoStlHjySTge4sy1RsVTHYfD
hRLiKAgSVvmNxQ3I/viRt+9h0fyOM8gPF7vHhcU7EyJUUh8Fbnh3NCqf3oBr3dMr
dLrCuGWIyKQVdopVv63hJ+O4TU4WxIHeydaViIXTr/pEeRc8A1e1d21zcCfKQdHx
R0Xe44lD1Qj0qtMeJqNyJ3nakdc9RExF5x6uKsLwEZmRsoukOEOPCtqLGTYUxnO7
WyCErOy4SL1SdWjmImfjlqTPv7ACWxBzoqvZIwLhYJlOWxA1lbBlZrINq9ZdL9MJ
TqzaZkZzqUygGz9e/yIspyLVctaatDQwgF1+WRaGF+hkqsBwkvESG6uWYx2MrOeQ
JRmm2PIfuG/E25TLE1giBkM8uYuQvv9smgQozVzv9BjRYsK8shaZ2aWj4hq4gqhA
Ple2bQAADMEVv4/yRXimYOhYCiw0WxSKPfuetdWUzuEKuKi5lWYEdZlk/9AbbTJw
yvisPAiIjjeTi1qdRbkYtPmZOsWN0TccYlq0uZLhx7871aHZpumo6gYp0aGr+NFB
0kqHDBvW1PfwfFp6rkoupl7i4CE2SmZ8+lJDcBH/DN6vcrLy/8Gqzhtwu+jsKMti
W18kBn+yKcFLoWFa2d0TMc8CaWCVpZk3V73AZe4/B8JhT6KYDKYFy516E879f0M/
BGkaW3Srl78CVsC2m6x78qEXSG5Nlkjd6uOXn6aVlNtPqN0yXOwQVJHzGy7L9vfj
V7BWanAN2LbGDMf5vFzEZ7u5Bs4n9IO4iArYgwr1fPcap4Q9nuoBDtLVUAY0ZQlj
8yJZWSlS8hPqeHfoK+zhe4D6oDq+wRNdoCBRSEY9swzDUmPlEaq5BxOj3llJG+jp
UGNBVN5/+qXiN5pY3HsL1/7uyA9bL9B9YdQa1+FMKpdm39J7/7T+KQVvFwLdyjG8
Xk4Y5uz6yWl+I4/65CskuLnwRP1J/scZKBCixDJN6w/QoCdWiLfVMomULT8SeO/b
lyZ3bEuk8G5v9lemeAosJngSWXkyA8IvAJqJA1XyQUbT9NIvMNtBdO4I54zIvMd8
4u8H/rUDX+6DwrSqG1KXhjFm/rsbqkaHcIaSmDJBjuKgQZ/zJuM15doD+eIw1wMR
QF7HXQL9EpMZPlXvomnSHqIz0Zk84bbcaQLNmFriXdjT/FHayOx4WrmYI7YBBlcV
Dn6lYIKtS6qiChzsX2m/a+ZrwvaVuLR1miZm2vpa3M72dQ1IUFG2zoycXxrFO7tR
qeKHgw2rdA9wrVS1tHVEpXZmc+7HdQ2fhv5/8q15abhX7syQoebFKQNYyrszEOmI
7prwtOJvlcs00IEcAwU0GDfUfapzjkPtJxindNNg/FHKSTyLWKDKDnBY9n+dMbro
psbZ0/NAbb3qBoYs2L/B5y/x/VrwJj5bdkuIEleDV6XSHCxNOjpB4P63vCZSlvSG
8S4cMqmGhepJat4QtEM/oUbZdXTcE083YPR5foOV/Kz8tQzLD1EB/HXRjidr6/nI
lB6ZNz3Yia+S9wYrPHpuablLBXQ6vENjuWmt2Ht6tkZOtx1POnt6Ry6xu2shJdrF
lFynH25uMei4TIYg5nAUnC2kFCZy1J3131d9YDmmGuQZcIFxsfzbVERECDuOjB/1
TL126PwRhUTfNBsXyoJ5791wENPbeMa5OPq3hk8tb7hFuTfdI6OCyZha/PCEHKFR
BuWPlipT2fvEdiBFgTX1KUataZcQId7vw33pMR8XJ9xgVVBHpwTp2GregfzQZunk
mbv+48hJ7D/W6pzO3WH76x2oNr9Mr0IlvG4n90//qtusJsyxNxZ3EWXy8mmw5+Kp
E73ceBvcDoT/ZlecigXiMTycjU+6+uH8Av3kKgrpbFJiINa8lMjzu9bHCRJS2E6x
2RwytUOdUFo/9sZKb7GHTyYTGgzMltaxz/UCkNRQAlIsN96Cyaq0aCA9R3kGjzke
Kvi7NLeS4Xy4hFS3PpnddLxEme5DumuX53ahdIyYRPuAW6rJsWukUnpF3B0jkMwW
Q/3D0HT2GoDua2wAFCPfbaxsXduksHYJA2fIC7YxgD6iEIglK1PAeVFAvvp5THp/
mMvxhOMaxx80+FVvYKwmu4kBEROGSr231NnpMjLzv6U1eDvQ4XaJkUSod24u+K9N
/uhRERkbw6lV2gHrrpoKfvTxKflX7DWIBWdrp4Zg85366i0s+fg3YW9VegqLfBtq
1+bL4gqnHKAsG3nd4C8QNDEU1vhFc8Htmyek7kVM2To2Km9liY0Ao863m7G6vlg6
WyBpNAC7SlRdJ7oXGDgWeXqFo+ym4j+9SyXvim8XBUyIDjAgwbpnnsuEwLmQuCGM
OYuYkgjcClELAx/jylrbi5jMPf4DVnAvFkOywIVXkdCRgXLrgNw4bqlNUPcm/Kk1
D2YXhjih+830meX9sOfkPy/wJaUqvXM+o4HyqhQtcQZTL1dFSnQ814fXpyxy3bJI
8AHTq46ikQkgdUb9WgQoFw9F2JYRiUXhcDZVkHKYVAo0ylolOOb0hRZfkl7s11jj
+L9FLjBrrL/kgNis2YNccLWtyOfvnMN8Tbed3i3zNRDsG1fIh9yq6dzBsK1TJCE7
dflEwveosJzm4eE/P8NQH0htPSVec06VCp5U8YonPWotI7R7JnOHERehheT/OXeC
cRHGgdgGkQDRSSK9z9oezT4RFFtGZdAKs/BxYKygTRJdvjlIEfPLULZ8+UTiKLJ1
7RsZL3ZL2ulvzyMvgDV/pBmH++qEm6mSdOVZ9IOqkc8n9bkz9Kh2xFR1e3xj7M8r
rRUDyw2D5rqMvvbvVgQxjYy+DQ6oiPVEVi5p1WxAymDQLymM5+7xXhIw8wChWx69
Gk4hZ07QWTny55AMYkBuVM3W7h8QvX5HmpHmDRLLSnvF1iS/5LAu2b7FT25KKkyg
UA1R3l8ZUXzh2FLb4zJfm3JdSsrJuvB3ITzTqJuBvtbxdUhln+lwWZ6LN/wMgzyv
/Pgk5d6P77l1nC2WjRAoFBTugiTj3vD0B8/dxWWrpviOtZLloHqF1CDPkEcbjcP2
jwHH3pLRQBd+E64ao0jClvk/Ygj35tV8FUYP5MvInYR3xSheeYC+ICklmy0RdgjM
SYv1fz+fB7+BebIofIT/fXLmhlccTgObDmSHWI/hZYEuJZ0If+1NOTanZHX3mSiF
O/1G+9UJvPyxmvUfRkDcXyJA8txVB9+iYADSMUi30IwsitCmkP6248Vb6fl9P0SS
/vhWmZTKGPJfbLnDhADQ7NmpyT3mevW2K/IGQ1oMerZB52g6+aQhCJViJ7Qw5SPf
bPTFgR0laHztlhDgm6/ao7n9y68M2qQwKCe6J0W9hLdhXmiYaqAMLqga+mg/mbSw
vRZfGOMRUFdS7izHs13rTw/sFV6rjM9L2B6DkrftVXi3GSzbWnyNtQquiI40ocRQ
10VeWtoeI07MPZGkXTaoXI8FtBUeMUHXHaMVtt88DlfTok4ALGC52f/O0j3wMbJv
4g++FAvqcrV/IjCchX+A0coN7PIX0i/trW42BrOsG5PtbptuktJ2O8VlAJKoGjL7
Du0oD8W+L87Io135yL+rxU+ett9ImKdYIH5UkDcbeus//SN4TO47kdv8hh48Vp65
zjGYGfvBjdBbCicX9raJ9C/eN9eexKrLebAmhC+uo83N+uaIQkHzYTzHD0stcuTX
n7hSjNCOKAEAg8v6UeSE4K9WyFIarVkTSg9Zbtaz5zd1iMfv7oxCrOrqOIJjL4vN
TFLy/iork2W8nT/3/blBS3DJ9fGX5yEMyGSrQggOu0MYhc7BkrdSsLv4TWO2F8RV
iRYu/LgFXyk0wzm7B6ADUwP6REXHUEQr2N+7dHkHJEvBTBUVkb3xEQfa+ykPDnTD
B88wFQaCq3ZhTR1i4kT3wqjOZtkLJL8f026HAp3xlJ3vPKRYzh3+PnBUPqC2CL6o
km+UiCj3MasAx7WnmwmB3ywyysWwf5JvkYBfxN6Fsrj3Jj+WqBUgMXdaIJO1gUHx
HX2jlmMAnEOG/qSr5EKNGvxNP9ayfjo25ZvF5w6NzR8/DRvy9RdR5yg1fw1FPbAV
UvpalKPF6QfErfjBo6OjKaLH5dwRN+3eLxpxxuP6H6gYLE7PPQiygkn7oEMvV/t8
blf2Q8zWD9QMtTHQZexjXnb3m9DL6d5AClWoL64qW+PjWtrDbaZqW+Jy4Hu+nNDj
bm+VTSVC5FsLJaqAljLcSd/4gjKReQNgEUDINxIghvguZafi9OPO+VerbCM9GtS3
G81BbeJPM+BI8xr/yywaoHlHXJv8EajqFcw33oT4xaYs1U3tWkMvHS/SNZ5vXtRZ
S1Fn+5IiQ63p4z+VLKI3TtKP891qyJehUqvwyQBhFogG4SMGyYhW0Mb/GmgOZi2w
GsEgmQ5GZfqrR7xuTOjg60nPI5qR6S/wzTLkgR6caPmYNeCSWG8k9YJ22thnDbEL
Wws7ZYXcLFc+7OcjHh3r42jiUCTSdX+Qa7dzK41teQeICh+DKyC/yBl7MTO9XXfp
iUt6HX3JsM6jYWciDOgbeZmbjGAHe7SV+/9/WeVvPimNvU/1/B6sciBr6rTzZiae
eTyosNHco/nKH2IvcvieMY98O9KTsS7rug9S2kBMGaQALSckOV9eTmlLBXE2NqiG
XouIV92O8IuRuka7uqH1ceuOuQd6EmnjRU5PQG/0q+l+y4zQX4P1XFMHpLrLAB3T
O/HIEoHsUjOy95HDB4Zo9dYQlh8UzytA7aDEMmvHOXEv/SNNYMc3CKNO8BQ+ocKI
YEWkgI/g4r+RoKOSNGiRP7KHzY5gHgofG3SV8f84YssG2aNFvrQt56lpqBANiEXj
WAaThULpgVJ4ZNDJRMtOs9ycXfjVaFjLTVKGxHay0X18p2wjlEGnVy8NJqq4YsWQ
xVlIIw4YRR2PLqaS5jLV4otkHJfSQ7eiujWP+QWKV30CybX//JavsqGQ+g6cJ0v5
0RTuXPe3kYD+PyyBwBz0i3HAnWzF1XQxd3Vu3yk8aEBPjl+n4IWHxtjzXJsGmhGm
/e3nj0StfAbe3kIiwjegLs96mOpysstqi1tcc+A07oDzPEYzfE7sG2TjJFJx/DSd
V2c98b8tF/ybN5rFTERGSsmoxP8c10tb/AKXZ0ME16uYNb55OC4KGMnPqf6040hG
YmXgOfcATWjhCilZ82K8VFB3PYYNi9vxsbOkT2fikHMeXyeCvUSmVUjPZE2X/tyt
wtokMd5bExyp0qIHUzbGVBwEGreyXuVZHPpwqs2ZdXIBVkOkIUboqUZXenYBY98E
14DLnJPpKnleMrsLVxbk1FLbRhxuwRcr4rDpOmgKNRHUfxEMWr4OExguE9tqy1eY
c+9MY01p60mJ67gp3a815Erq3/y+9ix+djDZ8OvMKNF7efrpCqlp6fsMvADGDMB0
QETUnX7UNd86rZ2g8KBANwN1VpxtJNyJYaaYp+0s5eVkMuyRcoWIASzDjNDlqbj+
oXB37QNfRubKB/6PSmWkyXysiIT4sCTc1Dss5B3fvP7pfTtrGX3Sk+X1kepQHJCs
ZhcEBlq9HFIBCB3fXzkDjNVO+F604vsRbDpNGJIhFUzDkLb6O9yPeU0wyIh4O4SD
nxJD6ghI0GTAOh2Z4SoZnMoZrLnGw0DElRO4mpJSqxdkWibjbtVOCeW/ieSr3Qit
G2evXUC9IT7XPvJIwJXpa4gVBXZY9yQK9sQ1mcPcur1t/huDPmxbwIw9UN4ZO/ao
aVkZi/IeKZyF32vfes4kqwVBdanI28fTOp6IHBWzdBzJVXkPcWOhXM8nGGfMgEGX
QwjoHRIiR7O00NF3oPk+MfLGu+HX5NFRMAB5eduMlFEMhWf7d6nBlhh0Kugf4R4C
tMyjG7tYbWHKrpnq+mhhUU4zW4zC+zJ14e0K3dnxahQJ1LgccsPUJfuLKGwja0qv
3Cu4Fh/lEm44Br+s4njJAT2BhmDrIaFz7ZDsdqnvYGUNiWdPC68ElxXivMtWQvM4
fSnYDzlUXyWJXYcqh90istuQkkc4ZfyWkJblJyHDlRvxt6GHhaMPEtUyoR6NT6Lt
cPAgfH4asABdlbJfPM3PThmL2FoJo7G90wQATf+NHPJo2Ze79qQIcHXgz3d/P7QW
S/zIdVhXSDx+R1erbi76D7bdPT8C5SyoQrOpluRL/y1iE58Yp/AiS//KSpxxHeXd
3XhxZluoMpcblZMj0a4eIN70dUGsXsGKPFwKVRPRaMWzdnsdqEqpEd+IcEZcLdyT
dAmX7JO/F1VAmuQX6QBCKFrwWUd/xYqPsMitdzX9UAJWeXpMf8Lizk2EJZ8Dlv8w
psUMhyh2j5Nyo//hTwxXA4yhkIQMYJwdpPZaqk/DdPYZ9H9JMX8J2cUALNKE+fyZ
Y8CzlRVIKNQtBEtzUj+MdujP3AcpM8KBAKURus9o2TSId9XeNbxIxQJWAl8ex+RC
kSyj8c/8Iftjnclb3QtUwDm24uKRgsi7O6D1uHLqI1fYPEVL5iTgOnUz6/qrNeHR
r177bgpIrr61tx5nY0wBDfOLzc9kM9Law1SnFpBw0bCCi9n2LgL/aKUa/GBWLWXq
kIGPgQG57lhRXAwghYK+QcXxmJTclFcyzgpCav1hkD270fvoMFguagNnjENp95WJ
gTg8HEsKH1OO6byq0ZjoNDDUsrbjZMMX+a3q/0XHHXQx4r1Zsyxth0eWxCZMpope
ArTFqLtBxqt394skp6GGn/ozcKNwSZB8ifLWNmLsa1XEx4qnaxTCnkF2QPOH5qqF
j5+jnbw0rZCQJFnlGGbOG8VIu0oEWI81/WaGR1lCTNqJzJdjCLzoM0Q4BqpfNZ4b
b0J1R9j6Qd32vLveyZMxEOdJ49q2NFSHO07MhY2mH52b7PExof7TQ6WPoVZ301Tl
4uuPjFqR/+LryyrKSQN4JZ7g3f3Vn9OtgUdrMngCmU5HWqTNQp4PkjYMUWNRY71/
E4rZlNgpu0jxpKfRQllLghpO7gOCJXP4V18g7lgbzJEe1cER8scLzB2r5DDqxH/S
rjNGQ0B1QPpGiPsDN22rd88PBk++On9zHtAfXGTooi7sCvXbuyDKOXooibr+vePf
LqTMaGBqDFDctO5Ihw335gF45ysuAbgl96CBkF4QOgdRnENgMhi7BG+kfqgSu2Bb
nezFg6dHcKDTbJPJPy3rDMAJoItXovoY2dQKlwNPMR9xFG09/d8AH49Mj4eSs16U
Krthls9ALfptjwAqHonb3l9gwyw1KsKHSb+O/BqIpbZimWftd8QiIYlHqWdTj/y3
bjihbYV90FdJMMwsYycJGongrwrad5oA5YL2Yx9SmfBCy7lNL0mrAVOLC71xEllM
ZEOaCiSKRNSrfkXVCM4XvjMRB5dq3QxubtJdzBSkkT4U4Q9gigTjrSYzXoOod5Ii
f3JWv9y1/gGwpYrPs0tEsklwBWD2oP5DWZE/umh1PdIEoP205eUJsamvLwbkpLfs
irCu8b2MFAlZwWGS62Uw6UxdPAX/VQIcSVm2pRMGj+41QeAFlAu6MtDIPWJNQP5z
JgfJmJfUnmBo8WMiY8wgcnWkdZpQwz8DZCwzb4+ak0C05IMuvjOZ/0IZdxk+Jn1j
1yZr5Sz/4EYUWIalSfzn33+/xKVZj0N0q5SLoO2vHTBbJTE1B2ipxg2gO0/Ptmvg
ALSWyeVSxoTR8rgSdElHjocMx6/FL5lud45gdeea8/+TgxXvfSxgAFwH7huKBpK5
TNTaQ6Q8sIMegG8ReIOman69vASKgjvs9Yx64+BZDW5BWk3npR916fgO6CYqlvTY
kOj77+YWbZ2xIDKJ0xmxPZt+Uq4g7k7sLhQipLGyIKTbYsiGnxSQNSU8LJ/UqulU
Xo9f/0auo4h09r5+FEYIn5ybWFMiLomc3b5OQL/J8Fg62I3N4Gp7eh6jgNYAkqHi
6RJqf+OJTitEbNdo5HJOsAlL1L8X4mmkOZFkV/+4dfRUNRfvhggtazOuf3QAbJ2W
gFL8vxEkhdz8piklNDGaWi6azGrgkxyh9I6kJTQ1zpyKwGol7mxP+KXf4kmq1/7I
qNquhXkZT/3oKbPUhXkgVExxe3uFld9QhoWwSrsLFQsTitZfc1w6V89h//m7y2E4
0ex2CKhcpx1WK+t/YXXDnuLnWLoeHw+W9iNzg2ZSV0pw59xqV6cJxjdOpzT8/lpL
QGM9MhvC3MjlXqyGd+ErbHEUJJQrVbwHOMYlVIDLSTG0gTnEWGruHIMF6IwxQX9q
hL7IPidldEO+S6ld9HKMLWEMc1R9nf6RLkoKt7WyDHZ1m9kDqjwb3M7SBEsgHEiU
QthpzThaKq93gm5/z6ze0OQ56njubgXSx0eqgHuQC0FWuwXpAytpJ0VemPMu6iJt
x5U33A3xwj7soo6UD+SRqSIbFK/NVCS8J1/PcoOW9k1BUfprVz5Pmi+/nnY0NZWl
FM76wBFjDl1Ayh86xMIUEEcJaUAr/dgPXOkOSbWb1/ix3/S0KBkWGpG2JuIV/dsy
OUyWZ2j111CMPvmdyITHtqqcKine2OYow/w1dLqDtiNjZ1/loQcgSJy8+ZOh3X/1
apIC9yO4DHvCyDH63LCTueN/7Ag6OeZ7QnXxu6VM+cIeugH+PuErFbk5krbdcAJm
iE+Ib97TTm3PRwlZjqDfpynwDowRvUB0iT+Pakr34Vcx3Z002P92o7Qo/X9QtONZ
fSblJe9DCK6tEvVHstJCIN/Ym8liYBgWoVaI94+qab1Kfdl7agstvk5mKoANdMXX
cDsI1Oms601zzV6E1IKhAdFyN2MpEBTh+giG2JL3Boyt3W9JMI5bTKtv7Y27A0O6
C/qIQUPFsrdvKd8iNk+Jh+jcdsBBVknFq6kWW1K1oOApdpEjRf+mZvSX3uHZYIwE
ErnVVfD/NBxkd33zEsdJclM4FbflJP5FKpLqXii8VCRa+uhUVYGlfATGssMI9F/a
dJmS5jcJjUKXxBUsxzRO/8Qbn2NZvB6sgLl2fwzBF53t6v8rrb14RDWAw0Dd7TTw
Uy4nqW94i7H6u5Uq2ba3IkpRiS/SP4ZwJso+qazkw1ST2hfWYlMrvmOzKvI379wW
E5olV0pat4ImUmD65FXf44qc7AD1fAc1mXYZKCsXo6+iHy9q5jseD149m8qbhH9P
nOkWPzbZ2WmG9Fo0Dbc4x5Q8gyOVymhlpDn5kSguF4UFQls4QdULLuk6Nx3gTWla
LKWx/CvtvlhlVA6d23YLerDbm2Ngk0e/U2ZL//YgamrkTNzdiuadTKxB5RqJRtBS
ZjRwuIws9U+IOHspcKNlRn91+zy3Fp3cscqaLbIj+023pKCgo/nswriHfmZSsWqx
v3kGkGsQJhpZqLKRCNuLwZ91tAgFH0yePoixkcx96CzXkL+eU62LoD/FDTGcdE+1
tynBbsoSLtuEyLuKs+dqLaNs40/k9yCyMuexUdagbi+mVn7rONwoDWP1OGfMj/Yk
3p9OmwQ51UXg5+ax+/SmZWGLw0iEwtB7yNvPEyue34pesq53twHcYpQMO4oGndtQ
GoH3fmCJ2mBWjfTE8rKKpaDXdgF2jvyipdEBZnw9n9pUJbBGXOJ98/aOCB1l+RYl
JGe3jdZSmtu/6o/Yd9gWwxNT4AtlQnyNQ12uDYD2ZWfoHmOezjpljw1332ZuFttG
m1P+44Cu9cYXGjnsiL//J3SiPuYMQKVllxuek5zsPl0Nutm5ygQo6an3Oe1EAEBs
kSkwczE7cmRKECHmnopda9Hz01Py7Kii/mVJckW7FyWjCe4OXYQEnJQQ7RHrYR/8
dcbzb6Q2uBZ862AmgQMewKHJ6AK5b7Y7I5FNdAnCnnepF/nev6kBNvbKN0hMSIMK
A3930TFVe9kJEr9U02GS2FAoHUgPwbjrfD+gIAAyIvmAQH1tVXhhr3fvCDPTYiGD
NeIGzjj9D5i/WzADWkPdZjdzd9htNz8WwZyJ17id+oB9XmtNJl/vNF/5QXDF721R
PTx9YRkRAvOUDhdHglIfndUOw1rx/2T4EzQ4rGiziqb/3nunwzXpupQ54v9pVtGF
vkhdzksYv+jdlmoBrW7JxT7r4wB/5qrmVhy9MxB8aEF0Qx3MhNDq0XfX/2qXnhD+
93Kyb2XQaC+DJkAuciJ9FNpEMqx4N81tUw8iNbnnHOPUjP2FL+rKcKQFxXhGFCUh
wbSZGCW5Vpe32HZAN5QQMcJczjCfQx6ExluI6WJP5m3Z02zspE6Nb/ys6PLtBJqq
LeosznCS9ja0gEUdRoP8PN/FJzVzRHH8e8S9RJOntAyqDy0JcEXc9p9wqRnoiMcE
fHVeaEGMJE5dS1Cb23+8PCfKnK8bsvYau/WV7Fuz6r2OrLTFYoGxwMUrUvETfH94
iQ+/ch+zKbAHCqNPUgoxevL1MiRF3/5PENKYKMFyTgUwDUqy5SqEFjJ4KRytLeEr
lpw9Zr8fsug45g+skt8ulnfFKfILZAWPtvmuoXqrizFeCJ6TNxL2dgGmuPr9QgE3
Oji+UaVJijdFCdttXgVvc14T/ZXXSoGruufXw4b5As3bPkpGcdlhcJyFALTFYImI
IvfPBHxB24OCLmAzch/FcMtvuFcGtW1iJMn0qhyZ3iInX/retBS2HCN1BqBzTYpx
QUjbAVzV6M9u8U0yhylzyZsy+xzUnPGEuXfQdQC6/xOnkLCQ64GfkHyNWnmNLo92
cTwDZkU+5AeC0o8FCr90c28i4lamko/+bKI+gsuqIZ4selKFbqK5qe6ZPj6WKTQH
9s1RXBleDFuy5qzHCILffO52wXyzcr88dQWyaFEct4riblT4BqIHMPAfG/TwYdNp
pdmucAiOm+ZoGUV1C2V2ftZv5WVwwYKwp3Jij01eWkqMCbcumfSAa6y67SyES/rs
ku/GrosfQrbzZE/4I3w2CWt2RjrA45mHquW2ZWdm87dfreLg4jFK/8sZ3YfWCy1V
6+KW3vxwVNj1HiHYqBeVeYZph7nsbsatIUxJSHkUqhPVY9aXYtgrTq971eUTJjgD
Z7westkQMVFHmzrr82gzqt3XOi6VHGutUTHMZmhBVEOPAhGbUqMg4WRwbqL1RyKP
jJVPdnJcIr1ZhR5sEem8JjhIPburolbEfKGQxRMeq2H8qxUtf6QYVJbgZzd85sMU
2jc4OPWhGEBazYSofiKD+iCi3QTNd9oYKx8FXkcvTV38pK8iVY8XLHH/1Gn6xwe4
lRbFvduBoISVMMUphf/D46dAKfNyuxmlPmyHBL3qo7RQa3mP3K9EuKpA/VtQYu6Q
XLYIQ+ZkEccPRGHLIURmtUKbyRV5/07RHssKngne7zvkOIygqiFRJt7BOtsVwdPk
gmELSmQbo7A1a2XSgu/nVnN7Cs5Ws8BQPgDQvuDXNORY9/NaD98ENjRNdQfGKe4R
2SRBPTO0GCEZ5dvrkuQEo3FCQtXeon+xnRwNvfg114lnhyamoEBSahl3C7DiGaKy
XciGIozB4i7vBJyGDhZXUP+1hqZ8clnL5vGqdWR9hp73HdX7jI3gJc/26C6m7JhF
3kfVVoeX7Nf9vGYJQgTJ4k10tVk/JGkdU8fLCD/5L8JRbU5WTE8EdHbeX5xOqjFG
FsU8+hyqDHrvyfioC62p/tqha2FdqaAM1WfLdGLA2fNFBcSCdE4TKiXb+RjiDaDp
ZJCGHpU/4OoPccqfseBzv0OP8QTNQh2b2f8DWuj+IWHtuv6HBrg+nDWzKCBMkGij
dza8/AcqDgzSYst/0qy5FkHTcfOA1K5bTsayiKrvkbHaoohkcmfcfh9Xx+Rd9JXN
zOGICORCQwF7WQiLbimDVaT3m3/5toMzN3Z/9QCGALcC4aicOImmf7NUTeiOAw6p
SV1y3iQpGrefReplWALnIECDAtf9pR479tpDA5Na1DpjyPYTidOmONwcm/eQ3dds
s1Si9aFFFHnxPcKHHSkvGDnc5ItdbSombyQN6/haQUx3/lPhc/wkOWzM74PRm7A4
nAVPsC/hVjvCBXnjiuPgQEA7xzLFo+c3AO+ZZaNVQEYAyWg6Cdr91eIMNPfC5c5V
nkj5arEEo6T8kuBw1OtCrfYtJJZ2dbr9gqRCC09Tcs7xvXzq+6kYyHRVYGgHrJ5y
2tvmsMpJRpS+2JXQQEDoM41vNJLRLUuJ53nKUNetXVqzDhMpujHeGQp3guS8k6Nd
7gj05Ao/WhEg3Bx7IJ548IsDyoE0egH98f25SMRCLJuXG76pye4TaNuJkulZUaFO
YEvsDS/hYtL9qhGttCw23EI7WSxze92LlW0Db0YBkHSq3YazDEwz7XIYueD4mIkJ
jeFU5N2vOAD+P3mBVHG3hHrUFQHVgspZe/dzUtH/CMRHb2C/0tIShxAIQL/zq3gd
zYeABrAieCX95caSkUoEBl5kmVsfcYqco0pgKdRgTi6hKbrx7zLsbGpsacXS39eZ
bijyYMFdgto1iVnEcfhpWG/uwS05uO6yAqTDip6Umf0cx1yTIMoJxaImZf0/2fMi
MrpQUQJUlficZQ+oTLiENBnWB2HvsWir5sgpXxHRwY5RByjMnGPjuZtD6cSfY/x6
30TSOMQga5uD+GTrMjkpJxOHm55u0YT/s/3PU0wwMUVGl2/UPRFW5OUg/Z98FAqq
ByuQeKbzvPqma3SmVAfPIUKg7CnEeX1fhxH2vohayWvibkFb75VVmkrvhhBgjTX+
J714LvWXj6PN4bKXJjAMoLkqAFV/cNCAnyNYdL9IXxNYym5yhoo1nbejxXIpobnX
nTncoB+0JwQGQ4ySJYuZdVQY58koJZDrQSzGYauyqm2+RiOKmF1ItcpSmXk2h2ag
nTHWOrQP12l5/M1mqV7dSXFWB/KqaFnZtzcd6/Th3hQZ8+h7aUOXFKKy/0gTZhdZ
8gm7BhL+B6PIj4BlBWu76QutetGxoCPNCC8PSTuQI44AGV9KD/QPaDzkE5PNTZhL
RZ2fDrw+ZzcLakJ4TL5zUuacMonMyLndClv8Mao7x8H0mnq66lxVgtXrV70gBOkx
p9yZnB7EIwHnRDm4tJ95WVnXJnVnJ8vuUEIEvDfgk38DQeIdXcIbuxawG1RTHjqm
PjhaDkV4CUE1ax/H1KluhyBl3bcpAhA6iMX0afMvkjvaLoBh6vQmDAKEfihiG9Lh
t+Ymt6oW+f1OJjxsEQyoB3uTVZ641HtT9DkmfWAj6D9k/yJvUD6FI5IEXSajURZL
OAD+yECJdQtWmjRDi2uBfNAokKKcIVbl50E4ipBXgNb8YlIX2Y4hJ81T5EjhlO+Y
9w+mZp5N8Vy9VWaGPPT11lddsz19Bd/aLzpjO60cieC00BQJpg5Ne4kkJgpVit6B
BBo5PaedTP5Qb7wKnh5Lbj1PXOcntovQxL+1FnCpwrWFv5+90Ggzr4qVHDM+gW6O
ai4z3teZwL2PNC955pEIsc4qlW9OTVNBUAeP8SOltfuTLBn4nJpcm3Phm1fbrGIY
f+vS575hbji59l/5gPfOo//bJopyXlYakxfcE+rcP1bQu2p6c8eYguKdPrU/AURi
STz4RSch5qoFzoE2h5XZvltS+gr+oGZ4kA8nDvivBaHCfjPZSAqmCS5qAodpmFM8
livkE6nEfMqKxpxUWe0kzc4zpuuhZWkGhXmO6nSARvu2tQa/M+1qUU86CVwOgnph
5iM41GWiqDuhM3idfvDKZWELfCfva46kkkykvnAgQrY4JsGQPE/dhszFp7kdDhCR
euGPrcQ2hx1544OiPgUXgvjytHghFa1o4V2j8ln8UNcyRYPatx8DWAjOhXScTr0z
3EV00kjF4KZX0stw8eFaNKHpkQH/eR3f++vPyuPgL8mrKoqHNf+g1A+G2kWZABWf
foBaFRxYddGVJs9vkFoivCqRutHtdtW3VfJ9D6DH9t9omNou+jfPbFCwA3x+IdnA
i88IDzybth3PbFrHZw5o3JoII7i9uo5BPvt5cxlI2vtwzcJef5G/dt4iQrU+dV+G
It6GqExe9tStw+DNMuXIOj9A75E/mgYY6xVR3EYZLuuRllaguF7XG/KMvH0YKnnT
/UyMECIUdbfU4UMeDN0EW3j4/Ipj7JRVFeTG8tjJQoD31Rv2iztwyfEfvTnldcFp
8yTkTNB8rXa5sjOZjDOWtotnmv3Ix3JVGXPpj+YvMY8KZaolKx/+73kmvm5EjURG
JUwsqT3PaGJ/NlGcPlXc8kNHeX5Csw10TbWGBMweoSmo1iz7dUEJs6GGYqlC4M9y
LDjoM8jjqSAIE8OMirIKG4Kv4wOY0Hv+ei8r82Fibq2KG4OgEa/1kH7615n1UDxt
Ud3R9WsQTGcf8ywCzhwfYk8Lq/TwrmYBC+yhX0pvaXVerkhFWCBLnIauyG/rYGXE
MorjRYl+/mSg56YFWQyXvDIEL/9VX8/X7W/3kszUbT+hBNUM8rxr7kSZPavcWIys
B03MJZL6Vu4WhnMnrq2yTeMh1KOGlb15uyoHwhVz3TXWvedHNn1d+QwrelvFxSPZ
DO9Y8EhHxBWffZxPn2/UIrH4/CmdNzCMNAEOLLrg5NLe2Z8bUOui6kyZmPEiDT8z
2qGZ21Y6NoySDgN8ESIXDT1l4NYTQhHaFFH/y5S2a0ZQH2qB4hoWwAmbOpkoGASg
EX1+GkhOPblpDlBURQQgk9jevrQNGsPP7DSjLnwoKvHFq8Tzy0iCyoVj4uouywS2
MbW5ybWnT1rFYU4oC8zCZ157vvPUGTWh9TJ0jQNxdtT+lejO4bOVT2Kzu6UQQz94
DgM2WItYOY0iOKqbPK7YvYShn4DOsHUPQlkw/jiLXKlrnJoNIiI7+FwFZniFPrjD
nx7R6MckRS1sT1OJcbsJ02tbRtH6+W38bcLCCdT6TzhJlQkORDStY4l7jFpnX9rm
Ak3MJqb1vycNW6oL3BnHBZcBdMzG5iuevBh3U9IB10o8M06IeK3geboVTQVKT8jM
g2HMCFcJPs60QvvKVJyOhssVIFACZEGcBGBuWuh7lj1mN6gCmtdAXiIL+lWTjtT5
TCGbfCivAtR88E6InpWWF3kTZ/tBudPSA3UtLA+ngd2nCA6/TYl2lZukv5nnbnBt
lX64K8eyro7uSvyT2byM48AhbP8Cq5dMXUis+TMQwRScxEWDtK+k+fYckuPy9wvH
vXpNk00hnyE6Sl+k1fHd9jr/ta6rR7OYdE6IpvDhMvGWHNDYO2hyeRGEIZc/tJG1
tHv6XC3tLWIpxdEI1SfMExJCt00QlCHCtWi/0+aRtnJY+ZVVfh7spVseLIXlprJM
Gb2R4C7jDe9/jzLxKkEaGr6gpkVkotnK16QANUOoSrzhoFVreDeIB3FFwk2dc31X
O9C3co64tZsfS7qL6rluHRT3KELXV0WdU8EakknstvD9997vKFnLU4a+bSBrlSyq
lY0lLpgxlWlQdYB21TUtwhFCuzoppcIT3BcS9o1j3U3thoQ/SHZQVyGz2n/wOD8O
os5p100VOU4bmyxBHTvg+mveeNVPwPYQS/+tFk1BkA63cCb/sbyDBaB78TtZ/AXM
FssGeyCxpJtwK4RNI5Aehbhvx+2xM3wSrVkLH/7H8O7RrbpKuwzeULNT5Gk0yIgx
kSDU48EMsbY8iPlEjEq57/K5k/vR8a+jnss04mFW1lnCzsZ4uqEg9q6TaepFLewh
8EXlMA32sql+LqHK/gz6q1nXKLXIDQTBg19qdh+AxGyfIkirt8wbynHCAcoWPW7p
Z1y22GcldX5yz22dJHZyf49mHxvLpgTo/uV0gt/UKMhD/1KKcYv8bglWoPo3KEqG
/IJWLc/gjj/bRN0tc8OHF8As1sYINM9mgB+kBKvmp4o1IUpnihSYSx5sVnG2kUDh
YrWHhNvDvth3JCuMwGe8dM8g4LwzV0jhO04gjmX2MD0N8NDelmteX85aUAYP3iTR
uIa2RUlbZcOxj7AkHvFWgGjBXTcZRjX9iuCjmKRD1+uV83VdKetgmMnOUw9+jh7N
B8NQoFq5lmkUBdJWJU6kex+EsBeNVat+CEwu/CKYTH2VALzk5NNSE34UNVebyH0/
Dkt89jggumGOoVj/yiUGqwEzyUZmTLgZ3uYeKtp9MfiffcHhuZXVnWPaUiFl05F4
gKumC5HPcJ12MzYAdB4gmvl9jpX1dhHV3q6t/vF1lkBJYCgpo2dPCrxikR14cxw5
iGibXZeA9dhXAp+PzCq5naJbSiViQ2I7V5K0xxwaMtOA9CUbtA9IDjrAjU8xx5Ov
/iSyt6ck9ttoU8wQPY7NWnjR0RDaBA0nTZZTGkYthLUdncxXeuJYLG8h+loIZCuR
nOzijxMKqDxcUQd+lxfv5dpOfpoWUSH/pkrSkK5+E62yVZlbJAFvFF0X91PH99yM
vmk4Nrs3zBM46Dz9BTuuxhyP3Omg+OTETIaoOHklR9S/XFDxn0nWQyG/cUwtiZgH
K8kqXKWRVVBK7myWyJRhG18qf4zCPgVopzJQ/PzIdGggOEANIGFfNO12pq23OFFi
90x6pZYUFYZmKvuVrVEHzVhN9EGiUKNdsmx2zx/Kc87khAj+O/rf3WIjilH8ceb3
4NYBxoWhpwVD8C54je8x4QRiqGtuZ2ZqBr/5FyrP8qmrCDMekXNqbv9j2MBYDgLp
TsIXwMyvYl+e+2Ed4Ig2b2IJiP51uxkTeUskW/lqhs2uSilG2P7AHuBriZQDIxSh
yrW7FWHQwEsMnWoj0pFXHUO69bp9B4vSTnodh/7PZhanz/qhYBwbA2I5YoUSugm9
1lUrwh8+1WC3eEMloeEPCVPj7UMo/zj1uJE6/I9QACqCFK0wqy2NDhnbY44CEjpt
90dbxo5uZY42zDrf7Nj96tubjn2qZnRzdHOXNn4BIc6Bb6KlwYKLOHHgrx24ZRxI
Mf7vJqyPD27qawjmg9cJIyDC9syA2AFitrVDj3TQgP73oZfg3YOHjg9WrLE00dZu
nI0R2X0/xgI1FFW4BcYCteQhH6KLqol0gllUGivRxT/Z+H0CGDD7quOyPXtivwrW
caey4T8tWbMly0ZDcbJlXQHK0TfBBbeXkq4VjsUWR7A/euAJMkCL2+pqjxMVLI6Q
gF+CQSeNAT8+spjptkiso3r6sO1dE9O33a4BIo1vDp+e1tPKTD8xPiuocyxHEbgm
I9pTCJqYGtkqMw/itcGrNobjIiiccTMtcCqQwKBJSIGBKYtvnxfzPQFLB4DtlLn3
rmwon3QylCJ4O/uA8resXASVlJ6MEf8jKAB8bM3+ktNmzkX5ox3jS+5RA9f7PHuk
31tJKJzy5Q81v3d+ajxtgy2C0rLOWwtMV7zZgfUHcCQ+/d/p9/c15Fx5FPnHwt6g
WARiEfF3w9h+NzgjydNALPBq6FEVciUlFMMvq/4d1M3hxjFcTSi66PdX+2wsff2W
UPNAN1Oa1yhtghWJFuJG5HxtDUWlzj6DeeD9ZgeISkBM1Q8CN/XLzoFCf5VvYy36
KisHIcZCM3b7tDi2IVQNcBPsLFrtZXe03g/14N6WGAdeT95Bjh5jXqa3Kk5xWgrf
LbUKbTTXFfIe3pRRmdgRHpZnSuY9mNmglRdnmtzmnAoxZ73mL0rF163OoLf/sVnm
NRXVnrrb9oi5taVhM4kksiuwq9UxOR5YAQ5ED3CEyLywruevsOWpi+XzuC1OoMYn
TWG4T8eUZXPcC3X/AcPNIOoCb4n+KGBCKTUubn8lKz4LV/NninjCZYKVFVUFTf+f
MkOQpF4I0bVzamOV5eQhkPTcfRMvx8rX4ArD7Amu0n+0+s7ZZYyKWP6wsr5PekJh
J+/uFnZuT3hQOi0iFm8GsktwDAxqK8qHaUsX8ksDapIJdwY8F1jQ1Eu+acjY2qHz
C4/UEhZfJH365Y7IQVjpwrBDLXgs0quqeMZY07+wyy2UkjfzQc1kVoJMzaQ1xDPW
zjqBN4uS+Gf+xSyovb+DlGaZ3eLxQJVLMEPjrJ7XKrLeTmDp7CjfhjZ5scFxHW+O
L5YZ9VwI4b7bJgldiYu8Q+xn/Qf0NUbCnm8gi+mfpB/Z5nadItBJnORaJhlOEfMp
Sfo4nqvfL0wn8WOuPix/QeoMdEPh23loPUGKsICO8ZoimvqbERFehy3J3R6bXErS
3CAzmTnUFNl6l6o0l9AoHoW8AhrBvTAHgL+zoyPYhO/9qqVJRRQJvBdfDj+2pGPC
hMsyI3dCD7B4qH8qqXdbo66qbbT3LllEIR04jKN2StQdPy8VJUP50kmwf5ZCg+wn
LfIKIervCpTtz7Us3Hb4NuOfTNhuva6vb3HMS6yFybOcsZcxFYxMEVw42Mii4lhH
MARncinfzQNiikXfCAN1phCmN6vrpdFoGdu3NrPsfPkjUc/otaJ0vWaudfGV1NKa
4wvHIcvtFKtyUqkpCooismZySs+IkSQnIXBjOAbsoxHn7ZHfljryF+fG2PG9W1pM
zTvlZ7uxCMJyhGGscPxd8enct6c+GPqNoCcKCdk2YlwiGeitwZzUkKmnL0kgwl3W
xZWcBL7YKjAwYO2s8JynHRPPc4G0KapIEclut0ZGqBSp0Pn2UnHYH1n2kRRjt+IV
PFZ0Xbyfec3Nes189E+k3oRNJOCR63zk2Yy349BriKE3Edh1qLpjwRnc2dnOsN0l
hMwTXBAhXXPoJBDhGrtp9M0MsWbiGpQmejv7qDjvuOnK6DKuqlWS2HD+BLnGGp1l
9+J+uHnnLqGujZj5ehpvWcB7qt/D+e+D7Xc4bnMEm2mSdteprG3WDDCXKmJIwTkq
WTGQsDgcMr30+cNVCjX4VJXi7I0i0sNgUqsL6g7q73asSrPoIbHtGVw7p6afPCgc
9AQz4ZfRaL98YYhB2sTjUa7Mz4dYw5cQpyk5M0HSMQ3CVYc6BpNzfqDJ6S9l8CzL
6dMPs5MeGw2mzyxy7TaJi+0/6u+7oU1HPJDlfaS06zi9o4wsfrpTt0LAHE/GSplM
yeWkGXqDgy+S13NBc5J4LBWd2NQnfRgrINTpL0wVrXS+reiil9ry0hlJ5eonUaca
1oSqq/OJSlfdQj4huOVpYqWTgtl4hBqHDgw6Wbx66FGI8E+tcahCRb91abAeCtfm
ySUgJF1Btwl7gU8jzVr0j/0A1XRvhYe/nCTDhk78GzUxNYHH3NhvIK88/NF4tOJw
TV4KctR+PILxkSZl/Zah9yWCD/Ob98ff+ST4Ktoi5hqWvLbc7M4DQ2xMZXXA9yDJ
RErWbj5zMQQ/lIj3W9g+tHX6pfqEpOWPRAhBMtQmfbp6Lms8Y2pdSPENqYV96Cqw
OofDtO6O7uH3mXLadiBnw0dBR3hnPrREkBCcsXlaZMDrFv+Z1L11ZQXOI2byIPLD
qDgOt+4kPm0FfKU1zi3qfaRK8xYuNcuuxqigE1ofOZoxs5XHBrwL30i8O0AOR45W
mSVNE2jyCyV9qIxy37wpx3S6+p04d2B3vLr47zSMFbWZIe/GtESm4V+qcTu65pBl
rXceXEaOhPXi20INeZ2GYSIjjyqMtiXSnSbSQ4ORM1h2mNZPPQFeitBkPFgh90k5
7CDvyU5WVC689V/hvCYGlJtQscfvKr6wMDxnZsBoOHI6EeoKlAJ9t6kBPYyjlb0T
EXJAc860u1qY8Zx+OQtY/g9zuMw+S7APF7ciuf8FPTDs12ReRGF/ZRaQbgX9Tw3W
V6h7z73t0OkHeF6gVb4nIojT4FxNMD5LgundUdVIuv3oWUHvkFs+gW79pajxNhP0
wAtXTmj4PPaYIkzDoJJWLoBmzwCrhKoCPK9Bc0smdoss7Y1na5QbjSUV6USvweuH
llc600t23EHcuNilaGNmHpzOS/MJ/sztwmr8LIgwvKlcNhEdMyUfcUcD5Y9jDk7J
fiWB9iVKW5S9xuvgsEVIqOn3sQEPvFwK2DJqxNzfAR6077z8pH1HyzhdGQNrm+Z6
CgafBPtPatuulOHHYOAPLbw6zKie5Z9oiE69keklzm8V7jr0XL5Imq2MjI7KgSJi
KpMC+RjUErm146EyApkY8HntmlcUg8BWhNZiKAjoJ3Tc7HM7pzJKrvV3mbtk86tc
3Lzd25pAkHKnLuX4dsYj87X8yBqPMKOqjrJJgaecDPiW6dc3l082fMM6LMv+n5aq
4d7iGPmwW6Eq+V0mnHwDkl3va8S4s0CqK2X2eNPnpUEZ5E+HMsU7dwl2nobnPUvi
KfLzAJh+EmrFxXryn2v5IR799uA0vdiOuvzb52ee/hqb+W90KgkpQKFF/55yMZFL
pp2X+fqH36dMe5qsQq879Ja8wo7vK5p3Xe54Hwnauej+K+MEAiK8GmYz6F4hblwi
F7AOU39tJ+6jYR3rV+Bl/xXF/B8j5Y1lzSs+O0dFB4jVKkkf4FO825RDfhOhw358
g4lzTTCxYqSCIVM5oZmBp/ukEbGqL9BhNIwJyRKVcjVn2++Pz0T+jpVebJp7kyJz
poyef8af7u3saSKjZj+f3/05sJskW8mpZkb8xVh6cxEFCK/LqEGGmnWKu4UNc1/p
1dr47da0fnTugKjzh5NeVTRt6YMfCp8nVY9/S1pSAyk5TD6Kt1Lg7BB1H5bOoA+X
qBLxAR+AvkjB1etjn18njRxfSi8RZdCj2JK+V+g1Zi5UxgSTuPARbWssDP5DVnaz
XRj6aSLkAWaFizt7AYybbI6Geq8KKOUlP6ChutR2ndzDmyQQR7BozVcF221GURsr
OWBs29e9FoVoSPDdECZQli4uaZvi/vN5FjKhRLiM7PhYSWDxlgKkLQAUJ3RwzL0G
kTYJbBKZoYMCt+ZNMM2Z1DED92QDLZhJ36YFkEX65ytxSybSIg3LTdZSkUmwLqt0
qhGU9UeVFVzeJrPahjWwLUfdNtLFvCEFHhmT9y8jBUuBPbkkAP9tBCAhdID2noHT
dUoQIRjqgCexgnI/xeg7Y6+UW6kvphnelnIutSnrCI1iZKW49DebrwzXwntsnirW
eoLFDM78amDkTbX3H48UPmiPyC6G3HQ1u+XHYGqPOEJ3FtI2fHjDkiXBhLum0ygB
5u1rqYzoxk5RCQFu9MxESVlgQU6Mgwptxyx/oJAgd44ulXzjJfk/5Kex0cdtafJO
LJHVBV66vzs3xAtott0M3BJXeXYm0Afba2wx4f9fbj/7UuVuA7k38mFrnqtaneJE
f1z2gjU+ODlN+bykOCui3X8KjXGg/BhyhFgL4ILMrVUzQvD8P5jTHLB8MW3J7Z2f
aZZf4dw+GL9y3zllBgiMNGhCbTz14Cq437MrfO2AqPqP5AlsIBOtYNmBiWRNxnLl
mVGIPVzyCEcum6efbVkf3Mx2xpHXL+HS5cAkhdh5p1A7okFVkgnzwWBHsr23BRe7
q9wRYoqCmPdTKfRHRVL5JemSUMKG08c6Fh/vGmG34ePXP8tbqwv8ByZI0aDaLDk1
eL5wOEq2qjh9oaKrWOVkVJKk2pSrdthvSR0FengEHG5U0zwG5Tc5v7xxBkQatCMY
dmz9R9fFbOBh4baQw8ldBD1cl65ssbRobiTt/5gaEn0NDviZ0fE74h9+z7LyLOGH
qAuo7e2tJWpLeQR3nH0j2ur1wK+XWEfK5NPq+Qb8yJt2IMxqFHj0cxyUDW+IShAW
00lWFpHOEvmQZntho0mdo6+523iK0AwGTcNIGf4cwB4G8j3frV448U692+B8jwIW
AbJh5weSYCmakLvs4bz+0MXkuFPxl6QiFccNWBoY6Ix86vA/cUUyt+dhmBMA9VzB
cmF3YiVMu8d88887Oh3GGOZiI2mKhgBbHU9nVd2HTHBPJqfS9xpl+Yljwd/kPJbQ
Nq4EV1861pnrKQOIXJTcplBQsX79yX9Tna7b6pAnr51UwsqYay5/oEpgldnjK84n
48aPM7bP51tafaMQ+SOb24updHfGXzRA1mkCGR2TeSUEVHS8nJemAnmaTivGzaOx
Y3yiGitN8vk0U7a2y1MjOA6Pk/GCkgfERM3oRJ+uG5CrCJFS+jkC0DAMUW3Q4Mow
wU+QACEB1VO+AERiepg/VuNZrJAkEcYjTEOxnCcixJtIeohAwkl/J/kUUNAzlWd2
Lje8m62q/OgKMMSSYSqjENZXuXa2c8p6QXoPXOyel73Q7vPk9fMYoUemMQLjNwvn
RVSi/WHacP1pIbW7FSKJu5hsonmq0PUWiza8imh8rEik1ZNfXdz7A+pKuzZYfMpU
Zw28jPcsMHVX74bVMZxp87Aaru+SAXGrvVAbXUV3hJ0APk8HAgYXqlYIrlopVREV
jwFI3M02EvN0/5JdB1+M4VrBxnMfJKRVY6VrvII4VJjFAFVlntRfH5p4OT3oiK51
2psCIkCWk/hU0BN7q90lFXnoFtQ3PUzVDw0Y1CikP4tg7NnHepms3IYcVMJB5c+8
7s8+dttbP507vWmYBkH1FixnbMez63agF6CN796Q+e5EN9g5zAVj9bP51bHByKja
RZLm/hxgEJqQpBppI//TNzgZCButYjsuzpsrrnO2RnRuxV4lhH4Tlh3GrKAmZJbv
e6BbaPt3v1FZ7WXG3ieYOh1w62m0Hf9J+j2E+KiwIeJpli5+ZeTHiV/ZXeG+gtfx
vN4Cehun/2CnGCCRS81qfEVqBV/FEf4RL5iFtLz5A4BJR7DZneecGgsASw2v8pJC
Ht5brRBtfzd9PT6BGQqubrzZQDpOvzx9vF+1ffhHI1yBNEDlPiUR2eBTy4knR/6E
5WJ2JvbSZXC1owIRqHDa5DhTEaTWKTHIb0bKmdqbuV3+ltdcDl0KeiEgLjTLpKI5
/pFq3Mk+rfu9uoxA0mH+BZJqBGccv5eYCXjk9QWpLpJfATTJsOavp367AZNT3kq9
RLKPWUOjARmfl9nXVXUHkWZRziwsemp3byP+uS3Lko3OJmJMI8CP/TAFuzgbTrOV
c53htf1tVZH/YBUpVj9pij2ABg0BJmjjuwhsunQODH1VVowBa76pgtWuTdZR3u8m
eNvKbiqgatbZHUygzOAtlTcdAQA/eaYsekhcSSjHuRHWjCqflH1i5clyr5j8QLk4
tNcVIQa4Tl/g8cRNV3gJx5OdO9XTTO+Jb0VUK3+zquAObvPpUp1pkgCcz3m56gtc
TZdIa5g/gNQScG8NSGtPZS0MiaRgLw6GtCtPYQHhJ2A1qC9AgKWDZZEkHqTNPD2e
4AqVEBhP/hOncLj7siFd6cQZh8003Yfps7jJ7TAgSXFj7wrKrd1OGhg6szJPcGU3
e8+++EDRYsPd1aD+tbdDGpXVEF29BGa5QGHWKAAxNO9lWsPtsfjKgr+De7rEwggb
IHwZrz826K3yG3nuvc3z1ASdrJMJDBNNKVDM1ACCs2aoVDB7Cfof3MSJ2qHVeCMK
oH1BkuAgtPVTI7jcQgVhxxc8bWM9caIpKM0R959UKHtsH9uMSJIINCRFFj4dbMiT
7qF6T8M0CwHi9u9jPKCBWIARWZYPXWydbB+Lh6nWUFbw26R/M5T+WjUXOWSTSL3E
Vghsj/zcLzGBgd3ofYfHiSrmvp5NeLw77ycAkKTIGJ8WQxZE3h08sksDaraAIeLi
UhcoFlY0EdwKDLWdbEAjmJbxQtiWXqAhPg5zqc2C4deFvg6TrwleTSa0NzACfjxK
gc0Fi+rdnEeOsLgmkte/8gHxaFaX5mjqbOrvTcKxCBH1qlxMsSCplXWsxlPgpwvm
G+YAA7p2nJfvmYXMQqhByg5vhDd++qoewcDr4ZVSvlAAX3H8JRiH8rbTu1f4BAQu
S1rhoEGaXGzWUhDnvo+Ed8A0vKvokSjEM1RMJQQoUIIrUL2ay9Ek4JGbDodZlrIS
y5bAqjU5KUW16cBKrpSWRdj8MLefb/nceqDBW6ObMIMXspoa62vNCzasaLT9880y
yW/+AwDDGhVyY8O1w55bf2uzd0xeijuuWQBz9mpwyVPpsYTRugk75Wsm4Nl68BFF
l0IaAKSph80V2tnk99yQSb4kL2AhFNMr+DajpVYiBDplnM+ZuEoCQa/1PLmpDgRG
BUSRuTnStcjc2cH0mb2P+HXQQjm8eU9tzg4fmtxeM28lufF9SIdUaKMu3LhTv8WX
+UAcDpmdWMhxYvZSQISF6xsfyjxXZlk0fQa5HN9dzQTYlqD5boKRWPv9tFeTJMp2
TEEhTWku+xj2ZcLIIPv3FJy6vZvFRgnWSZUxos7sVeGD24pDWKh3d/zd+FMylFec
z+tbrnPSdPW9emYWu1Q9LwbXIGY74dZZLAtJBiCzk6P0dwN+Ecb4ifieYJuonDUo
fgEvpVp9ahZZsSQ7jS+OvKhEmHU3cqyrdIghrRiH5kG9ckbqdSS4XpnbK9XDC6+E
QFG5Ecm1teS50h7vWAEdTDzsA4U6e78gAH2Jp1kQnPvQ3g0S/h1XtjKExjMgX832
7Md5mhdGwS6hl7xueLXiIpDzBAPDkRhuA2ebsuRHo5Q3lBa4ht1RBFgwnrXuxqwA
NTeE842cH5gBcmj4CCQ6Odx98qowDje2eEJFXNU6rsjoNZN9Vlp/y9/z5iyleClB
WsiqsRrmuvxt2c23GHvxwaaN5Q2vi8qSDDRijM3Ekv8nnhAnpHGk4Qfuh2ui1vJM
NLvgp8O9co6/My/POYH884JWrN2kqlsEP+2jFzxlrjHxqYBr0aYzvBvVOhkgDBfd
Cy+v0IhwkxAFuMZSFvQqYUoFPABmUHkIWLiZfC/nuVAyWsgvrvbV52aFMTTvgfdU
7zpVRxagxAcfmcuz3TP+LzQ0g3amaFvM6rJXC1LNJWvgniSi0amOCuX4rl6Cx42J
Dvx6NMAfwVpRqQEop+4AMWZhNfTxTQxE8NSQ4rdAwgnfjVY1vl4uEtVd3eTfoNxa
R5JUuIeh5iQAPEHRTsE+ItwF8zO1XGZ5IQ0+aZufpjjB9A8Y48+jTnYAGbk+bnTv
IvnMxbpLfhYUKi6iNcL3Qru89Gf8S3+UoZfCjwMw3aaw+L6SFZQUr3XdzoW0UyOl
RXlEUm5WzMbOTN7wtKtGyTzC0QatXKnT0rU6JDdXE2TT9Q3V3VeeB1WZ+TyZ0rRF
WmZSO9N3K7DETYcUlbgoqRzM6OlYw7q7/O7TgLj4UG/957UhhfmOIDiEvGj8yU0J
9k08Jgz8hPcIgmiSPlol/mmZgVGOtECGOF0JXFapXIhfyRPc2yVlo0ndspFVzgKz
yYkMhrY0q4P+M+0XZPv5Vu2Y4CbCPTe2uXBsLftaCwiup6KP0USYQwNW189igZFq
0e9nXuGMBS5y5nNInUYvEn/GKsxRDtuCPDAMX5JOhGyVCCCDDjN5mAM+vynzmce1
dRm4+iAJrwgeWlhm2NKASxjheejb5OAX5ESciQKa006ahBf8fsJ9pVpPREUkb4hF
QQKC8FI7bVCWKq6qWX1QhDOkO+FZbBZ+FT+UtKdjg0MKhRvsQxHVbrsRsktXPDaR
K9jNWi8HUHEGuf+WEd+5CNRYCgnc73f1Nz6v1N1/31Q8deWsovKp7YqBvop7WK+d
PBqYq60NgW+8F3MybpE/5bDDVzjRGT+6oRYJT39YpGOJ3U9fY4TVJ1vPZVFSqlof
v7otTX9kJyYCH2MlsECeXz2MBoCOqyjyfV+y5OvCFom6/x3mtnO7P/FuGpuF4oQY
Clt1HID4pxDPWP//pPHgkDpvS3FB7QCpRqnbQKT2hOOPNopjXGPUIE1bHt5DzwI3
CeMQvdkACVI+wsatENPWed1MhGi66Fw7IcG8+wrQW6SSAsT64CiKWqNMzGsF101D
WGOtL46f59vcBSFxWl7quDv3zjr9AEHAPfCtXPZyoQNlKTUY+Hs/dY5stnQC+KUt
ySxzZLA1J0JtVgc3sPbKy5dfq92hwdLHFCIR1S4F0Jg4JdaZbWcmPd660OkGyqxF
URH8NaNKfzf8jstXTD5YKZS9gsZaRHNWDRbUU/wOPnGaUJTjPpyFtD2JNbnI7UEQ
5nWEmjegq2zOOrKyVqkpwtxYdWBaI4deNa0W+g4jpKGYJiLQhJEcF7ofSDk9e17s
Ji/uGZZKmXRSRb3nIiMhS8BHDzTumyUOo2QdKoBnuMH5poA6P8MyTRayyBZu8Hvo
w4i+fdjbgtSRy9bM/qsnAKEMdDgHw57SfoeuEAYsZOa5hpjYoYmxnlXDSo/pqjnm
GtDiAgjzvZJjtTJQMapv1BCrkNDVBLdoUJdLt0xR499KILFnrM3IsHVxNgju69Av
vWI/fDkW0NRHD7q2LSg/PJM3e21E1tgBsrxeKIEJwGqwjQkNPZ9JEVOQXKN6xkA0
IGTVKCkwb5vV6y0Ggg7s4eiNWoSVCLkB5E1jgfP0RRJ1XXRHqblWllLeUXUNOd0b
//9TraWLGloGClChZW/MDBwUDUluDqCMo/U72tihuMrGKU4Mg4IwbNu0M+AbPqQ/
S3z+iD2ylXdwh0nEO1HXjZ9ynpQQGVJ2STGvMSIks8FQW7GHRWKYT4cyxKjz5Wfj
W2N5u6ITcGdVma5Fe4yssRNI+jU+bhPrQl8k7xST9N8K02ktS9xKGdEgGenhNHZP
HOFAbs4O2vDWgISdAApFc/HhtYkWitRsZL0PhB+fQobTx/WThEB8GS6QDgNDVAfg
ttC0dgTKKuO1pzhGltmWSJpgozGfv/QzbRK9V19Micj7HK5Ir8MHoReWo9O+Uoei
3e+jA5EOPsdJUE+cNzX8etRVB9A5MuXzH8tquB95BaX1CrC2FxZKWjQcekJClTcP
lhwzbnDk9GGX8ShURSg7WcvAuc3gNLI9rN9wNQh0hcEVuyf869UlgKfLG4ii8MXV
rACqRK7a1SP4GuzNVPrHepfRLdqtGD/hwYXOUDEOUer97eVuACMz14axfSz2qbrr
l05hOKMjlgNkNJ6wigc19IgbhUxgCUXfQFxcSo9DyyW0tPHTVApXes95zkYLryxT
KvmgqMY4viAc5Ui7kbKRcf6FxrPOSKX0Wte7hukb0TnTztNdQoWkpZ9sAq1CSBIN
+H1ZCAHzvsS7OtF7+hqhCmDSsZ3ZEo70VZoZJ3NMwBnQ2qOylfS3s9tJCq+EfvUw
Z69ao94L4YWFeFMNm96tKA5Bpjz7DA2pwaiXWAGweDTh74L21t16xqKbVEwfgTcN
h3JqEx7FrBKCugWSl0hZcRHtxVNPrVx2w1I4mEFl7e7pMVYSHoshzvNfUCgjolXw
1Sz7+/lUGZCzzOSpNY0M7K4A2K5nTiiHCNi1xXG23Tq3dZfq8ISy1I5x3Sp99V/x
YCnwEkR9qD2mI1AAozfnAIXfWjfur3gT7/RMco8AdDFLGgxtmGg2qAO2BTOHThCv
INbyNt4ALqdRZO++K6/EhIy4gFX8L8RL59rJITPSTJnmLQc6fLxL840DkIf9w610
7yNndGkvsmREtU3iJ1Rbzpuu/Qco6jzeSC+UMh14GdQ/Nd/gQm8z9mlwTZ0H7AYA
0L4bhvbkSflc60uCUKGg7TfdfFlBAbIflYsXhQQvn98zv9LU+qaXqndD/mdCzSOH
HrmrEx1S7pUNCC0AHoQpePUE63t6c52ufzvogi21JdM2AW5CrOj0Hj5JSAsF1xd4
yFZjNvG6uPW+N8AzB73fSYtAKw1GqGULr07dqk/Efsr3U2C9ZrLJm1hU37LQbuhe
EgeUlpGxiUU/OgDkpU7+jwtZ85Ndn3uNNYcH9Ot3A5qiOBWFep1gCZaXYu2yQCc/
nSeHGhv/TG1wkNU6j2Cuc2m20oyqExLK3L17qCwP9CRK1uauTjLCT7zkCJB3ElEl
85RWh2DK7FgNz8G59lriIT4cjwfpwcw/QKBDVZPpNq2RB3CIpkq6Ixw6vTqF2Fy6
Mbx4iCMJ/uc3gzZD/vl2a/nBMS4u5kO3Srd3C16t6+ousRv98X6NzOovti8m65bf
7lzeBpiycdKNSXNUBDOcVe0Rm8EIAVwTx9TSIW4cbPKN03DPSoR/BWeZ75opEGtM
bJqPmEG03rI7XdqmyCDfAyYyCEayRaLwsMm1OPAp4RA3yQePwEwaomij292pt64A
Tk3nPnqOUgjAcjsi0yGjM9WolGasSRHYzIzuG4CykH25KtyydztpXz5cc8iAhTqe
psdqG1nuT/cuhi69JoU8WDKwFh2ta1Y9siL4e1SQmmeQ5yj4yig7M7Ysb5fGXrtu
hpaq6z0miDv0K/b56V1AfqnvAyRWrf19VNwCYmlXLM0W0LQVK+IIWLKGu6PJfLDd
5VFFlq5s8obWxC79gdMsQufUtbAuMIt8+YzCrPrZjyvzJnGJDTU84UvJZMtfEC/9
W0K3vSgXt/dcNuuhvR/IEo7CVis0U2pk8FG1YsSc8Vk8EOosEW2NM3p/73NAj0h/
ZsgSanSIWpNwiPtDBoVGGv6jS5KOWQjwQfW8jDv2jFMgBc8OJ5OIoEdqftfZnmVL
VvtPbSe95NkFOQ59mnysZ7vPASJRi4VDFYyY5gULzTQZpk8RkByOFZVgPlt0ppsg
nCxvxSqmbA3PmzTH8FSQp6BIGPmfke02HT6aaZoedXzw7QrTXXaNEBRfnC+yAjsK
OesGXsUF/sTKI2EJKKHcdkXdxB/lIwEFL7+66TgqYGcD7/1s/J1yiMX5EadP+05W
e7YNbBXmC39wbWZlZpz/bIzuDDb/vhPAVbuQLK9ADtnkjlWcHvVvABIZ0P2EIcQD
DsZCRnB/jb1zhlSjbHf6Y8UeaZpKqRc7bAmkMEa/N+6049TulFi4SXXTszFQgx3p
xRfIRim/PDqg8Ag+CnlEdegfWY57WgtzBnFCIoQ09z6jrwWFDCg5O83X6tSCo2Ob
LyOfP1l8b+45ELAiFdxB5xP1Yw0gMV8D19Ch9j9/rvDyEN5p9PtqJ6g+BY+wmKoq
qlMTZJO513117alFXPgG6u2vUiQynHpd4eT7zUUKXpQYK4Q4A4djbNi+C/gKgg+c
616poL4W3R8p0r8QUz1fTQ9PzubjtL2CWGpcc70XaZiyI9ZaGF5oqhgF2S4j6/1s
ZjjbkI3uuOUNRPLD5HFNgxexl84wj3cZboA7LF2JuNFkOtYEyYU6CNJMVeBrK4Gn
7nIMtoJiyv9Du3K0i4CPnUFgfKhvgGHcawD20fRknFr4MjvhZfNJHKybuXXQ4HYP
5eVkwHVZNox8E+xZkX9XSKSypzlMbhF+vwb7eGxggdXBOJZ357Fnu+zYVOQqgR7P
GvPwIWxrM8YhJJ4k0Yh7yxFiYS0/5K5QhPpZa0tmG/Y5Z+HOrnqcfaOLOATTRs9V
QuvCau1SHXFo8+5JdfdxBraHVlJSNWhPZ3kZb4GZvBIQ+x6gtaLRGzT/I0WkgZtj
cK5dvpPE4egp4kC9gORTGeuRYRa+4xkLtUCUi/B8+41yqLCTXusWSk9Frm1w+Mk4
S8Fjn4FOWbWMvXj5U7Q/ru516DRBlDgwfgPMwyEr0aLMziLJR091haOwAVHzMo0K
XJzJgu6Je3znpjevtyRSunJvNKHMyq616ipayWlQhS19ctEO75M/toJQuW2U9MO3
NlRfZpStfMULLJbLnMye/OTcrlJ7j1B19nU/pUoqP9j9ptwGYKEUng867wUk1NYv
KszlIaG3lkHJe7/boEMPBlQ2E7vn2+AvsJ+daF/25rvZnMGc6OvyutG6SU+RAxDM
HTgQKKRU/msdHFUPfr3l9TBWY9wxy9fEkoAiDDnW6sd+cktrdxoewvZRYFoR49Ez
8SMd3VNw5w5TCXoXBwFWiIjQ7hSVV6lZjX4M6b4aCuGw5OcrVu9K7kwN8f7t3L5Q
9sQACia3zjKV2WTziVZmfkspWRCe8r5iM6AP1++15c5K17Xn5pljrK1yi7m/5QJM
43/Qu2cE8S1NvwQJmIeQrSm7cJB8MY0Oxyq9E/v+5NMLX/kCSCqUT2vyGLORm5Ba
pv0y2uPR9suDzy/u9wOT8n/qSHyph8dVKlfrn1f1ikJ0Ig77zwviV06X/6xZQJDO
sgR9/QWYZKIgw9dJfYIOL2m8rsHuL26J/SayJ1wnOCpc4zGzQYNFmw32C8G2btEE
U/utkRLAYnRj173yDq8tAO20W6AWCCz1rFpitkuoa4bGCMZZkOrf+2k4w7BsqRkh
MoG6p8kZv0/suP/HApnzCJvhO2jCIY+vfFgnLQAcXZB4F6nF0rc3tSOcdldboeij
QU0253sSuOEBRiY5WysB2+EW3gUo1ZpBqw+H+VY9vlrbcKm9ZZIUHZ2o0VQs2bLe
B/zqe42jFgGnmRynWLODo0jHLhmp5JjpNCOZybDm3Wq7WtLeLkI6HUqfeZnznJIz
xTX3FyCOnpwaEd9dlpJ0R01xpFrcSYRZmCI74pRjL1pfPGEufFdReYsg9UspJQPx
9jCoDhoVE6PJHSrw2ywzKiw6RI2TDZhMlq2SMYBDzsf8I02klt5n4JfLRrCsoRjC
pER24X/Zb9vuxN+88I4sqAuRqytv40NOJIvKSZ096cNudCDSwOSpHFZykMeBRjXu
UfSGN8ZZVnApgTLI2SPheOiaRt0oG1OB8gOqtiamrsduAt8AvIpaMrpYLESk8Qn4
Dt7lAptdwsC4YHirV7ekgtH4y01/lLTj0sT3/xjt8lOSrQrhR3xQsYAL+vzPBUYa
Z0Z7ZStmXCa0v2KDq6P5zvThCozjHzl0WvQXK9kNMT5fjB4rESqxjobls0LGDBG/
7ZAgMc7W+mGCOoqIFay1aLIiVQ7f+rhhp87qPeR8gqIEH257rlKDOWGhAuKl3qDh
JBJNOvU201UkYOMVCytOinJiRbDKVCnYmBIybPyKpVJWHz5qjyiE5g8wWgnU9+Xi
qNKgQx/uBSlf8ggVU0hhQ58ttr2s7m2oR6hLog72I4RbRP/1dpwK4yaujG7MHJgC
S4gXf9ICJqKJFqdcd/kMc6vl+23IliZLaLe5/tUQxlBEsjO5nJaQ9mbJZQEX9IqG
+EoPU6HiyJSA4nYRwPloUTkOuB9dNZF5hLJ//74RjRNsgXjnKk2dc5kNvWz89ubr
MFDeh+2v34J1ID+UDeRZfAHe3a2enWgYsur9qo8zfNTq0f1H6ePssS9ajS06+5sU
OrE4M2LHuFWAIwqmzRPUHocB3Trb0NxJ0wicRrdPJPh9FevGxYmxbOJjZEwmABVZ
be8ff/t5/J7I/ZA2o2JvW5d59mtEA7g6Yb45ko6xVnHJ+KsSgcZBNosIJv4gFZ2b
0pfJlGMUl41vVvs+fhhnW8DWJSiyzf4Bh421NUo4ye8uLJsToFTvCYMj5C72MIZJ
JeYlSXLkKectSSPGAIP5cR084jgnLMd94DmWF1pSciRCcGGX2QPgB3wxfcUrYv1G
zslj8ukjECiv/poZJcr3PSE5x/cRKDIunaH2GfBgBpQFmYgPG/ltQaoDzYQGgzPy
yPUHO1aJeH8m50a73R48u5s253hHFmne6avshFNc/7NPB3xpUZc/h/tsJPGkXgUV
qtICByClqXrjWBOIm6m/4UcWmpYGDFV6cABLiETD5Q3RT8+3MqfiGaZqLXdr6Xdt
vxFPag6nDo4sq12TwbANODhTUQ1dDdcRuRMHbIKk7zJAxmY6vZCxqv/C9wk6TgDs
sMFm2fpuVDMd7eVb5VEg2mKKHqYZ+tt6Y6MIThhlF5i0dfcsq0D1Q4uyC0mCRAGf
1+lR35GA6Dc9PjkqcjrBPu63hjx9+1HF+S5ah9ZD1PBOnl4eZFesqkqfFezjP9pu
DfzHePGPznV6qRP4qU36Ylle7OTqcoNogjBsOn/uRxtofPm2LwDcSzArsw9/uQIe
KkChKizdpDwoqWy8LBEH52shMQe43KYBrR3o2r1I1OX1qUTELz0jV4c7od83SCPo
wH5huBVnUbUJwrbY9dXw7D2NmekFS5yRSUePMnEFpxtSbqvk3na6IePuaN0MVH6k
MKUrBtKutcLEY8YMdgw6JInPhDxlkPy1n1UhjqBSwRHpYS6+FnrEg3RWJZnk/gKI
5g0kGJUmPQRne3g8PP90BZ1GXlzZkV5qj5Jxo4ZHV9xtlWZrv93uxffhSrMIH+Ru
XBDLJZIEwfWfy4AgddcQbbizUTfzzPXurj7uvgxZQvLz6+iLciNJydnJpPfUT58n
vQ6PN0vWdGb46YfAnFpNK9h70G3zRRyR2ITe/gXv3KJNI6cAIgG4k8Nu3u2EbXjO
qpKBUGuFwqoofUZX2HfQ4eSRKXlWvQHhV92JltVnBIrTE6/GsMiU1Z721lakg9iS
8pWF/dQKMOcAoKR0WE080c1wRgDb0Kp0hbuOp0r223gs6WopXRfITm174OlO8rqe
PUaB8UtvaRv/d8sng1MWbcztrZD264UoXt07X7ChVwP9s0T6/AVOMn2s1hmYvlJl
N6q0gp58GN5sygnp9oFGyIGMFoi7i3MFwN6E+YZkeybmxfj/JPQFkJwlofjEC9NM
iY83vbEi5qgTZSKz3PbJMbXAy3+0gmbjd6Hy+DXRZhd8IOsElR0PoJwfL57HWR5A
6aqv5XBoU52Dh8UhvqwWwMqeKmIYVNz8rnuoHL0LEAjEaX3Xd3uoybeIXXhlr7ZB
dUufMdFVtloxWwcxcib21hmetYH9HWlbxbpKoPDUDFY0N1bIixejLUszBMl/RstO
Doa8E2WLyAzjAik6GM8ZqLKxFO0ljAA3FNbr4rVXboWjIE39YlSygZEoE+Cb1n/M
QBvbEPd4gPYdYRAy3Y+JHxf4AeKcddOLIMYv+Xwoo8arO0ThsSDZUbFFEGcSPa+f
oMMkuiRgn+B1zDwwf40BwuSQiUt/IPtrOJgxec3QNUq2IU8E5TFQGVNCvlPhD/Aa
Cb5vwlpn0miTbwMtfSZaILSFu9v5VraNEbHIDtH7ixMD+6q7BnapIooNU3lK69Ih
8Iy4KTy0gTK2Klrgie2UsiDduZdCaaEwz0Qul5hQXgRAbU14U+7gu5ViNMRpHmTl
xyXSA+G7ik0xHNIX8PAYg6l8fbUCHvVVisxOhbNjUP+ej7Db7jzYIJqcPNPn0/wF
QEEeytGS/msuLmmgOA7oqcGv48uk3RTIpfJcEtMxaYC5qPTYZUNWq5zl6TQess7M
7FcZci5eZvq4OVWYq6oK4dCuvBXGPQqA+7cmxkwi/T+WCJd5HmC1rL5ZzN7vlx/T
ERTuTxh7j0TfDrKqskG1pxKYnYJ5Jm8QE2SjXDfVp9hYnqmv1zunzTwGzT+owSH0
bTbXv0YQfhgSDWTEuUHsAYZm38bYDCogB5bcuZh3O0OfY185/kYPVpSVb1fLno/m
slvXGY//+7Fn/YyCMlprvETlHa+uOuYmHx12ievhYrFiMuqsgM6OXD6GVT0rwBKU
bC+32gKFyTmEfGVk5vTAbh8NVi+E4QgkiSg3u+PI6I2/95zFV0vGYmNBPc+0tXnv
G9sEsXsxjSEhAYY+wRkQCdx5q7KzP3wGxCP1qEmShRGZoftqCae5UzPl+J0R7xRf
lGPEqOubETk06hEYZeEyces9Jui20NziLG+AWoqTEtn1xs/l7cjBnmcmV7lCpTCe
2C9uT+r+Mob3sBwYJxYJk89sMivE8Qdq7aa4HWnA0luj1ICZSZvsaGX8EwsKLc5E
y/Lj/4LVCRlmUjJwEnY9I8RVCvQkj9muBa8p8K0/oVbVw7isLnzjNQe3MdZICiq4
yciKlVPzgcFPKqGPW1WB4ixRNDTVp/ges85ZTOwV77tqp/0tZXYl1Ps+Qok/kxLQ
s5VztFOQ695kGQpU3zLASNjxJ7pVqP4na7M6x87T77VPpvyXxFhlejYUSVT/6Gbz
jafq4hLyDzmyARBbcjg/hPvcsznY0HvG20rQY5YTo3MGYX/DftEvAbJQOVWkyh0B
TCFgybnp3vqHJc+Dn/AgrGbkERhKtOHmIlJS3H20lYeHzJbSKSWDX21JWLtG3Z+n
mCp7IFoHoRbYW4kMyuG6pXjiEtr+/SUEtpy/TTMEqyfEEouhufyQk9nrS+1EEScm
ISKkogT80IXb4i3Mb33TkSMMq3mWYRlk0c89YKeP12jDouAYv4pu2VloVIcBnRb9
ucgYk+KmFuQZhmeUtUozbKJZPPhyPtUmOQrOQ6DACruMNJ6vF1W3QefakW/uOlWu
3oSiqngZ+4lA9WqdOxVEJZFvyk0cxJA/zkoUcy3hmYOxUH4QeZ0cbBUAu+CUDdrv
wh5KVRdqtiMRDyRLiA/uH4RuO1WNZ3Xy9ArXglx9E3n2QK64CUu+d+u4wwcpG7bY
1ijd+gBVd6hm3StgQuOn8IDB//KRR6+ziTx5WRP+xwSVxtU4yBPFSUeAlAnTXvk+
w6gecYMkdRzJoZxsWkeWFGoO1fpiKHLoTWEztQhIus7ZdJwCLlZT0+0Vaw3e4sxS
WYKM5A14wbLqINyTXWL5ydoKHqhWRdd+dKnl1xXY9P3ZuphlK04ztw6YlPP/zTyl
U6TZdr43IEURuD5HGEJDHK6iNix2Myw5br26JCml0gAoZrMugPlruT7VzPT33zzO
I0O8zVo/Qrvk4jUueCe/IE87Z63V7W1v6MarN+jqtKkff2hFq195WMHDdHNWOrJZ
onaDxXVj6dZF7mdSIcPUSPJBTuf/JgDdIudyk1Pkw/IM/RWvFUk5XBf4q3pLVJrH
HMBTF3TMTfaL7qYtxfb0T8oE+uSCDyqO4C9tQSKGP8pRpjg5HS9fIb9b9oxjDvWO
nFRJYBHelZGWP4m2jBJFf3RueuCusr2onCPEsOlEfSLgXX4+VWIRfCTbGJUyfxem
mTcdPf4ftG1NFwjVy7PbjmijliHgqzLaTpcEiBroI+CeRTYwqAeMt+xFr/gzuEfe
v/vfQXc/spQOCJxQtNvvGHSHR2GwEALAekhiSaTCAhDEInrYqRJwSO3mdSXzzEMW
/lQJyZdsclHBmIBszUG+Onu5oUPNM1BBKbGY3ZyH/PBNN2MWSBklKahIkBgJ/rBS
5DlMfnFdwRjVGeE84OPV+ziTYh8ygQzziilKwq1n+CNkwjtxAv8/eLPFU4hNi2D8
lNTOZVn6XGLknzV0Aj5PwsiJGty09J7lH/ParUzVcZKr9ymv5H7qi8I51W/Wh9qh
NLX7Hh+GCM3CtODtNS2Vz0AMn8eqlol9tix/vus5yBb5u1wPD8jW7Gg2Lwet8KqQ
SxVvEC1fOV8FrI0fGXDMV+CZZatqDyY1567LRHqhpbPYcHavMiTlZiLiWXPhb3m8
U3xCcUGyUcQ+unAPKkPnqm6s1/geQDk9LNpyXEL+D2ndPee2Y/zRE+r3RV3gVdY9
spsq5t2OHWU4T+rBwrCHzs2pCBQFHqkA3/n4BgYs99hYXZH7uj92QL8uMeIicXrA
hHYQ9+hsf9QENFKl5hiwOONk2iN1If5tSBu4/8dOHkKqa9wsof6suAEdoVfehjtd
MyzAU8OWndq/ESuA0SNjldBMgrTU/EWxFl7rEmZJxnCYZHZ8jtGqXZ66gdJ3oVkp
UM6aHcrN4slmUOct2xTuWt7lyy57UV4XV34rmQLzZQ3EgrdxCVjoC2m4auyRyLBR
+bfirYXp9PgPqYzbnir62pDaPRxe+ssulDz00er+j/p7ZpDgSUuQfKayoczAYix+
RaYxtpz4edkI07lTwgBqZ5qHzvpiy8bqT1aPlODSqkrwUBDCZYQDzMkw1EX748Y5
bkcN67VnDZxF4r9Jl805/M+c5058r0CkLN47jZZ6vyVwNOR4jnMypWIJfuCgqU7v
2BKkbon0ntrUJcCievBsvFKWTcVocA0BiB5n/8LIXVCFCsBJXsILn7jOfXq3+2RD
WZl8OjVcCmu3WSOsY3uEUHa9gDU9LV16qr6Z86rBsDqaQ8SJrtvueMvaxOUMkzVT
n87bkiOS5nA+Sl8etRV5krIOhXKvxTQlp8MeaFrCgTlMPbm33jzkDt1i0ldFEzJ2
zijvUU5CwLN9Ck71UU6ikLMeCJPUq2d0RMyPlWsEz5U2YnLHj59V/v7/+b98ggcK
reYzid7bOkhhCJ1hfok7F0/4pf2xC5ucKwkCtsN070/6+G4Os7nPMV+qfKKAPdiS
o305EMFgiTzyN6NdRHUs9zmzRzWi1p1WvdtuiQkFjP0YuolBH1dbSvk+HBcDsTS6
qUceT3a8d+qePKlOeJ5sTUFc4pvSWZ1jWuB/LCSW+Gmjo13aQiO4kSTM9qN/IuCv
c7ylCffSewTZ59rEp041Vf+y5aUdYMgTf7n1o+y4KOQ2yLQRmY6wxF3OeN0ZGK5k
uFMCJ8PLFLdhMOV4K0sORIrJcQR3NU7+nKkmIvK010BRwePvGdlOfN6Hk05ziIuo
SvEwen3fktZq+wJV8M+pPOPOEVX6Ly+vABcbAws2JEVjk9gbCBcLGPFCDJAiAP1y
YAeH/fwGGf2ky1zDbRyCkQeRQv3rKGwp3bGBPY1oysjb8IPK95+Tk0GGlh24JSbr
6VJtOv1q/wjPPgCRQtHiG4PTFenbsbdi+Fem0+8v6EwMXHeOX+XI/6okbaBFnFeK
gw8eiN+EaInyvtVjzYA/i6yc8EQpikVoOrq9VI0L6eaoTJpHmX9mZkCR7/XWo4+m
qQTDQWDFNWFH2eU3oeOI1j2uJ5rY34XmTaBxMsMlZwwqWMIGOuL+EM1dNjsPQwh3
kTr0mXzJvQS5nkQjyxGErf2qKGhXpXuG//c0dYZ/U58PmATfXAtK+DpWax8Ch/wY
5UroUzuvq9P0MFje7ez7ub/Rh2eKoTDsvlV6xSPqTudA39bVY8n0t3k9M5SeaHa7
Wpwnq241f0iDdbmK5fGFsbvGLDg+9rYn32CxJJPW83IRCyx6ShUxi+5yKhVy4Rqo
A2cOq9MIXnFx+mXrB8/MkUgTRZqztUf0DCneiVoNzB8adhkAuPPqqopZZdsc0UGx
GHiwM3sEdN3DgYTsLjqjCcZ2bjkNfanIC3Zm0UCDAYKtuRl6lUMwnitGDxKZrdWf
Fqrr6IEqegRyWNzuoYgy7aBLvrVOD0hKdZnbYnpORCrLiDjDdSU61Sh59WjkSBmP
lX16J7aq9yKTpw2KOxrFKrC4Kph9PvG1y1zf4lsoBj3lQJehCsFPwQKJuKgiuen2
mrSlHCT3Agk7ForsrW4lV5AlkLfGmL57nIsm45CEh4T05YA27fU6Kj03cBY2P4PU
KfXPjUyoZu52ErxLJEyMGrXlBsKVNi0tpkCA8MWM65qA9qyDDdlew+t+YgK0VWUp
7xV8GDv4a9Fuyo8gNASgk51kWcZ3weuk1Em0qZIUIGml/TP3yPnOhLwtdkUZCtuM
P1Damp5LdMK63A6cecyRCWtC67QynC+Uk92PHA7A+Z9kzxyPjEQNqpwUoiNnOMYO
vcEIowdK9b6We08rcxZlqPgM8xZ+MJyUjQTYr9WI6eHPD9Rg7suGuyDJ43Irsk41
wLFCXS3CwJWF8zQU6UeDyi5SwxB9kkV2PUvfZcrYADhcp1di+cbFmhWNebtG5uwa
j+J6pFvpfq/U+D9u3unPYS9GhXndB1mH5clmDtXvsjvke1UIFvbH8EtZ5tsjIObp
MRaPo5iTWzbrSIVMDKOSMd9Cx6UUh86jIPv61awD77vYGkF8idsbC7GyW6M3asy7
T5vFBMuQvAcmU5LHR+jipkDtMWJZPl/Zoh4zZCh78fDEedvDeTr3OHfV1Bk6VTqu
pJOMJosgM2LNeWCIEOpwWrB3U/50zpSRAxQe4RaXFKu3czrL95ih+i8GRriM+0XS
BhCMmLM3ZCvhx/XNMLkDWey3Mdacjg3xA/o2nczgbzr2kkxsrIIw3NVatsuwEIQI
uC0bXayfKwjqn2vexV4M+zLfTVuN7CFmnXumY3c5F8GlWCXfM1P/7i8ClNZrnQ1f
dmcpHjyf9M5l5Pq6yJAo7b6vyYZQ+RCaDiZXUWQOPkI8gZsMnh3hSlzcsYeITOeb
hWuVm5h4THDjoXim2xb4ohBpUsPZ9a4hNl0ym90tchnr5hjF7dsyj78sy7V3KpW8
DkOE1jqmX3tw2oyvhf+3PcFBLixS05u3oIcsy+y2VPsIJ2SiBdoehbejIlOGMYD9
JoDMO/cYP9UtLrh7+mexSKYLK01XLPS0T/sC72gakHfJqIMcBzZKZsukPJKenCru
Ac+14E00LKaiiBjcAsoJzmm1gW1U5jDJEqk4FQTnyKaEXrSrBdGYOqDAGQR76KSx
+Rxy2PgTCfMw1DpAwE7f+2eKbm8N5tihDNKCGq57ge/0iOJ1oHKnPUheMWOCfBna
HdS9UPCQWaXRT48y20L4QfIJewBNfDSXMc2GezRBYSQM7gsMoNi9bhxZLhgUsfU+
X04NVRXROnAw+qNMbfri9tNLj8jZWVIuceM3/bOl6YTo8vUHNDK+4ZwAjSSGQuAW
CN0DzEHiIi5A17hyq5rewIbY7q1l+jjipTcQZVKe7Mtxbe+1A7Yb0qs3TOBx7upE
vXGpj6CPiUCciIPY6UMyHtJVBWot9nxfgAHMWyjVi1jm47Kybx/1BiZg5y/StOxr
mAjQfR7vqboJRNL9kyXL3ri4/vECWuMue6vXZT8qv/02Kgp3jmLq3gO1F+gpZl69
9+/yThwD0zfHKtCOY3hL3nY8oPkVwdbjkkk74nttjH3KOilM/8wOe1QwmV64bmKd
oV6oQ3tPhfVYxMtSkz46EPZjOpjPuI50xdigASO24kbMZQ/NOSgs973edXrH4qlQ
KfdJo6EZvlkPt0zHKkn+l5UmVn5IUwHEzJoGCXNzYzYxS4RcD/cV6tMTSvGfs/Ut
x1pWF5ub8KrTGvKkIcUazfOyfWMYOduXoCV1mFxfEe9H1f6Z04W7cgzsfgnQCkL0
9mXCkQEJd0TzM/OIg3zA3pcAKcZ1U7gw+EcvBD5JMYuCfc9ttV6gAFVXlgWqkc2s
v9oDoIQY/x854Pl6+Cq05FkZQFDilv7kcZwk6xjMqKqN5eP4kD+TwdJv2IkIwXXc
EOJh8sx+mChHhYOVWhx5tNeEA5r5VgxZMZDhsHJ/NN54W+ErbGLBshZzU3q69z55
MlbP0YMp/yq5f9wKLdSOK0GRJljUS56xaXq5I7zdK01Jup71jlFNnoeiHCzy1IAC
x7ffV85KXSrwI90RbYOdkknOaiN39O90gUB8aogVmZu7DkYq5mD76AaqNHj8sFT6
cNbhn/4a4aHgKCNgAbyX9yOYpBuuSQS3ntMMjXfMNKdLH+edLRUcwgrABx2fX06Z
iiaCsqXSfpNj9B+ujDUr2I3koMi7Q40k+JjEA0ASMNlAI9mABTX3xdHsli0zRYvU
LKiiIrkcQyWHnfdpBYwntCZscaWBdkH6xKgL+DBo/mnXD20zov7foJvLroQ8RSt4
lYSJV4eoxJdg4UG+rPosLwDFdmFxwKlb7YUNWxLE8bIQRrIKawWFMJaSaOMNalSR
EOGZN6e15XE8wSmXyOBGx0inLf9rxL3nIlFlUnS33XbNtboVqWB3y7RiGl+U0pUs
NASoiZghCyYoJ13O7TxYasrdtV4WJ680hb4poVoVHoeHwmsfT+hDSYClws5H2eFJ
j9vO7YiGDeGvvJ3RKXFAqeBfVl0Mr9+SOEVe3OD18M8v7zLgGRG8S4VVz38OJ2Jz
EdMHhsmToRo7Vw9o0EowRHp0jN/5XRyTxQ4SUNsjbly6eDXNPNYAnH2J615BQuBZ
0E53PYDWstQQ+9Fx9greW9rXuvitJObGWKSgeugiSjsMQKZDvnh60KOzqTUP4D8F
gYFsCEhF9nevFyH1kRbUnZBO1WUPGELAXbDGAC+GMJ5y96wTjx2+/VM2KLyJPjHI
8MxWN43qZXdcq4Evxrcng5mfdxVnI7ft2LZQSTHrgfRqsmpEG2uyMEn5vY99QoV8
SzpoHSA46uWcq7P6tAM1W58ODAAlGwhQgrROELsMXMVXybxUq/Xwww2laNx23/iF
vE/rIQ8yKm8FeUoIWsAHiukVsdHxB2EwHnIwtO2/cGS9yTbvaGs4Z4ZENYFBMJwD
V29sJbAV9CA/9/ZtVvj9VVShPMlRyC0UtrBixJKUp0lP3/eMMWYPYtuzzguBIaOb
KR0YO4NEqhtNEnIQTiL3S3m3RH0YB6EUSQovHdj9JzpzaL3bLBrKbWEKW8O7ys7a
/R8KvncgXe05JiJDEAZff/nwgivo2za1olCYB0tZwnx0dH9a70ioHUCUwf3MVN5O
/2gvwpo2PrUxoWg1LUjcU927h+W0O0HIzu/MUCFqs53vJjrp4kzNoJDqMtralZx7
FlZViq/2j9Z7m3FgKGgeN3RPzN/6GLys6v0TF8f9nEqYSgPiupflx3Gh9YzSVEkQ
iaeh1GfFH3jhAfOQ6k1QsPbRAkjWZg8/DuUALy3tmlZfaht41z1NvApCYHPvSsew
6paJcpY0NWQbCinyqnku6JYyjirbBdv/Hggmr3kmYc+pcG6/RzV+PbIAcqKSfJI2
CwAQ/z3OT0+XmdF5uQtTzTSvKinwIGQn0cCu1T1+FNElJeNJ5U5v2Sc26Qn8uX1b
jsI4ZGWM58qBSYcZbtZ0GPXMb3Iwsy8GXg1LXRht6+P3tKEUJi2GOn9MM7xf5CPw
YSKL5Zg4BKOe+CQnHC9tcqxxCSFwWn9TnJd/BR/UABMFu2qwMpXo/08Upys/7/EW
0iCpBzKsjvGHnsV2VkOfH7zKsz82eecRgRlPPrqUawD5Phc22gCoXhvAiUkVpQKK
wiOFd9Xvv1nc+O5qGdSPwF0F3N4nn2vqs50B/msGbVj+SP4inkfWjCyPhZieEhxY
yLljwvxTJy1Z4liB9J066DkzpN0JB2vQcdc3EGkWjA2HRRv19wYNDBH9xyxoC2jw
8SsS923hIb2ASbyPGJs0PJjsCZBvZ0aVK69/FYCipqWLpc+VxeycbpDnMmIIeUYx
3IWwfec/rNmNJyPuKlOwRRc+QMEbcLXo1Tr308UWEwkgtvjlr2Q0a/G5PEiFnMrM
z1maAuRLo6iLMjvCn2Bt50RAsnb4x1LTrkLuQF513H2fHyZTIxHa1/W2pwIA6haF
QYsQOr5WTr6m8QYYXHXWujtisvrwMN0Eq/vpUgE99RjONhpx9xNfXT9GoVCyLy25
0jGwA1nM8j+Tz+3qq0kReFkS/Mp+g8Ak/tvEbXkUIDLT20G0AOrnABbHIqb0BDxg
SB+dXHqH7GIHkkHQy70eJiUDeovQlJbJ78Yry1QfWmXVgeNwuCscVhhbA9OzMK+6
rW2avbyint2GCoF+gaRNB48G/gITZAeswbHWeVlH6vCb4eQK5MeSTWntpkWi4XZJ
O/HfFdKiln8zL/AwydBTYj/Gk+A8h06FYYUv6fccg8p2PtF1R1EfIlGYPWRKWzNy
+fOVDVYsL/dCE3kIV8LEgpI3Msfb7/rRz/IRYCRTB+pFu0YOSe3fZQEVGUJ3iDTE
VCGphe+iwiAiw9QBRkE+bKiQN3HInEL3Wj4SxK/VTvs9z5xxAogzJwBjNxjA//fv
rOkXOcCld3bLA/zEJaJ4iPok/VoO8wdhmsXAt0UXFNLOg9usbC3ZdaH+uGDDHMii
eMWUgZvri9AlgchLxKCubRJPp5t5K+t4U+2hH/QVX7lwsdrZemeqpY7dcVQfv/JE
dDCs6rimy2lYi9LPkEGpysWaD6z/Q9rz0Vkdrb+lUHqdf5iX7HrV0csxTbnbVaSm
lmRjaLoyZTTTyJvEhx5AvgmBb1Gxn1sfexzA90idPfHIQzyvcnDFgeotBsCvtiWl
RpWTCkNW1PP4jEBaWR8u61nR0FrTBmdO80pEH1SzIltCuTIQ2OQF5QCYIU7aVPP6
NKQKl8mw41QoWzkRlN6pmNs/6Akxs83f6olA5Twc83Xt/pzUFgI50FZNhPq9Ik//
Mgnq89LbPRjht4YbMR9vzJZyouM5/dbJ5qBPoPG3JdJzGCBX6Mo0AT2OTrHGhbe5
qiNYGYpywpJCKtC5jl68Yo8Z8SBJrzRImJBCf9KYKffSUIJkrIkECIB/mYptOH4K
6mvFULOtZN/ySkREXLl9HyMkG/N+4U51MdG409ZjXOV8j0/14OFy/eoMy01c4b37
90IcF23t1KRXT0aqOWx2+yDNYn08CrEtKxhGrPkUx7Pj4gkTWx39z56seqN4mMJ+
wQGT+gG+2NJPtUTauF9kP6PYxJHK+iD67yz6AhJ6jMAODnVk1RlgiIolQ6DB8Loo
xB7ePopoi1fRZPqfH+GDe6tsC4VeetMcMbDOEZI3Xqfz/OQ305VDDdw/brKhuCZg
vCYZ6pR7zVGMhoab5WjJHxV5hjsWWLhRtn6EPLksjwVDbIBX8OfZdPGjcy7kPSux
cS4HhNIYj6jnHuWo0sB2JBLhWJk1l0Au+GWJSQWXFaNcpWDfYID4UZ6t49aTNo0P
5A1ndi4n0zR+dsiFDGikraE/gf0dznq/UI/g/COOjrJeA+/JpCGgbhWQ0SQasF77
y3LUUdqlByKeFZaUWZajAb/rrxvR6CEih5ctleLOnNUpFxL9Aj9ApWuWTikAZwok
XrBCAvSsXPoUMoakTjirkMxsjA5wrbmwHTeyUFPAkjYVPjOYQfKtOcJSWnWEVAKC
h06qqZHGS1w1/O2yOHaauKGXAge3yjnkLQSRsn0TtnYwXj7Rzjl71OiLwH+Khw0q
/h4GbsYvwoqaKuFtKVRdm/nDBae0BOvbQe8QLU0V22zan6Zg1iIZZ8mvcRn3Wp/P
5Yqo2cj1byc14p32d+Aw3qxPSZ8lzo9BSjgnutdYWMsWbvoa0ePX7aDmmn+f91W6
bv1mlCK1yZc6pMAxT7fK+GmYsLHbnHnKekvZC8lUyU33Tl23Lr+uAkUmFJ91fZpK
OdR6rmPGBAN68S+eSmpzI0t73+GHRuTNQ9eW/u4M3EmIqT+cDjf1PtJ1/rrXMW5y
/s4LjYpCopYy+3pQmLNVJdgLzcoVI756RERAEpSSaMsiVVGJvGyOgcOzwFSvOGug
ML8fHltk7flnt/njoRdQzCmwP3lZbt46PpYIuQjyeVIccXSo0+nNbmrJVnKvk5d4
rmmqdKRgGiDuoL0gJ3NSlx6KGg6VKK8n7cgJr8LH2gJaXl8glXFB6TgHUxSRJynu
pPFcPz0n7Ayr//qHSgh2rKWrxcrtPtnTypb53HPDk5nyPpOKStcAMNwVg+VuqOcx
36H3A6IxgPdH/v9deBS9N5hzeTF7ask89m3/9ScwXJwDtBQhseiTbSkKZj+mLQO4
U6gIlBF68CbVMEAxGT/aTHYSyLUn8VsejL763be73WK9Dv6W7HzhXTf/i9s+QvkR
d+5Bl0S2q33p9MGfXSooM7mboKXSRiWi7iFk0JUU9Kr8bxmdQvsXPbIwJfB4+Fq4
dhsZ2mng3mMZUCCgV3l4KzAxz/Ase2DerHEdrOMOir6+eL5vgyUQ5ewqEMLQFX7x
QQGhpM+KYWTSDnbGovNdo6e0wIsrGHg9YvC88h+zVoK/b5QOsBWs1fM0EkepzIYS
ZNmUWRvbL4B34060u1sj/wIRPngvNIn/XjNMJ+bgYYXL4Bm3jVhwD48YgA4iPiqD
3tZOcUKqXwVBtLelbu88UtExVMQdQL5RTw5j3Jas4BCKusmdLcTTiKMBkcZH/j8L
0SbQcnsMQjLaAfR7diSUdRSU6wEPO6xe58ogoAN5KrF5NR8rAsjja5dir5O3pU20
Gb5c4d3C8MbikPUqn0zyv+NKnwuduuAlgnkJk7WCrMwbHOmQQDkOy8aKrv7pIIkU
HKgPyQ75MSzvLxugiNBkJxi1XkWHAlQ1HsimbaaXt+1k5rOl3CjkyUDlW/MfKmBz
SJmo0yupkzx3nDd9P1PiM/PWVUuDPUf4pccQvgiTjz3rz7EQGj7tAj2Le3o0bjiy
Cg4zMB01fcutV85v1389v5Ll2iIl+oJawcfXFCMBl9IWUjTjuP2rAx3Z6yruK5yy
0UYipDAUGMXAg3mRx+OPbSStTzEYRFsN8fVd+OQht97g9LvqvL8SKecs7I3n8QWc
5a0YP5B+1bCexh+fvRfYpfNWj0ISfAc9rHJpgS3M2HYZ6EQK++17PXUtf6joXJbW
XDDUMicKkSr7YUAmgJBoA4srymQ6L7iGrSpoMJWlYgC7MxOdCGTHtHUJvGlmTkvJ
IDtst8OhVCEeQN+hmHcBqShfPE5vXd/N1zuOegi/X1xb3lqI2OYlPA7Ub3l5tb30
AcN8s0+GkoXuwgrhUWMvFkXsOuhgp8y8rZEgKOaiJgSklZURCN53SVm6AtmJlNOM
FqaIgALJ7wEtxkyS3DQOs9ozzLUa2/C2K0wMr66STB9887cx2Qj9pKuA/HpRSR4m
ozn0PJfm9rQXqPPzBu1xAes4Lp8R7et7dg/9qm5KAzbWDO9ZWb4XnR2+Tc7r1yUR
HCjeG2wuKAiGnqV+RcMpaeylwsOv1O6hxWomPaYiiN1Y2hqNiAvQw4jnslj3T9/3
gt2kJJXSv+OTn0HuzgHWxmZw0s5yfpe0bEYRv7/P+5mEWEtk8kHBVMsawdmDk0Bf
5aYcjvJwMKoxfkAlZbg+84EBwQAqk41IRqaBFgKX28n3uoW7q5hljalksSNhq4T9
+HmBwyTTpwsV3oB++Q6HoBFQM8wdU5ZczUIO1cnriK8mFc6QO0LNsuyCQ04skuyS
lCN9z5YaC/Z6PJEsAPJQWLxvDodGF0lUP8bKF9AaoSfI6vkStSaNDvFBQS4vLCKg
+6eMG2Ko4J1jlSCXzKNr8Ew2PWl7WRN2HuGhSN+nccFfle2Yg/zR0swEdGlMbiuG
qm9mF3qDvxfGKOLvSTb4FAH//F+8sUJF3NJ3mRFllsTGHezeivQBQSRRB2gtvrGz
/ZXr7HsR6YOZ4WzeoL0fO2uzvMXEJ7IiNz11I9kCEYa6AUfGZL/wcWkgTzYkxqrb
iAr+WaJGV4WNX2SWp/NDN68jghWHxQDOZedf/lmVGydu35p8m5k8/8PqJSw4o23w
UNPomRCOJHJvFVV4jEWXZj4A/n6v0IS3kel/2TorTV+4zTMJc+wOPDOU6aYaAPGM
kUNmFg/JUoepDLrXEgC9P6lkrm50GfcbDOQl/OkrzakxWL/51A3xGNPkeaFSyELQ
/WQBGob9mlFEHfzyb0DmcHXIFozEfx63knwSQ+VM1g/bg0OfMzRBEMHKkRl6d7l1
uUwcmBTvA1rurI1AIpasWRCsb7qgVyEl9twMYBkaOIwyzEQjFDFkSyTqogebGCWX
DK6RXUkgJFRR2/n3zmvLpzr6sjkbXBFhlhOnEDjb1Ho3SdIwNyHFgikro830XUjK
5obaR9WoFeZXEeDJicLi4+2I0Bd3rBLh0eMAkl7u5nscHul3XUIHMIsm+5Flr3Mi
Zd9dMXHbV9ard+B4OPA0T3nXyoupY6Nx3A2DqE9+qdcbFPnAIgnCAMdrlvzf+Fq2
zDjVE14zAKJJNStXx417IMLsfpQqaYpeUS53XQ1VChHATWdREupcHy9D5D99wdm/
9tqw+zJMd2V1FaitPyD5ogYJ6KfY01oEnmPYu6WgqQU=
`pragma protect end_protected
