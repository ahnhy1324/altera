// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fFqU6J2ZNNFMPDbxZ3GVn8zy+vGEgYONGp87LPHzxtaQPKxY7SaZH8fIbP4xQN50
Hvp8A+hh66baWNqM2VR7gvhR0rwfIECDDMdna8HG/cspwfkR6hClm3XKBzSUJ3EL
RKOFsaZmam4Yq7YVXDsxIC+8LHWS1CoRQvYnCC1N1lc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24768)
n7yWFQdbpdBc0UW4o6HHcyjTLWFGy3sA2Bb93VnHjK4L90XXmSQEO1wUHRl1REAX
WZEe+VpQSWJoD8lBD5ob/cWLBIp/UrNfxE8K9M3laSuA4iaphVbdkMHntSJMuQCb
QnjoUEYE27HHFXXJdD/M91Z1MmOo+n18NAzR59mdxZ7U1p7SBjwcnKGzyA+m8XxG
NwVdrnHrXwCoC4snABoDyPDi4Dg2Ym+KklajGB/zT4fn+xk7oUOO2w0iaM7/xrnD
LABF4dH4zwVzV4ld4fCOFRvl9RqlDE3YZrD2SgIih4tyQej0E28hlweClBzNdihN
vEaILrG68FALeKZGDyP/wvD5tFiNp7vkXyCCtzet+GPbdW8vAp/xbJ+to7t1stR/
6KTfvTWzrGpyPbjICI/xgaLAn/BJS/HxDC4JxQOk0+bCHsTtXJ9ecgbof7bpSbDl
zWOavD11uUJfOGdQy/G9kg420sYl+vnNhAIL1Q1b31pA0CKC7j2O1iZb3NGbYx/b
nhbiGU5SP4mOUxnmRDv6zuiysTpMcRZPNbHp9/hqntaLiayGA+jeSaWkDbp+JCLE
t7jgg9PWlf4NJCe3Du5bCV0D9PsSNw3lqsdqX7CRolbH3wg+AiEcT3OFk8fi4o8I
VnRDFg4vQBANEnZV/Xb8WuMEKTTWcRRdBmysyHbJ2ywArZ7SCVPeQtlBgHddCHA0
hmPveTzVK4ukfVk6X+iiWBBU35tIy17SRnLUOGY0NjzEp3qdVe/kVx/9mTDWuBVm
I+NbOhqBnx4nl48x9Ztm3GDZKHVibqp7/lPYyyuZWz52kUvrKH0qjKI58QD5qxNG
BmwgtWazx5KpIepKQfMqUbuWpCoMJMvmiY8f/ReJuxGa26k9qaNsD4aQrwPCj4/P
++i8fUqBV8FocKK0oQ8ZQjLZQdBM7F8mw7k4GaaHhYKjfPgXwpWDclLDTXFOhau5
9whxX6vMP9FuC75RFvtV7x2BXZ2S8XHt436UD8OiusgsNHMWKdDD7YzdgSYpLslL
8K6VNuHR7TAZscT6+LuYqvdhwpWaQMDut4u9JsKj7o4a3fdjdlxZddDnxdyQ2u6y
F5ermx0brWLmFQaSFE1SUT/WjgKldTvWJFPwO9C66D6Fo1qtYL3Xb+Jx5wt93oO3
SHIPag+Fk4MiQ9+ciGGrjnucdMG8sKa0wEI4XYyNaFK/9I680q25g46CNrhVUJVn
Qbv9a5cUXpuYu8qtXum03C+00qkLH6EaMgL+vZpZCpwAIS/uzTBToqbGyK231DwL
4XraH2c7i7AKCC2mMea32yehtXdb+ILfgXkjK03ErhYEjMeItFaBojUU3nDFuVfl
CsLQ62tOlUgGYFPAR/6jTPQRdzVOsnPuN+L3xCNpFmhHmLSZzAxKSEJp7vY8QDn2
SBkIZHanzEbQG9/mvJ/dLUuKmswP1+tYdv4cOJhTGSGnJcQNKJF8CY5tYRUo6drO
9qIXac/Qs27FfIZTsyOvL27MdIZWZ0omDd5zNu/gdUGhJgOl5YunTQYBoaBEMA4T
y7IqVvW7Rbum36cjBrS2visPZRCvpiAOi6n1fd6ybzeBRSneYFzkPk3TEciMvY/1
iA7+rtMMdZ4PpHDRnqLgIHenFMYLjz8OHFNg7Gkw3OcXuwVwSyO/uRPN6L9gfMGG
7c9o0h/gmTO42bIqNvzb+bx9lEjng/FWz/joEJ+xgLDN7nmdRdB3tzWQhIHyAkZM
H0r7YcoR9X7g4gEp3PrMvwPf+/5rgkqPpnWvv8mbuCbCu1JkB/2d8rSG5qVYGRPo
qv+UQUQyEV3t9bp/r7TOg+d/8NnlwzfoA53PNOpyI563dSSRksAEPatuiEuhUkue
6oOwJb9G0c9l0nA+O+Ax9aXofiKZJH+XyxIhQVZ4K/lrwQTLYKSrXu+YrQvkJvHA
VDZ9krVnszGWkVqFiOsB3g5iKGOP1sajDzHmcJCZhRfgx8+JtTvPnpEx7cjMD5mz
aFv/wpkGKLoQzhI+wzgw9kxyWsRHPPUZ8bN8eRHuVroqL0IniG0nZ6Xko20rolTg
mf8ZFl0AhXtOwCJtRt7L46JgohDkKv4CYdU1RCzp7cAInTsN8Gc3fK9eJwnI3Ebg
F0D0wI3fObX/igvMsHCGtoeRO85a6GYR9smeeK326ndNDYgCEZVG2IbCqn3RSUv0
mExdvvbNH4rppmvhaya4htvWG28nRv3E5LOfv78xQAAEIijLQ+IAwlGda985Ib/x
6IPU3zAVM+ofjC/BcJ+sSD1ZM5bBdb606tvzMdMMsvbjBYLrnjxZvPrtDGDZRTKN
MrB1k+ptKbMRNPiQk6xt6AijmO0ZC7O9aZ+Ly/MJW8DDhZR9XHDujBz43xCchNsy
Wdmj0mlcWevTTVIZ0/o6OkhICbG2bBiUZolgeuneDN7U7DWDw7nMLLakV3yuPOoi
gwPCffj2QacbThhXJRXqcdhEHwNUMbgD17iBpHhqFknRA4fxsN7SchCnzlULWt7f
Ahco/3LmM8hD9sFAcw28q0KTuth1AKb91J8RM8gEZT+3Q9rVudOpPS6ude3aWS0X
tmUexjC8hDw018ibwu0Fy15JSc72I2s4MJT9qL8nNLOsPfUDvKfyMbcBSust0Kjr
Khk+cbMU4Q2XokkWBWRtB5I9JRhm1lgHzyZE3TbjJrLbOMxBjgf+DfSxIQG6nUFg
lkI8LkzvU1EEfkcnIGkPyoRoZgDeSegMo4pViUu4vm9P2ppjlImoy6MtRIlz6R0i
kozMMyq4hGd/mZ4A2Z/Do8Cxa5LESyaYudElx6o0dP+KKhdIHXjQ7uXaOlSyDIWr
SP0Vl22JDO9FsGViZW514w51JGPgz4Ow7kg9OPSbbuqpI7Acw2SK7xY/BYvmscyI
40OeA/yHFvljQf89Pck1pEMehiEn2W2RFkZWG2O5LQI+7PoidxwO7DY22cp41nl8
kXZAFgwouzIOneOTWS2w02zgJhob8C4B+5M7L4bas6HjeZaZ7RVp3uZdJ3XxIAcl
nWq4AAP54SDSoRATdzF4sBrPsPBhigDDTvBdizY2RSuGqUHScnjQFm4ou8qV7Ex+
JRPU3ndfAGOH4xRHKBoccyn/G4ytVMdwT4MyiNOyGijJVwTC+fQZwkLmrVOAXG01
dUw1NnAGYzgBQ0puhmP7PERsCTPt0Zd0DcZSmUb/wYaRgzeoLRD0iaWwj4FRmHdr
ng8DcvxfsiSnhVz9Y0xnZsr1UX30SyzLVpQSANR/u3yvJt/0BMqT6RSl9Na012si
zJnK21lGZ6wne4elXsCdMn1tlfi35Cc4NXJyrxO795YXcTwka/bAhkN7BKKkxTDr
bgiENCIa+emow966LBYZRv9XQ6ANVHj99ISOTi3o+b/z8JdSpE+muvkQWweeh6iN
vPcP7S0H9aWWqHQMw5ArqOVhRPAueBC7YDusWz14mKAyNeqpGfFTIzS6JZfX8OM5
z/ka7d5VGnXkQpGZAMdnNRKulmycy0NHz4/M+NzBqtqAvsloPXNF2LDStG0Hd0sf
jSJchYCBbbXxixjA1sW9MFeWWkqC8txJ4oQ9rUGx49Lm8K8eCxT99QJA4MzJK8w4
7rpqpDOcnLhE8jx7xGiM64j/knL2Q/C8rUTZPxVVety+0JsrCU4M48c2sgkRzV5T
fuOdEh5bDoKdWH1aPkcLQ7ERmAgv4lo2xvfa/cidIQujWJSfTVXd2csXutyzr1wa
FFZ10GO6bbV375Ukp9X4zhtidEWYfYY4cl0PHAxGd9gLWLsBxOng04ffgZMHyoV5
o3wLsCjaQChbZAqTCjmhOMC+b3URjP706XOdifADGs5ZuwMzj7q/COcQZVbLV/BX
C5Ku5UY0AyEZXhgmMtNMSDmkM6pGDf4VnMypOft0YFakEEq2N6FPHJTDGecrSNGe
q1ohn0yyrnftcoZCDrRZgLG+3ONaBKs9VhCS1rsY71iWtHc+wxKnv5bwIpsdxKgU
EDqnRgMCWabNWGDDONFwfm3PbaKi18WYdH1K3st4w3hRkIKMwndMPNkPpKRcHwQw
cw3HlBCNu95HhHE8OhAMWydeeZLTzs1BG92GxAjmy7HLqrNItXlMyeCWgvN4bRYO
mrC3O8cia2eui1UekKmoEX9O8l03/S/NoJXwX60a08a0dvLFwsYn/rkEA5qlsU4i
dmjR5ksy4AF/uQ7NGCqAuRBz/C8U75DXIlCl6LVdSVwhxkSFnwy5ZdAulhvYmMwb
WHbZN//iDSRd/Tx27yakC3FagI1VWDTdL3hTBL2pUC36WEBQ0MuNIAR0vLGDS1W/
Zuw10Wqk2tLgDJqwVZE/PZcRZFkUASWpJKPcyBLdw8xNHWV1h3heXgke2Q8UQwQB
VGDyewh+D1gvLo9le6GJ4DuSTh0wGNtgbXiFuDJFT3Xf7D84oCtvkaQxXFtSW3Jw
alj3l6x08OzrQ4GZeNuIbJKPbCAv85dz2GCeuDVUrMGNYT9mAqy6vdzEw2GGoKtQ
KOQElqtPi63lH66b661tsmmaDOhRw9gaeFOSk52XE5sBiGwVcRmd/wP/TCLaz5SU
aOprbmleJ480ZcYp3pKn7pGw8s0vYJGqXnfMxKRd5Y6JMfyh4Nyf2DFLPJ+r8Brp
/bFm//K6ZJ0Q9KyWPiIKMVegtPT0fut1tYaV5ZMadvXM+YZCbnc8C8uaYVsJa00p
fSSEw/STK6iA+92vOwPI5OEJ/1MrcrSlu8dN5YAjIqh9q4WkyMqYKfgO8xqbEbqS
sYHYnc6RPSoXmGm8At+ezh6aJeq6eBNv6VXY2/HfX552/IcShN8T3vnWK4X2RlGZ
D/pxnxjSPCWG4l8jaHjVVYpXzl0kabsbyDWcOP71D1nMIC9+NgtNGR+PFtDZCyc4
qbSoBUcxN/zcsPcdZuR6C2exaVH91QmubR6CagXkWTNwk1+ji/x7CWnkgfRIjq2k
1/o/faKFVYU2dgpIbSWb0kpyPjGrT9uKXPMwq/3p1HrCNeavYLoj7WJcddjOhEWn
D76zCfPc6JXWjLIi+TVcLiHG3x/hrXqsLIqIncr4es2JXmgGx1+R2R0o8zCscTzk
em+JBmWLs/gqVz61oV42UfOKzLA9sSJNgJV9Bi817cRQnE102pGetz98O/2tSWHn
S+dLvgFn2uuAi0GLd1QxrnmRKp2bkRivBMqv/MfRFS1anCaY077cKT9qEt0Qzz42
1ICWUyU4rztyzXG0X8gUbmNTUtTwGIP6akfzkhuU0aO58oowY1H1BEV0jj7nyjNV
+Hvv+6f3H1lu2WbIlKObztQDGtWG5LqAGXr/QsT/PMOCvEMzduV8zTEDnpzX8NCd
hVlhOaBuhS41DCNgyb/I2duQ20vvhLg0iLBnPOlCYD6yrDTg1W8EsSYKmwhF6vEc
S8O0H79g9L5YZdc0g/MUTkAApDkeCZAfANiDxd272N+zPrJZyIhZcwROZhwz+ixH
TS0cGciUJ+j8uAvBzMHmFO4yipEgZY4MW6PDGgM0BM1Vz2WRTp8o/FLQSdRbGiLO
DvcT3pzb5u9+qE5F/4+Mocp1wz3ogDsJc2RXTj07T7lpRk81nSuBfLrFFNfAgE0R
iIVilMEl0KqxMa/qYnGboLeb/Is3D7XxYREgC3YQzs/CvqZKLZQLxHfmsRTv1VDG
5A0Lp8C7jNEKq8KUYxUYa04CWlEnP7NgAJfEJkQvpHGRfEtwRTbIPu4dunV7t7JK
lSwlU8AvwxX77mECCG/svSjij7SIJ/pDvTGdwcIufB9HqHKuAiTirXIRpEKDvpks
Npfkyqg+aSRe8pZxWMhsSmA2w+WLnYVCeA7jUgrwZDV78rslbDg89bRCJO741tq8
gHxQPFc5slUdsEFRyVY6qU+txmSXl1dLuF/PU+lQo+vy1ffZujdqFja7YRKxmLji
ZVYS6AhKiiMSDRXaRhKhEr2c6ttXTsSFuWaa18nc9Tw+LvqF+y2sk3BbUwkVLxyS
Meo+7ygMK0zQQw6Y+iKlnHxH38FcPmISXHOWFMMq4XLsH6wxJ9WYjhXm4bYSfsy2
+iaHr+LR3gALsIzXraTZeM9LJSysaeGaA/VjBll2NI0VqUNtyvfHTQ46wJU7BI2j
M5AYAcAOM4XYo2WX3UadKKQlZOJUpjvcgfoIgJcmELCNx995PQhzGSqx2PqW4Bln
RJwVsqi1hw4yKzlbRJGrcmBWFqQxuPs4JaZSllADdirgehFKGFd/7FqDVBuIGoQR
drbwlktWXHYu5bI4jYvNTwYaD7amO4Aw6SzgTU78EUv3ybRDYUcVaEGPEtIWsMGo
wToOh0GNOU7ibYjSoGa6PD170mtypVPV/TVHwtLqPye9RVBN8HQVUHG1HF8HZV3j
v0GWTF4QXbIPyy6w5YMAkZnby/h2C1vJZsujUevbUCVTk8hZuFHARHAbEAfRPdcY
8toTEauSCZmvngfyuX4trNtu+1UIHBSiogqBplNjv4nxMnxrXHcNQO9mot+Lv115
VOT+wF7atfJpQbSTJteptCyrRmgcLn/2E8tfzFNIAmKoi4UCwc5KgmlIoA/Yb+w9
kMMeoMZ8prZDnYoz83A4pz+eS3IzfCIXKP08r4U9mazVPnNCSFDZpM63dlO12Zad
sTspDlzd6Au+ak3avG2iUegFOHle7pTQLdlJTImNXniBk6Jv8VOc6Up3s9YxhDPw
406XKuiIxwbixFsz3j803eGZPYPu7UPj5dXK1jzWgPABmDHLLPZt7nE/P3iJdPlc
hJG6jB2ztMINf5LczaFzelgEWbCaf4YpvsCPlTM4y/MQWXzasp2EFUJ9xquwLZCA
Gbp0OrrIfAGMkzI8blpjODERnWrUPaN6ig99s/Q6RIKzk96rR8Fgb+YN3u0sHCJl
7OELnxYASVWwAGiXrWUoCck8fPmX3bRvwkHKNhL5pxaTZXjMEHigEadre+keLOda
UV6q6EzbYxQXgZFdd/glpwBYNDvvF6FXuQxGFgqTbSRNKD6hwj8BUm3SV2UETMzW
N5XtB0GUoWL4pbATQUcmPUHWkhYniTYh/EJb4l9jUCWyH5IGdyLFjPv6kXHHoG9m
9pzF7rjkg5DygFoAMsG5JoV53/nKKER/TQB92EfVeFQMlMAk1R+eT41wtToYsQ3h
GawC0OA0qs8vyeV6W2wf4DvDVNSo/IupmDUQjhDVY2jTKlx4VRxiLfkyVCN3nvMX
vD/531gDtERd2mblPdPVUYcEGmWShjKZhPkCpoRVgQOlzd22cJeKWeU+Yv3gLD74
G3+99/kXjtYRb8QdhAy8RNci0UTpA1QloXNpeGQ2Tm2kDAE6TH7P93LMs8bN8+l8
l9WAa/KG92yOUoMGtNNLGnBwX+38s5Xa8x7AM5Q4DcMxWXU8fdu0Me1qHGv4iFXy
YGFUGdszGr0AbySNv7oxw2CEjdObx+sdKCL7AolsX28xSFjblFRIu4kEHLDsx5D7
kBkxiDFQjWyLebEg8A+LIYO4kQfXgozUo9DMMz9uztQJE2UGv6eICBtyv2AcwdHV
PsR6PC6XtMnNnHwix81MAXfd38pHwwe3WLJyTvGIDuSAJYMcWV2ICGNJP8zedhzK
fAGwQLb+aCqdZRsqnrhafnsXg1HmQx9JNfCoLfkIl8qm+U8GCBWS3KAa6e8wlcsS
c88KmJ+DbskDBUJ5be9kkA4dec4S2atIEWFxg3sxCVYtCzn1UAJQoetDJunDJ4WW
d6Ffo2A8Gp3bcjccMOTJOaIVPiUC0w8/gdxB922NMrarB4gMdnv0n232FrNDtaBw
jxXJUXo1DAxS50aLWLrkfUZ/hDPIHDjkORr5qCQbOgY4ejhaAPxZCIIiciDl/Hu6
ziJIytice01yvYL/ibGO4SOcnhKz7B3qGxms1ngcm5IVFP9oLLyxvXX8U0tfhXGP
kZwUvTAyjfETafxBNveBCotUAjp3+jcVZ2nBfyb3oSX8ToOSI1fV5P2gNMR5MU+I
Diq76XIN7dDzV7BG0uKA0j5XhGI0zFzM6RKYvpRrUsGszXbd7C54ZHNMmj9q83ne
nT4YqQeIB/Y7l1F220wPWJ/RHqVE0zcFhoNzXpK2zxPXhv+WDk/hahW47RXbvohN
xXvshqaT+NPoNAKVtc3Qtz0lzqKbeSEmjAGscF7IDcZXHnWlspxY7alFZ8z+ROlm
AlQnNLwxJKv3H9Cium9eI6MjYcyKcxYY9xphx39/Y4AWcvydVmI2igheJ5cCIIg0
qc5YymRN8gGxZ0A3dUJfRBWnwTwBAvlJlFSNoxLnQGQ/zWiHKqoEbIfM8jS2iWvp
WDs7hO2GL0TvuuJ3yO/NZW7+teXPdjuXHrKBFGa+nkOOcI8ttMIxQzQVZipJaG4v
9ZSrXz470JocG9MqNhsPTBCJbElY0GMG9R2Q2hor8joj5Q6jL60J32iHJ5Q84b9D
ad/rLKJLr5dk/fJWm22cUirhdhwTLKF+x3n3OJkZXCKWNXMkxu3zCfvj2MkyBBpq
E2ran7fncSxcYwD2QD/KzKEL3Dir+haPXRbkhe0WgoO24eoaaeK+A1qAJGuEqhhW
tidFrdUwjnp6J5f68A1Oc8BKRcdpd8RL9kgv70FBCqOTo9xkUKqB+B/+DBATsdrI
dJ1JJ5qmmcvWnPZ4Og6VDibDYUIEKhj3OBn7Q0KmDgkfbrsu5Pso0WBCPh8I/0HR
OeVnSFwvgVG9ZcOe76cbyp1M+cTOBR73eCF65FlxZ4dPjUX4LKBIey++fGYKG6pv
8LjUv+DVToeDY7SLpTm7e/+oiP8k9pggEj8f/8ATryLu6MqI6wuMZ0z2fDqqKamV
cMi0x7vFbdSQy2Ko2ZAPjQiV4ubjsb+rfC01tlDYcwLs2bzMOl+apYq5Fg2KEosr
KGaAby0K9BJCduSM3IfkS7p306hLIf+4Dlbox5LZdq8RzE1TPO5AVRC14xSe3Aw2
jpGtpj1tYXl4eoQx2Uf76nOwWQQkxtP5GImWGmuztiYofajWWauFRv8m1eYLDuy2
7OeZBeuTQ0EIw6vaYiAzSLu25p0eVOHgV+Ie0tT+zBuESTDBPTGWqDlH5hHIcRtc
3+d5n5t09u8q7TvAXCjl1rBQ0CBsKb3tzrthfuPHDsdc1FvEPLCmltT2rkTa0Tew
m4LClQe/YOqP3kmdKYfe5DeDz0Z4uXeEB1ERwCupFYGfbsFW4TSYHQg6/j+QWxFk
WqHmNwGFZzJueMcmQuAVpKyU8U34urA6dVSykehaXVI+tEqBsRZFnwxq/dJbHFWU
IRSmRkc4XHlIX58ruGbS1fX7a4pnQjkQ/5RfWbFDDWQTbSENxhigMivvxaTLoo8h
dinJpfemoAqAae/7t3Ych6BEbhFVHp12IbQ0iO+Mu1lpzwQTHyQJAgYaEcY7a0B1
SXcl9LVmxklEYbvMQ/F+DrO20RClWD6cFCiMRrkUStTbVZQAs8COsp4l7m923dJ7
nTGmqDKFK1BOG8aew9V5qqtYioZB+U5M6C1QhmaVfB+JhS1lZKhrbjzZXn8Yr3TR
qZuJ/Df6WaHxkzqOx7179U05X9sT7a+5hrqYS9e95A1c2ogbHJ7DCjfB3u6MxOkh
dnQSQCGaubQc1+QIK9DkRWcut6hTZ5nWiMRAdwomCJS3hCeXCAi63cJvv2/jwVWo
jn9eaqJ59e2DujBl0GnyQn1DiLAlcBIkwfi52P95/2n4juQIsEpVhPI6fQmU6XMb
8ktGxCmnwnun+gkajy+g/hmTB2pOweUuft3n/vbo8J61L0r9YFCwUbjpocelWtza
YVetcdGGd0djDUwci16UAsGu+REmmrZmHnBe4jeUfgP/p0QKaWe6gwUNyEzJqfu3
sKgRqDKbwxBMLwYkqa8k3KxMM/o49/Pd7inCOfFbXWR3TgBfFWo/a4Dw4FuAMcvr
Dd3VkB1y0ID3Vc4T1lLQsfJ7Tg3f6hk/1ibvxONLLjmbcK62ErFf8x6PKWI/h0sj
GMV66bj4S5tCusr8wrbshnamSR8d8fhkNFU9tpop0fKy4NoPKqr15l2Geiz/EqFV
YSzzg00xaL1XXlScxmSTHE1CVn4n3G5Zd8bebCqrmgFbzv0NfonA+f+fdPBHkp64
EcALHju0THxRSE1RFCqmKMbgXTmaeioQNYNzxWuk2u9fvqUGwnxL7FiHYig7Cpu1
VIK/d/m5AZwjvT4pMuShHHgZxmxtvecC4VW9obUvkk+x7jonVh556wcNGtRRNVt+
51vDZoFU40kNUpeHpisceI2N84Z9Ko3Zxu0Q33uYGlCAx17w/fO+BCqBGF0JLK60
m6IuBR6+Vy1+cWBeJKl/GQDXElAv6tatO8uSBvvQjZsLOsDDzIzie10ce8ORrEat
9uQgU/5WztNDrsCsFhQxnAd66JKdAslZ8awx/iCyN3jVnUG9KlUeTGfKQLsZozF7
1Pprnxiu83sgsKAIudgTaUWgZpV5a4AGQu7VP70oIr8Q5V5dpqv9oyAuaXfFqzrf
S5FhOWsv0aHYWkda3JhFzVnN7+mDqDpesnlRwmj3cxkMqGtsZbRbuSLu9kOlk/Gr
uunIrjNP//kKkhkgYzKNcpx6DsS/I+CVzXvQui0K7JUYrzx/ayWgfeR5x+jEcTDY
J7aanYquEG1zU/vvlODBHsHwllaBoDoJPjzteokJ/cOg+/hfE0eymqPBUWs4cUfa
1I6S0LZ7dchofSjw122zWFmJ/8qD+ePTM1EJVuRkQbkqRJVDt2WEaNgEJJxbizLw
0mkk/p1kw1Kr2Kjn17ZOQSR5acP6iDJjtSlmaVpASBNCnY47p9OPSgE0ulF0AKWW
OI6K6WL93yNNrO31RihwJ11aRZBWsfU0MGgh+JtOKDGYLj1dIOqsQJR9cLkELXKq
igY00rfGIPwAyIQcS6R3PK5f7PJjIIKYpPaDQZ93cVchyf90wt2T3gmCDm5OVOwa
uLnQA2oqf1OVm9pYlVwvzIjcaB+A7YHjZHUb80SZj8G2DXzFwuKKj+fUv2/kULPD
KCWqORmfAShkarHH6QR5I2qcIpXqqyJ8PjHGf317PD9e2R+JGFevWwcXe8GG57mc
UxZRmJuzV6q3Rv+aZxrs2F+P2M9U5l3LlOv0KiaXC0n1DwYu0weUqlAdurkcOQJh
zlcc/TmiGs/GbJ40vZr3hJ79MwpBJ732bDxO2Zrtrw3bxg267RrT+1ZlejqifH6W
g1WSXS4DdTA9s6HuUKksmRZ0Xu8Q2m14N92yPQ9tAgu96JODWHwTXmOBlG2xqG6w
oUhBb90G1O+xxhI/2TbntuY5QJYm065a/1q966Zio81p6suLuZZJNLw3+YsT2NfA
qsMo/ZbaaqpThv5cwN5iUKBso4SFNmOMvO2IIXrJ3i0fS9d2dE2OHOPtSlUj6RHL
tNCsSG1zaOuTSPZviyN5E55/IqK3mWr1KJMc/WmlFtEm44gY/ElVL31+2IBGRMdB
kKDm3uewW3DvIz68UA0hAVxoTgABx5rtTqrwFHl49KzBOCw8UAF+xHE66kKIlDpr
3OmVno7DVyoxMLpTQBG8UTIoVzKTGrw/XSOY89BbdntAZyQba9b0/AMf6eXWMPSO
KcuN+1igsVOdoiG03szfoxKY3fd+jHDFJedTBSz17mB0kWADgJE4smkVI4wdLMtR
DcvctHf7vALQQ/KjQA2/q2MjZR7/Tx/CvOokZtXYsp3bGJcOoJPqYvrkLpqMsoF/
7l4pQD8xrOz810U54xWut7e3VXN07iladwZNEqHi5XUTGUj9cqA9H/NtjpbL82Ld
TjUrjzrUtDR6yVlCUwxBNEcPCkVXT4GMsJ1eur95GFcQN/F1O429CqgfLt9NVPmQ
bHf923uMAc/SLiXbuZiRUHCgunaWRlFEJ/GC7qTdfufDBuRAxIsXo84wE3c6H1Ul
5eyQcB4lDRbTFL5rCRnpvHm38E126c6GHc5pO10VpynhWJW+TPB52N98oBqyVa9h
d/p2myPs1OMhS/57IXGKmVymudgstN5jIfekC2dd+kY/67h6yYfnoaun9uCCnm1z
svRRZEni3lFoOLIPXoc919jTdzwSazidtl1ANj5NpJMESqv5o2K4YD9GTpJwNupv
9MMf6Xj5E05NwshoEUHxJZkxV3K+E57lAvSZ1WlOEDBFf1JbAKjA6/HzEiAPyqbA
kU3yl3qjXPoeyCixEHOg8LQNBMPrQ/xdl7hsMYbrPAPY6tFSnwUEINfEufYVLBdn
i3asbIL9uXZERGLBmNcAdWfE2gXb8abzFgITEufJWGE9vj1LJxHJVqNpvFSGmYH2
l4E5SMv7Yd92pKOPZKzqQwIhndl4ZlPRIz+T/k11R74z0OjgYtyw1v9L/UJPBf2f
GcH9PJYdMmu9r4rUVF2vWDc+XeGd0lFb0P74NDhRhH45SvD47LlepdJYw0gIA3yo
FFXWcRfThb5zv24xkXY5TcI8SXpUXRJzDqPbo0Bs84/ADX+/kHU0BjJPFyByQq82
Elsjcemiu7pnirka0r21LZm6jDWo90isZBiv391MPjymGcWtFzUFzJ6v9uEgaTdU
8FFb1bPa5/uyIqhmwLLVR9fYwtCmXpCqhR3VqkRw9FScGzGRMWzLFl96JbTqifCa
2/FmQ7SSq0vrWtXr30Ipt/dSfEYKhohLAsSfGl8Bmlv9kfVb3XCB72+pBT5Y5bMa
l4X/IvcND+kv3wyKQLeM5WQ9ZKj3l9xuWSOPZAYcCKKot3WPpBIwBg0TV4FoCf5F
wOxiTw7e0HnjsyUp8TH6zNiJXbKVQXNB6QqBprJK8FJkiCBYL8T4SQuost+HeAb9
Kq4JjD0+pq9t9otxufbfkOvxt81F/AffMfiHgKgyrd0WC/7903xjjimqAIRGi725
P/roliyGIDl/c8OhOQZjmWg3cetPTdAs9klHrQoeQro4viEKzOivgGqUpzObJIy9
8R+jcygNkOQ3qoxPSpf4mPY5skOGDZ3Rq9pTz3BwdwVJqeSQKhx5Bf8Cl4yxNdUF
4sazQh4vV55jNpULJ/J/ev21fBlXO7te+IZlNZI2D0R9lo42ZyE88Y//mS+4g5Zp
t2yk0PRlGqnTauqRdenAT8xE+igqB9jcG6f6iM9Nc07V/FO6Y07DxmGgZt48sgb/
M41mdJqX5GMW5JgR3nN5ZzqUqOBRhSUrQhHnzuq0OS7cMjNlVfH3lALVs4sWjdFl
262ITT5UBiBbedVIYs4eG9h/hwNU9xVm5ASmhDWRsF1IXU8Fn9yZeGfT2uNo2fmU
CJ7G8vDnAXJ8KWgqU4LqWUfpaU2OIvskRYEfXEBr3+xjeXx842orCKM83MT4OjUp
j5SAKPyEjp0djMmt3VqoCved11lpDxd1m42p9iVoxYKarH1ISE3gxSqyW6U7ty8z
vv3FvaJGme2ndt1cQ/v7ZEiJG/U2Q1VyrOOMedl5E2IsquVRzIUHTm53cuUUVLvM
xeNDCMeAlEGDBnQpvV7UBL+LVUOIvfBiw7XcJxDZ/Mxv6tYUFLFIj1Pnt9OqEw5z
8YC6SDUti9deOs6Z6PXAa3gtUR3FHc9CFO52HEo4YHPOp7HREB1E3vZTQA9QU8px
BfM3I8zAm3DrlGwVT4wBzOj0/MHtVynVCivwQFE6ItN42eCF6J5vDNAk+e3577TY
8rHPJ+L6q79cz4ggpnWAH8ck9+4ehNen6TAxMTdLWZZdX9edGxl/q4FjIY+7gcP8
N6qx+f6vOjk6NUf/2AKaceh25ifHdVikYhZl7qXSXIzuO8IOXX8ThKSXxwDule2Z
T4VYxIZ1bO7aRbDKYqCmhjen1Q3GlarRK/hyz2IwpnAHUETdpvU7y113gtz/aMlM
j7PSHf/3b8tx/gMD98Psl8lJnEmP8LGW6fAIB0TR8fCP1CSi666DOnbxdLJ4E2FC
pXFaw7z+FEWpKWbNovqYay5o1eJGfdz1oszjP3SgoLGv8IFSobg2xIvWpyNtyU1i
HcyOp9vLVrDIgnmIOvw93nX+DwsbZprPfUQLbM6vnV2RUCBXZbHb9pgZbLrEVTLR
N5HmXxHbT1sA+ooQzPMjqL6jAHT9rCyjCDmSVYEh03Wd8d4MINDuwijV/6yFc0CH
cKUjOEGVyhzRPyUbok9eiWbjVf5Fscx7T3fHS9HyXhKrrPaDNMVVRaBuVZ8qxhGv
RDcrKHYUvJbf1dbb330RN4336lLImCWA/vVmQhNMkpnZzItLPLj0VH/8ZUeaAYZg
A0q1pKFwb7HGjkRDmFagAKp+o79ZKCBVmK/rVTDSYpR03K9UJS7r/6xb6gerZqo6
WV/GrtdcUDzBnsb8/raXN2M6Y7SJp6Xrebs9CK7+xVkIUfE+eZhbcK5ApORkYK0j
nQsxeihsHd8HQzTPgyHZBLoib1rtlLy52dy7gvPy9OPQY8bHIaVOHSeIiNDwQmal
ToVKd8xoUZU/0L9OvvTZMlrpj7xWdSBbpFj626t7M3acFIx6983llIg3tEaHpfIa
9UwNrzLWehX72qwRivZOXb1xbtzQ/KJ/5DM8VLFPW0cef6lAPcOzYfmXw8G28NlD
GMyxzjsyTZEuF1O56MggnIm5bI13H82Zy6a65jF0GkY39f+SHN0oO7Lxwhhy8q1p
njbog7cLsbAM4X/LMS1T6UZzcZxjgn75356vaYFPoUGCf2NmKaZJI9QR5Wg2VPVI
fCGJwf8ns7nZ0szecl+HB3/E/K2wL0WpOAAIFboQS4XZ4Vqk/HB5DAc9oymoAFyk
tfWYrQa7DP9lh1YKFKQNr9eBsyE5RL7szIdBO/yYlumx7DUcWyt+idCYGVr0agMr
S2RYeuzaUKzm0+FewTKdXswEKnbOOW4afJ8WWd4/tI5FwCOlFDTYqxvmBUIAyuby
jHmBmlYvkuhJ7iLJUrXZ1ASPCsaSglUK2zwpQRAgXYvulyAm+YCr1ToMj+PmXUEM
I5zToMPB+b54m6JIHipD7esllHQOKPh8vPo3z/WiTo9Gae0XIxfAdbX9KDg5VZ7g
Isuyortx08QV07q6wLcBwgn5Ec8+2hF96IfjZhPyCYMNY4cxUEU/yDEeGRj/9V5M
Oi9udvvvdCqm6w03Ayhx9jOAsaLIxB5CEN/yOW6jnbzzgqzk2OtPfK2AmWTueJYI
NvLmYwloBWFs4F5cLfgU5vo9AY6CxdDjvQMQ18xytR4KyA1GATSf4c8E4NpnSnhV
HPo9xKqikPfGMwuBJvpLs+bPpDHUHbv0pbdne2mgat6JKgquSLs/6AJt3nkXV29P
yKVyxZhWgdp2SdkOmwHtkMb6yc9OwphHYNxyjHVkJ8YGBqzsXbv1kof82pl31tWb
TCWpEgXptDiDRzyDe8DdpdXzzCiRn4LVb6wSbOPubyO/3yd7b6Iko5Lvd4+DEfLM
q8nx86wOS6fKh/xXfH0GHYJdWvgcUe0+BfNMBRLRPlQdTcoEYcyK6e79ZtvvMkUm
OnsSkzHXdkDv24ZGJaXFiBUAuZWLl6zGASttzPdPqDVQh2WEQ0AbKgQtd7WN6Z5+
4XYCsCWQHPqZIdYhmZDmEijJnZ4wyAqAwJBhdBIjonbs/3xPHTK+k7REyJ44OAT5
Z7NlS1Gv0vZ+jM4khbGxCtNYxbMAbSmJ+4Qy4gVlTVktUcv164GfuBrmz6JBZ8O3
66Lz6AQ+27yiHUSMTlPlLLUIzBYDVi4W35ZRLIl3FbcafvAP/wcXrMPCs43AdP2r
0Me9rTxLkkORCNo0uYuuZF/LZO12tHHH1n3FB2iq0IFuXRcG2Tm7CWPumwnXEyvo
2jFIeRWTJgLPaYgQeT5nU2WBIt40tSRAL/7cUV4ze5WN9mIfaR6IIUk7bt/EywE6
ZRnKdxff2Vm4PmyC+dsPPnF+wPfY2wHDr7+culWOPUZj37JgV8ra4STPCP69X5Zs
YQz6ciknYKcoCt5hCoK/TWewcf6LimtfUrP7MYETdQ/oP6uh2pQ7Tl+e5dSR8piv
Xo0ePLndDz/82Z95rVs6N6aoAiLBdWSWvVNB903eTYVLnoD/4NrZTbiGPk9s4itm
URk3OE8dcIYzfZ4pRMrrhA7yS+VwkMxzYZuDv3y+aRVh7BfHAGqVRBI+jcafoPCd
IR+7ZIB2Z2nd0q4lk0Aw6AYwdGg59I5d8l9wpPxJlETw/LRHKA9D0Wzg/6qJdaZf
4bezhBwT35ISd8ZaAPkc1sRsjQiO51CBGkGKPd2RQm9Ow/TMu241cvAWvBZpT3jf
Fkk39bIAG6guTvjTRHYsTABpawVEAE7RzOxGkBQGPt0Su2N7kDefBYbIMTJCT9Sz
KGbhlYoUuV25E1WIwiry5We3+lbFPAfCgTVgQd3sb2/bnt9iRzbDOO8r8BDJN4r9
jm7EX93aM7pDC2D0kSQnkLyI3QLpidh8sM3OYrsv/IMNVc3dM0r9+lzf/7ZtXc6p
bwn9fGVtq3axyh7jEfBdJQ//R4hShTyIHxbwxlKFsuEEhT8LKP8vAIphfcfR1UkL
/GJOpyUbyIr6VqA3VADpoR/qiAkYhAs+KZzlxw8ybmtDdyFvkoxwo/4vW+bsKVVg
PHl6gjNS/aK1mPsMLtzDZsm1iz0RMqCcd0VmiKRpPBOkMz9O4QhLug6wve7l3ldp
XErjUX10gtcLGY8OQVFTcj9Ye/9aOhm4C6muinmvPU+1KkAWNy+W1UXS0YCOCsPX
BkpKfIc3iWbXEvFqDBtEgdWgUxmmgCJCvsnk5yEsiFBVPswazD6aJFzabuD0YxsG
vxEpeD0Ztcy3vyizXfkEc9RLJmyoMbXdnzdX9M5rF3bIuMadRpf/G7tVO9OE39Ef
Y96p0iGckiKLYaPJTavr81Q3/DGi347MdumqEIFNaxiqOiboK4pzDWgnSaEeFj9J
8r95tBe64o9u0HkEZlbt7ioJDZfLSv4Fo3PedkRVtlY+66FXioLE370GwYfwQwxk
dfxrd+sWElH0DE4wsjrt+DrnYlxrVlefynktHzaw4mSVa+AhfwuhKkvH6+XHjJlG
hdmDiMNWUcBQHkrGkb1Zc5djyuC9Vs0o5/M88PthR9NMcse5P343pyw3Qbe+I2Xw
15Mi4Q05caCmMMhwNRjfzfwJLuNjdCxOQObBWSC9trQ/gzOIPbzpzrC4/USnTh/a
5w0v6LhZ/kEjNHZipev9a7wss43C1WO32grOhwyHXyx0bVh2PTa3DpDSCuJA347N
taQ52hTZU6bb/2dYUo2rUNB2buZSKlfGsPk9shan93AKIE29fqPhu+z3XsWM4tCR
71Rt0Cq1pYUrKXHzr7WVEBYwIPPesrqLHej/1ZOxuJJflkNOww/qJaiL7wFm+/vO
3fz5iKgN1JJblxnWtC/Z7aXc5DdhCLcJfjwuuJE+uLZBeexSI9MPJoJkGzd1BDl0
aZoS8pVsal7tdBgZ5qb9Qt2E3x/m7mVS8Lt0pW+CajHNr927p+xzHMCEXaTPyP5B
Q9ZKwoW5/wsGgTYKUtnYbfpH3smlD2FEi0BmMgO3vAZswTa9vAUAplSx0foQi6mI
nvDnmIY4obqnaUJJMNOylf8T+GBvLIqsKEUG+KEag5Iix4xcrEyf8fkjPSHDPi6t
8SvndvcpkzCQluktjyzq1k7kaFXL9EyoaSGdFFebKZChzjdS5+bBzBLMfE5q0cjZ
FV/39F4pO2JKwQ8fFMFfHKh8MMHyExb7V0c4AnNIv3KqCKMs4O0WzV6tGCv6DseD
1yHdeNH0xxPOK3F1dkVwCXMFSsFEI+y4d8LviFLDtJNkCZr8SEk2OpCs7zFkC054
0Ex9i4SJ6KN3IDgeeu+jZvj4B/3uKeCzVea1/j+9oHjyfQtzwgBNOUw0M4/u4TQ4
EW9n6iOhNSkKAAa5kOyE8NVBS/ePbj2E3pt8cFRgtoSvTkqnYFn7OocJUkZpcIZu
4SfGc+7TbClYhhGsjI+L+gok+A4rU/iWURpFap4Ig+3CEj3Bd85rBvL57mpqmsDk
DeKtS1wZguro2s/XnVOGTGY2pSAxwTKlM1/1SYqM2+qlHAtrh0EArZxHgURLSVjR
SRda7uyvaFzDjhcj0hEVOi9+414Jy4zVYoDeudxuh77T48IykRczgUMjbOJx6qkO
/gBTxEJ9IpUH5iDpPwPtx6geqf/cQ7r4nTR2KBmOeeCEURgkUFvLnMfvH8bzg/+S
myMMhVbxbXBCEqkAtADgOoqQpa4/6hNd3KTRvSQ5HOTIXjCc02/rxWvYq0ChZWYh
WvPASYgOhT3N5ur/rUqTCJvTs09+Dqlx01YHYGnJKDazdZApfssmsbHk6V+lVZUq
s4L5jwTN/fiLrX2AT+hVxqrrfxEAS4AeOWq3TMzeNGMitCrUyePg/J/sQHjOyMXV
8CnC0+Shz+MeAw1iyfHjSgQinNxxRgHYPS8OyhqSKsBZ4DWXMLKaXJAoj+Bcdbh4
qHvMKJMdAcWC85sgon8oQfPxh/GNK8i14L4tmUr2SQdBlCShwYiGVvo/INd0psAA
qJw2EQYCdaDuQceJKFDuw/l3AsYGwqmIzfZzTFHln5ABrlOJf88aYDjh8+9PMyZX
fHSbdLo4NuBnux1FhCn+bOwVI2NHjumouBJUZjfgP/f+573TMCCt0OvxPGVgYn80
AoyAMUFpi+LBWflNU6VsF2BucW+wKo0itZX8EetN6DQcwcXoIQNqMupXwnEUzbjC
Z8vKy2mV/qEcfYed/OAEPl4jdea0n2VqTk4UElpaq+Jg/groImpIlHAGu1RRAoTQ
GNFBzBs+xOlgFeISEqFA3aNx9dfl6KTsPNT2/YSdeU1QNpap49qXQnvmGd1NU14a
b47xq0C2IOfzIF6rXzx2N+uUclROESvCK3rZAVoOwmZzVjFQGWpqcyJC85pZvp7M
0spcuIUxasD8RdEJQ4X4+1VSJZpq5AaM8Bo7oFwkTcZR4PPBX9AuA29ahWGPuLIg
JTdB1LNWFWtYG3GcUpl/DjirC2xEgD9TRtmNhM7QGmZu8fb6dGiR6S7IWDkY0brR
gSBIQx7DJkmPhA+MNN2cRv1KcJOB/uPUzNwqK4dlfYlILrAiCfHMq9sJpGyDDi6r
FvhGUE7lCPQJVICCbNQ2aqg56ERPlHkFTzd4M8jGkhVmjqQjMnbayqKV6AvdTBir
vOhHbJ+B5GU2CSP40bUdcikGegBWjS95O/gKEDF5+PH8iK8kL7tQHl2uifsQSnh7
+1/JzPxiJEvLn/5T3yCvJstqH2yB0ZMvr4hlVu+i7oUbacuTXnPUejpE5wMSqKiX
FACDMb3cSHWSDmj8AtNre7vqoofzn8Pp04zq7N7Nml1sbpgnugpkTWAIvUb9fJta
wA6HyfHn15PP32vYowPyzfiWY6FjtsrGTlMG/ngtjq7/tmHHbKgeMFyQ5S2pdT+B
EYIyu3mXgqYjjxOm5KVnAehH4SR3NXdCbxVXiQPpunvYWOgbhGF/dujrKg+shRU/
N8fT2vn/TIGwz2b32lHDQPX9cK/QI0uG5r1gWP2PbLBTOtmNCVNMQ14WopycTwtF
p4DOU0qR1fdM62DP6C4lCTkIWwg1kbNbveTL5IrZxmqwNgkLeFY2aJjoxG2P4A1n
Y6Te9TGxcFyoS6GTLFWbOPDanw3M9iDrDauvbeHOc53DwJceW2nD1ZkepKPcp4BJ
gZbnnblJZJB0YKSGe0kdYXu+edZW+tPs0iTrMcpzbGPZ2MGXpwW2WICehWav8mSi
vYVUwiN0gLZw2r9P+vT7SlpacfevpgWPQLVDt/gr6435T24RjfhsC9NBX+Z4QBsJ
KG0pXyj5BREKoOOkd2q/bWrsQTVprkFyu/Dvw4vmaLv2/hiw8aPXAmmBXlyuMK0H
jKNLeocOOvcmTJP1IVAByibwOBCG4tIZEQNuAff4Q36p2Y1r+QnbpDG2ahzYTaEk
Co47IoNsd2wVXqqnmIDgfUndziAOCTRJha4l2m2ELpRsUTeUwDlhllY1bg2J0a7b
e9lFqm5QOucWzqyyL4uL5ZtAn6dAKVCbhn83K3RJ78hEC9+fBoWt9dcTuREUBxu6
4Br/RAsRqHm4HJDzA9plZ6JIASjk92CqKljf1ah/mMfrHF9U6bTAuwpL4JTHvdeD
h9/Wt+T01Y2c159IMyjXxhqLaciCsKyHAzkNTRxzt4GhBYt4Qi+jSODuCDCkrdZB
MTPKr1QmUrPh5UlqZpiHPrxG6nmWbHZ4hPtIsI/Qchk1sSS/i7lG8Jd10ZJqAl/+
bDQ4ZfUbg3pryzI0KhBfUmBjRKRgsuX+m3C+0yXjcJjZjGroXPPZbeDtoIWWqJqG
0vl+ohZi0up7vcIETpm9JPg2YjzB8A2+FwAgcfcECCYhr61tgEcyZIfrdfw0Qirc
RQhiVFf+DYSHmYcHvUYhG9mZuMC1nj6QhM9385N/4Zy3znIVMLo/JyGdKPHNhpJ1
zJ3jqs68o9njy0NbkPGdgzKJzVlmLGPU5DaXtv4YFNAoDHnsKJTzcIolgC9yge9Y
eiZmr3MXQuS4u6npRv7iakchMfCz4r2PhBy9ZDopfuoDWMFPGZhMNxgOgfiwsSPN
b6viFJNFfi44zkLqONeuDAiIT7b31wtweYAsTI87Sg7wA3dJcusy3vtTr7IaznB0
aoiHPxF7nGO62NNp/W5hGysM9PFk3AiydQEt88Ns+hYg9qlQahoSAo09JbPsywM4
NQUBYrfs8Pc8ZD4Qm7TMmozIl9NVJ/ewNaaITGngZKJJAR2MD95x4Xy8gGrbWUSa
1FziCcldEhDW4P/0L6n+s2NUs5ThBK0BiaMrDs3KLuAZ2rKmBiLRy0WcSdIdapjt
vxJAU97FXzzRFKWt6aMFIGBNA0dd/NWSr09aHtWpfT23xfgN5TvDr0jA+G1QO8DE
KskbjCfNVH/bxtgbPKNw1kAKC5ga4K5Y4Tz9tfEqIVdGx5jZc698NYtJcIsOx2RZ
pffmH5vmE1x+OG7q+nApXaeLrAVKQeRPdJhG8p7K08+UJ4k2VGfwrPtZNXyzLXu3
ckFdk9Q+XZT0Bh2hg6/QP+Bpr/ckrLcesPPzO3pGxr9bis2Vin0pPTq9px2Zo/fz
VuABMcs4J+12nmk0Bg/CJPuv2XUgoWLKGiG9OUWKRze0px+HxovLhrSl1XEMntdc
nQ3LSB7WakPtrQ0jXdlDBpDusVwnTlWZN9aG1wxK0x+PRU3otjQPIwBbBvmsMtmK
YQx6rePmGhmTUdJbtcbIWVt8oKTCcbeT1LiE4OF13AQSc2QTQpFeMqcHRGFSEMvb
piBVfqNxezWTD2ZYX92RwHXkYquusrniTMxNnXtY9ygfQwKtlgo87v7JK8U8n18D
rPOqs7mZPaSGbdr0RhmBGgzeCAvvYbVtvLp4BYFDZuqPkDOlS4f76Bxb+cfTDQGI
S5DazmOpYbQeiXR4+gv5nxWkipcMTG7xhxF2F0tCZbNqg/fXq9QKI35S2poKQA3V
nCrVeKjW/k/CwFBIUycZBnxxwQJTjMBXFB6IISIH72cR5OsIDoD1cBkwCvt6W52/
S/s7HYQ4IH9374rvkiCyDsJiNhSUimBhOmn2X5yRef2j0vpqwpnleZgN0DR4IHCK
WKemscStNBVTbdzhFO3OFH4NOESwedbux2CEHJNP7oxKVx1mktqY7+BdpI1Xu7AV
rcNCO3PtH7Uxjkdmfi7+rs7yPOV3Qln4GlE1ymyrsRyZrX4ufNHJ7Pja0DRCHa6T
iRfZAwMIYh7U5n053QlqmrDs8t3SEdrejpKRH5Kb1E/Z09RVQWejITYXhQ9o8j+L
/3VKOvJNMPxRxMBr6NaLGmpS9hHaFGNp57xqZHBZnJ1V4D86VPJJMD0aTqOfza+r
wVxns1shJREwyoEXm2zVewIOl1aJkFXDGzmdrw6+lepWb6zDv6LTXM86qDm8AQgr
I+6Zr9ouey9bPN8MyEnuRyQ0+jZSDKRSp/ndfJb/4tcXsBvhg64sVrufKcnjlONJ
BvrDKJ9poTf+JErrrkZVjC8AQSGA21hgKd5SXv+Jfeot0E/DQpiYoj1068qsaF+V
U2pNK/HN/ZaIX9bW0FMRZ2Z2lXgw20ncAZDlA+fiC2fHZ+CVu4nHoDpxWCmNYDDO
8bx8flNkYGX11ac/f9aftBQ+ZVWB6VvVzgkPHaSdxlFf8BTLp+TEabmwxicSDEEe
1hsriUovYkf/x9BzcnkMdbpncd8TTIdNL+aK3ZBojLDIBpygmDbnNW9xR0wIa4SF
Wcs6YmISz54jbRiHrpqML9iW+fsxU3Plsv1dkvC/w4fayNUHQzhKbIGVoY8awJo5
2ZNhsc63+VjwHHgZSmxjeRmSgCL7aKBhH01tBsCsKGyOOzahPTYg+KuK1aX/tPXm
wC5MbkvG887uHC3PESfdDL2/LIW/EHDlZrMVqJIj8Lz0bVSyCsSzbytK2oioy3xh
KlMHH7QS5Qi2dfN6Z9QcBCCH5EKQ/zyy+N2E4+bhUCDeN50E2863eFxHB4q4q4HD
Ee3VlpFGN3O9mhUyTwoEsN2UASXxzquPQxz6GDTOy/nGd8Lf/Q5I7L/bruTWdYOK
M07XbkK7J+MbHDfpo54bPKtkaprKeLGElJclKEzAhW2U/trHB5acw64Hmw0GnBGw
eWbp+4szo5aNIHe0WaxQfFkPueloSnRYwTw1sdJduEhnzGH5dTVZe0NL9DHYXVzE
ltgSx8nsFVctVmW0Fowlxmh0Q+Nm8DLkUsBlAVz5jLmJHxq6gdI1jBZ0XxeqEaPN
fyo8kfBJFURVfga3w53ZGtXm8lw8RwWTjiRelcHkI9k0ZGQbPp1dFb0Wg3hwYwLC
8XaeGH3Vldpp6yPtf0a3qw72PczBuuRK1Uk945bOk+bu4RJ14nGBYE8f12aBBvp+
O5DHRXD9J7qewGgaIR00FDWiuPbjk7Ywm1vxXtRR8Rm6QTIGRiOBC7oQMOocP7Zl
CuaYx3P+FXFLI7Xsj1rh85xSr+Qt4yjBYUeHLHcRU79NMVC6KKdgVdSlXquttDpx
0QiAC7H9gcyWTdPo9N2Pe7curoe/bDljGlYWKSm2P0S0ZAPbovFzhoKUIJYpFHZs
xKU85D84awvlCfXxzBMlhxrfzCCuyrgd7VFwQWAzh/szMiUDHFQWi0mf695ESCfg
/kYLlb6D8znzx4Fi5JIYyG99qxgaW+qqI4xTnqOkfeDImBEaVG5/JIi9VtKER2Ee
gtsAMcoYLlJNx/Hi52ftL9+HzX8ImrrJFTfpDzC0bypVihIYiQJmPUcIz73we5rQ
QPNdZJIxbjd+8Xy6pJchGGBTf1Yz2dmEeWFkgP6XXKKa3zkuABg9FBCNf42wyU9e
7bhlv0Pnf/3ekcyxds60uUoEkGNFw9fCQX5VuEnqmSQ+dxJTvXFrVbZzfzrlhdF8
/pMwFe/MPQjjI3dN8mU4yqyMVXGs7UWz1Sj/fpIsy1bo7aRj8woatGKbFf2+vMv6
7MxiP5UftwsZfg+QeVfbtoPj6jFpvLMTN5dPqGDdxBDF+RtDP5Soba1sJEQDOm2d
5Oc5d5tfM42loWYp87eH+iHGMYGTGhk/Cn/59cs7sblihohdcSTd//4xZJvG9Sza
9QdPfrLxsXrapzPr/sMoJbkDbyf8qewJ1d/PaHDmzMJJ+od5N29OzjF02qRGO47Y
PDAPmKKFIgLHXJ2EUgKNj2kpB2vYTQMfFt5L8zyTr8mgSmP1oxxxxA+3VtS4Ze0Y
7E+t6fKc+B3Wbd/Ehi7KfgDgmvMDkDqxkIxMgAyVoKJFK8YrgsbzHfV2VbdyFQH9
I7DH1h14sqqyMOnrvs3E7yjwB/maB2NnStGVAhf1fF/o7pEXwxQ1nnHU/OFb6ck4
Iq41NGGCX6Cp1GnIWuqAVGJeJ7ma1rfpOzN5RJX+K3z9C66MMfhAtoZFPv5svFbj
zeQyCQgh/AxiC7nhQwZl9aN7+PjZVVAOD/x3h3lBJF/vgtXlRS8ZvZf54lzEUwWC
sLVOXOUWH5lp0xXBud5QbqnkL1n2nNqQHckQQYAYVpp6nIT3wHVXY96TaipmqYoF
+Y/rzyOHRF5rsLD8fwr2Q0Xz2OKJbOUr0VUdrAS6PiL9FBZEcYTkXRUgDDxl7RPO
+FgJvSKraHfTiohC8rpy/QFpvHm9RIdOSjVq0x3uIFbiVtCqFRlZz++3IvA3hKbf
yNLDqwZBww3Bf3I5W7BYAUSITpDxV3td+lsE09M5S7PakW2LjGtgZbxA4ZzpPBlL
ogsReUWRaiyVl/P4PFPidwxDHdk5xNdqwYq8gH1Z661HJpy/8CLK+vKqQ8EyZU0S
9fVnxwQFv0iqOknP+9JPTgNHvRWLue6+uGJ3q0t9fDgFMzDGpEzNyBspk7zoHrsj
NdtWAyJ4zNsntrxP7QTxmPrdqD4Y6J7Hu9mlZkTjC3fLom+bz43A3ncSog/cV+pO
P23CTv6ZzgbOLKnaRazXWHE9bJ6etgYhsAroP4S5ywsjyzcp91PYUlx5LQomVnvA
H0wqI7ezqrNwU4eK06TQzgeQiKPuy5DeHZ5MhY5C/knEZIY2+XkZ6QIAgMpD+Qd5
OQO4FvtYi5dVUs/1Qb7Gpv6KuT/+/CDi8bFwQG6FgCxpsVxhhRd/OFcVaIRDh3XE
kE4qs8T94Gair17dycbpWfMyWWfylDF+jKtKnvGEmi7mEwECFK9NcZ6OeuA17C5l
XxIufg44WR3uDGZEUxvwPchidCWBDbp7fz7sJ5fotLUUHwZmxSNRd4bdJzmR/7ry
6mhvtt1FxzrveMaESSho4ce+v1TTJHRU5PwzocZTaQO3R8EdaDeeq2wn5Zr7Tfoh
bEXi7oXHc2N29TawwKb8DQh20d1D3P7zAgdKGYAw8pxKYIqccb04y0YUUyivdDtH
Fiw8bsPNU7OFdkReHKagYl+AUpxO/eaW71aDO3+ILijWIgT49mJf1ZB9o4/cFQQK
NVMQ06THfjXRzJ/1vkM3sNdwvip1EWNsPuAdHSbvCO94vS2yrwV3TXhdkHK6ryOw
+PxUrIK3fmmzl0i4hhwgJCY0kp8bzbvNAz9RXng9AVanci4/7lADUlA1KbZnp6nd
bQsgOacLvdXzVd5NjiUsa/3kTi3c5Kdn5rvbXgUbIlVhukzDBaHo5q5iQmZ3H18B
E7EZl5J/qK3HwTLr7CsJ7Xl2QWCI/0/S2arnX64+QDmHnP10ar/xFixzw/pXRy51
lDwfKtN7RoNICBPQxuaka+1mwW+t8L2EqU0EyRzvn3vKbDBcpMb++7m0N+XD39F2
oClEtmE6Ghu3nTgeNlaMOkxTkEKNcY5e6VBFjhUWAhj6ujxYMX02lzf7sJCHfCD9
znMZPNEY5KdObcNhTRPn/WuefyByIa9Hvt+RpuTBiJQhxXffe+BQ5GQt5p3J13co
Py4u/w7eNLq+pI9fb9BzNhwajC0iIJPLTZ7b54BId2gbeSO62WvpTlj8spJbJyAp
dU1a9vJ2RM/kF9ReJL6ZMeivO1d3Y6N7iqPcyM7hEbKyFlOw2Ot6Bg7tiOqizpyK
KODLX+gOWVwrO/6CsiqE0zcOgJ8zXjixcZG3yKcJ1HbYW2FQmSrHfrbG+6yrPfl6
DFTJZhqridQ1cSG9veSoVASvkCe4oWmTeTO5L7sdEfkRj+46J4PqhwrcWUknSNHp
lcWS81hk3FdBa2kuhp6dhu34BaUcxrP5r/TVxu9cRzFX378dRWQ0dLt1dELK3G18
VPckwQzSIW+ea6Yz+bdXmPUaMV6DGOM0Yes2xf+rVl7j9V3JPMTnjVw00PHcia7Q
L20TwyAsiCJRheG/0uoiliMURk/kqEuBvlVU78+3/aOPHM0X44lN1nj9wtbf6x/X
skBoPNaQy3LqCP39dEx4gBgBqdBwL4M0/0MEOmoA4AjtLZH/dBOPCRHt3W/yFJ4P
f0R7HFDaWgSxwYM3aiacc6zUWlQzgAmGzTCs0Fdqyua3CS4LyMLPf7WUYz+m0OEB
mV7Qdt3u5eNUDbHeMHj3BYNuH6BFyIR74C3ZrZLgF7Uz2EZPqtNg31Hr8ryrxPMe
a8xLjvNRPROKjGM6L4KhgJaRzx01acobIXdyCR681k4fvRLpNr5RPw/elY9N4AoF
jcgckvjOcDMO+kFXFb/mUORuqJpGoC/LEp8Cv+AF4W3uY4wYJNFbONMUDN4RGMOi
iEn4qdtZlCDcDzmR8gKnd6Hvt9M+rPAxNf40c+sbch2absJKZHroMipQKDithr1v
6ORJ7B6B6/9UyM5AFRT4B8Gb0zpfFpEZhkI7fpu6WJQ5nwGq6Fb1BPD6ximgIM4X
6pMfMlLdmgn3yJCZKpAzaufpVvg20VH/q9KRxXdk6SF1Q9XehfmuTxzizXLf+yPp
+/WJTlcYyjma24d0zJk/X5LW8oSRXJVSn49VCEK+Tah6c69spcsNISOdBUUnB3DA
kxSacQ8WMVAqoV34wJbQf+RIM/0v5Vx+hs6Myb6nCijbwAslq8DzePGECUTjoUKx
wDUaGL1NcdjEZ1wwLiDBNnYuc+pASWpZWj/oCdROL5u69R2BOkxuSW/4aj0ABQmZ
NbPK1EKK0ZFOxoGOG26Ei8EG0BpSF+F/DbDLtzh0OglhNXMsbnA1JlwZGtyttwm0
342Y2POAb9f59ooFRahS0C0whrt31IkIESsV1YvxvGOzdAkcwPc5WuDQvIl3Q4B9
+TU3GS62xzCbzwkmSkcWttrmOMfWzoZ67abAJcvJ9EQIhL8Zf5SPUOAkURv/p0NY
3s1WaIzfisosXrcT72mS9iSM2k5mUgKArjJzJ5holgvFlAssOT4bvaUWVyW/Nsji
AQTq0rc8fooxQ66HvJA2ThUMTyI7oj58SesHj53Uemd51UpaeLWsnIxEULGE/TtX
gdBAT42VPBLOte1YfupYhT4g1fbeteOBtJgWmqov5AiJ3d9IeibX88YdveB23bF2
7FRT042BMb6x5rdSmQhcRZz2FcY+AsUQiprNRX4NTTx0Uze2YEt8jeAEbMHiS2lS
FNVG02V6uKzI6S2s+xFEnwq3fiM0NV9CeNGIi+9FEWmv9CGxWtJgctiRrzJoEe3q
UAgqL+NCPvzgwfyV7dsIH7Urs3M0BLBmlxzvhVnaqesGJ9yJYtLNL7PC+uXmmUwR
6O7takCHwcI+NPWLoUlCdk8MPl8JQGvLdXOiwNO67IbTZdlLH7cvxtrIGXax5aBL
kXjSGjt4lOfeLVac+QtqwHE8IRzwdSAtTngOdHLm6Cn2m0c9Yt0+xRSuUHLEBCwT
pp/uA5svS7Ye6s8Aczv14T2SR+qdAoM4vkpVNw4kDEV/v3oJ2pDrXO0e9r1DOFRE
YbvaOGgva8pyonuRf+zYxpM1+JeF2pxk3zpSq+PT4EOwnyD42oMlxdmEXpUf070t
ywdP6ZV8ntBaJCoedWTHdF2i/hhcY5QRtqZQnvHNBnpfpnX+r2RwY6hiAEepl3Zm
L/1i4aYBevYXIJYfYIkNnKiFYISZDauET6La1yIWdwKBjtu6o2uOm9My71x83za6
/Sa+SvOGKGX8mQ+9oocu5pmQARfD6gDn0TSB0IhYAEqnd3N4sgbQkQh/+P3sY/n7
+KZSJ9mbHaYW80pnk2YiWVPH/cPHTo0blHWZJ/0K3lqVsHnyERm7EhCipVY6UKJd
9+NcI9WaH8CwtxwgaCH8a87QoUS1bVadKASm3s+pudQPF26vd/GdBN3v8Z02C1A3
vWVlAL2lB0fdA9olZQSg3yD9EMG6FDnNi7nEQUSH7PDRa659yRCP9LtqwH+KZVP2
jCoFLfWfn1V0eLhcSfhzGDMgfdGTxoBOMHirl9fFRncXvjn60C9zDLpDp3YogE+T
8MgnP5/vwcU1Mo5qXzdEfJZBEB4Pw8h5GTH/7JRDX4j49IhicyyQvOCtfuPhYdyy
QNNnkBliIVKLRNqiQT4XgG/F5/U5yKRI9heX4Zyt4QakMAyzOZrtTveP+MYuqrc6
NS8jdTyn6sHiXgoF/BsincxNa1ItH6T97ur91IEVGe2P5wwimVDKQc6DxLR6XwLG
cdH6LTj2t0eTe01lq+Y5v2tSOgZdjjI0DY9P1pUSkA1hafYSXz4ayFlhrYba36Lj
6IHhHDpg5yQYvln9mZqgk3n02UWEPlbOi5RV7HigzCjI6rbpFT8O54BDuVrMz8fj
nW+CDt8iDUi116WOa1GSLySE5bTZT/Ej3VQ5JhALvxdmaNTN8cpkIXKgSo/hPGv/
a8eAgPtrvbyAbJLbEtYeNyuKd/DyymTn+JY8/btiqUzkiV8HNdHHRbQ3h/afi+aj
1wVAe62X7FAfOs/JxpJGS/80qBR6vW+1dXRLf5nxdwk6/yQevc6XX1ckLPntH5cl
T6m2lRHFZuV7BBFKdiSp3MqZn+PSuLJDLa112N3sorFnxjzU0C4M3Z3K8iPdVBSK
7TM5GneCKnp0gyr2fDlWh27EjZegwkPpKa2omlJCXXSrHWKpZkCO4u5UAbJE5C7O
nu1YnSHh+aP6KoRgWzrCSuXX8qLaHoRf0mMy7K0+kYp1qk6dUCSQsCViWejFDWu1
/TZmOZHyU+fVtegg/whQ+dRGJ7skIwFSpYA8br6opwfwcZap+0Wt8uL18H6R0upb
53eNR4FDYpjsYi60LxcLH6S/HhBPW95qX8IPxUCnqG3uS2VYlkyHZkjEIQh/JdiD
/A7MyBOr3odh2/f794Gkq4R0n2EMGfpWsscEU8EEaEQWLM5WDQjs4Cz7H9sUKpIm
DFgVFQ86P2N5iGJewFbvpvjkf3FdpVxIn5Uw7OzJk/s+yexXZGi+tDfp/VxC6Dnp
x6pEnjX6LyuHRo6+a32gvW5xaPoanzjumjbScc5PMDyhvmamcCLm8m0iuJvSYXGY
PhU0SnXOHAvmgU62/3xxoDw7sAU7xvuWp6sPdz+euEyLwjORIkN2mrxAN45ArWv6
SwToAXPqjf1ri+xqy3dck+grTkyKI0a8YP78S/8zQupMPq0L2H9SsMf6790Gee8B
cCZ7NireFTMDuuIvrmQnvjhrDqx9AG9el9CERIRgneShIlrEWqByqWd1EtL3YE8/
8HhrJyVU0P3DewGBvNN+mc22v4lS0OMdBuAAZngexz9DkQqWc7ns0bWXZJqNknze
7Y3vwZiN8XNE/N8KdE6ED+rk16wGsduEaF1MicoXeblwFFXCJsCqXiXbg73UZtxO
PlcDMeWpMakCXdcMHBHPEKGgYxQVZXLr2x02KAWrFJ2Ck46+cUs7kyapwD8MaRHG
TmD8DnMgM82iwpQTNcpgrSbbPXEGvLhf+Bgi5G/G2UwAvhwfLjMTKiTXlWwO+dZi
IP1leJ77+kQL+IpZ2ISjKxWQvTCb1GJxYrnnjIZARZB4VvcOfeKUCEJZI5e3OCqN
lQgOl/HmjZXrUTEUFupiiV6HoiocPhIGFPdy3oQd6AyVBW6gDpCWHtvKJPlJPRbM
Dp+ZfzvaNA3Ui51ApMpdePUnogQ0ZjvvE10GR9JmraLPZyl9kUV+HBLTD9SGMNu3
x1Dlyck9YWmmZFZ40P3zanTKnMQuK+2BXtUHqhiOlfCGYLO8/cDgpFM1YP0SzgYl
Dath8MpfbdPEOowe+03lr/FLDBagyrEZgX1009W9FB+eWY30dGXpdmAQMOqiR+TT
GlkwW4lImcM5MbQlOBRv7al7Ha/oggvGTjCE6Nip5sbFADdHYD7beAIgSq8FUPDe
cIeqe83N6m+uX7N3DGnAyPUxix0uvtr3R3Ln+qQLUKcXCAHOhJk6ixdR1cj3RydR
M/HqwFnO7W4bOigMs5qrwSimA241XbT8cLEVSElP27qi0ccTTNRc7rhCaUmsRNpg
gFZ04ExEllQnu1Z0nQpcb/ti0rp3wUsamp9VoiDwv+7qwlAdmmu2Bq57zT0a9DZd
hc2ijKZz/0fD76MsiKfTiJeSUcMI7B+DhJWM1eeyPmjwMZFBC1733yuZWt0soWVg
chW4hLdv/GOeT2g2tbaMl/fLhguohSJXSDYbVtDI25CT/3Efe1NIBIwsEvEMQudd
sk3INT3iC/Riv/mDwu3v+I+i7drv/ja4OaukoLwXK3SbgLouARN4dvVbTg98azzA
iklgq1Uz923mNsbIskRNvs8zinUSXytxlGDoyqU8FCd4BNtH+qAHcFXhbuIGssM0
Pui/WIxf5vXD9IU7gZvzxlDD3y3Q1QfgcJhWYSsYkedeBKrf5ayGoX48JKkF8YSX
b2+HJi8tjWXULbnKXYLWtmkcJvUEcekkjk1W1JXcG45SDT1eEmiHlUewIcOMTpiy
ty0S0vN1EG7im/yEPT6kcwq5P7dDmfBI/ZrLLt2yK8UuYNpIk2Mw563fOxqPSwON
6v/iW+9vdaJw/3pO+PHnJFcna5bGwIaB0hcOVNtWuYvvpUrhfRxiwwzvlWiqfZ33
gnssh1thtee0AZV+VG3VGed5nsVqeztcM2zdnC3wX2nf3R99i+ayjmM8DZxu/p3L
ORn5sa9ips2fTDeuBGdkDr+ewirfYqPH/6Tp4gTUC8WJg/Dl0tzH1IZiySuZ613d
KmvB0PwpiI+Q2y8AgwsW4sPQ7Rz9u0fOC3xBQv77sf2FZx3874sYI7EXiBe59GF2
F/7jNrzL1nizgeltspfhTb5a+skB+oW5ANVZI9vimrqY5mKKyZdcUAKptvPk6Xqv
jeTRl7jfVRr4tiwo+k/GWO6hBPiInDrJw/R4TAtZmflLeKFany5i7VdVZGqS4Iyp
kLWCQCrMEek1I8u82Iu59Al5vhs+l9x0sZGVxJV78GaoJC76R5mP7BTVQ5NCT+F5
opv0YZmkisSmL2wGKUbC1NDFuLtOZBC5t0L1J6osZ1rP2XE/BS4XRLX9LEX0KRI6
F9cmAZ5LZhwfahBljRXJLfpsjeKe0FUCwcSts4ZcWLSz00zVoCNZLlklPmd0MiW0
DqxIotJiiYJObgl9GB19hyE040iayH4lI7zmF63Uf2/5rbBWW87CiiwUXXwihhYT
mioKRcz6PFIcGFAc1GqmeNr/6C1hqWjdW7quZAN0Um2PKzeXMc8/k1HZvSXYDVv+
ksrJptgZPNm7kpAXZYHWJAGtTM8zHJaKXSUH+o4W6z1IkCwBn3cpQYT64hN9ip3V
+EGFT9eWa6IKn1L1KLOnqG8lLgNVeu2k0bNNpLKcEGtff9/YDZyA+M7yjnzwbtkF
OIcKzy4ZZWrV3ho17ZGTQv6pg+h8sIq7Y0ci11h2TKV+8uIIXwDXhZd7gApizAXC
lOZNrpl6j8OySO2KSXPbC0n5SQpDvQJLLHD2ul1LT+JLUZLhMCM0BfTC1Sl2A6FG
nPqzrnxTV+iTiMzQnLHP3XQlVpt5EyK1JU/jcVR8oJOUi0HfqNT2t1awn4bzYRlf
TXvotmklJ1xxi5j9LbFQwcMdnEeG9d7joyAapu9YkHXpV59cCQO9XNeMq7n1Dc1c
ZxNyKjlhHJ4iIUwyqLQfPCiCk96VL9MlpxZCxDJcISXUltMG8Xa0hgdNRdc+pKW+
nqcGkLTMbB6iRIpr1kwQ8auJsdyt9afrH+iLfHRkvtTdbabOQ9l0M5bRQz2vKHGM
ciiRLwB1eiRIZVwLnaRiTOjPdPcPrE07i/bth7KJ4HzUmWMuoBqNrQ+K+xh08+Ae
N+tYECHDIlpcGJNDMN5GnlTxKBmfDfVUEJvquws5mCid9pNIq3xPzXZYkc7TYgwL
LRokh4OD5KLAW/sNwyzBa5UzYew0itVvTuMzZDc17C2qWyEHVhO+zxYBVincEZ9h
u7/8d9Z3eo8hU6R6t35nZUDIQ0FDreIGOxKQ1zhi6gb1q7kBeVulRsVQbvKQr3Sd
1wK20osG3GtLOMz7DqJQQqWF/ATymyl+6vHD5VFLTWFed3QxET3CvgAgMeULFxvh
ewSF8L+2ixfKDr4tTa4Qu3THAVeU0aTH+nGWbFcKOVoQ9HMpgtRGTTA0pASfgckw
B7FwZzEBMx46jYxe82qxXZfihauFJ95A7xPkylEfKqzakywOcnfVfPRYG5XLjOhS
DtQx44/VbfaORyfNCmtd4niv2Sl40iPnSDj1i7SA3jITK14MJ74TthHwyvDCwBDg
UU38uoVbQ9J8pDRrGhmoo6H7MsSXXQj0YPTvy2WttSLDPuP/PsE4WqEPwTY8yq9Z
yL44OvIWb45UjZiFKj3IUU74mO1xF1FhHVDOltq5AeE//bSoWsgM7i+8deAJHpIx
6GHZRDt3KinFvwsPG1T6m25JuJMd394vgLV1lyJ0X+g2K9FZtxa+7mVH9kXrdwMA
yeb9HvvXRz0kHIJGBTAmhBRcFcaqCSKVdocTNWTaqqAq6FA7cR7eLcX9T/NTHoAm
jwYuZmvMMkEx5tRStJYXD0mAPx2ZsYk6AMHLAOItCs/ap8Z+9ix8eOM6WkEK2oO5
TLcf6F7v8WZkVRWjfbscE33aHktdm7RkkCDY4zOjkjEhgikAtDfZTbT07SFtzSOs
nzSfLtO7jkfufw3tWmjBuVgQYFYWfBwgkFm8nN+CxwsmZNndAZN1YvSSJXyTk/QD
x2SfBZxXbOGntF1xTSLoV+0tEoNEd8d+xKWcGLv5mBiynFNgH8tSeKUqIYzVYXNl
0cm1Tod6Oy5bLwD395D3C99e/cHoqYK45w4839YJkLD5tWduCuDvyRs53X22JIoS
stT1B6/kS57l1xNcJUb+yxfAxs66y2S1DX7fU/QZi3XsL28+rfnPHpMbaZVwe/JU
OAnqNeuxy4ZFYSVMRLQPsQYwF6/C2Xa5LtyWAIGM3ruHLIiy5hMvA/jSbQ+g9lVt
nSRJdz9q9NOVL0oX9NCqqTfVmlkjH/WtpozSbLEU3PamEgA9XRy9RaUmpZa2rfqD
r+sJOiRxiM4gKIeKoxG4WBNq1120CDjRuY0NMVFbAA1z8zpJc5GkadRg3KXcwC7i
BdMZyL4or7NpZHqNHBhaVenf0jZMg8GQbWhFoKU+7xVaG9571EDk/HoU4ViMZTaL
5WP44f61/7OtduBoZY335MeTAn8YGRU+4b+E7FO0jScGXmxOuRIGU1CzUs5jpLOO
9Iv6vWb1QlF3kC9u7q+yUMu/nNkfptGzb5SiEehsBXXZmIzXCJEBpbujhy+/hRa+
JrjR/rRmOdDMfrT7O2IHM0qyoruKs3rhdBXXY0PwQlddeuNjw5jzrHi8GjgHkbJq
kIOJxzRG0v3812xWTfsdufNqOGmJIR8lAhDvfLT2gUzcAHfGrnLgO/5Fc1WSwnOx
`pragma protect end_protected
