// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:54 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LWo3JQZeymUBy3mK+JVSxWMvrb0V0lPaKKXSZgE7xyZpaa6wqw79Fopre+qBwYrO
0EvbvQ2qOwK0zMeyAsRk+3xdR5ZRsspaL0W+Rz5DzOtlx+N4VrZbmrjYXuA1M1+c
N6NYJzVoMD7KAiYk1fpci+7/5nxXmiE/kC3FfOJNoM8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6096)
e7RGj2edcxF9oNLxayq2w+RzgsS1iBv/nADtoxnBJ0JijHPIdigvhqYQZ/WmujMo
F0nSt6RLXOcABw4rUbDqJKUXTsNhDXhZ89KbWskxWbArtIdbCeGzjJvC6G0ywlul
1p1BEYpncAXxYTsyPX3e4dQa9yJWg7PEo2LLFlqJ12OLAQ9J/ego0vaWTrWEOnsf
wkHgPvp1WiLvLnMJ7+Yt05mTasXEw9Rhyw3OsxoYddyTY53kEzM3s7wu2ct2BufU
/YbXNbsEFBepRTBNScFPpHHsgUS7KVlhnp/PiGphJdjnreOIK0IubJwk1Ev9T8ax
2grhniAl8Ik+RMlSblP0M+tPjftlnEWicp7nPchv8mLsg0MUsM2RfPKEvarnmRWk
+DLos43yYRixaDQkdwyScE9a9bm2waaLo5bODLDq4zE7BIKmkugNvVeG/jVQV8qU
N+ayeHcj3XIsIm8ScK5MKcbFoC8kqbSdXTFFIJ/nnDF8cBGDSKA6IViczdc3eJs0
CmR1dvLLnpxezcWDVm3o3PpT3Ghzv7YDhksXSPk88u1OsifDg4vq2oCT88zQ8iQ3
OSflUHQHqJIfVIr9aTOpuf47+rrVY5n6SxN2/hvZCbLox/73BTfY7ROCRCsCdAi4
dA05Emkb+F0ItFwgvZmc3bRqkLZ8ABRAVhlADIWZkEvTlAVfBh+NMv5kbmQtyw27
eMzz1cA0TKTKDyjPjVv7aQFSJ9REQ2/+TQzhyT5CxJbPyTGFeCZ3j8el2oASlIY0
z85R6NASTu1r/XMDMBHJn7h5e3grj/4l+qhqBWzi8Xe3Jq9D1mV0JIMgHYGzTkFD
DMoyCpqd1Oki+L+afyaHkM/CYwXYWhpiPaCh2ksk1I+rENWZbE0a0YDGdDLJDM1s
S2MrPXOQnMV72KOuXlRzHRdMRatzdM32ELPeyXpFDue3+8PIE3Ut8mdt/bAvVt0D
jZjkJYqCcItbMPUFl022l2bca85ZNd4ptCC/NOYmxuv1jbN0u2ICvljTMsNOpc9B
Qp+W4oIwA3T3Xzf8oa5yuaKGjmjzuoZ0Y/GYjZwhs49dNXChlZ3nFlEp6n35a6jC
lFQPHQZl2dgvmTTAic+6X+O4L/k+EAFoAkbUQdqQ6RsFFtxqRtzW2kuosAjpQXzl
BzhQ9kUlWintmuXayYY8PrI3I/lEvsAMKms+091t+WzfBjvny2tKRBzvTVgNjLc/
0RO+j+Mw1s5YhEQT2YhvBGTmxhbMxMSLD7cLA8xEw1gE7b55dXozvw5vhAUM4lLe
P7+9wufYAeg56Z5skErr2Xka/j5oo1j6hKDy8xHr9jcrKq3quHaeZwop6Pwbs/xC
IZ2KtOipzmN+GItYcesvVjlpbfvfqmYSHlbVBbn788Q3r9a4IMQTarWRjt+7L+f4
wMG1eI610E4cIGmnPw0oqxvhWaPN+1l4XswENhEMbYCE23Jb2QeiCa7LhObGkGMk
bjz3zWbnVq9fOuMNWAM7SggbMkx0j5sT605U5/nJnSr6ryDlo4CZGWDjFtSuZ4V+
KABpCx3zFIf2SSZi2CV+MXDakySBjvOMxSY9ji7fap7BRmFU9RNHp4rp0NDhRqwB
hF3dJQz7TaVaSA3OCeuPbXXmfmnWxyHBWkFyCLePLjErwbiQM9jjFRNK4BLDMWr3
IQX3I0ozNtaWGNDIouM4ObeVxOFcZ3YF8d6CRYB+qaCbenTH4yCQKCPCTlf5od98
22aJFFdLJbR6nyRlamd6QOh7SAjXZ1mAdX4+ZJn92/OGFYR7IcZ5ulf4Myk35BzI
wC6Vn8Y+pp7l93/17o0KowgOqlBwz7LMWePW/x6qvVJwmSApkrVc7iNARiebnTYC
cm6lu/IvX3ViTLRphBqPVYEH953xLSpKl7bABtLGjAWj6+JEv+foG9Oec0QCBWcV
25wved1MDjT1zAkWI0Jo622Z8LjchyDhBD7TIZ79grRmqmaHZFR8shRJtfeK9RmF
ovXvFEI84vepvyAHRiCzvFsqV5qzHYMlIsrwb6BrqEgUzO3fqBPa91Zz6URsPpkQ
VSTvjzI370T7vbR8H5fNOFUWjqStYKkw14LLfIVTuUSugxHpxXvdq0pTpmVK62lS
fURWu+XRQ2fNF/k768uJ6T7s5GEwVeLXIaIeN5n+4AqH+II2y8zhpyJOxkHNBHAB
s205sNU5G+Id2EipUzrX5rP2m3l9gsjYmwSwoazgOA6D+SYyaw2v5SIkY7//hfPx
mgR2tgea+JuWyVFXM2H9AC4lWcqmM28vMusZOFBPc9t/Td/XCyzRKfDVCM034iwl
MgP+u3Bf0JimC6isXOF5oeVNkSldSgfydBYAaj/WClhZv8L8HiUibtL16j3YPNUs
i/o+3okqJbmKVC0skE5M+c3q2N7Jm3sLcINxPZQ3G4uwTi2iyVdwkilsgAi/DEwk
WE52D7Cvo42PSmdmHmDxeCz9QFN3uzHktXE98wJE/ggnOpBnzQcDtQqW0FaC0Xwd
QqBpWfN5cJm33BCidT6SSFeaAJ9iCjkQZcBF4Kw/WQJEUUasTxTa7UvrX0Ya5m9A
vm2z+8Um8cef92wLmFrmovwtRWG8m+7Y2oCRhwSfIrUogpCbQQAh8js6yK/zuzVo
yK5VEGhixnsHpIXneCGRZeEUhg/r3hi7fD2yfXMWwzXqg6WG6jt/iugsKiNxcnQb
v259HS8yefKkFsOIIkSr4nrD2iHrsamuUd1NezCH5R8B8w5qW562adTdZHVUol7j
zepsiuHjiMzU5KPGpVE3KHgajMGV/BUjdp7XV4w0jriomyOGQSu8gYERzDD4jxVY
yCIpW5XWs2S391wr45XSeehL1QvqYjc1NVQn3BU6NL4vrN38mDgcPICYMlYBTlLz
5syl4D1EPO3qlNsErON0rboyKLTcw4fGwJhtlyao4TRk8dcVoEu8CHkrsLX4SQBr
JUdXsipKC1TGnJ32DHHXxvW9zTzaTDS3mFaO5UcveOe5Z4Y7/h6z1z9ZHmx1qa5V
qLvDrKgRK8Qrz0rdLLw8LBCaIY1a8++b3GWloPF2j7KGhWLKyIqiKevMkR7TCYhI
8bTPfb35n6cMzHpSu6U6lJVoSmOkAEbbAJNNdBu2SM0O7/Wr6dzkVbbPf8Eg/t2j
rG3l0OEnqztgWRQy6oQxk74oAzIKcezMprdWQuutkU6DJeUDiAfHs9GMnaV7auLf
rslDSmgdgD38UMq2ZN8X2DGIC+qwIEy0c0/fz0UQIeS4GkO79Uy43bEbI8s4jIKM
CtLiVO1Q/EANX+wetYIVphwzacpc9MvFPPmR+OgcBzh3rnfmQudjx0bn0aCWttvZ
k043avc76m9yl18w8fMpL0QjpDN4a3VpE2b/yPWnVaRd0DL0wiJ2QfDt7YYABFhS
dTqlf1wBu/OeDrpuVCWKGd5lmJ4xGyNFHRx4ycpZa666bvBBSU4LXDaGXllF8n5D
Om8ka0eyeCdabyFDqS/F79LJ8DolPi2w89/gUm4z8eHPnMoJgK0ztsMx8xPnjmF1
mN5gLrH5Ufo9uXK3pcX6SpV2XVr8zUBMQrEoQl3FJztwWc3doNisEcE07hoNa85H
tRE1Pq6wIcmXpS5M9zP1l/XoYb4/eT5vPhcAlKdVJv9j3UfTzXkMzwC9JZE3R60v
PdSau5lTPL1nzcWDMhJ4du97SqrwgI2PXK64QqdRcbHYYqyToBmMf9bMxV1P7vpd
JgjwJ+NoKfogXH7Jvd6Brkb5dKCgLyfIDKyNzIi7FsQA41RTAvseOixHxfekNHAW
eqdDLiA7nr4pg9dbCLrF+ZiUj6FjMmk+VKq70mbgBdRHnhVaBRHlAY+WxTbPVkfE
x2wrFeiSNmvu+QCeUJafM3EJMEj9Y7bKFTmhXqpkdQtJAIWXn7CI1BTidI5Btt0C
xmvNrcdFwZ66ptWvNj2pCdvpGRq7f6sBIDBQ+U9gZz9BgR95ii81NFqx8uONAGm7
EbnOJMBjhTYpOxH26twLtSLMe65ZVVpj8ebXKYACkHftN9tMLiV+JAT1tOuKU6f4
1+1iKlMI75FLungA8JBXP5voNqHQigZlUqJ8BWgX6Qx8m2buOSSYnFDWHHq3n321
hLJHAgNw/Wj+8zyPnmH5bAGorraGLIVCYtU5bWD/qMqZq3CjFG7j7M6j+vTxiqHJ
i4/LZRVRXwldYkI19mRN0NgCPHRtExH73NGT8A+rtPeMEQa+2RDDI0iSZzft5Ed1
b5I2wF2+n3RnjC0/N92WwSDwrM5U0OImP2HHiDRaJ900hJRaz6Y1pkc7n83aMXvp
ClqLR1qb7GJriBVMz3+DHimMXSIJnrRz85djoFLv3N5NjPazqYrPOewcW+yQ2vuA
TZLPGAzX3ENi66GVOjdJzz5IK7oGOPPhIM3TBzgLWdz6aV1kkAEPM1SZCFKkSg/E
yC2WVVfDCImq01NAIdvhkC7FtEuUYbFoSPR5imtzb63FNii2+FIuCY/lAgAB1jKA
acRqNnAkSS9wzPfKWsuq0V8yhtctPcOv09DFMExBmeubYnVeD4CCd4QFq72LIZci
ceVQxpaPiTozhgZgKY0ANFY7GuodBisPrnWgk1iWZN5hxutF9rt3eo9s7jTtaPIK
EqM1RRqhIV0/8vcxqO/rwPY/kVPYMWy/qy+IVSlcG2fyOgLM2zalekpB0jMPotyR
lsdMSuIgW+Q3zpskZTTSp2lyVZpFn9R5X/ht8NzZrKCELmywiXhWIFUOgqf8iCwj
5bHZEXJ4A5L7oQhpQNlRpUeXsnersUEqCs594Ax6JeG8b9nN24HC1Ot6D9BgHg7e
oIkN4e8vkPAhALeBpq4oFyUVFu7IPiSfFkDUYSPmVfaRHB0UUGzxvI4jWesATxBc
iOOkbrjGdommM6hCHeT9iLx2/RAwmY1BtgzH4zbgBrBnteX9GHVRtPpXdf0xY3PS
Y8MBgBvJUfZW2Xq//AcNGW1R4YWfW+srOyoBFy+fphS5T41E2cNYeVLfKrOYEvmQ
GQBJCaKaf/52+hUplxagOMdLh1Ouowg6GgD3+I8oN88boOHEokExZPi4KIeGR5d9
Sb9fZAgir7qlHSFlXBMJuOaY71sEBHplR5aE9V6PJsTlX7nEX17czoPxMUWXhtWn
WhOI+UZvET8pc6WChuXJvtLL0xPl5Hoyrgu5goiBaHeW+bGXAsmObz4KDpLq1OVP
zIelCSDlNOzUV9ciAN8kX8fZCSf6g7cAQ0oVHK3JmbSrFHh8p1yMhmedrUMfEwze
/oHL8/KuOUPW6/axTLbloLaNZnsICfkxjwYXU6OpGjxXt+3A8/+mClA4HUBREICZ
03++TbTtzMEhk9uO6y77ETe2CBlOreNf9WtoJauKUFzXLZaQC/WYhShdxTzwHwKX
o/SA0zEMtaxo/H7i52E0D7WlpIaQ22WHhNP0FlLVXIHC7dVlMDTdZ+fsZ7gJPr54
9Yq6eyRaiprvGXPHrMs8x8glBPvBnZZRutewFRP5XLcr5Mu+l/M9BpS9XECU1Xm3
0OSBlLkhjabM75PqxaddDoXFZsuSHzWFolDyGFCZ7lDHBfUA09o3YgtwbD4MqLno
y5cFopsyo9kgkSISBzWHsXkUeeY/IUe83wdndd+A3pYoZKPuMhoipdDRJ2MxOa1Y
XALcqWE7hcNcpY6oa206BRbMaHxVU4sBJeJqUT8lL1gCh1PZYjbSuL/KtzveLVKR
vwHoQwbK/r35ljDLVef82K/agkrixTji2bYDoLQLdhhkhCGRAKm3EMFjDHsQDnQN
cFGUsCjpW5jyUbBmkKIsUH4/qqYORZE9ep42U+glEzYjyIbAh+9DjWLJDvjoNl2g
wwPjDd/vUEHVkKai5HdC+s5JhgKbvDHyjNUx/3cbOl323TmL7TJHz/YCa6ZYvbjd
wXDcrejtTNfL1oPELEYC6T6jdK93pHNTB4pSfmMeJJ9dCcJIZN2bGS7C9a+akTJc
23eEmrP4323nf2Fdze/dSmXCffLlT767O7uRvKH1v+Xpv+HgYbVQdZfQHvlg6F3G
WReGprELdCBV9H09R3e7CxB2ENpfOjLYNtYCTnpSqz2YOAIWSEACE9UZRign2Y5t
1WGe6XKAqK4mFytygby7QUmc6HpbQCrwIV8K2+WU3SotBrg7evKFbSxHw3zrODDS
3BNzFZy1gqcUZpKf+AiplpgiIsDXa3BAw09iXYj/Jtrl3rxuNosMT4biqnPgbOZB
WQk/cQk0MNn9o3rt2ovOY5SQm0J92AWiWptiCWMwEGdOHTRSE3BVSx803Vi1lN8A
gRSLgvlbJzZ40j6LV9O6KWpSdDaDDCHiTk340lBCJPgiJdlP+ZYXnGvrLxyKSrfc
X1LOhJfuPX+WkeUdJ6hhbBbIsClSok5Q3/TmDZozp3Q85pJrG+8BHk6o0PJoD67P
8By5P0eXtbfD1mWuN1yOGJMCKvPa45u9d5ngnnZm+CpJHXSgyZUdRmFsSAjaJsxH
HPES1R4IPD3Ri4RGQqWArPr04fKUt0Y20f2SVEY2qCiW3/RUzXzp2bfhBbfgMg6i
tGXTvm8YQFFooRLEpRKQELu7S0WUIkShxs/eHmIV4nLOehqcC9OZoaCvwWimZmKE
NZyJJhbShbcbbdFgMOCLBcUaDAnU8GeEyD+7tk5Z7kzjayPtMF1W6EoIUH85a4xR
QWs/hlmgbHyQeKdWr3Yji3ZD1DeUYjb7Y/szSF0w+LqmFolMOHUSS0d8/Go5wVcu
+pMMiw4aQAJ54UcrTZQHOYtUzFyPk8aH7MFJMAYMOllXqPzdvNHvuZ7ZGv3nIegM
RxwCyyaYyThraflMDd7dJBleNJRPEK2ZKlX1ja+8cWcE+tTHI7A8zXS+ybo3ORlq
ygmi/QqwRgLTYmJwt4JbLX54jliC2n+mOGX/eXqyN3G3ESI+OYxVP5siPps10we8
cRkIPhwEv4poInWqBOdF3kLB1ckDSC1Wo2y5nWbWwGo94/+mHARn4Fwniyr/kT0G
ikmEuV8R+wkCuWwZ3/qXePDgiR/q3Xx7KxDEh6bmltAoQvv/tJ7I89aO4RbR4N4y
RCl+T4EupIeW+fBTccazDeiDIC2IkVSEIWk7ESrYWOIwOZpoIYpXWIVBUWyW72ao
scI9My09uxOfj/b8uNUHN5W9kQPtU/zzt7Nylq7B7Vu7P4mx0TiwVGOw9ubChAaB
CU2vkoMQbfTLIj4dqm6JOSiSB0d30PsfTTHE8Gr2Yzq4c0L7MYiyoAjwEjZNHepY
ZidoJ7A3o1/Z41e5+HsjDiiEOxCIla4BE0Qd1XmMlrycRDlfYv+b0cb5SBRajyfV
hRFVJXUrh3gPTljNTU9PPLkLX3PtVyAPacx5cTzRp27kAroOke4WEYyUZqz9H8Kz
Ki+SguAK0ShaYwVeTvMaK/C5gfkWHGfH+MeFgXbB+qlHRhKZiMNsMBbkgIc7zY+5
HWhJGIYwbsM4MePyzZFlJJD8oy7banDadIVzeRCTDO1dcoigFIEOpBEx3EKaOv7h
Xf4Xowj35YeWntejTm/esoRmbA5VVuIF7As1vViHCkMUgp9PiFraez1p0F5EA0SU
kVMR+O5sYu3xTG6/kheQmoHdDup1l6ibnOZpvl7tDptApakrIADlRQYdUnSjS/mr
9J3i9A4iY2Xt9PNgCLU2N6YZv790T2nX6/IbspWCs8QlfqQ+IyaDy66FmbDTLx33
Fp5iU3BmyNIiQny1ZanW7Xjro3dZHq3n/VQvb7jmH/385xx8VOxaDA/N9YOT7FF6
+zICc/oja3jJkZAXud/odgyK5MByTcNwHW8NzWhC4llcMW5SRo7XeOJh6w+BpZ6s
5XPgMuQN8tak6ZDAgK1MWBqQWHcyQZRCHwZSio+kr3PYFxqVeKw1XNHbN6JG+JxK
w0EEfrJN52lV8SCdIv/PmvPipQeA+Ldd2QDhfDd87e7Qqgpai9Hjk7C66A4LgHKz
D9l+fGpzMrqS7+JKjMfeTBfksv4o9BndiBj0dbaR9IGwoXKHPQezwBzqffP1nPa6
G5SX/U36AtTsv75DrjAqvIc8zzwvQ0BreR/HsxhuEwLZuL5NoCxw1TbdKPkiLqZ1
diyxJFKPY8J67BONRf0+LJySK0qNNC/KXgZivsI0Xgcni8c06/9q4AwaSQPpWhkA
`pragma protect end_protected
