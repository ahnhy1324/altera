��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O����w��0�R�;��s`�D�MKk$�6/�"��I^*K�4o�~t{������1����f	l��>����� M/��
'�TO��zŸ����+��B��L �;���r�� Z`f񪘽D�^��bI�'�s��p�'>����M=��@� W��Nf�82$�g��v�K@�&&*T�u�����KHS�m
��0D΅LK�c��9�?���W}�f�7�8���6[3��H�lQ	}� �en�Ѓ7"���
�����0�j=(�>��.ޕ��g��v%����`9mݶu��9�_+�S��I���qA�z�\��YD|4!a�/�hKZ����>_'-(��m�>H)���Y���G��6��g�S�dZ2�>�[{G��Ht_������4�)"
zߔ�C2�u{)�d�r->��{�m��v&���b�&s�Pn ��������EB�11�5x��Iy����ѥ��5�J��}�}G���>��	T,X�vm�6�f��q?�V�YzSս����l����U�&K���h�5����C\��+y��x�I�qQA�O�� ͩi,��=�?�k�O�n���s>�����cۄ�|e��b�.�gts7"]��yh���-v�F0i���Ymf������m�C�8Q���	��G��!$߸9O���[�:��z(f�:���1&�}aMv�-����E�k��x4L�Rx���T#���2��B��ɦԟ���_�D��6�eˇ�����炢��ΎDPn�ܱX`�Z;����׺8�'�H��;�����Yć�w��^Tt�����U�z8�ť��~J�'�t�2Sp�	'��c�ɂ��"%���=O��m��Shնo0ݜ/H9m��Ob��|��~Omϝ���Q�'	���F`�F�eX�雡���\�z��N3��p�;=�����W��E/)ֽ?-���?)�.�~����u�f4V�A]F7�oӆ��2��$YG��&���Wظ�Q�x�	��+�Gk�EN����9��e�5w��=ȅ�����/>Gu�u*��}���#��w�L�2O�n|y������,��ꐎ}�2W�-~P���Ҝ���U����_n��J��J����$H
��TO�Nh��x�#Ą!�Nv\z��>C�d$�(��rp]F���]�k�5����|��7K����/�[�����)�V���M��71'$o�MdJ�1��q�Ivf� ^�Џ�ߤ��:��Ps�K�HSV�����1�o�j���Qx�"��nKDaScc
��[9��龚�I����k�F��<�_���e7A�=�w��Zc
�a[`T��m��ߌ@��>�,Itu8���h�����n-�y���z�	�C3�b�*�kǻ��  rMr��¤���t�5��7g����=7y�R��/����P�K��/�8q]�h,�u|l�U�c�Ē���c	i��O����N��4W|S�.�Y��O�@Y���j�B7%+�dz^��(Z���}�7h�F�DM'��r������ư�r8�e��h��s�K
Ԝ����;��U��HhҺr��IT�Y��l��VIm����8��(��i!p銲͈��ʳ㗨f ��襅W���Y��m`ɵ�g���T%����I9}˨�؈F���o��:aGY��w�(!QJ��S$��Bgˆ���%�H���hhe"�e�ݣ��ߦ9 "˴�N)�[w�ٓl�	y4/0v|}'��s�ѓz�2���'�>x+Ҹ�X��u���%�~��u>&���iO�hB�0��}���R$)n�%���z�%�����'r��и1@���@��
�zBC������X���O�Qʔ�����afު��2(G��X
..�b������<�2���ٚ�߲�QA�����U"i+�4Y�O3�Zn}��F3�8%��'W�h���7�u��^���&�?]�#�0L'Yp��׫|"&4Dj3���F��욆]� t�	���;6�}�3�����RJ�����h�yЍ�8�X��Q� �x�J��t���{0�ɜ���3����χ���Gͣ�H���%�"d�y��*<�AHԴX�_fKy�Q�z��A��dj��~(~�4��'wZ��@�i��$�M�!'��`l*� �sS��tz����e�hS)q�#���֡E��)�� �5���H�5YR��#�O�'P�
�'�C"����?���w˵�j���*t��s�=�?�П0h���;}�਼�����c�t��N6X(xMΦ)�M�޳x��g����4E/����]�
@��UвV}h�%D3-��.�����i MH��HB'W0M��46�����s�I��'���݌�r;5�� ^�m����,��#�[L�4�/�u�~5k"��CC�.�f��Ր[eH���ƨ��K5�O�;�ݠ���B�D�{|��@����Ũ8;��ߵZ�s��M7�/���ˠ	��He,k�U�V�El�ϖw��V�W�;�rH=�������vJ��Iڟ�l��m��5����IX����
xP���)|�<�%�����ײ�xnX���'	�"�:���?CT_Y����ӏ�v�ѽᾊp�XK��wo���t�Q\1�7�|�or@
g!:r�3)g(g��o���z�C�0!��\h\�aԼ��K���H���s���]Ơ� �5�s��]^�^A��^pU�I�{'��:0p�!ԿR΄��9�nB/���3�-F��T9$ӓ�!�P�Z��^�n�y�A�7�����'�n�g��}� ����n��:�9��Ky
%+ظ�Ox4H��V��|D�.���;��:��N��!�F�3���
�����mȕ�����(��"��"�0�Ag� ���KS4�j�4!g��$�����Ƴ2B9�M"X3D]�N�\�U(�-�^f%`��6p8r:dR��;���d ٽ~J��Kn&�4=τ�{%Xr���~�;��N:c9(��QuRb��*E�=��7�G��Rs\{���d2������u.2Y��3ES�wp�+�1�\'jU@Tv>P�tХ�.�5F�eX�Lړ�g��}&����r��3g�X��7���TOmT�T�^�P�_4�|A�Y鋬A/�cdϡ9�X�n��ik��C|����j~%�W�}�x"G�L��伧�](?��"$��x}?�s��>D6�6�!��P���_��K1(3|��$���.#i܃Zq����ѥ4zW��]V�c3t)���d蔳[�����;$��G#�N8��@4 s�P��ܡ������֩v��c�p�z��q�K�E��1�ú#d�}�Pr�s/q�����}��I�Z��D-����4�r�=Oכ ~��Cׁ5���hA�oҬ�7��dr�umһ�Ƿko0{=?gc����?�h�\$��^��R�q=$���iEd2*F���\M�����Yk���o������������sJ-�e@F��}{���'��nJ+Q���l;���&�l[ ��r�Ao>gMw5���{�3��Ayڢ��y�LI��c�S�-��C<DKP�]f!R�9)Vʽ����R��26G�����JK[���`5���aK����SJ �z��hfS��?3�����F {�5���=�7��)g:�9�DgQ�sd5�����S���I<�
7W���O-K�XS�����]��L�R�H��qҟڋ��) �%B-��,5)x�%bG��̽��+P��D����
5�(���w4R�׹���r��d�r�*�y�ߐq�u�3p���bK��`�҈0�p g�������	I�1���Dv$%�˰������EL�;8�ɯo��v8G�	1e
�[ɜmZ�xkN����F�l��?���C,T��*V&�e�=�E������� �cѨ�޸�Ia/�~n��Rl]Ue9��L���{E����h��]�^6	��g̥±(I��1+�j6�7���t��1����/����/Ϯ��6-n�o�DQ��Ɗ��iYYȫ7;�`:�V���M���t�pS��9s���F�p�^f���������ڣ69�۰K��n��|Q z!��zh�[{CfD1b�y�|!�PB�Ƽ�#'������h��)��;���>���X>5��^�ȼ��uP�`����o��6����
)
�Q�Z~���z�^��^Է�U�O�C�`����ݳ*���+��u쥣��W�ɩcV���Yw��$Br�C~
NƖBU��^޻�e�����9�X0_N���������Ű�p��e}Y)�[X���[_J�0bh��6�m_7����f�`n�8��q�]|�j�un���~��A]����uX�oDKnf&y>��ʵ��޲��m�I{���w����PiE�:]A��
�V�s-e�y6�L��Q�N�X)N��ƨL�A�N�xj�[�]7�;G�@�: >w�Y|�v����ԓ�뻣����.�4���������ZF�MM$�\o��Bv!�����fήA�p]��@|�Eܸ�z�fG'G�R�z�����i�T��J]�ϼakܼ�S���2lޫ�SPѺ���/s8��+\�)���	��:�,}^�A���z�/������$��`ënhiO�s\R�0�<��@���o�в��Jأ{��vRq���d�UWU����xt0.x{<$~�jNzJ���6K'�����]�G�h�wHN)_��J�"�+�%��@N$�%�o��䩾CB]إJn.P* 8^�x�t�:"5�'���Bq �8���tL
P���W"�޾�PZ��A���r�
:h"3ťfk��\;���V��פGm&�ݡ�GZ�٪�ټ�t�y!����l���V���c��X��q��/���Njvq��mџ��;�
/����QtƱh/\f;����ٵ���qPo�����B�����`������l6���H���y���8$H�~�ډ�nxpNB��6�5|���1ɠA��.�T/�B%	�w���L�����)1� �Ģȯ�J��+�$�с��}i�Q����5=jp&���u�G�D��ǚ�o� ��M�L_�������
�o
8�1㜰?�ݘ��t�6��`^T��� �7+�ןg�hQ���G?@oD�}SJ�q��I�4�*�=,j��,�輔�����n(u��� �O��;���I�*�CP� 1��'*x�pʱBq�g�1�<,��mFPs���f�����m�	?�[`�y�4�����I�8��r����@Y}�]���w�C��A�sձ''�n�s}�����Uv�-�PEB�e��@�+F�1Q[{X�*��,8���5���E��P�`3�B��$�}'�(\c���lƒ��L�������q��*]R2a�0Ϣl�Md�mF2�$��dTq'�?��Y��F܇Q��|��n#e�����LQ���&뺽�M
��p�<iř�cN���7ܬ6�?$��C�	�X�I�W�xN�Z���">��Z�4!U>Ε��K�9��Q9�
�'�H0AށXl��a&��z?��r��R#b��jڪz|�@�A>��]����5<Z��,���)��� �v�x^�����u���/g��D�� X ��F�  `N3���@ϯ�l���s�^K:d-M ���j��J����qD1{�`�_�
"��8����X��8�c���V�x���T;�CfJ�7Ɉ��LK\�%��`�V��j�0�LJ��ݬp|�w���`)l#�)�B��A|��7T�j����ϳA'0|�n	�j�;����~�Ou܁Pj��(�omh��l"[��w]ZFe閇�}!�Z��(����c��i�/�~������g�@>{M�!s�R���>��M��N��D�BM=Ҁ����g�Mc�w��uؚ570Vb���;w0W$	9�"�/��ND#��C���'\\��?R�IʄA|`�����K���������wp`y�,O'	T�.F4�U:2�*���	s��R3++\ٓ�S�~4'H�Z�	f�ɴP��Q4�B��ǂ�>,���� �\ćCY�������8M^���^C"�g��}U���',�녡}���4����GhK
CB��dM攜^ ��y�#쩼=v+��
�%mr>	�]`�aQR�?V� ]�;�F(S�>�(�zrA4|਋ަ�!
�v�:8�|R��������6�dI���{�ɳ��9�ksN�JBGV��<�g��x���$��5�_��h�R�8r*���hȂ���nJ�/gQ����?��E8%��*�cL@a�}v��E��0?�gʄj�Q�e6�F�lc�l��G���LK*�Mҿ��N_�ߞ*�%V�iR�����ޕ�RK#��~j�_���o�[br��k��jx��:t�Z�2�-�ET���3��)�K�t�e����"!������$W%a|K�{s��im�6�w��Ҍ��/���4���ǽ��~	��ܬ	�q��ؤ͋���0�j��|��:?���-K�V��O�-�i��8es�;-y ��N���+Nё��u�y ���G}�M�W@w#���2R1��p�sZL���nL�Ț�L����k��J��u�f�B�Y�$�i�ne��� �&�sSԏ��v�qj'���/��K�e��v�|f�Py�7���d�|����{D
:J��d=�8l
�"6Q`⃮��'$ye��MC��/,ޣ�3x��SVX�p!Qk��{�v�B��M�>iT�Y��:U2�b���&�~��Ab�;AU�(�͢%�e���H[�ͯZ	�0+�f"�_�ީs`�K�y�65,߆��F�"���9HҚ�����`��
��|wzyj���,$���C���g��d��)i?���4�0e� �����5�=�(�78<@� [َ�_���t�O~�~-�,,I�y�/��h��Щ�J!2�F)Q�k��������a:���K�u�7,��}t�9�0�S8`�nABƆt�
e&Rq���c�i0na~���`<�1�Q#)���˶�7��̅?�y�0��Ͻ����Ȩ��J�Y��C��*��B���uyÞ�9 ��<��LĻp���s�Ƚ����J��