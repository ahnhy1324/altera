// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WLgatME7R9T0ZWTzQHLD1nmmM1m47Qoo7m2IzVETo9qoKp9TxeM7px8jJ2wnSMv4
I8J+WKcUk5C6kwymqCDCU5u/a9v05X9P4BDzd7/QPmXbsQ1tG7NBiS90X4UVBQiN
YmJDFNgJT77d+kEvz3G0GKud7G8rnRWNK44F4oU+mtw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11696)
UUxwPSXLyv0q5D0xhT+nVdSxAWj4iCo2m+WPEof/W0vw/LabrAjTmfZ16RulIBXQ
rzmDnDVEmMcPCk9X7Le7rtKmLXQzc6U8d8Q4pOfKRNWtO9ud8egucbzygz2BIgSv
f0F2z9+LVOlqkVq/2C0QQyL5p4Ynq/bGmr+HUxNIeYcl1XUs2MDtDhCMFODQNGXz
bamzDzEDaUUaJSzB4JPNy6hmUBtAA/AWFd7zGjLtlA2xfdH3OF60bFxzV2eqhtnL
H++Mz+wJP1jrIboLZ7HmxhX3YG870xrOIuWpEEw5cTYmGCWLa6s7+tSYtoRAOdJ+
wLqf1YfY69tEBZLIKxKx5jYpVZdz7qFQ+3+NA8WPQEbeKNdhAajShiRFwLLLUQap
bjrc3FGH84QPAe1EDCDM2vyx5ZhY4EpVK3PqQppgHlwHNp56I7tfGpAoOOuZn3Ic
Rst59ESjHV/GK7VVXwfUMv7ZpOdV4Z5rYG/yqnOcuOykWeUhfNoex1hl3lbcimpf
tDUj9vpne2tNFEhiNNPl638p8dkqMq5CbGyq//2EQsGMwxxiNyzqRj9EcNTskuT2
eQsAVNfN5bp/wUp0RihA82FKd58ekRhLUSXQiafav+UK97pxrWjhLTBhxoAW0T32
vNq/SGTg1xeJKf167GTphFCvRERoaTJ1yupjh/ab/tjEB6h2eETniNuc2lvi5gaf
5iAl4RJCAmGqxPN9+Cga2Xc4ETL4L1kLsb9VY3GRTBXpRMHF6eSDr3YzEak8YGze
BswNRQL0JZwKZ69xzZI++ESt7ydRBa276CtV5UkEMazQMCjd7TI6yyrT7admCNG9
rJpyUqsVZ97fIeZBTXWEHcvN1gE7mTMTKoLzckA6jdMERAfq4VUvjzn+9TZexg/k
+3tByRr/6uvAC8f+It2j8If1sVv4Z2WQJm6Yknd8dhalIs1eLH9v9quOa9awBiAy
kPJhTM6dc51294YaL+QtvrIJfTcWZXLXWP6jNZ+VqNyT8gO1/NjCjOjkO7BxY3KK
hScOTQapH2wq+zdWTuvNlYSXprociRJxeJW4/WGcs+NclfHBywW08bj/tSHAT9h9
IhmQVZjgdijOZ6eGDuVM+30+g82m+t87sUeBmWQ1qHOV2TkoAdJSOiBiUJUrixcw
zADPvSrnxkgVlj1sxDgVsX4vyrTezl3egX+P/brb4362kw2Ux7SLBUwjW7aZ3M6X
Tg7PqfVgwgOKOIzEB2vaTEUDgtvtA7RJDzx4EhKhgnIhR+parTqsZFkOOae7bCt4
SHPTKa+bmp8kdzSuZ3wRzCTkVnvEWJcxXWB1kBwtlirriDGqiCaz7ZNDk4+LORoY
V9Rl9UNfXjChebC+SrptQHY2emGxQiC/0sIW52tmwzRPBIt4zfU5YBeJM/s/FOK8
/ZTPEt1cpPSXFwNn2/SjueN4/1qiiuFqQqF2yPYNAXiUENYAgF8p+ueOlWGVBEVb
UNt50fBk2ig6NWhdfL1iCnfsJtJrRLZk6c2GlQt4IPGMMt8QrRjOQ5v5DUZ8RBKR
4Kh63OCy15EF/7RM0zc3/9QPekReeTSbmpTONVC7E79GH2Aw6PKhCE8hvtmhOj7n
Xvw5H+301pXN8yDiG68srZhb9ulKTNofAUigplA/T2Ct2SgF1NxFiEr90OzT4nAK
XJnw7KCUtTuV0PxpbGOyGmX+sVLYhvd62TMz0SP4oAJhuAUFH1kgTm32Z86Vq7fF
vj5E0grt4sQEPrkQCE53wP9MYvdwekhx6FXKtvTzNA2AQYZ4ARnYmzsEyN3Kegn4
zVEbMVbZ16SP2kS30TltaQNKqkvYSM8f56DE4FoCOa6mpLIUjuV2KaU26qDhDME6
Salv1nlCIPEXBAnE2Rf2ePSN1jy4YGa6rIZil0I74OdhpAJeTtkYZ0AAHyyoxzGu
pjTNQE8NCIhLfbhgCCqJp8OE7TK6yV64n29ySpAi5JM3RAvVcwC5Lmgw8yD1FmG0
PDXF2Wc7OCVKiqz31rFEVxKX0rxdyQqMa0LR1URMzvNHkEnjZO6S31hONImWx+VX
vSQupo8M31HrVqxIJaSUzSyKR9vxN0Y3Bd3q/4KJLVN+aIOG89veVnVii66YxNfg
9Fk06RUOrdLeMUOWbssgYkFp0iaiKzus+2Ajg02oc+4wqJ7jsWi/9asVWvyqdznN
SteJG8uRzn/biCPeMkrFXJuzGJUijB8L9eqlWhGfci5VKBJcSpKtqRx+4L4D8j6N
LxQC8jYEUKeRlYpvDpmm5AQjdzYTNdRMcTCRuTFlVFOXGR4rCb4TGDJ5YgxO4TP8
HIWvEpUtitUSANz8TmuX20qXI+MNf8foXytTdL7DzvttrZ3yI/KqIl3ojoyoRXZe
0O5DOrlm0/iUMOGm2yEUc2DiK79zz3VO5LYV4ZtnHoiFnhKTSwISoGDw4YrfrJKM
iIPTJ7eeSGxt+3hIqLq5MBXlI5g2QwPnbYd6VwbaQa/NNQoPab0AKvBrRI2fy7/c
6abPWY+zrM0imxDmpuHhxI/a/wQ4PxWvbGTiyeih8LVteSVWEmcIKs3qH0y8j497
cvIsJEtcqoXZGviTjHJ94jk7qIm4+i7pUtnRxiCTMtcpD3vWJc12HHFc3I9LdD0o
LfiDFp6sJ2jPSex5qgmV4hAvGCdmmc+cPyCRuZUdz9zWyq50sL3ixDyhXIasKSH0
qeR2FIUNbbxJfWUCFpj/JQ4jDwHFpDp2GARdomxnOtrk30xLGtnorFvjarBhVEpg
e00rdgufgOj1fPIjXspvBwJkOmgmtWIiNSasb5mCKB/8p9O8gwmJB/rP6qbgAo64
SQOOS29Q0gSL7VDcdjZ6QCEIQe77HabOEpzNG4RHOwMTf8mmhL0DAg2kkpv8p/oZ
NQmbx/yueLBd++KI7qgmj7sHKBkBXZNmAu9jneqXau0pM5Udr1cB+27KmbQ6vxxL
X2Wp+pGshOBC4P3zk0YDGkYtuPy/Ok70Zf6Ymqw0E58VCo+dp2jB5o3uKse3qOC/
nEYUQd47XZ6JDvO0b0jD40Fdnk6jtuCrhYfZb/7SoHvSta4Fr2B5n5IDt0JJuC/0
4qF5PNRzly3vKKyYvFqExp1Ujhl8gnXyQoqz4eRmFNc6tBuUWHEt1PJm3clqLtqH
Hbg/ztrDMbt/kEF0KN3aeUdCFJ2RSHScisf0SAOlpElyl2a2N7FSlDSKot0r47y7
LPT39jHEYPY2MU+y5/5Le6jD/UndsHrnvmD0yMxZXczBO0VkJbBPRUG1w1UtRXcS
/3nBFqjIkhHuQ6tpTRHcwshA+fh/ew4yOd/ZRQXanAF6KPMf9oMGeMkFSwygR61M
40hF83e7tQS8URUrf2SNq63OtMlEwZaq1md3dU+GXvmsNUp/xJRwjcQEjqDmVruJ
4fnUWjR1milbFWducD+yLykPm9OVWAkZ7FC2QXVsiYyULbG1tst/VEe006EtsV2d
GtF+zgU7r2ME1gTWqZaCGGCFCIgidQV8XXjJHyr8GUqf53mKNXwF6+ueK631ShnU
+5oER04q/yvbui+JfQ037vftRcn0+Vf90fZZwKyi/LiTbA2Tb3d0adI9SBz5Uu7O
vs6YaRZGxxi/f4r+vKqXjJic65a0FoT7sRsaf+c/dCQ59UB6goy6iu2ixQ6KcVk2
NFg3AlgeQTr+8gUaJwkbaF8y2OWNc3clWLsVe03TLGYQYrth+LMsQyH+TBbiEXcb
H9GZRbpQYfkMyWMfmE03fwmZnTZ1qUf0/5ELt5nAzrY6u9YaHkQq19BUiPqo6vn6
M+koTv2g6NJ5sELpDE1PcqjBlXHnJifFL/ATd6FYD91vxqg1f7/3FttGHgYDaamF
pP2sn+uhaot57pWAnFYmZFhGaiy5e4s7YRAQ/U1VLRqkk6yGbmfL8PXdidFiA+6P
dyBeaxAnDSgoaKbioZVuo2iMYj2cH28tK//aLr6YbPSaTqQ/ATRgPWT52luMNVva
t8yM4y8bElG1u5xdQKqVx+jkp+mFNSsWjrDsqxbntUPo5OoUeIO/QlkjRnynAPrE
jJprcSEa1TdYPkLRBAf1nDU6xCdoBmmLl+7l8loksvEnstFN7z1rsjGpFS3UdBVW
uiO1Hbz1C49a7sXg2kAQ+0prttG9zgn36YPZTy1tlnJtOrThsCXsx9ylYp0nRQzc
/RvvT7KfNLiF+PwpS9MhxpaG/lNTSjGiIG2wjTacJs2OnH0dm4V1mTvm7hBo+RjO
ZOcdBgxuiwK14ja0fPai7okMhY9W40iySSo/eCHsgZL+c8Vatt5lJ6tre7NgaIv+
Iv2FA2rNRkvGe4xET398ohSErAWRi8hzhO0JCefABaOS4BcXFzSIO9FQjqP6/FBo
2GBeu356wzqIaNHtlSWV9TUj3qcggBDUjrZWML1pGe1lHI0FMdEnPZ4zNmBNrY8W
no9+/pk0dbdvKLm9Llj95807Mx81j1jUQq4yyCipEe63CsO6RSo8Dkgd12+vgjPz
84XWYpJurXIs/eXogNL2707wLunLvMgmsiqH6XNhhUwFyh6wwmuWwbZ3q/TFQyc/
pkT/XpYwjbwtK1nNntXijyy6zxqR7DI2yEtwMQyW1yW8DYj1U+Dw268rnMPdTcZ8
SpU20yTTwtwvYXtsCH2zPpHqX2BMqTIk4anAGo1HV152ZBI63jsHamBVqH/V8ZDd
1AHsd3hCTlsJQ0ryX8Fr7Q6AN8fDZB4G1Mgv7h64QKHXCgQMFGY+0Qp6MCHvq1IX
3bWTws9JLkBoz752TdV0e3MqLCw0E6XR3EjHeKzl+dwBdXKPgaF/zTEvw/hHhDU/
MY+fHh97XWVqkJSxpW/eiWR34NwXKEPw9nnizyjp0DeVlO3tnmU6OyPRRR6WDoKR
XWtZfOBYybUiYwAXzujbhZnc4SF+8GP+fyaDDLTWIZ5G3rHXCETFndjCkeVAGqNb
ESEEJ3cbfi8m4LerIFkf9K0M80xmZRZK1FGPHmXWy1wwuK4KbNbMMnZWSiTx06wM
TSOsJVDf5Ae6p/M9t5UI0D5eKBv0rWkifXI7GF7SrN6DA+EMOdZc25CIzDXOyK21
wQe7+rWB6pzV0Cdfz+i4ml33ZqJ6OyHMuJ8f4VTaCE3cOe1hT4M050t57qlLF2dO
zzWniZorKqXWjVnFQabSXwGjNXwSRYKhqXDnEDqjc281N0vnsGLLyFsL0kh4pty7
EKHxC3P6GEL9QKLFaBIQNSNegNOmeuFDYeuAX9zxjOPHjRO7Jbfmw3cFldqzaZfy
QRMsMwaBozD4ND3TT5UhMUb9rsTIjmoHyZclpx4dtm9zVkSrmVumpttLrRANEWmQ
gRxprz9A0OLAjSB+Fu16CDNkZIObbeLG163bNlA+NPK8JxJDOyUlQsFpGH89KLy4
3k8yML9o08TC9UTu5cafrjBg5YUNywwP+0D9nCgmNMZGXzkOF8oTRWjgIrFlOQIJ
BtCcVOeZdz+Nf7sZLI++gk2okNut3RchkTikOOaC23McByaTtKiAwia0unqOjil9
Y8p3ASnewOTns2dmkt/ARKwnvUrIRxKS66aRYHyXd/YftfXYNx1DW933HZUPoNLh
dKSHFdBANbMg3LO/qxra2IhQ6xEYoqU5EQLhqmfoxuNDuD0YckENPnMcqSds9SD+
oW1EK0ZqMmDBO75+1HGO1E752Iww1V/iljqUCFKsPsm96e5ABFA34eqTKZlQqEDs
PNVk8c9tuLcfHuwpV3bfGWwQli1356WSY2mWvvVdJ8V6nXzKd3g20dT8gbdQmYh6
Z6ARO/mQyzRoXZNTnNLsOwy5Qm0WRYNzdJkqUeKfRpzJkNvyaNnAKG0N7tle6BUP
C57P8895waDMpU2PXFSG54zq0/aNc6iGFEW+MXc56UnKw/A3Ixs2rwqonxsoLuC0
4pcgLnGdYr7JZui4vyWs56xOk6BUlqezT94XMHOUTLc0yCoYqL7CX6+bnbBagb9+
weNVbVhA76CD8hDcNxQIuhsOmJwcp3X4H/SvOn1hklhLMMJodEIxxhS45UOISbEO
uCKbynFvR0Zy2Ew456GmE3TiX4tPA5nBmTqPv3EVf1vnHgmqQmU2ukASvlfuaKGn
quwdiXc6X9e7PkN/TMRhyKiTtsgV7JWfOu7PVgA5lYSBYkDxZ1UkS3qhZCWafUyb
AXcQPtyPZb8iMOh3Wy7CNJ/KUovAPb1/Ii6FMA+THRH/775SpMtIOxUdVrRlqumA
2fAc/txZjdNQ6IeM+KZGpvskMChAFKGSd1BOwXVLnwBI9hcwxZXSvSq6YQvXXbCu
FzA9SAedCezVdX3nO8XWj6CClqCngF5t6wXWlKzo9aDquqbzqLaKmnwoRvi0e8Go
ve0gquJx+vJALC0BeBhojM80ZcFyA/fjOWKjq9RmgGVVxvqpE+GFBRaPb0gBYkDG
2UwO4f1Ku3TiwAq1+MbOhxwFGP7wF2eJ9jLFZ8a8jGZbrAWFxpZIsTVvGm0Nw5Qf
0QW6gRYGQs7NLGa2aS0YEk0xq1eAh7BRK90XEsgIBj7DSx8EGdu0QbL+1hqezr6g
EaD4JuXV5//1oRPkuYc/BxpX10ZjvOhwxc/yVuXEt7UVEHbXqKpjxz+gKJ3ONGST
UqO5DUqNguSccShzhG7rfalg1ieO5uVPykHThIlWEYu89nT5gLZN09EA9oXlUO7T
6R2t2xS5qdxVHmDPS5xVzMsK2Lp8rZkE+LpTQco/m3i+ZKSUYhGHoo2HPxvUYuoF
Ae5OBjERb6zRS9nEqfjEYsjerlJdQOc4ESiJraWCLMWnpX/9c2zzAPOvYYMFDaZa
3H2VemRjy9kzkyEZCcQ2ccqp8w/+NYIDxig10vZnmLmg9oFNwq+VQZWl9sy1cF46
clWt8mAV7XbTs97X9IK+LnSCh6AktHHghAKPOx1CvxwEY9s1viwmjwc2INzefjqf
Wabok+Tnn5+f9WDj5hW4T25Q90mM8Y87ejtuRASSoo7wq3fIynu1SThZ3zU7B9T6
igSepoRp0RhAtTWqMNmiDgbkJdgKaBo1DJcnicxjOumWdm+29sYI7gw/0NHu3/DT
XR2QqDjkR3nlJKg0EbNGo2csXlvZuOd7THTc3j5jmDOTYhJk/L5L1Siy90bJRt5f
J2V9vxc4ZLJ9jgRIp/epgoWkB/iuSlH2FtRkNOjpYsqTZhFBGyyF6v7GMZTQtCgo
KFMO8wo/Qcv5qcZ4q9b1SvMSSrRJatYpZQJeX8wEjMKZmbygk7lQfuKJcx6bv035
OtNEbClr/efH9Nx1lT0+4tVBy3ur/uMbmP8obj+Kr9WaVCoUopLjIMny1GV3PTbE
fpKWXhXt9y6H7MiqmdYGfKDiXxXSNIheMWXZRVhJSEDn67226jwLni7KMAgag7dx
mcwX66pmoTAxxq4dImPVYByuel4SGzjXQcl/1NLBs2cBcTkJHAX5nz2MpJ1iIVYY
ew4UDZIqOQOEhKikTcmdvpnNBgsratJwDCNkl0czBSxcPf5WH6A9cR0lCUaqBNoB
kW9tDCGO48hHifcVo8AracMuR6b8w1o/TvkR8eyc01TozLwWVt7StGfki7F5toTD
Fj6moEfCJrBmi3jJkea6eTDbclWqgMcM8L4ZkD+SDT2s5pY7s776NueAeqg+OrNx
UCUygQv60htEPeAIkb/UsO7/QfsNICTqZi5D+ae9e0N+s1x6U5efzWekdlkPhz5x
t1h6eS5BdyRyAOQUHNc4MwiCS8y1PYYl/B9n4AbKBd1V/gHdlXOpoqWMZskTl85H
ic6FEChForliiYq5rOjZZWH6Fe577m+B8t2cSRDUbe69Tz04vHxpcQPNglDPzaJ3
NhB2PCE1SOhvBdNglG6Wf1tJg++2NYO9Xe4TOw/X86cmsRXOdDJ2tPwIWjtIgjPL
qKBzNcdkvcsFG1UO9rOo5x1oftrVQJw1Rqi8wFd31wn4Toi3WD9DGvILaOum5hyL
umJc6KfwRcS3KIGYI1sf2ZZuKduyUxjDqVe1NXHjTBJP3WWfdgPbp5JAYMxucGA5
LWc2B6P/Qva0MMoNzHA2ytZo9b5ijlEsTii2ZtjfHCkuarSlm6q6Vn1Xsj+UcNCg
lIPfgt7NVLXbluEbHoG+1+dLR9gPqKIwQQwGYsJ/l/Mw/otHwFh43j9D/7/6RZXK
WBzpronc4jgNS7St/7xiue6RPDh3ges3YJMf5d2RDTrIWsInQDKol1BiCR+dOQ3D
ac8zO6bNksvUNbuaHlRO4UxwlqIYmtmNvPZ/ITwuaeg7F1p26yHVNhP190JSwrTS
oRB/oXLx9ol8cAvaWIQvYrKQ19JOpWCpW1lv8VYueQNauX+n4eBNpG3j/ZKdU1C6
c5gM1lPUAb+r6Vi1SioBytgoCmOCLsA7EkCuUZRiTKqnN4sw6objegHm0MmhLNcc
L8umwG1zXMNpKavD5WGYiYqLAEWmGupm4jxs4y5ATuSa5H0xKrc7RplWCq8ae5GQ
iY8ll/4O+OjrtuTRrL3ZGXLYZdNjOnnleL6d94AMSD+g8IRPQbRRVY60Tj3J8aqw
f3hwEICbexkY5AISJkS7ZKUGncq8t7KEdJGrK0AtQ8RVxw1nsbxHV9i1J01mtmo1
iMk3cjbbIWhu8FKgEVKGFT9AVyf61MWG/Cub2u7fyTxfvCGQ/GYnQxD5l8di2I+/
5XPZ5byYnIkhJvq4wSuSiiB57WwMZB7EzqPexAyemaLk9XMeFsH5GY9ci2KgFMBj
yw7tW7BL62MN6CN1AlvE6QagkjjJEy5OQMeB4SvrGIQ2N7w1fIxZNOxyJ/9FjWmx
i0P9w2ncktaxajGhGlqwNnz1V73XYX0hQD6p4TLsbwsRCqxl0+u3zKJdiS9fG3WK
R582Z2ukhe6sg28tce90dUp5ouN+DOSVPLw+66ejwA9bLPkCLXDKs29cCnnWLntR
LM67LJsZfbCL2yvP771atd0dZ35J276rkmwXkTabWbn5K8zaIAHrQwyFcgfyhq+8
Gcv1aGJWCz6wTjGBT1SnbR+/th4IWTv3UHPn6Z0t3qvFWQ+eaIpZAwtrMGcwGO7j
6l+8ZUGxRamLj1COWE4bR4El9RQeIvT+owBZNcyVFpY4il7xqm8wuAGgSrhqABL0
kU/rn/qsCcmF1T885pk4oblhVDgVOrfvjBxn8Mwy6OXlKGFmcKViBK2NZ8ZyYdLp
R3RErxXEJi4DqX23SQReIMR4N8b65TxYQcgN+O4Erb30IK2T9p+AIjo9Y8ot/qMQ
oJ6GiKxMa4yC8nyXQ45wrCvjpfipzbjbMKcDQ7BB9SxwYISHMC2omM7arfJONHMZ
dGfpQZbtWeR4F55loY9g34VH3XlVJixsqAwuphnczVgdjp/sgbWpDLYfNONgPdG5
mKM2vsByZRYpnDJbd5Mglz1RA8BwRo2kxccSK8goSK5Kpm7cphMuMsuVIrBf7tKA
a0IMDX4pIZa7EOow8nreOgvyZd8hqKOWm+kc11jKOIvAcjQRtgHNfGDHGKf5X+dg
gZCl2qJKFLPQFpPQlTA7jImk8CtrCPfDXQLJyysUqAywTwQME00+dUoUL1BM7HnR
SJbRDa9rx4+yE98Le1Izxctd+8uzPmQWq1s1RYVIjUmJH0XNnnUSKyefB4ewNg/Q
+BsuLxuJxHTe+f6MhkbMFXCrkEbRlhCqxYja9GYaLwa4BWKmRmgh9kA+cCsB/7yE
fGDCz8AEkFVnxfJaaBhjMh6jxGhuttpK+3G9QtQg54cci5LrtqBwd/lae0N+0h4i
EgctMrpFJ+S+4XqnV6ImjNkYf8h/exhNqpPShXaMdLVNXwtcLQt4FFYp3PsHKUe/
Wpdz+0hsC7iqqwyFJc5qxX5+W7lDaIMBcOPVSUU+/76gZ8PP/DH+NU9xHcUf/0G4
3Uq/pbZOSb7XBKiSNuR5M/cV8xyKWpq6PGHaOb5j2aG2okqkV/eie8Y439mTpLxh
5pG6bdGXKC1ShofflXFRvaNLy8Yvp69FbMoie7LJ2VIjkr/8k/W/g/aNDDMBbxh1
mL5jwQUuzkT0A9sH1DxuVczFEuEmTU7SLBIeXdzcbtq/P+J4rHPwVeDw6LLvyE98
1kbL/08uKU0LFA7Y7FWy0ptsdNs/V/lSFw7KRiAJ0IxT3heZUFpyuu97FcB8zxV8
biI05+OZ7QRKfcFII7OisVHcpRcHDN2aEG+0x4cr6IKXjDBLBzdttk6MvvgMUfId
+R+EDJId6h8WBCITd/vxd8IdycUMgc99V2FUWHlrl0ninFfu+P2LO8o/lkrxEsWl
MGU7wVM+QrFiqfaGB/ydb7ozwY7iZ/34Kpa7yu3VmNkrSAc/Tw+H20kAVJCuuDLz
+hf8+XAa4/F5kajQ8JROYB0jcxq3w8HwJTUA3CgLfGyo0/iOu2UM18bOA8DRtmMs
/LXipASPqg1nNKnIg2osArybgb8pX34SLtpxShyp7Foq8z6BiWJWvYGvSqBDfkJo
5UPcpk9mc43TpgTKzLk4di/9dn/k1K2WBIX3xUbVEM2eWzqS1nMSEz+rdyB4Hht6
GcdIq75HtkTPZ/hhE653tsY70f2+1MZ9ypDzJcJGWwZqVokvDxGQLF/1B2Fbvgze
kC5W7gk6pj2rTUbZ4pyD0V/lnSAaKRWhT9V9Eah4B9o71tl9mmjatf8ASBl4Id8i
c1s9z7LmOaOJzodeUfpYUHzssq9sfR/TxG4jF8WkTgSnJ59j2LWmsYTOajqWCSv0
4S7VcVvz23orcaM6/KTIElu0YBW8GzqXKQ4atVrDCQgk7ZJmUVogKFWXNPW4SWtG
h4tnxRSIldJWptOpEVeKGKXc8HBnOlgMRXqsrjw75yq1wO6eJPu7F97sIdbFx0NL
QSppExkwu6nPu1AsBB30IPL9987OTNzUEAyHmdJetLXEldvMLo9XcE0F431W8nE6
2DAcZThJCBQmYGtb1n6Kuex6y/N/wpYetFUO8fogD8CLHWOJA7/ZNBAAbbpYl2BL
BDmRP/UsYS8edfHSs2OgZXAQwl//jF0dgiRmDl6MlEQk8uigXvRy14YpL9/TFmj7
1NXqhvoZeHexhlRJkCeDgIGJhQB0LabMV42h2SPxDvg7RFfJSCIMTXq0rCYVWfF6
XjM1traRYxAXuI65C4KT3GQpfEdJRQ2IJTGI8/jb/gxMD1cwxjE+ARrMKuWbD8tA
PX0h/40K1HAiIXln7ykG4y+g2Ep1FWrt4ieFr/2vneAP1q6q5DjVrcbjM3+rDtkr
H/aPmRHtg0XHnc7/I7kZ1W7sxnu18wGlRiDZpFJyIcK23c7NJcJhcef5x2HAXo4G
jTv1o+MgCDANUW3wuoSZia4gwmTL1rFdTmVEhCkrQDn7rkCbGHDRNTy7ocxvsVns
ei1jSK0pgi9naB3rhlXcr39jpQ2elcnl1/2ZLy9STKJb8+yR4g/yUXBtxdIT4cbq
1ut3H4ClPxByJxpV8oIjqnKPxBu7BCNv0bCYlrOc39/WA9RJhHQizuxJNqqccN7p
OjCDxhE1X+bBABqDuecSDRjDj578a7Cb909RklCRLgggukg+77BLHahKNJ9TdvzV
M7Zi7fwm+PHRGupxvwQfSB7ehmTzLPREbYJzszr9CzQ9cU7+T1b+xVoRBzRhF52z
9oRAKoC2+2FzhBa2mwG7uZG9mt/cGRvm/MJPY2GO03yxy1qX6ysM8lh0Ngu14CTm
C0JExnWWuIBsK11tWLJn5Z3mC+W/4kqyEFFoy0wU3yH7nSdWtAO71kfUqTa+ss9F
4GN9L9S6vAaVLKRSZ0iTyQPL2aBOepo2QPvW2fkSHuxqzxBmsn/gR7FqhMwKwIad
Wi8OVTh+XDz8l28rSBpyeZUu2qKR53N7GuqL4YmllXtFGBgg2Q/771UzHne1RZE+
Y2Rdu6Ekdqif+Xnjdb0etTL8BYpK38AXXnbUma0XZHh62R+MNTQtcrYqyeD/KNhm
XL45+WcFNNqv5Wy13tqpb58DrU6i0pbDhvaP5R6O9X446VUhUhvxxYMnoZ8sS379
8nb+Zc2UOTy/AD8UL389+Vq/gDcQQQ9pq7qwp5kM2TSu6D+MN82MEQC8dVYvZMeb
aHmRR6eygGVDGMqmU0qybgqvIj3RduRs8S92nqsh7bAekbyDb8LdrlmcEnpv1rAU
QYOwCmlPEzD9gN0m6YratcS8A/j0mgXUG9aK7SV6YymU1ln2NXF8z5Fy8g4pBnA1
Y5dI9By2x2NuJVu2m6gCnE6JIJonY1c6IZbgml4XAdtzG2Zzs+XiVqmWBChCBSxW
F12xIzm5yHIcsUZob3X9lqdsRNCxqbyV/g7oFJFwPWVsmTxahNE3yegnli8g3T3V
M2+4z9fCcj4CB/gfp5ht1yrydrGUOnsqBuvudPD7GJeCLlBSGDf5Qeks94MD9V+6
2T2J6lDQJVSogE5ar3MuhLEZTT0dASGURgRLU0s6IFE113cgWRrqIPa3y8Art8L6
OvkOPwYdHsXydlLUPtQedhAD3tttdlwdykbrIfeSR6paSm97fPexU25vmV//Gtwd
2n0Bg5bE0jHQgD7p4iYTAp5UVfcCNzwrbIhqpbOhXmdWwj5+MPziXApMexhU73G5
6kGSnI57pdtgkaNvjKutVNjvXC5BCzdU1Cp6cPCqtcZotkLzoxuyuPxT29AYwoUH
FwxTYUbgEvN29k1Wrwi7DkOrX3eWN/tviA2Of3ZlSDbQ6aIafJrNdlbVu3aXOjHl
HIgotUn3+Ea4o3xRlSfjadnb+5tMv8+BZ2X3TfYF9P7KFDtIIWqISY6S87mWyQK4
DRnUREAcnOvavoMsoxmN0Z00iW/uQll/Rf0wKeFOerV2lQlnOd3USXw8GEl3Cy9/
hVob9dyfO9vPSvhgGdglMNmGGaYI07BrqJLRy3fCW2c9Vah6RouOAPwetkTP5dd9
/Ri9us1gpuUtuW3acqZuLsuBxxbINW2x7yuWFh6uM8UZX+RXWz88TaaeumsfMjlv
o5A6PniAlBIVIRBGrZ4jTHUcE8uH8L/PMZYgS0Mk3PUOAGVr560SgWuSCgz3Bc+6
g6VvVIY+7lDqmW+zIHabR+T9vqW0sSUx/ymvtynbHoG6v4Z3R1Cmpt5RMWYrk9cE
dRnlgqL9OCeooxaKHIcSVh0UHar3pUUWbeq2gc7qtq9S19Hm/PDzK/mzrkPYsK2/
h9aLX5ft1teDbDkeYSqwcsZWiQUBuEyz9/kbHxJAk33BSSviNFNG+9e+RZ14T/HI
4Mf4lPEkngxvqGLKgoLDyoVXd1zxH55sU4yhIV5gwQUGfCJjzCf8m7Rv76S4QU0L
RzEjXzFBBvX7ZXpaAsV8U1aqVwY1uxfst6O0F+ZkjTpfAhH+Pg9mWX+Ep2l2LGmS
z8OrH8tUTxAoNQ3pBUjkttC+Z4qAVch3st2TfEM7jg39RL6Psz8xwGuywbNnXXPu
+nfI3v7EGTrxwm37iSESepE2nemyYpDiDLYkMqvAIVWGJRw4yWYzzz0VNh+RUAxq
2p/ZsGAmT6Yg974NdIH/hIhylcCrkwvwx4LLo/GJ/bQVEveyEM6FFxPBO94bmHxe
dRwzzpsWXFNtNCMKOGI7nYzHeT1570+TfUYqJdKaGqtrfftPFI04p3JLSv0DeJwA
Htd+cMsqY55woBogk3wBJD3Y7PBJh5swqxaj2vsVxVa/i8j8o+/b9dsenkiCLsMo
wCfEgCJ1U6aJ3C3Z+EIEGy1b0VPDCTrgarC8IcoiyiHPUnSNmpQZgFPFyBsKuA/U
K0Hl/y7Cj+lkApG+G5j69JN6vRClYu8ELcs7EgDJGqqDij20RjRkhQkPujHRAQtq
JUCloC6KcmcFBIOdDetxMGAzysswgd8+dZLkIwK9LfOCulaOeIGTGatUIzJGPIiJ
aDJaiBaHpxRA4q2iRiLg0tX7Jcc/HDE93hdJDr/zb2SI8PngBYMOeEvV3H0nyVmp
3uZIPliCdH13dAc/lnCvy1kXHnxNbs2CC0xGZBn5CIx3m6U9pFNXULaCAXLaNfbN
OD4yWFuQb+bSF4rRgTKkqkSEFJkKS+1fBTynybCmT2YCNz24JJdxGTOBcBf/lA+C
X06gCMHdrkz96R3d7hyHyUfSFOEzUtYoYGl1Wlgy3ko7AZUT6O5+VIhzt2WrHRJ+
+azVBYV2kOUgvJnYXVdXSjVab34EpKuALN+yEWvV80DqaDhX6tLEoSwy5ukgYaTr
eJrbZtIYaYY7K6JKDa7B/xKdSTA59bhDTSuGDvpvLcI5RUKRNsZJvXXPiNlOO2GI
iRYlJGhD+hQQMPQ6tNrktxDO8sjlTf2vNbKD6Po/fMEGoeTI5RW0REhUauk2Ntap
CPir+ZB+TmyKdGKU1CSijGD+bycNNZGnxIK1yLyBwNft8CCdgVUxDQ1+RIArpAtD
B8hXk7lz0XH8IIA73H22NAp5J1RdXkesT+8y0BZZtXqDxtJ6cg5UzEoqWPG9Fw6S
Ogubgl8/XkahYNx5VbbkW/NbNyNHpYlZL29gj+W13JaAQDdhTcmyYJIaVCTcPSj8
CMSC9VzL3PQyJo7gg8nRi49QZsPDoH/C0QZx5Omrc2J0SPEsuFO3s4NM3YsjTybV
FKpniXGhYZj8tubQTiSqXeuNnbgkO03vex44cLAVAahNkUOyEGUalaK/9QHQwk+J
uCyYFdk+McjmisUNPFG7WIiQiJa+5CE4aJlsq/kpyLmWa/KgLduMHMNuC+4gom6w
2ut0eXcRfzcOlMb2iUDQNJlacmEecTcf02cyvGnigsuLajQhFi4PrKVEY3qjWC5w
SCt4JrNAw5FwFmqrVEUzvKaMuqvqdV+9iY6q/G/syxloG/wLKot2iTNd9B2rGqTS
JEiXhrazR3LjyxFa36DvofMFCLyG0NUGhP7UnijamXNJYju/oN+f1QmlSCBiaQWX
Vpr1Ez60DKkaebvkPeIzWl0xtEMscvtGiMo6jrv2LoXpcxXhvQyLWR/FW9XNkCDs
GloErlDcyq0uFkEJ1OBG3VJxm2Zoqr/CWTCzSnMf+dJ3XBO8bjOJXKR2Gmv27JyA
874s41k2SaKdnBDeC5nKpR5Hmsxzv/1ccXN5JwMFToSBZJZMLpTw8jUet1zgBP20
URyv5VRNJ09M5QnXC6PICclJ8kyIs23xKPGHbPU7z9ltNXws1FhDesc4P2GG9vd1
OyjQkrOJH5tZ6s2PNQPEnxJNWacsatGDnrBfa85OUp+6CSbq0tUCecwvJrcjdXMV
FsoqNLPhvj1qnrtkhXeByKiFkeRfReqShklqbwi8ljYenkOMW7BHAB+l52eDonJH
y0SSH/vBivzN8jdJGMtukQtZinnCEDdqx2Eu96eXHEbxfYvdKNoQ8Yv01msXegW1
vvN3oIcnEpB0dUXVKidjqzF5hpy0OjL2ke3E7VTN+w0sBnk5EoJIZp6VgOQUL+RE
2FX+n4aaFovNF7RTSE2WluoqcRfBA0JaIi0HBN+GxpnOeaiZHa7J6WLq09DnbMCW
ggOML1jbhqQdF/Y/VcgLwKDHZYIDIHF4NQGlcZSIpfcIbAClSOUSNUIiugX7oGap
vni98ZoJ4gzP65h3GGtJkzMu/HRI/BjL/8mfwR+NpaDH1+vdtjxqdWpwOtaFBrvt
EFQOVARY1liucYCgj3tALe1Ujocz4P4fLN7XjroscFo=
`pragma protect end_protected
