// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MdM1JN3bOfZgMreNN82mJmaFE9sUOpRjEBdwoMeKQgD30SpZNsKtS6JeMw5lPtYq
TDFZs1y/1g92pwmNnLYH8bVR5ITKUWkN/Aa8PwXeiEu3m0KwNyM5qSxdN9nggMnl
273W5Zu4m5yiZFI1Aao/GfuXjxMWV6oiVu5eAGBVbQ4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25216)
joffFm5MHhKWgoAAUTT9lKZ8IwS2CP2wZ7GWJdJGTAi+Pyr/gP4Fu4i5506w5gnR
Th6FFSRxYE3xt7Q/KNeT8pKYqHk4uE13AHYyJcFSVQHV6G7dRjJeYbQlhCwKBH+6
ZT+buY9KtCY08UyxcOrT1qbY0xx0kkeaP0htT7VQ4aJy22ToKCSZSdepO+pJD2Nu
wfjIRut2+Tgzg+aUSPQTXZss6UPepIIg9QmrmgZ+GQbwCzAfW3Sd5qIVT+G0bn0p
29yzGjqKi1jHZLcPzo26OJTIdQmpWWi8w2TMZyb2Lz//h8DgN068u4HZYiHqNmcv
1NsN8B4RoZJMN2eGZWE9yE22Qc/nPuNpNYe96nqCnghFZK7ArC/UeHwFINdfgvDZ
Jv3LuTIFVg+Y9XpFw8lNiFdGyA2Ti6shKR/hK7DQCx508PJgwhAvwrzACq18twzE
542lDmfyevguH/m6XSQO2WrlTgOMaf+rRaonTVVuRWE3GXW5aaK9+Yn+XDVFsNnX
JwCYf0XmoCdAWDDBig/YCbd7HhFuQgxbnkAx8swOUDsi/ZllDETbbx77NcYzmXHk
7YHqpf+zFF0jMbBbxJlvAAeBTswDhTHsmbOLuDVTOy1o1fAhWBgBhf81/cJZ4Y6v
eQhqwjk50UqlmMhVj86TIzljJZnGCHtUiRRgRK5MhWLUHDQgYvD9kPsfG+qrnI+u
aM2fFWZYkGOuyhsPE/subFUb1H9N4IMcwA1DubQ6v8DnBtmA6ib0jZl9U91j12Ia
7q2Z/25LEAG0+DS0lg3PtU5HX24jSp/os4KL0BX0xCDa4gT1ZbhQCbeO4z5H6QFb
q4VmYl235G7vjKmhV9ZM+mCagrOeRTBS/HHqJR/72YDofVCBPqScKRaiDFVc25Ru
gJ4RAUYGTq4guBYFy8Li4jze5NdQRWkf2Otz1GsV+bL7EzFASvzV+L+oA/l1E39b
kqZFHJAQiA/t1Hgb2i5WPpi2VB1md7sQ+aQHtYPHDS8cLjfQEkXX6NDOiSPvjhxL
3gr69iYVUb0CvgPEN2UWII56y+xk1oQGz0gF8yfidfQcO8NU6MvZJ/hHluJsXN0d
sEiO4d8CrJR7A3of1uqgxZA5f1+rQKUv4pj3bE44XNNAoLbja7ruwvBESEHMcIkj
LJmvsz4tnUWoQDScN3hjgjPs9YN2Y+UfyAONiUispmCjXlUdqfSBYGRCP56A1CvF
mDtD/HCT96zuj71c9bAjLX/IU+WL5srLl7fCnllynjp03G/uixG3f3vDsgDEqobY
Eb0ninNhIzxGL1auQY67jIPeOxDgMIIz92E0Lj0y5QvhwEU8Ow2YB/JVkiLGVLa6
RzUMY/WHOIeQPdXUBqo55PcgeVhA6MVHNV8/zsp0xQ57kNU1ZQtQNW7YtJtkIFZZ
PtNBWuThb6umzPcrqz+w2b/MTaro992qeWm/tmTJh8rj+lVAZNchJKeBCpYzglOK
vWF7koUPdgTGAFPHhuO6kV9AMVnveUCePBuwkoCgp3cKwNTdip9+QLzZNNqzh2eh
zYSwkMbHLICg7bsRRLVcQ0OtFoPMJVo9cezSJXFAh/QNS86HAuSSJbPLrbJFVxnR
JoUbU9zNCdMTaUnHifj1B5Voxu3+xwhiF0Ml48BcHKxop419isiRv51R8jFlDf79
hMwyRFuzG9ikw+QhcpPEPy8hsgvdWJTGzPYUZByxj+gOWOzWFlDDzzfAiqmAZaoG
v93b+3NFoLCr2GbXc2PNj9uyq+ISX07fkT6H51tQBJVg7IBhWu6SPGerEY+30Ugd
wqI4JATXE8XmrzebvYvNSvjnFbGDRNMR/C2M8P2LVBbeOt708XG8iRAYyspXaz6q
vbHkMz8SnXRvs6oV+k2diOS7OZJBXNWk9mtXh5jm6Zm8/t3AN7ZZS33I3sUQvlKD
mh6xF7r3aBCfMYC8zJ4+DssQYsqKEUZHe1DkHtNuH0bD8LuBRm8ZD2NXIfcIp5T4
RoECiYsH7iPnQClTd8tzD0b4RUGFimJw1H6ZQFBtWX/vQADzAQN+YstwOzMuEhYV
e3XtnabIZl1Lp2jU7AwehTXcxeStj7DbGHwy3AvfHoYLJjoWuPRvzmOVlUBA7ZGA
7/r060lEGc7DkmrX40mKdiHSypddOuGXGpYYeV4DeXMQT0Q6mwktS9G540vsfO+H
8JqRdWlK0eptDKxspr44OZcOxm8x0LI9TTz9vitM3kLy+uzKVzrJKOIhajDqnFWA
GWSOwxQ63RIT992G9l+5661PqwIDpGkfr8kPs+Kre/302nkynzIux5iuEuImKhP6
CMyavIKvUk9RrXFqVrBV/dO6fJujMK2DYJfHRdBADMGMTAHaWv51cvl6B2pi+4Kh
FpO/9TTTzaUAbOEoV0VkhRe5p/+MhGHP+HNX02OiedkIv58/IbUZGbzhuIuhKUFQ
RX4uoRYaCniNT5b99eUnIfSwaCZWHuZ6WfLoyKk8LLkXfp4YjYU6+4ZavnaisQS0
XcGRyCs2dpFXRsEErv0qVE3//UCOPvVQ5Ub0H9t91d6VfAvx0Sll3FDA1l7ZemBY
aL0TelTT6RIx3wMA8djKUb/lgvIl0G3zDPTWfjX4sAmrS+k1g+g4x5bkWt/p86S6
QjM3rqK2oFlYYuXW4qrkqVOrbC0sEg5J/CzlNK8wzaBbmn54zfSCDz1edLY4YREd
zRSCknzEVdLCP7FRMS4U61CveMKA4Dw4CoD1dlAnaqQz8/uBU76Lrpk9YB3RQbFg
Bc+cNSYD0Tr9Dc+Up3XabXhKm7VhtA+ie4BUYRDt+cfbrhNUGMTyGDMvbHvgOjDq
6WkyV6dfOMZ+oeKBr0LXYFMLMf5GVCVTpwsUuZgMqFdfoaGcIW9unE+cC+gzO8re
jiMjxUmaVhCoq18yM1xkFiXd3H42pleV8FZDzOIOAZ5QBiGt3fcpEtPJL/yHcCMi
/MuFutAH6z51CAgp3uh0xb66n+LnfjPlYvgCA2mrN0joD2BlUGUoBiEcLFwFainD
MZqbKeGCLa0Yc79LT7ndob3WhxReJNbckkP2XEyH3dVFL0xH4CQIk9hGRwwCvT1b
YvxaJgvKw5H4oWWQNyQviXqQz+9yr1mxC37RjP6oYXQ8L7sZpHVqA547Gelv8dWZ
YEkGDDSwciy2ERjBShbT+FUEqwqyseLvOY0AZaCcFk+h/0Ma+KDW5FU7prM8stiy
8mCHBgTr2cLxq+xnvMWWoBhFa5+pFUBiDQTL5cjx0S/SEHtcjUcrilmqHK8hsSU8
RSTxnJTS+/UkHCyo296H+HNF+5TENc19mrBpAjpA64Cq6bNaM/jv8Ff+XulVKxzL
cv0Gl4kI0A5WUHS/zuBlrFWu4f2sdvIXSSjbG3mXim137b9HZsBkUOQtyHF5jJ81
Q3Ygs4oz63KSEir6Sf+mJWxCiK+k6h69iYhsjxaJcGjkZ04JesCQL0MVeYI4W00C
soT54T39uVD8JntVEcisFUB+00F1DdXkXG9zIwxavfu6gO56C6t558TAqjColQRT
NdFSsrUe9ov47DY/XDUjhiXzi90U4mjPwdkFf+73dsak7gIvo5vLl2MinYsxMI6T
v8rNdcJQnzCb/8UAtH0JC3SbJ6bN2RY9T4DLxdTHC00hk6IGvaooRVy3Ot9hxaoj
eCSfacTL7isFiXUOQLzc9FIDCN6PzpLNvAwvZuzoW80utDD8/55KZrvJzVHXJBUA
FyGYCQCFbh1EpXH6hsr62fnEjh7wqAyeyAZ2pdzBX2CUrJERW1+zbr4+J7pO5lBG
iUXg2GioCFObf8VYLufJcqRPZ60xFkn/wEfFX3MbcW5yWndgo4tDo1xWF5hnznRU
BCZH4s+FIpnguROf6oan3u1jBEONOmzywu4Cv+5ew8i/EQwwHKkelceo3hzE3W9e
WUIpiN0DGFkKQVZRLV+zc0TX3GB4h+vpTCaRokIdq51YHI35Qla8qtpv3TtRUWJO
uRVcylNdVn5cwZoBb6DCzbL58oWXE0Fm0H5VYo/CGvo01DgLd5vWgzTlKoGGuiKt
8y1gerTZ/DqEiOjzP0nkrVJyJ/TCygECn+mfMd2BravYxC/4xmpUZtUK4ZLBX0xF
lZLNzPBVwJ8zTfCsShkIUOR8yyoAZwVRstrMpCp8AHB7UnLYjKlnhYP72pCt8Ji2
u3ZQ6bSHKxv8n2AXi9aM2DXq5JeecsjGnpGjk2MU8nUlhVjrw+sa6WbW/UEjKGi0
ZUHZgU71Q+hydDgR1LUV1Kx8MXa+pb0E8pk5rHQiJ1ImN2T3HuOf6kjqPcyAV4QX
EWZozKltXwxSLivtOyFXUQNmoXj9M+6KGLwNY7RdzolfCFFFVt1bVuLlJVBiYmgT
NMxRC5vqF1fQLz+jx3bsFE9wuGpunO6N+TBWSwpCVp4Req5Gz5BNpjYnXr+P+OYL
g/gCrw9TNfmeBdc8Ybqc9wJjo1r0LZktwjT3lhA2NJfGhMaIGAHpNFde9t3qDBTH
oSAUqVtBp4wJAHWJavlVQFWRsUvIFtYFoO0TAtd0zFJo5t9/AH2ZCGD3TpptUKJW
G2Hcx+HcW2t2ZGiIbxGzCJYp4s7ekl1gldpSsM8cvfWU+EG5ZeU5rxppVCk9cpiR
w8nj62ndNoqI57iwBHFi80/0iVSSwKQ1Vb303u9Z93sKmehZpMBZMKybQs3Cvl52
FYkPOizs5oGDVVBG5kljlVW5UaR8JzFvWgyffXK8BSM8eJprMakHeHtHRr3UEJAb
f/buaLRMYJkZIcIasyJKXaDBZCfjvQknx1BPi9FHe5+4g6O1LPIjNx7CRtXuOvHm
pnEJJtnMeKg++MxpavJBxBkuShwQz1vtvM8sLvN/jb46q37+PrA9D5YUh9Ot72Rf
+J0fR5kaFGcxIyKQtSczxytpqaLLUBT4toTmjcwxZiBYXOFpYUXrY51A+LoE1H7z
fdx0gCiFB5U7Q/0HEXPP/A4ZVrV2FRywJtD27c4Y0df8FwA1MXkpLP7KsP3XL5Px
zkAJct10qWI9uKWB5k2MfXCDyT3WjVt+1aRbfGiYfv66X5j9fxmWkzq+wWroe83r
17GDY3hut7a6zFO+32dDGpJO/ORFONcKdCvCCzLfJkS3j0TTmkV2xodlXXOdZBLx
knHtLqK5DM1wCZ45d5SeMQ+ywwWEoPv4mS7d+eptdfeMIQLRbjU6zQdiFDGU+AMK
4s6GsrHKBrUFDfH9HEd1wdxbgZX2UJCw00fvNYWTr7esHRCF70zktkOTtR72BOz/
g2lNE4BbH82tpkbPE3DkWbxLA7+ZTd8G0pWgfL+eRkjBzzuCNY0bZQ8uKYrG2UW0
aGuTgxG1sOT3Xl/TFZmdzjyswhmNHgiRLYtKEGgPzjhhwvw0ZfdsHE/T+GrlAk1P
+nilvWbvvnrs2O0dtTxbRmvC8KIqBNbVXJAFyDG/51fbnuDqkKOH4wEZvIwED1IK
l1tM8fsCzNMvAi1lU8FVci604xR+xVbHphtwXQOy/CdLLX0BbuoESbo2dk8yOL9z
P+N7YqLWmJJxPUlW4dhx8UI/c9erQstMlLK7npvCOS/7QHINsXZOAwE2YgQC65rR
IAiY59HYvBAw+2Wcwzu1+sTyCTUBWOCnCpNZbGT8Lr45kf4ZRYdlGbthwY3vngYl
vSvUWe/DbZ7npgPjVtkncNwxKAynRQ1ReB+6WE2k2kN6umzo/XN9pBeIeZbe5J7J
7I2Pr0dQKTab+30us1i4zhkfFr2K1chiIt42mKnSGoscevpaKAYq3XIbb1gyFa70
ynRfnOpjrO20Af9xrQs2RVpg05pygDDOKOtgof0vhDx83vUCrHKSIxIXXpDC2pEi
Y0LPQFKsqC6qs0j/0hSf7u15RsrN/ORj/FMhmB87JM1C8Tny+//vxzC8Ww6ef+uP
EbkeWKaiBqcFhkt1gFYnmw/VyNv50qJTyIGr6SAt2OQ161Xsr9lAZEiZ/PFz4UKI
hoCV5Iq5zb4xQj7K1SVFw8WflGXG9nXE+Etv9PsgJazOxV2gE8b1u+rWA241E5Yv
zKZnSEt4upZ45YkTW9sQkB5YTVse1yYiuYiHcYPUEOr2EvwSb79I4zdnHbsIkvNJ
L3uXniDiWAU48Q6B4Fle2fxXaQgU0oRuzKYXWLGJFdlbH5FB7cSEX6NHmGRHyBZP
yzVxzeSP19EehBFKFC+Tgf0h7EPfTOe7t2e85QoBrNTTol7zUXwt75W2njzd8EIN
2ez5tIUzxf+m/lpM9pw0XXJ3dLStIFJSTSKPZSf3GNbIGMKLcnzIgRQ8RsxHFkXJ
rBIOmzwgVjPmKrRmfyQaJzAyKrrbwTEI/QIB/OHlUQRStUlXR3xWAzdpMjWI/zwl
3TZi9+rXi8pwGSnu1AWbw+FCz0Jw0XJ9TYsL3N8SgSqjGAPSYM+8CtzhVTCusP1V
CELijYkFOEAs2iIYivn/mvw97mil/UPvLAsttyb+cmtVbKI8Yae+MrETcBWgls7p
34Tz2uXW2obqzcW2mXkC1KH6z/Ef7KnEzihvvtfMorTncjZrpNfOYLf4ev2UZVDL
ADdFrO6bGQK2X1gucus5XwG1XThlaFJvD6v5Dm1o0G1MZYC9eJKCNexXsM0Z2qwi
rWOTtBMfPvAsorAgTtpmL67POfIV3H49bM7qw87N4OMT60btTLqpn2jprAQG3sBe
3S6Gtmms+3HnYsenI07VE5TWdqA22ZCT1aMpBF0RXxyF1eFmU6mxmL22ReYK9GRw
CJtNzLQLg/K0qddeq/fD6o0Zm+OBP03xFSFLuy1uliFUJpzwxa3hlIpbElS5E8T2
ThdVR4WAEaZ5oyEXDhpGHyB4zMqajG4W86krEAGRFaHzt97D6Mt6Ja8b1VhNum6o
ojKO74PAGmkg9f5pRVRtEpVcXzTaNWijSexjtpWacbln4d2thikaPTdhdEMtGiyc
EFwIMLapMd6yQvJQizqvDs1KPvyOjoJySy3yTykDpAs9i+VjlIqr7nYBnR/1+aYd
yiGO8cLKwRLyjQIB3BrLbc+dbs1wgxmKHZ0huGOjbtwhqgMvOPaGIc+GergZtakS
x/iKV9k0YVzSxh80lb6DRBqB8pfUcSTY2Wetsz4WFocDrhWFSMLrxVraDuHwY1BV
lquWTxTxUuiT6pD+gNHcWSAqLxsJqNHPpaEellzhHdfl08A00ONojJUP8IXC5Vdb
mP0EleByQXrQUvi0bV0vjUXK0wBpwQB5Fq41/T6HbyoxHJ1Ev4ubzHE8UpeHBVuj
EKywugomaW1TNye0BIn5IolRPiLkBwAJnNFbXavY6WsZvDZ46TZqdAe6SeqeWwJC
msWzzW2u1FfVX4D63v9r0SrpbVllnyZv5p8i9Amr40i8yQpfi5R0pfKOwpcWCBX1
tu5YRjWl6qGlD/b3BeD8QNt76RA0TyBKLEQ2QRxPeOBeg/3JErAydgVBiHIO2MLb
d6p1cHahaTgw/CB/7xJHrnTDs62/MhdaXZ4DEO5YW6rfypJDoNv7he2LLRrueIx6
o4vbsJnc38Ndjw1czEPArIMl9eyEWCEp6htPr4xclGitD+q5teYOklzJqndkrTei
VElJXx05IM8gHmEkzrhs2rO3+VJiBB+HNRLFwlVD9SeyPaJqqHXeAoPCma/AInB9
tCR3scoAsF1GdDSqQ503dWR/NpLH54CMeJJDgsje3LbFCCd1tlQS0MTdS+Du9SgJ
lwHM5An6Yb9IgKFn6gi/AMjNLKxPliMNAx9pw+4773lk4V1fmLe3zHcoHSGS/NrG
u03fjCaaXGFSq9fUw6RZSMe9s4nrztAO521z6P5oUMEunx3jJWK+O3E6lWPXTcR2
tjO7Oa1anrqxjyI8VrYlv5AdczW+gVfKd6ObW0IPRWgS1Wehg1gWAjncuHQcShvL
i3Zo8Mvxg+gFkDvO6eEPVAYqrtI1wRNAgjv62Ok5hwb/3vKO5BW2jBag7Qv4HyCT
q2JtDK8a4BnSzS9GZq4i/s5BHBW0BeQGKcbDrjX3fwKknP37/pXInARqW04tfeHN
zfMlDC0XND240HC+9xO21S5KONCThzqueUTC1xZLsJjEavyzU/53pCvZGxVEXGFz
0noOqU+B8pk/BGPU9p6xKQHr8THBqgWafmTv1oPLdcNdu28eSAcDFWAETJkmh2Am
u+MhdOi3NuMzFfEKn6F1eidWoczsrtAncGfxEVrgQAAaz4dcOVDnQ/LmgUnEbJUb
BJdFhfR54lP4iym0lOxAwsnr2UM1c8L3fPnD3+H3tKKBDRdOYXPtT0LjsdLH9Gcz
eebKMxwceazvk4WLt/vkXIIxGmgFurxJoaOtB6El0KrqcGABrlTssZb6a98/qf2j
J3HuYQ5TfiUBCKvE8zyAQJjNPbaJAuieXugEXCohKN+lHjL+muLwPXM+COsFoVSi
b1xsCq8rRpu7KmdP2Ol5h6LQUOqySYwSb5PF1JfkcxNDQQErUGeqCx163BN9lifx
AMWtjJbKSMVVSghKn2Wiv3+LzpW4zoaAo6csg/Vj1IiLlP2CwsUmueUlmaSXDkIv
Wh2zXF/0Bd/xouAan6piXjb+wiulzf++BchV4lx2CcCfYOYxR42YnsihzEJ4xjJr
X+HAK4WE66qynfUeprQHcCMauGPlWZpfg1TOIxLNz6zF4PlVr6J/MZcbm+gYHK62
qYbA/r4uR7YAyUJAXRSTScs+KJjah6bUYmYD12ygkZn6ldmSgYQKtWPj5lKWWQ+V
FLa8Yh7wnp38hf+A40C33zX4UHBzbLdXbSTkB4ni4jdMiFIiCBX9V1ZI19FRWned
LQcUVClJpoIj524oZ53d9pYG1YdFSkAPvg5dSNiCglu8XQs97NRCxqhB66qNFkwz
cMYWtuJuFwdpl9euHKQXlryTYAl3HjZjTlvKLwPasbQN76828g/V58z1Ng5s5Qis
WIiVKmOkG+//ze9yNDUFlr0dQmi7MvWT/Nzk3lslHoYz+WcDlAGznGecyKj7j/Ht
kzwQVTrKsPIw71eXZbyp3ZlT6Vi4DQsRY+eylxGIpk1uAeEZLEd6raMXQsbLZod6
MXvo/4P1NZR6YL0V9kp0GE00US8HBp/Jri7ThZcEQSf2NvYIa0FlGkLt64VlTJ8R
db1MA7HrUQDCzN/kvVJlp//FGUqc0jozFb062DhHhblNyYWACIUeJb/0f9j1tPh2
Gruj4cKPq1AcPAAQmBZ//+1FZHrMc8Nk2iErMOC61ZzUvNno+dCQ+SLmtKdQ1Hz5
woBd3pRJfXv0GkRrbpxXkRCdtDpkjSynOkeIZy6Pjda8nIuWe/H4GzG1ryX1oIRD
3vt+UqN/tYVEboCuExOMqfuCjH+UCdb6NMTtVo+ceuQZEP4bcCMoHslUEaWp4X9V
5nLGZUEgXvTLTbIlME55xC6G4kYFAvaxD6w0dPMkKttiZPuotcs8KZW0ypmbpK7r
YzMa7323eZ91ZzX5KXnqi+JFzA2BIZRyzF5v2shOlnS2YMZbNtC22Nid+tdUacmE
YMi1ckMv7Ak4Zx2dXoQjVwJl0A8aLe1hfmSSFEdyhVSLQNv11O66mHKFffInjA+W
eING4n2swtrEO8G0sLq7/iEeFrX3YcEKALzxLw5ZL7AynCN1nEPFzep6V0mkLG/I
babgICr5UN/M7r84OsYh0ZtW4CObiha4uLR8BdNCMxu1wYkLnIMPschash0CYc+h
jY5dh4t4jef0dXZkDcS0g4KR8ERMZnOqSG1uB5kOJhv2EVaHgjZcbE6UV0X2sEoL
p2My1vtT3INlI9xaMCZH2AgJK6z6XscGsWzwrFs3JTwJJEQjx0KNDJFmb+g2BS8H
D87mExMHIoWqvhJNGty7r99+faEs6usTjluMCQF/DL6h0vMiGgB8Ea7oZ6QT6/Jp
u/2UY3+HFSxdHzE1G7seuv4B0cx9AkRHiSIfiyCJElDqTrLQfB0pPNIr3MOsmOzk
nlNRW5WQxLUxb5LoSQQCLozvivLk6uGZLdpXqF3/SM9icqDNWl3fLQEl65v3H0fn
ou47MRcJ0Up/GdO9ml++P97+y8GDuwTmJEJSkWv+fGH6cC5G9MWQPbsK5PmmcdjP
alQ8m4Z4epNxx5uuCzjFb+8ULit/LMCFpcaAnkHVPhxH95zYURNdd+5SVfD+bZhF
QI1anPSXXHWFs+DDEE9mdMnPD4IwC+JRkbJxIRRVY6Hj1QVb2QE7q9xcEmwhmUxF
RNOvTyFLfQofdZF5TMWhJlnwZtrEzKALKuJuw0og/j73TOWPyHIHiDHZ2aBxjE99
enEwrwMdG0iijIULYGV134+ywot7LsrOnIHzTQDZdK1e3ieZ/2qJRZ7uPOJnNZnM
+Kc69WgJ32UDZqlYaRnWT3mpZJXjlsJFjMpKfV2T4vV5vSle0YC5/hp0A/P4D253
14bpr7loIVznk4FW3i4sR1/Ar1hMMtq75hLP+wu0v46oc7iqeCaHnUf1hglUKgC3
xRM18aZnKqkvGxIwnYq0tyxQnsoQ4bJawQLenVXVl0A93weIrLvsFaly2aKRcogM
cykM+cf6XVY4nNPyCQiCAi+Qd4C4bBoqEfHoouQsp2MAtw/3eHMNPuGL5Uj8E5yb
tHwHYQZQ1u67kHXpdk76wbWl3T3TaxZJoZZdrpG99kw+LQrn+o2E4Hpmcqfeg2dT
K4ObfyEKaGE7WTy+VkdOtz+xJwnHtzlyl9D/oBb6N8NojNz35/NeCoIJYIKKq1kg
iAAxh2GBUgue7/H/f21Nxm4GGxVV7IgpF1AqZIRKV1+n8jGBG63F3P2aVd68rxBW
vA3A00/DeW2VL58jBjUS69YbjEss1AnzyF0SQmzzx9PihzFpz+pfdLWegr2y0e1k
xIQb+wp3uzSFIOGLIiDbZWNzgk/655e7wYpxj26e04yCAVBohnEs3Qi/RwKqAmxe
8oF3m6DPw1jJMMdQmaYezsTeVhrGPDEYpQtWKfTvPPlFS9qXVLMY4UoB7gdUklpH
usNRmYDSgWPmh0ycs3SGctq3dVwDlsQWl/BhBrsmlmfXDa6jXHyPEeDZ00OuPj1S
aN4bsZbCAUwf/Ia/gAYSQj3qzBPL41bdExWPAjsJWcHPY+U15AOwekMSYVeSm9Jr
V7jiNiV+wsdHXlXCYUAYsxjs2JOErTykRKcpAE/xauSxca/ESNdsoojgnQg1lFvO
VmqkQjB8D4soEeZVQ79LTrghUWjjjEDLt5EN/rP6/whnHAUbpLkX27Uq1YzNl7f/
aUNjtaSHThCcC3HDSVLJnUC3ox8apr2/4O6kkPLbNHQAqFnQ9zL9WgMyV4/rNvqV
IXPa/ksUREDB+O8FJzc1HG6HgRrNky9+dEEkIEsXQTzzRyo8ghGjaEMkwZ4p0zNr
ZMPwKl2RAju+QdzWvI4JC8Ry5UJm5KQImglAdOSIm26lOutkyPKw8TT0ElhvcUgN
XR+xg7Ojl+Wi95lRH3QJGNtbA7NkhU6UAJybEEki+bFn6QFxkmrhAmhPgVeVpyjI
dSfeLc/v3VqL+LjDS0385phFj+Ly2u3z/sqWOfXLN7N1p7v8WP7JHay5nsUXsvIP
Z1hgIv8aDVL7icRvZGm3hRmAAyeTy9UtsF/3SM/q9PbbNCXmE7zv/VliJFD9NShL
SWSoVnxjnLcHw2Va15Anb7FHIDyQadxfd4zKxNisZeJih3e/jO7UrECK452LjSew
A+UdN5jQ6eC1UAUsBZvKK0tdOSzxu0sxB7mIpHxsN/Yla6F0VAoqPi1xZduEKTIl
veQVZHEWyQMkl7qL2ViEYn1ipOkmvDA/lu64iWy6BrKwfQOy5Afk6ObAdO3zibg3
4cOG/n3z1/hndlj5O1OXCZX2cfAp/BOApYs3kfzqoKmoNfM7iQmlCU6dvvJME8Hq
SbuCEtX77FayraCN9TEKKegv37SkfYDFi+R5Lb4Da93VkJLYs9m/O/y09ZGU3AzQ
vC/H6MKCce37Fg1WgkGMzt3mq1MXMNyiOTiT0pZFa/yJ9lZPSIOUuTpFVzOJpfOM
69qapXl1JGr5R01218YSNEpXtrGMzWFUBuLxIVO+EYzFnJXEZREZPMRCv7M2wR9G
ItUipTci85ulvVoRnylPFssNW0SwVNnhL6nel3JM/tV5QnWndsNbAHBV+cI67P3I
AUNYYOs6TOms4t1cAUoMsUjo4Ks/+iipLertLbip+NyxKySVTwVLGKl7zWYfhBz0
jkIm2DftTkIpcjD3HXeCjgWmBGwuL7/Z63N6m2SiFajzHde8W8Kfg2ELS562v4hA
+pGZeCUk1FTUfup8iaFAmOJKdn2JhS05kdBOF7aBBCYVxxofTv6m5KJ5rzVDbvdZ
K0EpHuaXfyWneJbUPUHA+0+ENpGL5D9b0mmYxXEl/lwLBiNPo5GideW85Ez3zOPP
G/yQ9/LjRGfegqokVQ5SRw1f1t6JlWtAtXe7Hepog7JHVLM65G1FC3j43GUTm0vI
19lNr9gX3M5DbKOe+UG1v90goMN5TPgeOu67cSdyQCoXhxQFm3J0F3ygRLkts+Z5
NTIh2rxXBddisWIpiyfZG35t3pe07iL8qBlui2sIHPeXclFNIxcWnWeehqpKvWRh
W31t1+Ew3reDEx2zwxUo8KRzG18MNbUL3LFacm0WdlXyUadrILn4xY1EDr92VUAV
8EnJvXG2J+PLN+jx8BtiQvAusxFyv8HRXlQ7t/qF40ctjIk1UhSBu6gV4koL7QPk
r1kHWMPMLaoeNE70XriTCGbpjrmKBv+x5UmhFopAFyBZVmnx7bp85iTJh0EcRlwT
6eeKohPWatDegmwZ2cInuEXu+3/YeMrp47n+SHcHlKC3OiDKZWmr67AB5I61Lj4G
zJ4yUJDpkIH3OSDrpewGnnzcevfCFkYZArNzbxucaFw4zdR5gFm8Se9uSxUlKd5z
MdQoDFN+bu062mu/pACUbVapZn+yifFjSHmlYd0NzvefHEWv8FQrWW3g9Yl0lfkD
L+qJaSLAMX9peqMT9acbNzOUiXU16SODvqL6B42rodzJ4czdwVWYwthK/sQMRTcA
YdI8GxhCWaHaa8pZ7P2Etec7SfEHvthAMLZHuoAi2GwFb3aMI90myp5B2jiEesKo
TKPnLs2iksK+vVmNrYhTtpyh7BiNeADMnJaqrOgJUUf0UCXfZ+torI/KesiOpLhi
Z1XgAkrB14ZY5CJTGGGeBIq6Ea65t9u2vuHnTd6Tu3on7C73cUDWwKCtVZBVAny3
ij4h+gZnPAG310u72WrO/PEpcS6aFNMILx62cOO6H+JIKdhawPb8eA5gThdQtwzp
INvjQzaGQw8VXl6BUMPNBJN1LhtZ2ayoQGysbSlZVw/ULDgLgdEI0mFn0TU1gsUD
SWxUf9xdJcLIDvxC7SMWuL3wVVQZe02dSbK1xpGbklKyK4JGQvGJSOSgU8l7yPRP
KrpH5azUNA9PrhZZYTCZUDsmlF5bYc6Mit2KlrPPI9mXLEGJ50PC7MIgD53FCOlv
J553yp+l4WjFgziavot9VwzZFaR2d9Yd8SN3Ugqkfy6Yzx4yNWrU+X1WA2C3iHvV
/juhm4lfI4VI4qP/Eqdq9sfBHvJOil9T/2N4zJmHz8mUI2R1unEwH30lf6GWo1Lw
YXx283qfE5UJ8kC1uRxSwhe7M3Cy5fV0liZqFAg9XcTSWrf35vzrfQajHojGtXEz
mUup5cceOaeQauM9ZWDKexWyn8KWG9skO3NPyDRWKGa9mk4BKKpSagdA6VmwCgNp
If2VU0otME74ydMRw/FgVavO0v15OZzGY0BCVZhz2Eg3rHuRvShw+r8jQINYaX8a
Qseiwfx6tpvpSJd0wLIx5dN3s82aA2pOyAT2qiHEF8AEI5CzpXcCXWdqOkgm5dj+
1Eu1FMA7Shv2LRUhjc+wbWulM6Dn/LZ8Wk9NeSA5LpO3LaHoXf59bMjWGCEHdVBu
ZoibhHgwqxWZvNzpNVRSNCG3YPTMeFPhaYnTMRD5dfqVQbyrz3hZ7ohKgJplEOnE
njf+7zgJ7l0S1VaP/uIVJLJWB3hoa3VtXGW3SmwIgRQu/TGhQftlsQ4ztfwvMj6w
b9TfMzqHYiCnvCGBaXFDi1Bu4XdLAZ00uZDzc4ClXrifPSQe3LbbbwLjyOYgqKld
JMK8aAbgIcMnx7ck2lI8xQ9/vQ5oIHNmfDc7hD75wE+fJszfB2HeiICbis32gziV
HpXfq9zbnj0GYRVsYN3/5eR1jtFkXv1DfgIiHY/VRtED2AIE01EVq5z4y02ZMLmE
QmiG2Hi/+QDK7TqgIQOXphDzvh9SUos+NFnSZ8KWim1q7zNPAvt1NuBAn/RtLWC/
TfkSM78fAxwaIOsTZeyNSF8QFdcubMJpbmMQyaxNGRLnR9mgxLE3gnFmPhukOJEa
V6wwaCVEtKtQ9QZbwfqZgwPVksn7LRQ0XYf3iJkqPVv+pFyPtUXTi73HTVuDd1pE
FdzQYFdvvOwxn09GKKF9WfU0gTPHob7llQDQRnI5XsWCz81BdAuu6oOtHtjbMYKs
O9XknrXgPWVsh7sV0c15ugfmfciNxkJe1uT14NK6osO6g8qIqgLYBEv8JKCeexxl
ztVOfh56rejKEu3xmMtGjoAZZF6aRl5tIb0k0uKtCp+/bticDINvHLew58c3q6F5
ghWI/s//L4yuYKRXYkNP9903LpixQJLwBfwTnhOka90zsnLy7MiV01vUKNhwrpx6
UL4vfNv1/UJ7dvvlTeV78nry4mc8VWKDjoRnFgyCnYVX8cRymzTnNrLduGSRwxlU
sqXcGwnS5Sv5o7XkEs7cde7yrLq/Oc69Riz0dmeLDkz99Yx1hg8RVkoMa1G16RiL
cLQaMJbT/d0DpLJlB1irn7FSQXqAx8GIrFd5JKbPbX7pjmpxrr21enaJ8yn/FNBl
mnE7ICnhbvlLKY2B3LSxsLy0jRRC7eWO9rXbeLqiBxz2H/jBh1OmgWwONSnoAm7H
bRuNvpqIjUitTYimkxtAGtJ6eV4MqmU1uwHVRcO1r4GL7D3+yrXKIn21dyLdNN1k
D8Xt9txzflmTSDMfqau1fX4BFD/JyuhEwXCyT99FYfQE9fKvqojyxViopQ1Qn2T4
PhoNOqS9RfBXWIszfP4hFyy2mWezAtCFflHHodwDDiPsIXCjXsExx9z0t4SLA/KO
wWwW2y9lCubeczgdG8BpwI4oPD6U8V1z5Ff2NSQCStu2cLFPuA0LbzARC1EsYwW+
5nLf3YdV0LCdmc2Vs+lds/03J6nRY675FYfuNXmKCz9IJ4su9/PpPy3VTy2nyn+K
MkiTjxP9G0kk4fycbDGJFgJbYH/BqKqekUW259ewhBW32gy0u5RHPjjZb8hGF7Pq
Kxl0sbiUoHCQWLZ0h1coC3I5mt4t/j1Zpq6vVaGR+NB+OvdyQpw/C635a8RaXyDj
7cwMXKBi6Mr+H9zBUFMdVaTNRpJX9WremgbRItwb342yE4DqIkRlBdaMvFyqKV9z
9vEFAlMYLm9BoaBvrhZ+1bD5QMBp2TNUmz8DQ0AQGDm3poZc4DroEbVIvIeTsQiD
Ok+U7LQTcnu01MyUHNzFZ9e/6KBKczFOj9HUTQ/N718XoAm2hf7K6yX682bsXEFR
tGxyfvURGDS+o99YcohN5cCcNdTvOLpd1TVjJpVu4cgYBXuMJBqPQitxcysOmFwx
MCsuvCRqtRSIaRGnCe+O28pFD7B17ZN93Cas0cgYw/z4Rk4xT5rVrFCCiy6AoetZ
n19jQQElzwcWiEOCS6DRTnv+pEyZ7Ri5FzUQrOVZyQ3iApB6xzQumpLjyRmlyaYC
dw1LnKKOpuEteRZswOvdmpnUKGFxEtJdn6kRmkneMvq9uXcAD/RdR9ljOCmHhxMP
uC9NwfTDCYxtgFzIn08B028CUKeuUYeN6Q7D5DjpvHwebpEYDcFwIkfK4G0VcEDy
T/0jdj0ZJMDMlwbnb/vdjI1NwV1Wq6LK8Jj084WZ1eg400W4fGhRUTYRDyDW5lOs
YupdtRKR99vpYOhPjyQ33E7LNFQahgoh9tzrLFYUd5327f8Vby3sVP/RFClN2lWx
Y3WzDEDMvUt+YS8NU7q1QaA/UWai2OkkXmD/z5lJJAgxVn1nRq5iUNJXDiZxxdGG
FMxR5GJifGCaFPU/eajOEcynnp94jsmsQK946T4D4sGmwWR4OkmTq3GxFyDRhWm7
fdSkUiecthEvbrg9V5vh124xya+zuK63xiS3wV+ucht10GWtX91G6VRmxK7YsMpd
oFxctoatanTH6iW8QCsmVC5sI6qx4HhJZc/uOy6QjJ7xLzXNEZCHl+QleKzK+p7m
A3yR/Z7yhiX7JSaJrBylnGj3e1S1cKgzyMNLPYsLEn2pcnXKGi7N/gfL/sKcZBo0
Vcxu8f+hDqKES096BWhzTaHwxM/bfY5iEmav/OpNGhXagXcWF94m1mcbp/o57EzE
hAYx62wPCXbGR4bwIUAn9JvLwx/mQ7SsCi0xhTnuq1NUtIt/wHKit3rwSI2pjkjp
5bFobBt8cqf/jSXIs3sBgdn3oCaP5fHMIai5B+lesnIALoGtMy8hK8Jym4Uy9To7
pqcrnTiAVsBe4vJ7jPty2FDjwr36mOto/i1A0PoOlTToEL4UH02WXIXnaCaMPuS/
hYS0eezwSojWfWLBaJHerAJMrV4CHRPJeUP0EvW+lzOQL4gsM6sHXFvbWUC+1fyC
zftqHKtjYpCyjTzlPNvEyJ0COq/ctth4jQ64KZ8eCASPfOqM07RJvteLz9Q9DVqD
xhR3wAmwjETENPzVKd10pIO53a+wNi9aMGxXdfwFj3E1cEhu/4l19sxeQUvMdtkO
fF2CY7aUuwkr6pvfKH4tl6i+shYSDi9D8FZd8Z6OesSvTl/0Ubd2lKwOiC87rE1R
l0tUNr2VIB/023BUn0/+YrFNNatcShRoD/ddDs9c929Xk9kjSAgQaxQX3LiEx4Sm
RpPE+HWq7azdNhDlXqG7dJFvnIXkPJmV9rwGnwzeQSIAo9MnHZEA/QYR+uZHsn8B
uBka21Dcugqy6nHNaoGCenbz27VcmzkQTeEitHhTZDw3JqSmagYDsbuTYnMZWeps
vykkrlbjKy14+CygYJahjt+kERHWAFWNWjI2QLYKISD/YheVdr18NYUsDLx7FGIG
M0XRRJgY4wdRek63uhomAvA6E/l9vsgS3ZMaIc81nsPwAfcxKCLVJQD8gHrJL2ki
wql6Dwr0mo9+25CxpN+7yd3pbFSKZtbzHoawrm6IDocG/RseTTewixiGcsVLLH1R
sLWWzlg6Rk4Wgd0CtUwKoPSzoTdAgML7AV/jgo9IOXHxHbzuQGPpP9Oi/pvEVWuZ
xTytSffs+1AvK46nH7gX50h3Ti7sDdmCk+1IMx2ZC/Rq9AdN7WxOn7zdVYJzeyOh
OJmzceH+YbmJAHMoIIFopAO9Gy+AgCIYsfMD2IelSGY50M3yPGXT8kQY0TA77h5Q
GPLQfvzaGtCwhkvA83AFv4SjCr7mntUPR92yPoBmwxVeload2XffNxUdf8sV+9m8
f5XzJmKVbMhSnURBbC8UOaHBMpb5rYlNMsfz7M+pqNAAS+/+popiCrRH5YxuNbNy
htD460IE9IbWQPTOzdDFnRNgZ/gUxnxaLgHmaCriz9xUZ7RBGLqBFjsVEoaJFj77
liB/2dmPoTLIPoeYbH78IbAq4ukR66SCc17Dom2zE295GoN70AuzF7zFZPPDPxrZ
R69QYZ1CZgEF3DBeFZvc0wWNu8EI5itTHCVr4CUay1kojoWRpn4wEuzOEQNHvm35
Op2Qj7Bo/fnqCPuugYQBTIHG/ki0qgzxuCSkVzYc0qKSb7tS5Hr1jI7CVeH+ISEr
7dpaZTBTyTeXMAs/PzFeJO7Q9RdMskq28DGwBew9AcgZ9LaVht/RbJ8LVWyEKD5P
gfUTKkkr/RcUvU2fHHdBS7pZV6kcrg2UI1E0sMSRA5PDAwx9FxervqP/Ei+pSchG
0AMnJmCu+Qr6PBgr+x5BDaXuVftqaDnfKMLOKH8fJsH4m0q5UzqXNUZOgt3Vw5Qz
tuG24T38ijO3ncflsHLX63pB7jQSvmy4QMhb64Aj2XVuXxS03TGUUxsuU84W2ytr
BLVim1a9dPwUKCEGxFfTDp3wKFMlcvNgRdZom0Y1SgQnmuhO/FGR/uDvBXVxp9o3
mVDOUW0XYaVBnFV695tdoIHRAe3xamcR+AcThESDPyb0LYzh4d7TScPs6M5DquvZ
9fV62x/zuYIGk99dr6L9h8Wm3C3JrPtD1u492qvnAM+n2c3by8fR2T/Nru4pbf0k
1BsIdoXUp39hZ3vuso461T43AYw/YB7JqrSgdMHoS4gHfUsQl+tOn1goHTUtf8Wr
ECYjU2LWUIUxiQn1WZt7LDlqh7bwYRG7/gCzUX9AhES6D4V2SF7mHDc8oh11wb2K
toqCP4NzuKyQiN7SoNZe20f8Jh7I+7aTh+LgofDClgbft+TO9a+7cpbtALDQ4KWm
C5UC53C+Ddzb2VYs6nHIXhxjCnoIDzRDyC40a6EcTCnt5M3Tpo77FJ0utDdqfnjJ
mJIr8E4fkHVlvlFvmCoIWVJ38Pzpaph5McE2OzObSum6A2KmFKXRWGeWC6B9swJr
qT8KxEKqx07N+Z2z/vp/LpVq2k9E7h4//USZvovhHsIV0FqKRyqXyCDzY9lsso8a
AcYdGw6V6vGBr0E++Nnb2GxBmW2EjYgGc15xdLMxU9s/bOLQLaQewKqtE1nUXFiE
s5cN9Zeg+5Z3HOJb26A/VXlbwVkWXBqYQugbZQ8IQfYAnGC+pRZ06y99lIFSLJbD
6uuTFmDzxwWc9GJzplvTvEQ4JeguWRJx0g5AILRobSdZ7zk34K3TZlZ/UOogPmBH
9zF62k6J2PX29fR8fPXv9tXnfxlNwEQ0W0rb3wncjeZ6oTmhIhLyvZ3mCnZ6TVzb
HG6xBpylQbiTQiYAngGPKA50uchq7hNrrXfsBksGxRE4JAbblcJ0NyhX6u5nvzZY
GLLFIkQ8MQMCDLY3ulpJkUjQqZGft++k1CJzvsVVAyRw6MY0vOjSFSjBUtWrcC2r
31qjW/u5OGtjUW3HLutezR0894M6CmGSKVzHumW9ke/3wgrEBMPjfbZyu9sQd44I
KzSiZjYmYjW83kOUQ6gZwDJmukVGNZiHS3ju4exGeAxiTlq/YmX9FylPpSWEReQI
iDqRuJD1p04C5hzWK5OzBrBYmsGOIHdwF2FKRMONPHPCsCSLckbExtt2aVFZgUVT
02I2hH+wRQQ7MG0oxe88m4MHK71c/bQZbxaUS4wTGVPpVXVVFyoH4aQerzcmmcY3
urEY80XKbXAWZ6pEMdcmsvaDU8SohXzROFw+wOXSgmHZMthbD3W4p7lob7IZCXwj
BfajI0C5vjBWhNsKBnlpTLnzAnbDp8eVORrqj/J36Zmt9ZSib5QlVcN4n+UIl004
XfqegypEqHLnNZMyYsZNtBCMvghLXm0NjDGRfwI6JjwRAmHA9PHpourVJyDWH2Vr
BN4ZNIQI3Fe0vZ6kiSmpyZdScViM0O80bdUA7lXSzY9Wf4vigTJbC5yUgc4lOohz
DyAWdzzmVDhDmIIq8Bnk6FfJWdFYCpbXIek5Uh0JFBb5Udcc1iVcQNl8aZntzHP9
oMIdXkXoNGyDNUgNLqQg7P2uAtcz48GjSAdjxG2YgzjQpjkNVJC/xU72RhiE+YD9
DkXmg8JAAV5j35ShnA0X7de8dEbLWhE7HYCAm0hIudhkWJwGORhPH9dZJEtLhZJF
5GfRvYzHagUH+e4sub8eoHhWR+7xfD8Ff1e84gTWa9FZ4zX/5o1JWTv/NDXh7eUA
jRHgFOcvxOHSdk/lnui/BEan8I1gv8TK1HFACR9MrtXWU6gOnIF6vFewrJJxIeu9
W9D9gaou25Y6dQL8qPlg1CD1pe+RBkXfzQm1Ci6K919RGsqH02o5DTSt86au1pVa
gi/dTtUtBWmKKMCCY+IwiBC7r2xB6FieIosoms3pLh1rnDs9NAksy/ul7otORTB6
XYpv8/IBbjqUU/LLCbzc/uynX8Jh1RpXIponI8FeXyzFuh2JpvyVThxIZXYey7cZ
fuof5cizcFczEMtv5SBrXIZ3ERgwySKxu3z0N+nuMgS2DDpA1IxKo1iOW4dpent0
HlsANCKxszAiK6sQWcIk9EvUazGXYqjnS9HTTqSt1eULceSMTfB0tUF/EVuomhEx
SpGjosMTlUL65GA+uqyLRu2An26IJrNqVlc9Dlxe1e8luMvA04Y8HrBrWxua1F6e
LKl+5uefXWjIEbhz2a2xep9IWHCQKfdg0qi+1ounCeUCSws/Wn4TEFUPU4FJtrku
emn0lqco0s7c3oIapekpd5YHpCF94d8KirYW5M4r43DVi1ZGDaR4aawUnNPN0Bu/
9rnIMEMNrKREUcTSMeJI0mVhwZIVWkBGVY6YlpgouynE5XyYNK6RNDaOpdUBhgOV
L8FcgbCSc04NJS5SyzJyE1qNeIBQB5uuJ06RUq8ruH642VZvJwg85M88/4wS+QGD
AhpOwJEYW8ntqF+gt7Ltba71HpN8D1wM1ZOobmwQzfnXQygb9g8+nsWECsZ4UScH
VLyWP5qi5uvroIVCE4kADW3C4rfttW+8MwvQhhDKqISMZbcYSpgyNZBg3lvyKwkq
rx0aNuSt7zZsej4fyXyIxYZzPD7Vwb9hOrdg2ceZ/PYWPwg44u+zv1gaJS4vJwhM
aCJjmdoxabRMJVWXQ1rNO5PeFjFV89OV5cCxyx2NlQb0qdax10DZ7hgXWMXc71NN
+dFImAL+hML3YPOrJKiPFJNIfK0HmZ0C1VHmOgG8mGpfI3b87Kp8cEuFvTn2t5qg
lSOdhQmCXmT+P1qK/odPVdnzFD6sUjE2G061pZ3GfJkJbTHVvtMSRU/WmuWZCd2n
VPuplmH1Y66q9sMdx3Gjuayj/6pNI5smiVrXR7Tdex41+Y/DmNqvqJiZ7Sec4VLs
fPLhy4NEV8K5ibPKv9jVTu7nmXzK3BjLxOI17BFQFH/fdJOdVwZyLHhJIAPwW+P0
zNsQOvdIFuuDyFduxBWP/NH2ilnDdQbVX2ZluDt2qvXSKmyqXzpNMRnofBXMXUjU
R5pHVmSp6kLQM1jUA+DtmafVMSN42E9EPIIMsIDvdszwP2JonzqUoco98RlepR4C
5cZmMaWiqDhru3JVGLhAp9JSmz2Hhw+u28K4MEyH+fX+GQbr1G7pEf1Vq+sMkkb4
a1q9WVvHpcMsUD5CQ3BZZxaq3B0AMnZ2xvlxtLBxjWtdqA7dG8aTXgpfZ1dH88tv
Qt58PcOZai8vxwG4BPlpfhGkPj1I9atelx2JqhuShWK1Dvlo35pAl43+kPriq6FP
IeoY7jKD44BCMXwFEeNVDDmaH/XsLT/+mcS3uh9iPErnVb0h0bs1S8xcpfF2qpRl
MtQcI/OjRgGCIiW+Pk2c4Z/cbVjNNxqhgWbxBUsLHnGQM/oj+Nz455ayu0rQ4wWV
A3FlOnWML33np8GqopDnj6q8hX9Cmt1YeGYb6KVaVa0RrLt7g3dl9uiNcrg5jSaN
r7L33KwpWmxD/uJojIiY5n3JRVHfE7uHmoNgt6PzAFTz6imM4P8xzoT+Zv7HCMKi
0HpbnwW58XG0znEL7T47idqVheV9oLjukS8CmKkcR0+xeAd0kDm4hNx4IabcmglB
SylYKGlC/27743+AhsM/lYbbp3AL+vPxLnr+2ArPmSdQG2iDAuiIcaIcf+x6Fg4Y
XE5za9sK4HD/u3lt/lLeppvkTbXh5RSV/tX5Uups5th3h0YSSv1sxl/uPanEA+N8
UMDHq/EXTkykFg5x5HHV2FKlvIdd7b9UgIJuk8KdWpMNnG2AgcGn6ps9HQu8TD30
lVrF179dOIiFBhGLttjomjdEmaqztRL2Z8u7BH39hlKYX3uRJttyNP8CAd/5R0tR
20UdSSsUQ/4b2pQ5TYkRiww05/350CsFTTBJrPmnCoSinBeortneBzpPa5eCqRw9
Ji/eSvaS4ujdiyTB8mRsXEs2QZJIl4EoBmZ7Gzp2tH9peqGcA3Snvok+oOoeATTa
OyAKug5j6Jn2M8aGjKpndmJw+FjYyilX1oaSVPnDbTmLUNiZl2tEHCGCo01f0wSd
CsNdcB46md6j8fnTjOq6HQXsINTvtypR5mR1feW0THKvESyXr6xwuQz2UR9HPkUR
sEttwSXfEpm2Y4reIIAQHg+KkYxcNxhFu2x/ppTL92gy+tDa+cxxypMcuZ0ltDbH
fCEndmqAmzjo/qzfr6VlyV4UkgooZfPX2WyHQPoM696hYN0YrP3rFClMMc9WcRYB
QCw9uoDrUqnWEjnTwCclraW2hwLYImIiazU9wrV1RSM8tVSl5BCN03wnB4w3KO8H
hyjYEsSf1At7EoHGhboHO9+NNhTy5gzYFM9I/ZVReyQ40K4qfOiWxrU/PR+hdLva
jA1nLnVIzdNEvOy0JVQxwevnjnX2Y/2pL18T4rqJLiEINjNjEll1DWeZvCXHpq2/
/UP/e/gauXDifMGgg2rXG4EWbTlelmZr2kZMiKeNlE5O3kw8n+MBIzHHPcmerQkV
VsCApC7dnY/EX6eD4xuroM0JtpjA71FQvOcPC3fynvrLHpr8I3xdVcD0pMt/GtPo
XBj8jgUvWtmu4lSWGdkfmGOPjVjX6HYoQfB9iAe1AXHFYOF5pgt+LS/TYqhooY7A
R1lrfUZHnKbF8v5evAfoywIdJsow09k1+KP8Id3T11HrwskNL6XP28oYxYv2d9Iu
/jL9elVeghJN3W7aLlil695qHYo9uGwwLeQBA3d5LH5V2HEeT6YlTH//MpgrlRzl
dS52Fg8ErRvpdhKRONrWWEdv6HVmW+fg+NQyMotqPKWyAtBxFMMKGC7bkS5EUPgT
kdIVXG2oczNgNFMLqbdFUUILm/lusp5URv6dZB8xd++2jo5KNgIBeEZCnb7X8A5O
YkLGvaQOOT96hLyDDcWrSB1eQUKcl539px74UDVsnhjAt37GCy/Cx59BYa5xM/7e
DmImupInZkn9QRpnFzIUGsGDIARVdC9AJfqWqJXfU0OBv4hKD4pYYtqqUvmfdOSL
hCOgEfQ7bDwnzWkpW4w6DyPk1tGPaQq47UOlaQomfIT2EB5DE10Bp+KN3saBAeTC
ffRL6+uS4CSTnNjUb6kAiMacyqhrRnktY/sH5Ig/w2T214KYbZ0r60d8slDHnRr2
o7Fn2WnZm6N1L8V52HjznzarALJydBvy5ZGz6rrLNGfPQ72vXUuk1wk4s+HLu9jg
rF5JMcK7KcIyYzFJmh3kFHmi4Ul+AdRf9gipCo7LJQ+yA+oAuE+MDWcv8Awts8dp
ulQLOh5wi9Vy1hhl+9X5851LeRIhLFy9IHjBzTpGL5OvUhdpAg490E5zPkZLSV9U
kfsyq/QdXWZrVHD5W23Jr8U3Y4+Lmae+l1/aw6F+4pusaHJNCVDKX0mx+Z1d/Ign
omctv2v1xbPdAYDZudhjm5zSVM0vHT4jCHy1IKWxFQq5vCXjI7eloLTacdKAuj8b
yBi9x9I3rZa5G+xxJ+NPYJQgrJ5vBtJt8YC3ykJNYQSlTY/c20sZYt2Cf3HgIL34
71BFau/A3B9JQOfCk2viv4UV0i40YkgnvgcT95wgUVRE5jd7JcOJTSHmVvn7R9R2
A7lqVrYn+Xklk0goluRNjCIcpgwlhIAL4EvcRQwfzmxwgh0D5SS4t0JnON/WNuXg
MA9AS1JRTlEzBpgPgGGt7NDjSsYRejmTx1n6hqtQIFiwClWnFFThSstse/To/3TQ
QSj61R4XUr/mS6K/F5t1MluWp3r0nDSpVzbTKTUkda6Juq7n4KcitXbg68M4A85I
0CNv96BpkZTaDxRnNW0rCaED7H08dGjNdc1pNoDmk7+ut05dGo3zYcfa+z9b85A4
P3PFJdCEraVJp7h+GrXVtUvrOd5EWeNLtHF7YLvyYb3Y4zClNF53p9VExLN4/tOr
pbwQg42bUuev7dATb4yt8gfFha8jbtl2WCfg7KKUiMQkCpb4gXkVXSU5sfLkVr5r
4V6hN4KBzsY4+ffmD3YGmKJUKGaBRHWqDvwoaElRarEOfNTgf4shO6LIk/wMEo8u
f2cy4cTmh4YCRbHHSO5uG7Jv0YO4UbidxGUP1pE+Q4VC5XJLtdFExn5yDpT6FmtM
7cKM8zaUf7Azfdpeq07dlw60Ki19qccPIXRF8XB8mjuFkISeXtIR9BL2f80fqEtN
+zb3rgxs8xSTJw1t1JNBIKE7Z7g++jD6xphq9xwliqoSwW3wOscO31KBmBDvRQrA
2ZVaBFhpYym/ge8fjcsStGViB0rJtGDq2xAyzPAgCRfVuhyNQaz1YkYg+sv7dkzO
sFj3yxjqOzekdcalBNmYalNo+Ly5jKDyuOVcv8IUIn8Axq7Lj/gGjPZcdGcmPSzy
t79ilaXwr9edM/vf/kLFLK2zfCLik0zuCFFyFQLUJpRhAoCKsczdmMDFusn/9k7l
E7/8OYoFKDm3o88HnmkEeiGNzNqVxiL01QxdI+ZXE/G5azB7lXrmYRvGEVEPepYT
D56tNGZvjyGyZRiIf/9huKL2d9JtvG9fwNZxpr3fO43W6Twdv4e4+eEtp7J80ND4
H281bIEEY0Iz1DByUsoJC7cHKHyxTFAw2gSMDkvY4VZLW2cX2slBFte455jEZ1mH
7arBDqYWgHSNkXEj2kV9Euc52n+htw7aWDwnjRCpljeeAIc0RXunrieUqx03gbMq
GI4Ck+y+HSOz1da3MBojisd/m/FB5SOEKSI+pTbf61lxwWHB7779hdulo3bME5RS
V264Gxd2jrn3H84a8ta3BWKBOWPa5/7l+DGqxH/GoNM9B5JNzP+EB5Zl1YlHSqzv
5YkyTvmosLFwOxtAAE5+dL3fHXJN7tIsbd+/gY//1Lurt2bI7qbQ5XvWPQvwKBv8
k+XepwAn+8KJnXxETPOVYEOWr66pcuin11Vpl1dfXhN32GVCpNJqJuIOmcdCT1ve
rZ4pqbcULaL7t5HVmRqGn0lLRJ4eDs9n8VhGve8PM8CeMMXrWDVJ7oeHzcDoVlLU
dHFakEZiizsEactmrwQ56nv48stQd/Rt6jV0mmxt3gbsVR8Yn9FeLL49dvQ2rZ70
Miy9u6NtcYiuIIXquN0NsA9P+kUIMtaXGRJ/1xqxwhqxwmPLtMtWlog+CXlliH+s
YIjCjVBvfO2OBHqyVQ7oXLEmSsEqXkkLnOM+eUvvyw+mfChkOJlT3j4EoqsSgcrg
JhWkubg+i6mxaejiggqtRwIEaND40MsgG3yi6DcwXhLWdJxxAZxPCyPTqiY4xqMc
EmiCxtw4vZRDLXPw80esBX5StGSTwtZl2XDjPTAqJJUDwVkgNFjKFDSoNsJHR4t9
PHvNXvABZEAyurv6OndrWrroSVN5kRD/vzJ3L3mvRsEyN8L9IN+RcVbB29n4itDE
4SY+e18F8fN60Q7vEkm05N2wC4BGTgcjhDDi/58bSbOOH8xbcM6LzVmEa77Pbnhc
o7TCcG19BgYYavOmRmO6PzGUA5WxHExfJY+9lZvVMAmWzfXzNrYLBthKxmP7Fe/j
70h8q5YAlJ1u+bNE2f8Gb6G4pKT2Vj5UStCnsZL0da/LK+q+7v4vQkjJx9AfmbIz
sFER/NwKpn3mfPuZ2xOE1TKXmhUgcPj8sy1XCOOBEfctF7fmB6sI2acUE/buOtP4
sP9lOh1bmprt2CKJmUqgLjfx3jqlCJSajyPx68MafnId5rPiKkjkMBZnz/G+5lGL
rVQao5LspUid8AUPoFOe0FDiLdTmakU/5594MvRxLAUovqDC75s2WVzFFdyAe+Ao
ZYqxgkfcnh7sb7Fi3aND1yOCRyIFPLmKXV67CPNLdFmJY47mk09+KZwh+UYqX1sk
f7bMtIz/71atNMjGTMRghwzDra8OvdiJDrxEDvSoqfcNZROlq/No3tU2WxHDKMaE
4J21JLVQ6nSmI5c6f7Lhnbx0S6ysa+Wku0krvK1A71ly+nWwJOuBT3aT0suF17CK
3gknCfo0ydchWIthBqqmo91DQF7ICRM1zdAj/mOJoeFcfUU4T2K1c76oPv6QDKl/
41QQFteYgNY8TGU4fEWGimonwlHNjfN0SXp2yKeeJ/o3+W+M0bL2BXtSvdccdgoF
RU2NuNgCznXCzPNbk8lpgg99820Q1V8Oas2Q0ADEb3Ufi3R4ST9IuCZaO7hvF79P
AG2ELvun7E/A01txjcNn4Xgw+VnvHJA4CAG7m6XVRbinwJ99770yXV8f4pB8fubk
aYjdQcbwuUn9ZnkmhT7QhIF5610bTqzz2ezp+n4Hr5Caq7klkB60jTcCI8LqbPa2
aYY23c5q0yhhTBfCNLHOotFGZ/1jrsAZCYUor3q2/k/JqnIZ3mNLaKrhlDQzH2mx
TyYswMzGNEtbp8x6p3MR7HmLPoF5Ir/7VqPWYH+hGXkcgQXLD4ifzTUOMFIf/zW/
jEAh/M53bxPQb4jKkloti7g4+0QiqRjntBl35NYJeg0K0g8Vb8iw1IsmqHUs+mEl
IKN+Usi2ffygSMIhFcuPH0J3K8e13JA7Yp49+1kg85/hOEngHmX1z+rfgTN16t+s
/W4ciThPlAsYCE4EZgY1lr5VU6TL7schvFH8qKCp8VhQyD9Hg34gNx9xZar291r5
w+kHrAuFvYny3F1Q0u0cbiLwziX+TjbEKenivClSGtTlFgZd6g0yAuy6UlrKu/o0
KJ2ujrOtmzGLXlTpI+wx/rtPe127OYH9lm+jtoJdSsTh7O+EZPaHY2KxLT0G3fdc
skiv1B+8RaJ+Cs+MLbF4JbGM1GsES85r5/jXBJe+oq18aq3TFZeTLUCsAsv7W/bc
ViZYY1Bxn6bQJewtCIYsuqglyM/qy/Z67J7Ii6TN0+qPBIhn/WSrN9WAD6HzCfxG
hyeqtiD04qKtU0bUgcJ9VZcg0yvq0ewRyQrkhS6v9YIEtJ9R5sO5DQ9IEdQtbb/3
vy6yKapg1EPMgZhVNkKTQ+04m+A8XwpxjQmlkuH6YzxUGrtcverCzJXa3WynYWFu
Fpmkz3qx4a/6GOEMvBGtBaKZjK2hT5uj2sdhsgj/rFH1QERqlq81unf24XTRTKLi
hIDIDSEsi4Wo8eG5MZ4CkrxCjs+seb8/82m/IjaJ5y8/sfrtAHthaZ272OAX4udR
E+ZelWXbp5rqYyW5SmfvzGS6tg1tXxHIXp7WidhTuzIFw6uz6rHbO32rM+2qQtaJ
r0rffAjmM56fCI5Unc+ue1Cw2OTk6djXLv7eSF7+HpTV+SSomCIDw51Rj2T/MHS3
bXdWcXJ4uAoC7XFvPDejcxkIeuCMCfyWz7armt7/cBcoRxCEA4VYdLBG6dC8BGXv
bjBNHI3Ym7lRm4/l7IbApujkbsTlYC9ZvHnYpG+alENRfvMWXnHneXeZlPmnxoKw
iBWpAlmEtmJZlE5uQ887dUmf2yRfkmwbit+sTG6b02k1Ra+aFou8iR4uphOsk/HC
dcv4GGonmIwelktqGRAsDLGJf3MNzFFIl7Mo86Uf0u0caVDUSeil9eCfGYgBF32g
vCOpVnVKefdqNUnDLD6jv0oWA3rluzX9Si5VSHj+kQuS/Gn8tpFfkpg77P+P2iUk
GIP2hvcgK6q1VIs55+r0V4mX5Aw7Oxja8oriPbJdtv3xyfsvpaYGphClR7Gc0LcY
pxrzvQyCO24nG7YEKdyRQ3Kt2Gj6PU80V5LK3JqcE6G1aVnlPwd2o9NEzuoULjDr
yL5yruGK9jJ5jF0PVFDlDRmD3EPTKkdHmt+W39Lao7k9JhnbcpcP2jpy/rvZ5eM7
HIgqbuziFrVjXAMh4OMv1OdxvkGNISIQksukz6EkpwrKQ/pVuVGo5NcF67/OYkNI
VrZ0swrnhC5gnk6t7qNHI2002IfYis25K9OgYF6WmCszK+ZcK9k4Nvc0MCW3xZEB
4wBQ1SFgHlDNXK/h3VOeUCGLcCtcTSDailWtJvD4GRfWqvtbQ8PQ0g3RN275Bp5/
SHX86eULzV1ioi16X6Y+HofD5cO4oOeaMUdHjFf0tdoMGYkxWEa0U4bxSzrHRll9
wxah938cZZcjD/q+o0odnofL6YnQIxgeiUzkp25jCX3I5XB/oelvvD3DNQStERQG
2AMeWasRp4BKNkg4mtW3TW5vIdaBnlKJ7GKbqwz/Yc3A8NCacEWll+mx+9Jkhtdk
fte09DLlXj1W/xq5h23XQ5TgTT8StY9N2TVxDFHN49BZ1rAq5tU5D22VmAfPS7ZP
GabW0qQdMS05JYHnkYtxNI658twhI4drBUF2BvDzI8CyCXv9mV0LvXjolg0Q9pk2
Z2iFqo7eY82mIC0okGjQKjHizZ3+0EOeahv9ocG25IAAV9ieqjWDj3eHfLKO8igw
3ijXLDMOVLEDrdrAnl85iQiRdnKupbzbCSDuYeQZ/pE05bDpHPbrrbGpgEiXsp9w
JTOUs75SpdoapREz0U/GZ3bI9fTbbv9Ha/E97oggSPfhyrv5LMQnksAHj17QMzC5
NnMDjdSnX+JziAJ/qzdJ3pQP9kcEvPUIDTumi7rtNqatlB/VAVPOrsMU6kXdTa+n
HYWt36SrsFWLs+NmpEUuPS2nEOHo7DPrItYQaRKWB326nDkf/JEF1MrEvWmlbH3N
wupVQfKOGpo0PoOx49f04Fc1D08TWCLfK8ywwAly1rFBrh2z7xoT/SmZJbdGuDeR
fiLQA6x5y0do7C7v7Tok3TTTakiwppmfMkFBVNKOOpb3Fh2U8v1LRk/JmKSkGeYS
wimQrOXDkrmKGs/fi4iuhi6s9ejgt+Ef2Kt1NM27TCnzSIMYkLMWyJc1HQPzVn1s
OWbAY57bvCwHQLs5fm2tDrKCW/vwV24BEBcGL7u2hz/sT7KK6E6SIiFusMH9CLXS
rCA5gXZN499xjoZQ5DRbPQ/oLtFzXjdt6Iqj8zkiUS9zxMJ1cKJapn48MzUJ3Wj3
f2i/5N/R4zizBY9hx/OaTe6bUMF2ce+KkdthqfXkfYZwu0JqEvKb1gIvZO0swiQS
8Q77Cmbv/LLS6e+yec3tti2oRWOFp2QdAzOu/BFypdb80EMcAzl1KceF+wvTSPLT
myf/xcSLqq4nQcqs5pEbELqXiYSnH4xrw3+TFHii7NaultYoCfixUHvk8QAk2p0r
lHRlt8fsTFvjWBU5ZW17ExUHb+9WBxIeH6preWcYcCuOMOsG+3QTrdv7Rjv1NkcW
uuK4DMwtTkn7a6R0MvhZbRzveDiXM+JcPHcEiIkA5/2ZNY0iU+sYl37VO1louQvl
ileBHXvPDE+SgfzLPSV18MBTR4vWuuI2f6lmo8gWQl0Zz0c71sTLS9BjwBx2/9X2
a7ymL7FQigo/BA5x/qBt3K7yJk0iUN4GwlgjRmmuij47UMSsK0ZM+A2B35PAtKTY
v1VuHq/ddC9+IsFKRVR2HXWvKiBL8vR75BdXSMBkXYV1ZcnNlJxfTCpUztM+2xzr
xuNKxo125wlkeuwcmTkAw+NsejdXEKwDIljiG/RP7iMfpbtKdOIWfWShGrgj96BT
g16ojYXyssPjpYkrpt7pdWqQWaUoGCnrfpW6feMy5V4sVvPh8Q8Y4g88LFxafUZQ
RksbAyT32C7DY3VjppYycoMah0GTfuS/H5HbsBXy86sfE9Hvz5zTWE0xDCxL9aCZ
swK7eOUmOvKIxpMWFelhgd/cN7i5Vkndj9GkvR55BrDCEOsCEMXUYdLHA8s0l8q6
5Vs/CH5XV9ay4hYYtc+JcYjQTz4wu16xcii70KIq6bZNYrI8FK8NkbPs+I5JoUR3
PTsDbDHZ2tfSXOk4xjv1gnkVHyqdpZV2FOoPDiTioCV0IncZ5FI1JBxZsbGCkGAu
jCY5ddiSZd7feogAd788onpzzUMQ4B1pKGyDgIYc0pq7dcWVoXCg2Ati8lbc17+j
URxAEMSpKKIn/iGXeyVyF0X7XbkV0WIypHGeZb6t3QgP34ivD8GobxNk9h4DMbDw
2s6QyR1sC3po4meeX0e6gWvg23a0T6cyIL1TEZLYRTrK4Zdif6jT944sMSBvpJCk
dC1CJQNj6UzmcfboX33se5EYcpWOodxllBaslRXxsOCc/qZelI0HHsR6ayolPJ99
g2I6WqfpNkscAfIIv+mm1SQVKfzEZ71rZBfLBxk4ozC1u4tLmJAsTO4F7Rae73IQ
n7uKPOUhJXqpnvMNe9JGUtvQbrBCiwdJWmj51p6bm0YZ8ttNYlVyfOzhMAMoIA9T
KYFAJI2Dre6/F0Z7ED/Q6SXIUJnM4os1EwVKdD2tNjXCBRv2C4Lg5jUwE/RjyM55
hBbktYwa7iSupXHFdRyYopILLRzX69JF4WHNEqVNr5aAbKBAmyk5ABw9zJA7m2EX
D2SX8arzILfv5hkhe405DfY0N3rnPYWsTgYuSDndOX723M40ZFtWJb7CSnw3Bnha
32Zw0Tu7UWg9nIWQPhyIfKFcToVN1dHYHVsV7jQm6+eD9iS+jgfHdg7H+1TS++ae
LdUnRyTESWMughMESrMsr3OOd7+bzXAWr8f7m7iSFM6JBzNAvz1ScHvXw0pVDycA
D4VNIHwjh4FW9bg3jBPMTYLq8GkqGb0vs9hT2THZOETG3bXFTu4oajwELJyCnTLx
ynQuR38e9uyTbo9lr10V9wPY8BZ3eJA3FEgrIVdGd67f7E8X77fKa7MIgH0tISZn
nTbdGRrGBtVRmsjuq2U2wuCPRTpAeFqYATtGHTBH56AvMUowYNZckUlXiPXUSwQo
99uQwmusgzPxUvosL0vEuzrY8nIdlKPiucqfhXb+aTikMs4l/985IZvhiQhmL6OS
poLNbYU+eGa2933W1xirX2iJgVJ7URGbcSQHixBCPsZk56EjWMqhKxeJLQ4/SsgM
rOwHQyD26tE7O6o233RUo84DqNwG7id5m/NLMdN5eCOifGZQzCjoxqEVHzUD8tyt
jPqU2kcgtTxQe/S8igLytptLjkpJNRQj8OLLISQyP3zSx21+lh0cvROILwDgbZcq
ttMFGZPtvyeqf/fOjQ5mtr9YPMpeZTM3+aFOAVlkNMmienUhqpknNvPS0H6LZ1Uh
il7AV2zGkI73yJYs0rmZeuOpp3/ZCOraFi4RCafF8s7o07rep7IJTVU0A6Hec8XU
KKPBEjg3t5RbDgeDqbVFHf2kFdbcUCnGYHxkMSbz2OdAy/Prvlyj85/t8Pt6nRWI
QwORgGg3lMvsNZAWR1NE4vvAazaNGgcuNtgD77OqVpocM4OASRI/fgf2GAygQex3
I7lnQmWEMzae2ZjYIMguQhX4YRkrIVFBXVHlI1F38EfoP25X9DKC5B1O4DXI68Ef
EZ0i1AdzEIYNlzDsjl8R5bqJaoKBJ23pFpYsppnkJFVxG5yUuE+I15plqarlPEEV
Ky5GJCF22M9tvxmet6ntBdvzn85SimjESFUVyHH5FreXhksfnzQ3R72cdRdUPTmX
/TrX74cz29IYqhFHiDT6tUMEDcBnv1NfnoJHaID/9rpX+uAmyu1heoEsa6lnK8Cf
JcWe+nWuLPlC4+/jvlJO3cwXcHmN9GedW/zS9CIqc3HhmBneKEOHpjN7H9S0XSQY
7I1K3zKbeDrLPCTPwyCTgQQhV07EhtrWjHhjimFa63PGNIFN8TsqwYHRxCY/fwYV
dM+WEqAD/4sLfWaa9q0vUEvb3dFk+KbrC2EsNUaXdGXzghfFPhMzUk+3T7d+3P4m
+oBZ8qxqFv3pAvrSv2W2qMJjivQ2KxuUhBZGopKjudyKpxYrliyi5O8PwXzfEzcr
YiTs27PBi7PZJov11YLP+GhUihDoS2PJs0vSbFnteASpKfAj60gHE9KhXjAlbLGs
u524x6AWa07q/7t4lCYGu6Bm3GK3b0MBaB6puJWag21Ao7p3RtLqJiyQBg9UiCi2
EiBXur5TJiBVahkwfbsNtnxCKDhkiHlTHEpGAnM5kY2iZHbO84pHGO9eC4JOCKJl
Q+GaT/CtRyoEBDadL4A1V5DmYQIQecPMGvCQcEWm5q5DHbTOA27iEb6X6dczogxs
ztzXxZMp7pB/tYZ9kYuuJqttbTpw38leWwlR5A5/8WxkwwZpWtA3jr6IAsiRMCPA
FP61Pyegn9I0FMsrHsN5aH7O0Qk9oRnPJE7jM28Or7V4dmSXK3pG4BUF8zIXh8K/
o8mFvhf3WSRoXaDFXAx7Nfayh1meqmOsESN4BAAN/X2Yui7QUyPLupzT9tu6AzDN
b3RjBIHBlyv26aTS9P5q4DGS7ArAYJdstKEWPDtbtkmKvq141m2xlyl/vlkaeC5j
0ojq+Chhu3bA6MHM98nNHnEIK5RoVJ0awKP6UOyrz/2tkxTtylXV8yFDXG3oiWcH
Y6z848IAwaA0/7LFFvkJxjkQe7xmvCGPfG64GKYy0sKFIRZDPSeKqJ4myi0kesam
7W8EIJbVGXMg1nZXPZcfzVt4lcRgpX7KsP2aXnol7n6OFL2Je+lygWm+5jH3ANgZ
SuXLNTg1/Lod05NMubzBALrb3YUMiTNexx1YJB7nP75r/qGCYGLL3IaWgZzloqod
5DqTgSe6VXv42Gee3fsbc5LMx+0OpSLOLOv4qWNHxOM1EjfyBW34id6NAYxS+DK3
mFGsC2TJXgtGvWbAZi5lDygUPlkTvKaV05YQDwyp/GRtJUrrhILDt7JuQHWFKoVL
wiA/gp3PyNV9/IYF97UF+bjMxMnYI7gMwNJbTpEKfhRCRpLKFTz+I5iQzSol9s2z
PGZIO4+PSb8BvswqN0CWCTcgMLtpqvHmCiQHtHFW8QC328QBYGCb6+hi/892WCoa
1m58mJMzi16EaBbU+UyqpRvlxYpTChG8MtSJKlOUa4CxUVOWVxtgjzlXpqBnGsCU
M3ILtZ43vwjie9WcCrom7YVrGWoOhFa/JGvG59ltnOqPuIQvXg7hRbncXRaCnThk
3rmuG/2ev9WUPQtBBtciJfRcoPcQO7+Gshf0bebRCUHVZ5iuqutgyL7IGTGUZ8Wj
nYmEZlOGgQKMYA+W8Vln/z/gWnC+FwovSjz+xzyy8JIPtNfUiW1rhYR6iG4tIqyz
S4phZujg0Lu6nH3fyMOOGRw+tDrlIEJMPdxdAKQkyzKBE5vhRFEfewJ0NL96FaWB
UCakGJuN62snLEQqNFrrL6KAvtZ41TReXhk4phRy3LwKTZpx94Q6tM7D8Ht509kG
br7ZXPld0lUAtqNAdUi2KY1oOa0ArvMTeDkGNRvxb/uxi51kid7jli2F7G84nqYx
ZoldHXRZcx3YNudSd1FcwbAALhMlT/xfcf60P1F7z1zX7v7O4VX7PK+TnMREGEtV
vtNzFbCTxksqa6k+PKW8LAHHUkcZaNmeSlsrRagtkZrUc/J+UfOSlLWXwSIFexJE
qT1KYQyKHrLb8AcaHJyHO17H/cDJ3gyDAzhkaUAOTb9UzmmXoy5L0iMO2gLFjgaH
ovGfqydjwI8oNFfhksOhEdSUqALhuiGiCj28xKWWmbomSoLO4SXIJoZTJTexMk3A
CT9nUP9JX0ovBQPmuaFFCvcsdP4OVwgJS5CuUhoF+EFkVhRjqqA5ZzU+gPP91Jcx
U4mE5H+YsgUm+qoVqf25/J59Yf6D1CCHitQ3z96bF8f0f8iM/UH2vQwMsqETl7Rp
A+pIZqsELp0rEufF+I/Xow==
`pragma protect end_protected
