// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:52 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OyqoSyQ3xq2mCjsk5GZKV0c2xy/hJUT9oIZZX2v3oyzsBVXRmCRSBIfKu19ees7f
ctQ2kFUcsLI79W+E0sjBOO1De3rIRr9atZHfL9GN4L4QARPDKLJuHYeAxQF0fN5G
c+cLwSzTmFLJ0tiHjY/6bPjQWq1w5kq4XURcwce+amo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5344)
efNMIMCcwwhdHQUZxmbja9dSEGSDSnpYN6fHr2jhTqIRbckxs6XqPSDqxOgWl2wB
YlHDxjzzwnBWC8pxejywW5r+c7jJcrkj/eshiXhnhRoqkz6DPieCacb3B3ptEjJE
BYX/pj+0G9qWAydOaOA90842/JCNNrVPmv3tAh3bA/NuWX7JfAHcUXT7Os9LnJCf
TeFl3moCeOc5d10QDkVRcIea4DRyUFp+ELC/fRrN+hJ8+aPRpAE70kekOQ3onz77
oI7piravDHBFBf1IFr+aZNq15aKxp0cAWJYMcufKDlzbzhJezIV/iWICa8Hu+yy/
5FkXwfrpgO2+hr0orKb3oDmd9+5JIZnvEN2fLqrXCHvAWrtoM5QV9EQf2LRnKzWN
TgIHdSJ6B3mX7J98exTIWgA2IujgNd96qeM3+fAs3YaAotFbaK5tKzwwbhCrm7oj
osXRVXXCiQmHwk6o1jRkKo6cqXKubsdwzDPy5YYzAleKkpW8lcbH6ueIlP8PrYkW
rUoDE2myHDcgifIgFlxz8OadRF+7aVUTofL5eaD+wmPqahWcZDkrn87TYE2xdt+8
lPOqeL1fUoNRdU69qndGDbz6ZEjYI32WhOV1URBeC6fxIKhAdlbDA5bAMhEbhrWf
aqYrDzmTg2FPNhcd14sb5Orc2280XRIMrTMZ4LXWtHg53aOoGZT7gBeB+QIKN4dn
nE+TurSSdALJhAqXKzjWWwoi83yJ3nFB7jorvUdmxOuk7o2V49Srnzl89oOz5C17
QkL1CcbfoV02OLgGnUc+AgzV8TWGU9awPiQRbExKLKI4CwJLdITFEpWQX5c/Yy09
Mjum3Uihd1qz2ITl9zJp6CHtucB5pC2JdoAYZIo72053/bb4PhW8a/imJQDYISNv
iw9vR6f5DBP9jr79CtbkssI55cVEc7129AorABVIWh9QrINpr0+RvQ4a3X0s+ObY
G3UQGPuiMnjR3eTlGPLlRIzyeFElPiw6Rb1tdKKlfzCaRFDsgZBv8VBQPrFOpbh9
SwVdd4bnGT0QyW+BjgQScuIuUpwbVOp/yXFNBThVkqzpl/2l7bSMbMUdf1PvF9L2
F/lUAHsmBC6OUwX37sZy/4PsMkrVxIC0/8TIE9QdTUNI3KT64WDU5Oke+Lq17P7x
z9Gp51dX6/7bnztoZ7Z2g74BfwWRmII1gB2QsYzywmHRvfSJ6N3nMbRGoHzoK8yb
JO0xXtNKyaXn0sgfwa6BcDge+7q6ACi2ebyTyHlH1HkQVajTBYmRYIKbthcr6PeY
m5gMk9CNtvJFQjkiI3n46hKzn7orfZv2DQ4LHTpy828xTJsXR/BSkRlY04yjvf6M
V1vsUw6ZpFhgbARHabuJE7zCoKtGpraGz8newaDiUgkgxmBUgCe9HvCadooE4PC/
j1CkAxRTTjx1NxQLFRSmuzfCSAuid8C4SUcPFPhzekIFAOWO0Dmj65vghBQQ1B1o
8BGuu+aU6L2muXRd8oQ1ICbHROaXXLlIdbAFsAhJwhJDvXH5CuldfGuTAVwteCVt
M/aE+EDlnVwzYCdebEBKv9bZnjIeGCzKC5DBnSUxu5ia49EEQVET6IIVb5eUgZSL
lf/lRuCyX1xkuIJsZuTYogAKuvzGT52A4KCitlKNKm7NZsYzXoWdKHlsCDv7ufMl
13BUqYhxRbeS205pFw/PEUQew5fkSXXORSWrxYZQXivPcaeEKqByPodQJjWHfmno
giZr/2mEOWtLNr+8Q9wuVJHbvd+ODVlBe/O3p5bgJqUdrYxgwklkYcz8lNNzrNrU
UrGCY1ut5cCXVBp9vlj9ji7O1gYzxCifKR5X4N2NjbjPXTFYA3rPvuhQ849eOo7P
APUW7ocKjZMo6OfTcBHBUfJWPqY4gGIVzC3P8k8IpnKBk16+T3iFjttp65mDpwL+
QpPQz74p/gIFMH/6dL/rpkThz3/KSc15AerbpOXXD5tKaFr/zsFOADv13Z+CCJOw
YQY3N1VHNsmdKTq1B8KR0eVUdWLyZn4lCpJxJfNncJae2SFacXQoVS92f8732nKB
ZbWOImpdz0Me+62AYQUo9b/y0Xe3CEhXLeC5brLujP4AFEi97ISX3+lHb30yfL+u
yZnbALAFbCLiCyMLVG7Yd9tv4OnliByhWh/YNeDmXYEppndhDuGw6l2KKuSRO26p
EjyjpGBUNhjHeodhuh6HH2EyF190fV4TlZpnYK6FIkEPwc6WtBBctYKxy/C8SLxy
i+mZGk4d91HpW/HFm4paTuKtKqe5fBLslbz7Ocf44YFGGrXVRS+K6PpLpQOYxwzk
3Vz0cTGIe4+PNcGnMMJUUKUWtvB82Taa7bbSdTHo9/24gYRQo76R7UNHq+IRyWtF
CLx1TzagIHyIPhvx2iz6cY3ErxhICostvCrzf9iW+XNDZ9T9hlJ+PyWXjurXYjsi
pc/Q3pxXHGqNAIyD8YbZGt19qCE6AFCuOArZXANi9EmcRQdt8P1CbAc3pjLdHfe4
EbNJQ16p2R5PRnt/5j2GyQwEFE8kihlyJV7s7DKRlb4/yeZn9ctOIWOG+mxmZaID
4i2zazqs1YKvmbWam76vyyl6J8L9XlJngjfkO2PGZCJQGElKfaRYpv6UXMjyrCC8
Bwp91qsIMtCDZs7uha9SPnvJAIIUvBmyubv0EKZUk3zcnyK6CbWoldC2kQddpNh2
M2JKVo23tZBtLZM30qTsPmehUYCXY+IJqCrT2Y84cpt+90I0LcuC3QeawqlkQPFz
mZ2LQgh0o8gtuX1Ibj/2Da9MgHGGfVO2MYgpNtWOdcriv76A7AyrJ9CT2CHyK6VR
/nwJ1lcMvhdU2lWcjwa3v3nDBE7/OSxrlDZvAMb1Fj8R8ygL/TG32ailPNfLs6Dv
wpakQTAasJX6w5HP2XUbnCoUIGkGMpM+qL1tHvnrszHDkkT3fvizl7vrJLn0jT/A
3yxiMG5duU0hW2EDaLTsLvcj2Ut0OiCMezRrKyeQONzwXz1ehS9qYm4S9r86uoHJ
KTfm6GdKrDldBdt2oVNLCZcj4nr5Z3z3s50ZIcVFRh/SmxoHFumqyYOUtLW8vSCB
pN0Hn3H6VwGLeybdmpSzbHobw5z6M0+5FQbC3esBfNQthqpYWBR+z5u+BdcQzREX
THTIY/6QC8TVnIQXSktkXkvZai7/Q4rX+E3yyYNXRAb9QTO/hw/NaFqiGZEV62AO
B08poU+ozPy8C0HN3KEqB4AFt54twKPG76KbqSJBGhvrI48t3GKXskk/6zH0vqWo
MBzK9bTlWEicroSWvSP+xsqgufL6FBe3P6lcXtFTWhK8i2AxUPvLFNO/It/2M298
zADP4YRjjdxmdyYHdLVfQt2nv5xoriynFb+KRRgFJptjeJnd9Mf+pM73CJlHuPUi
O1yoSE4IcZpjzzixrFFxdD209BkNo4g6uarygDthmPNAh0dOOFOjkPK2j+raQNuy
NuvNzUNLXyeKNRL+T9086RdhOqUSH5yAh8forO1n9ekLivErOwITMkShljG4KyxZ
2PqVTYUUf0YxICQK/4fqLxEHq9m0UFraVZ1ZeQzsV4F9BepskO5s8/vNTVmAv9by
Vu3vzV0ETPIs2rey7D4+M91ru3T7/WvkR+BVGND6jGZMsZrVV6CrEYeCD2FZAK4z
h6p0zO4e6PGLYsHPFlQz3uo/DiVj9k2aM4K848RfnCFWyJR3IS2tbZyOYHBjcTCK
YqBLa1LepzXSSdT0myIRF4F2H4Iv128QpPVSHp+SsM5s36pFMnXeGhyCHwMkBzCW
6YkaqQEr0ir4WXDnNJAd1pBuQqUqhtOTH6vU+k8S/6Zg+8xzuJb978VAYNrVzyTu
5excr8wGqW8vzTvBoYvhdvdobL6IORn9ORaeDGGdOVJrfZr/IkfPfCiCYpMEPa8f
nW66ZZ31dNLzvXd7wtBa0pCyJIG6h+GIDhfkWA29A8Uus4uFIZFT+cy6jk76qNH2
RAUKMhDEu4os+H1101cl61sDLs3mJTgQa3PBeN5V7tC5gfKPLKbBTC9PSbvXWgGy
AQrauhrXrJfq+iljzAWUDH+g47HlxE4AWVl2AkprSAUfZEIvscbAP+g97xued+t5
iqBZf0wuJImwVnW8olTurd1ykrAQdEBl+C01/XtU+wp226+sWPSIL/YYZahkkK86
oCjNLqZgiYIZFvQr8tqoUEveIb9NMvjqj/XRuepfu80N0jejV67Aurhxlz6iTTn2
WTTGhC4cquRTNs3IgT6aZLt8uvD9tGla1fENQjHJsFCFX/vYr4ESsXA+Nj/exjFu
r1arX4lDK9BcyppSsDONz/AgneL08QwkVagP6Ts68Ku9hhps0OHm2dsFzHuFu388
5PZHQtqFELB1wmsUbOmcRKYl7bhnUG1iOVEAa4D0/E5+wy6Ek/elgXZrzt8GzSjT
zZqp/F4kIvhZKRsmi4E+5rrqVjk5hSMywGXv8D8Kf70F37k4mOunVHcjap3iaACl
mcIuDe1X+t+h1CfoUAuhCY0jpVlMfip3VyBm2m9jLMDNJ942D3fQPiuj6whXhJol
yWN25z32wGCBC9er7wa7BrmnfF3vyPnMDsgrcb0UJ562o/97onqe5IJ6B2mWakh/
5CZ7SFUte2DSraLWYdAUF59eWpL7arm/hn9pHqagtRj4reLt2I0ex71NzgJa8puz
oivZKKcuZc3DEfbOaDmhqT1Y3EXQkx2O2NNmQb5cSCbG+ndkCVHhBez5z9NKfz/b
YUbsVxPGaEt4y0RxgD4Ljdy42HriyRc6xJ6onIn8DlT5qz2KSVIXLAyuhRJAp5i4
BUhR1o5TEndR2ozz+CD/etdx9sOuU0ru63LoXDHcofZmiV4kNhSqF4qs5YjB4VPy
hVkyy1Y9zsFX42HEJHO4oIdJ7Lm0Li0X7a8zqM7sZwLMvimY67Vwtg5sQxtUvo5a
7S0nNZWqk5Dkvrz/Gg5JLg/6Rk6DV9do8DR4uyWSuvaaRB4rV+rHhV1E6o16WCXu
jU7YLNnRdvBvaLLbySMe5cHfVizk0ExXGIrmqkSWO1DwuiEP3Gu+fLlwP7huZREc
r/811zj7QbUbRlttDjo/QXICbfplw7Xt3jHW4MhylauGPUb1bWLUbLQJVJx2c7LQ
/ju0XLu3Alu0yM9+U0JhOzkaCL41pX5Xhsb2rY0bZby4a1NXI/O+sxTt0Dvp1wMG
rmsFbYdIufw/MmAPy308Cmj90azgZft+60WWso7+nUtfnyv5+2HQshglBMWUdllO
MXbu+Qauteafyqh0yWnAKL01ckyChPmeUbvjnVcFLQFthdhAzYR4ZbsvdWjn5lby
Lx0wcuaJEn2vV9/iSiz1A6M+PvtQl7wYTLO2GXr1iFFppKwiNUB8+hSEcbfpi77S
GUarAPZn1l+7wGcz+939czsGXcLQFZVf+nukHdG75uQ7zB5nxcFME4hzy8VdjrhH
vvHUD1zRziVISIHC3YgdpwfjfIsNY7tSjq+zNVQGBMQQVxUwzFv6OfgdFg+Ci1NO
uLL8MN5InaAmJjqkhsREKwhuGiXdMUua5rzTBAhsBUxxOU+vh09qRvEpDkWFWrBV
jMZFR1mUZql1CZpalM/xnWsl0NT2DmLlBjl7kAHq2YfJdJg/2bptmtvqlNDj4KeO
8Bx6zVKqra9P2KK9lBlRU4QZp7s5KfnKgzYuCi7bPkV6HTkld2d2Ng7MO/5qx9Fb
bTBNtyIMViYZn3mMoIVL9srMMmCXaZM7OH+UdQuVqHuRYIz5tUpV8ixbgkZA2Igg
TNd9GMTzZbODzxC+3IE7C8kkNw6NRNEXCMDUAM7fwkhjo8AMHRG1BHPZ0FoBSqS+
uXEUw5fju6poplLIHrfQjy2TdkYTChaZrcTEakECeWgXVZ91fF5uQ96edh5yE4di
JxMAHjOnBh1BKwdhJggeEilOI8iPe9jim4D4+ix540FXENKxQvNLtOCU18nNrBuY
jEvi7ic0LOUznhUtvvaRe5LVHYwUzEZ66G2UCMtziM+qlek7UGAfdSILzeqwX0z0
LP0JLyfNthYNkemI8Wx1jWUmSb9sFN59HjkPSCuwVbrhoxweueTXcxKY/8jV6TAl
5IjdJROTbMV/CjWBxiCwbQBcp8rwyvGEjhpmJfbgzM2kgORwEr6yOfrb6F5kfOEN
cxOkWDQQzYOTrIQKPGP7YpDCEJAzVY8WQiCgWJbNHe5pAVt5aR1TBTngcca88wBZ
jrviqfwLTRvBT0L5a+B93d3ViTO0xOr1JOqXCTkDLJYFxLjsR4YuDGwpbGCUCfQB
Z+uqSbfr2Pk9aqDvfBq61SlNHsQv+ScXCH6qp3dJsYBNlyP0QglfvSIh41kPoDTk
HceKmtZJ5jthhrbTPDjouKk/uwM0SnSI2zfTqEAAMM4JGivyapvKg3xpHzYPGygC
w57WGvuAxEdo/Ic/54tl89TjIMjogVU25w7Ga/rOgYgPkYw9x1J7eIvQb9Gv5yEB
QiLPJcILFjGlI8Y5+Lz+SZFMBnJBYW/YH7XfOor5VdsVhJUK3qHXJwjwoex3uez1
z2k+ObgGq2+Bhdqmr6/lOq26U4B6K8JCsCHGli1NEQvhOTtX9sUCm+DE34atOyXA
/HPCFMyKhuIrgGEC1f6ELugEIA4DaPxip1w7cSFNFyAzWzzOSVzj5xlHOplQ/4bj
D2CRwmfTYXuTqZAR7Wx4fU4gz+C95gzUFDUmiQSepIdtSqRLS3KWpTXP0sW3CRcI
IiyD97kNUmWJidKMUjaV9YoZ+m5InfKwvDElgqhtBYrRnf25ckgFIPr2QGYjOLOP
byS9IKWvjmQN0vletYvkOuJ+o+FasIalnhNtB0h7zliB9CRxKX/4qzuFCx9fo5cN
xnAH/3uekHe9g4oD0NcsSya9Ugezs2ZtW/9PdyjTAIivrmUXCZVxgio2i0c/LIOu
PuWOGBkzOftl7VdHOhxvuBPU+59JiSN/z5SYORRFu11xdrxjPPX1+xzzU0RkCfAb
QFINNUVThoDkZgQJ9guQvzdC0uIaZGuG6jcOzvWUaJZpUoJDcopawpjpekjwsXx0
pDIHsIeZzXT4SsoszR0+cyiiIkCONNItMekZ8tG/MueC+yca5kKaO6BzJK5We0Io
PHec1tRBv4aVRR9Q89XgaA==
`pragma protect end_protected
