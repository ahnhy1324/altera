// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
T9u5Mnc/FAxHQsF9nggJsKTLduVdbFFrouTGIpRa1vGbL8+gewsNAHAT7BzWUqdrWpi+9rQjL0TA
xBYzKOUmWw+uA45yNS10kxcmSGFhLX7he4q+3nabdWZ8P0oIDFIOKEl0DxyCPw0usUOzgjFCdcuQ
x1Vo0azLHk7APwOIBPPpl8hOppjBkA1latEJzP16FZA0UVfe6YClEPNRQhrjWcEa5iv1TmbjzX/B
Ya859i1b5ftqn23gPFoV+5tcQfVwpBRzYwp1uiWlY6P8pHMA0ZDgQGzitmOwUuqdOhtd8VIhjwBx
tzZNLM7w5lKsjKQ7umvSeYh2/WC3ZdRjaK6ImA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
I9LeCOhZDLA4ieY8Y/M4nBicuAbfXjN0rwocb25+pw7D33d/XgDIu/qs3OYKf2oZAXz5V7FOBrXz
1U6H9DQW3krS2zr6Pf1dg00/OSMLPrDVgegEmuIbuCiCgxSntZDUH3Igtl/8tr6ZM5UmuAUmbst3
IgonuZRCuhCh/0wGk27xU1Tv7+X7JAhfFIYkoEru7Uzf4yN85MvQHnJeik74Ow8mZ6UjaYaKPyVe
GBS7C0RkOidH219Y8Hn4Y1e7Fc26m9yK2hfoWxkBDbOgPOrWTgMU1WFL6FbE/EtDWFXCguPFLPLM
6AVQvmQRlbZ1lou+SPcIcMqOPxg6bcYFe/vueE+eLmTbX6T0Wwdw7Mobh5Hq6aDuUOwqC+/4smzX
vPXn5h+RNR+pFN/mH4oLm/VJZopUleniruPfaCMfsi/Z4fDFVNc2aTNmpG2OYRhSKlfHlzz0wIM3
WTHSC52owSpV3WdNcGipDjXTYVksWOTpcwa/zjJIOXg4pdsoxrr1ueSBZhUU8K/SzuYpDJ1SfaYU
k1XIixSIzTABrMwA2hSTAxFivj8AwHPtGzsURGq/Jx2RUGtiySPujsN/E0mfzRXgUe9n0iCR0PbJ
C0YXVDrq3O/haxN/jywwqH7vAaNGN7y57Egev0VjELvOhqIk4KPQQ+bSDqL3Qbe1rl4wYV776R2G
D0AhJqIBK1PtF/CB+bvi9FzzVsIyTCrSq/2h4BAiCTVH8z2Fp0F2Gs7gCVcg19MWbGQCXf5bXRPF
P6cMAlho7FcA4fafvTKWGf+mbm4R8QfD4RSqehMdI7XlrEQtQIzoy17FRk/3caF6k5BqaFu+bgwk
LZqbFSsT/Djp0wPQiXCCTR8v/ok1Di7PD8/gPuqVOkC393dxDgrawjC6WwY/lV4Bz/mxER4zN+em
rLqjG9+qxy4xp0cEdv6uVeU3EjnailPQtB0XBKlc65alp1fXen/YoAfCtYC1D1bvP8jLZnZERShy
oe0BECJarCBPuKhNa1VwlS2UgTCGq4SV/cxbTQiiCgWyaO4pV3c1DY8k1SAWIgyjmG8Dw5Rbyx16
+dTVPnrgK3Uq8B4F/phxFMZ0O0nWVCRXevtpLtAVQPyR1+uZZnixQ5oO5cKnheu11uITktBaZlHX
6bz0ieizZwwjTSg2XyxDISC71K4K2krWPhmtm6Q8RrqZBv3ZG7YJFs6ftievoOZIwBdktlFfXuDW
G6g6w71FrfZfF3RJAEwdSmu+8n47qX1MLCK+LCoIwCA8H3SjLF3x6/c13Hx92I/TIoyD126jeF88
a13edEAp2o/b9nunlRdy5u1/+Jc1hx7Gow6eqd8Cny9SpL5eXiSjEaUE54LzZeEY4Qw73yEnoxy0
p1vRz+cDeXMhmvQr3wIDBWWhKZyfRrR+wC1oGu8xTafCh63i0yj9vSsffZzIpnLBPN1lfu/dDkTd
G7+rFgbm5jMGleRR/uqS9a3fi12YHhrHFD7+NjC4JnWB0VEo8e7yiOTxwkcv3kkQavadua7QLcDK
tel/oT3aBptj2sO/+HIOMnQCpsnjgQeYSFTA4CnqUcoQCbyKBwpcdpUOmKMiV3iTCb5FzZ/lFDCL
nualP3ufd5wJWwhwyo5CwKndKK4eZfiUSl0exGlPXvXw0d7t1/4eaC8T1049xVZl0+8twA50b2Kz
zbtVJMzi0EFcpcdSiru+FNas0oajy6zNIICbDZSqb8vreF+RTTxOEZZcinaNhGoEAsMeA+xZC2ed
CDwieBeqC2dymLiih2TItN6lt/XnfgxA1UyY+Yzn1ZXlVbmFdlbbyUggytgSlT10CTzL0AQVCDcd
ljwEANWDFug8aCKis07Zz/pNkvm6I/PBDxbO1wOpU1wKuCeXa6SM5QA3lXrgEHYuHWxwmFL4LFLo
9u5RuxQCjj7qCaGaNleJUMQkASZpoKWkx+KgYIb5gWSDU2TUnOxFdEdbgKeLYLyHvDR0GGiCxshF
E/znBv3LiHkmmFPBdRdVNxJ07M2TFmsglBAD+QyciVtr2Ed+APrdIU7vtrJ4rZz6LoRxSlgXTKJT
6f5aTW7yHimlghHo7VhM1PdgHeC/+4MBGr4ey8HNeH9acAEQoZlujUHOzvftrjz0AIiGDhKAJ/Pq
TE6EjUMEzyrynaNq8qoVA6RpyiD0RRI9NZSxhIhhu6weFagIFS2yPyp66kTFTRJFKp+ptfoKwk0O
+99N4N7jEiszD1ROz+rbKZzuq3cwpLCmoELaUOjX2qD20UldFea4dIY6D5q75W+uT1+vPa1aOpT5
ZFKzraGmxgrw1RF8FoFblUtJLiPufG4t4lMQGf7ldgkXVIlhKz3YsNMUWgjHToZj6PKkmXd7kexx
uEvaTlMfUOKOGxodqZUEL1wlIKELfqBtnNckVWN+Znu7LK31itr9+QT0QmPV4KJ7FVVwAPciNNwy
9VUwAEXpDifA19Vf/M66Q0kBPeP3D8LiqI4/naGbq5+ON6mbEUIErH/Nl/qf0Hfubt8rqyaGzn2u
DlnHKAYtO7mM1Kr8U+of+XtcPMN5LWPJjMVXBJ2ua1N6KSsAHg6Dh5TrjPIPy9FvMGn/HVsAT84E
/nXSDvn/ORhdfGMhbcEuUQssMohtMRGN9/VApATbuCznE+uHVdd4LTJ/NZtajlnEGC6zEu7/J0+i
52jflb9FBoz6e+C1vYvKOFSGEwPb8j+7BCQB3dlrWNpm698Lpv030MyX3+/cTjXPYxgsL+Cd+JzG
NSLmb4GHNX1s5+zhojgfvhV1mCf8WpfUyqtUFVeZiX3m9GUXxNaQfb99/FBxGIOTbLAOVpq4JpRW
juPsaj3OppXoS/mTaX1FP5mynlo0DXuPU6AutFmC1ahPXDySfdM+PW/xcQVmI0jK6DuK2NESEfFe
wJvWA+mTxk/503L1/UztjVwiLWZWw7iVX8kZ9p/v3NcWYGYWy4GuXjFPoCvwc5iOyEy3uhRNWSPS
ChRvGqJgXr4EqXbC99+7npqtvpHEX/n0uDbIl6gVQaO2MrdhUVwNfkYjAdYhESCUJWNwH8aU9xUB
c3Hl0bS2FBII3/IE/Pl7FJgPpw4dlj2wzixbIMaY++hBrpvKrvmieZsKKBojAYRv7kjpcIyCKkMN
tdjIoFi/WrtoXjdILddhSeE/cUO220C59lavCikr1k7F47TuukzuAM+jrFtJCMLcSmV8/m0aPFQU
0rFainA974uRzm8XMHws3AcL1jxgOjvLpgv09OAQUeV7nO3Quj3B+UKImczZDaL0veflErt1zCf0
pLEf0akrkBacRBqSL6pRTyV/TCJ3kwj0vZvEVRy2c/o+UwNegKwvP4LVEEKF5JlNHnBI1+ml8ide
EfMtVbmDJsEtthHdmFqq0quwkeySMXRDj7a0MQgssp1uO/J1RUETekhnuRFS/M6A1bdSif0VMlBH
Y6KSlaZL70avTpPHVFNmiScGjQTrjEid8kfVWYtQLzzrSiYVxBPsJrEGT+ipeWgJbhzko3/9rdgU
uKGf9ucv+CcFrE4P9tDAjZEwKvZwku9Ol36ZsrNp4hugGjzBl8an0pOXTb7xki0nSp7YzcSNg3a/
J3il2A/WHek4xfRAxL5wr+bNi7hrQJHa4Jm2pqC6mXTSreTKYmDZZKEdphaNwHh8ImbSceWFNyzh
PC6uRD4ogDDDob788AI3OYAl9Lz3w0aNPYpGpNlIjqDBwlAaupldTBJGaroGMqDj4+R0yitgvn2R
LEK5cV+mlOpdkm/FK6u662C5HGnlr50u36Y9An+8Gzz2yUdMJO5nvMrTM8piurNtjbxj3zWZtP2k
0t0IhbtJBUEKLTqcTrV7XehXdwzzohMCu4Y7teN/xKKgnZFHyXsRZccOS+KTVvqkUsqusJP1rxgM
nP0XfQZBId51ZCL+4TTvozrZbuC5The4O8U97w/VhvwwDVVNiiiQM2OrP1pS2Mbssva0nawqYmeO
G9o4v0Lr68wKuaLdhzWqEIfgbz898Q2wNWNsE9MuY1KrwozA5qb9gKcvQBtSE7SWL/N0a0lJe1py
z8GRBfobP6W1z/zKp5FeOEdu92+XWdSO0wDGVX16Q2K140lxpqzBg++J0+0Dp7qcq2+UY8Aj05lA
f4hWZmpwYAXKCgomX7KOXf+fMeLHATXGg2wQsU+qbOyY4KrTI6Q79GArks7SRyFw1e2Cg6vcJ3qi
pimMoO4m617pZihygERs8UT6OcZARxSNP9ii4/pC/S+XWtTa6QUG87659g53LvjXkjI71Yzq6RvM
RjmcNe84MHfRfTgHK3iz/Z+ZNFoUql2+Af8KsgEXFCMbAguIWFCZoK/5+Ya40ZwcuutuAvBI0ZsX
iSkgp7wWm0N8feqAGi4JL8BMkbpbvC3pYusSmpMlWxnX3eTO5ypTJHFJYwtzGHKtj07ZhLI+aFy9
vRN6rbE3LBllXU4CbDV9Z1CxPvARWCmEeY39ezsJnCeasMIgIM6qHnMjbyAmp0BbjuHt8tmk33Dt
p8vKYEtMu0kGR2vSQZyikyYcXAuGd1R7UjgRUlSetAcW6RHXh3ZD3SKMM0czbPfxgU9skeyuhKu5
4inPtMd6GvYf2sfavxjf03aEQEPaszz/YbBPBB7nqui8oYwTYJEUoTXRrk56dIpRPkOOAyxBquVm
T+4LaNYu+REB08Ouoa2gCL7cUmn4l5Tq+BVlJYUmLiDhsQHNjlBmkJPgCteXIZnEJgf70MAZ0tcm
uHux+leh04ti9FWLM6cWk+MxOztTYePskXzkkXO8n0MLvvBqvDJNBpOBtCLM7lb+YTqA/HipwW6j
Rr2NF0uByYz5RJYoTYUpSixPCKqxh1NdBk5/w6c+LIHbwL2DsDsXG1ic37WnHm+iMpJ/ACsU1xiM
y93QOEBA1Pc7RCOLMkoNIjVkbma7ZqFA7mhnQigACCBxa9C+Q3fG3YAYokKCrrlge+XWRLJnnAFa
eadHyqDp5KyZIoxsJ0WfKbMPF2uzK8guMI1n7zjDPDE5B4ofprWPPWCoOHUyRAwqcUSde02CX5Sh
983+FyQ96+/j1lLhCwDolhRMY0QeR/6RiED8983EfwkKlonxBEjG15j9C3toVH310yWCxQy46VUr
ETiCNrT7wBa4IH11MDo8QByHeIrYqnuWsiffom8lmfYXR2vyxOLeGoxJwiUczRTYXx4JADEjQM6T
47cBv8xjzGUYrwv/Wo3qni8RDqxRSHFsOQ7ZnQ/eB7bd0CE6xZDLO3pwhomo5aOhP6TJMTQL6gYE
rtLl4LezHKGJCrOnYM1zdRiVKMRWNWnj8alTUc8iuSg/eWXNdqbX5yaA2UazdZpXb3WSyWsiGUTi
Pv6DvTvR6SmaSvPGMNysC6c5wGpctkA0fzd23afwGzM8BcaPIgmUbwy9IsZw789vXKwURotl+f1S
66Rrnr9BVv95XYMzdbV21VTwj1+8bBfG7RiiGf6c4CuO7mqGnpT6/QfUIlTIumfeTFMqPM0G9RqH
HtgfVf2m8wJtBx8zUVADIskEzdyKVUW7JgD0LPAsixkVfshvFym41ibZ8YoTv2lai7Ga+aw3FLkS
btBOa30Xc3EhJJW8xcFxqZAeGmb6YeE0c5HlVaIwxtmosBBAv+/6+vo/bDRA/mpXT9fN5iwsYpeM
RuQ/t2wT1UyTbbSi88imTuUnKtK7EHw8bMzU0Puj1Ag861JVfCSYRZTTBQ/YG2RkRlZSwSFzF9rM
rQspOHjA1Un5zr+j5QGRItD4J7imLGz1O60ADp67iK4FjoHegm4ZKRVga4W8+O3P1Gc4ZDGyHEke
D6nH64HjNtKXyGPtbGusHkqrr6LOX/3vqmuCvJeQfDanukAlgbyxxcgVKylEcfAz6u9MQuvbnaIa
sY3KIjjv9ZRzSKqaAq9DFOttuI7861Usc9FpMwawe2vFJii751JKlJDeBHVuj50tyZMyxxOtOlXx
rLQvL4HqzDXKf8Ip1C8tR1obs31zvXZa3HLF3sxt9IyHqBxRzzqcFO9zRC2puaGV6ysb6HhNH6j+
Uy9fxosKgunz+CblbLHCE/u8TwUM6fYTUnizS+ryRDmatxGlon3sSeFcDOoluZ3yBoIv3m54ic8V
G7gBGYPgeeIu3NqyMXQ9fRs2N0XQ+odbUllo1Fbelwxz+dXSwAYADla1+Fd7bP14l9J6aqJ4E9dZ
CL46uqwN1wkzrO3RzmVjV0dR+5Rs56/OTne1mjCIc/4Zjga4HVddAJgYHztFDpoyfXt5KB/i1mam
CACEEB5DVgfiCQBR9VaviAzh3AlOcjzm8jp/Bx/skQ2k9LosrzdVMelmdxjq3HrqzWeU8CpRX087
MjpdfBCyTH3OGfmfNzl8Cb9F6X2H0zs7C9lqdwNY7WkZLoU50ke94/PbmHlnuvvyeDbjNzdWniMF
6aAu6bXfZMkM7Li3ATOz7pqDZC3TqI2119XehLSKd2djaer9AighNGc3as2+1qkNh6/saNCKxFzf
ZQEALT8YXG/2bgzfDRwnKRjFQRnSlJHYhcbrOEToGwR7ZaxeChpFcu7aD1xogNklT1+GV2m8juhO
qAF2IaAevSfAo55moDSWBkBRgVBSDLJ4P23GVMZI7MV8/4IftX0HR2x7DAOZPyoKZbRwJTtXgH2/
6/dDCYrRhi+9QFJKYMm50US5D2bnO5XNkcvBA5UTDW5F3HDpNXeLze/crwKeBCyKAmWo3mp/PaY4
sek6ajkKTQma29o+PGYeh+i/Man1Ub4OZS4Ow0sFFjluHoStJCZHhJgbLkU7YZk1003WttZ762nV
SUxjJXmbIay2C5Lo7dmtVKJRnhGTkdRZHPVmxLwcTlag8cuMFC0Nxj1aDF25aeuJ++HiMnJFmKhF
JkkMcSzEpsiYRaW/SCYJvNf9TYrUCONH+3+aLPUsNCvdEbfsFceUqrrFp+hCi9EW1IALVNR4thmU
Mg1XH8pfS5D0uTF8WB4Nk0HPaD1h1RpPVyHyVJSEPqy6LWm+ISqXipSz1Ron7tWx7t94v2FO9iAN
CYCyuUB+dKBmxkKvzLuQMu7z+BTUhIFDqbP57dyzioamuA8/JS0rMVDWypTJW/JKRhAcVAmiJOMH
mdbjYTaJnMLtdkszdLUabwH/vWZj9+HLNBiffEn40GuMff9Oa5PIk90TRbHIhwTCj9rMDRaDuDeW
kIKGVEP2vcssGbv451fAnlp2LOmdAFm7V1ZiJVTjDpwiKWnKQ2Oto5HLm/MF2gwApkC2lQj4rlFQ
gvXj4+fGG1KfucQ1ocbNalBBgVYbRIyTwJdLfqSMnqf8aKv1yzKkZgxjmlBcooCJ7kapwRuVRCGS
qqKVE0U+92NLdrGAy/FCI5i00Wed8ur6Znkxw0TTXFqcEZyhz3XM9YVB2ak9D4NC8IjNQMXhQuW4
Ldr8bmc8R3kVcNKFtR6upkpwBZoQ9ZWcCv/C9C179HsylSRzdhoeNjr+qlEhdg1DiZ+FI/RtHKvN
aHbKbOXhWfew8VEpmhD3XkegVTz6qkj+ICF5PYEQJdeWaMYB9yuk/ulFatn2efx0ky+GWGmnNB5o
Z6VcjX9uTRe0tokgwd1wjh/tWjdtPJgsX5WOKlmLoLPP5swECmP+DkwMpdDzPxB3+vW6uptrcDkw
2qfGhOtSa5D2Tug7q7L7ZGiX8aOukQ+sOCDcRPOMgExHicwAWWleVP7NuQSZG4cpy6Bs2jOnCAZh
1b1oHIstvNW3oiPgYIj4D6GfL1/u/mbAYeB1krmNZiZffI29kUKy/S26nPCkeW5WF+CEbIJIwCkt
4FA2b+TW5yHsg2ByuwX/RKBCLsDUoH0/Y8jcvIp3shmZYaJp/SguIwdMQT3tWRdOqcXPE/RUps04
P8AYeHjY67WJQ/zmGiuiwVpsCzgpiAG77AmjBSd7hbVD5RdbWXcbmxwkPxLn+wJW+FmY1Yh2tz6P
jmWk/n+n4tvo1ruf2zxI0BfY9LV6HyPN3LRmTDVn/1ykag1rcNlG08bc7fpY4eU3dViXfCTdUmj8
QlpU6PLU2Fyhd+BDe0TdJHcVeyXxC8SAiHHVyuR0c1iL84fGu5WP28JXT1mJbudZLlOhXopQ0Rpb
sXp/O+HoB41SbU58hLE16OHWN9Qsuid/KPDPc6UIbBifBzrRchR9/DpJhdZy1Ejv0Mm7D9a4C5m4
C6NkgVfNIQrnUmCoxF/MUfpm/RPl6TScx+E9JaCfmGSKCQ1Bz8QQQtyjwRKj1Q1lRqS5XEODCYND
ktNjI/gXZT+6rnLQlQMQqHGutA49IgFKqZXJCxFDeLEMQfvotmSs+PJrjbkad0moapqpaDHlQK7b
Rv2eZduShaNlyTaCPLHb2EicE+gX6tZGlXNKJsA4Jd//uSSni8m9W91Z9kaJc9cqwZPBVRQSlCk3
MJwGZpmBBLjBv0szVhQ4n5HRb1NaykrwT+HrVwEn2yNWAJIlfQzQYP/svWIFdhKp/cHAbPSFrdH7
MvWbIhsA+r5yaD5nenJLg4c1WkVg/B0W5nNuALmP+i0mz/rrSZ9p6OpGF8R9ISyhKdYH/dqesJeS
AI9AOd56zFYDtfifJ3zF2A0hpg/Iy11j24UGL8v4o8TbhUuYhs+X8K+SLrzZhgDK+y6Uz+/KjvBy
I4GAnLXR+G+MwQWNLyRLsGQ5CgEwc9LBw+pKdz46Hc8QyLoXzYLCfchA0192N9o3LF6TT3ytNUZl
2HeGEIuZ4Z77H6BhrcrgSb5IoQMi39a90iEkoNtxjFj6X1fDsZhQM/aRq/Gp170jhby5bCC6mcKu
8LOpSrwmHHb7tPbGwg9anLBZDU6JszBeU8oJyreGOVgwoCyj57nesZZlkfiDRF6DWGu5AJhDzIPJ
l2djRwshU48VdKcg3Y435D+CQaVMwgXAM/DCVS6dqw4UbrEAOJPuQUqbU8ed22x7IysT3fjUnBV0
6RxJ/4Y4YyB0rmIZDV3L0/p4DWCXmD6YdcmpxA45DlHxOScPWNI/rp3WSRLlsFf9ZoOLsrg2E05r
xbazHlVR7SJ24xXzDFwJxFAuis6m7VnfNA6kGoUkKY5qXlfdjBGXdmiSQBZoxeUOQyuBOhnEQoct
Dl8BcGKhGIBkkgyeqRz8I199KwO+z6lbXexmvv6iDqff+i64ewHb1WPgZ+7USsrw2GT9QxfnCvJq
yebFNVQs/2oyJ9KyqdkC1wH+f7eZ/MA5DNFaOJ0n+wi0aFpS0g1tkNdkErOXQOmehGt7PYWb5dUn
n9HWzHjSDPTjjau/Z8gRzR1iQL/XtW5NtLs3R+NC+OVq3b3M6tVNplExM03M7Z3iSqHosZCPDK65
CSTje2irlE49RPgEM075PqraCmdUlZOxWYifLHKYuNsTgKJA4542ezvGrDL1n96XC//sI46SnMrS
5rxtDK9fbldo8yPXVhAXe7AQVzUtWvHTmFMkGLf5F8D3+9YPeR7/Gu+dUSE9wzyV45hq81RZL9j1
bW4qmIVS+Bag4gCq394ulNGJsJhbRmAQQz4FXGibWiFJ7jzsG+GcHCMgv/t29MNSAIAWJWlY88g7
ZbJ6Z6khVa6oAtXtQAIfR7hslyA7yPZdODsSpF/A6DCuwbYvbcPWQKnLlA+cj5pS9R7aV9WpGy+0
dMsGBQv98dg7Napw5soaAmZ8jOrY4n79AdwSDKCYOMfn34V1R/m0wBL1I4xn4W5lH8XlvpfFUwGw
Em2nhe8aFijK9xSpl4xpqBonFEfWLZyhLGbahxCXc4amFT12PggH7xcpY6khxbMnC/fSt4RZdP5A
hvp27jfKvDPnlWh9JfL0DMzeIaWfkPy/xEr7AOadGFLODspfIzIk0jJaZJ4RRKRU9B8IyHku8wIW
hn4BQuEIKfAhFbIbthUurfwpv/JCbFNzhkSBr9y2xIk8ZZWA+4gQRNBgfopGYelq3K8qrHrBk+Il
zfYk1zAfSd3oHCDkM2XQxbXNYRoiOxRTBiVzLbosWWGsxy+AkmKEXa2ybuM1To9vImRPZvrqECEr
OeiJSLraHYaF+7YnY9PuquJw/j2WnFuNERNTXxIBMhgdnudgFzleORt1hKkXt0lbhinm3Kum59HE
nvJ+EMKLxHr/fOrp96mVM9B6h1bLIiQvRwLalo2ekGYmy6DASWzKWUzNfaZtQSkQh/+cJQj+G2HX
No4NJ/K63eciyqrnMFOEvDgUyHwtfdF7kRJWg+z9xWY4hTlad+TL4LJlrUfZ3I4BTxecBaPr8ruO
DWpfKAV2c8R0CkJriZVnZ8e0f56RmgYm8+w=
`pragma protect end_protected
