// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Z2Jkpb+UN6w/NUGtS+lKcjcf6XpibzOQ3BOnG3WCqsPOJVD7UCFJrFT4YSi39d4Y
fJeyG5vi8tdWpZtVSO4wRjx0x2iGShBKL0xdDtPfTzTvkV85Oss/t/s5H62dzYG7
sR06ObCrQmatU7qGL8aVC3PI7+3/ZVFfIDzbPhEAGdM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 63088)
7XGLDOvXium7Ik7XbZL/MLq//ExtjHsSkW2Tp0nokyTgk6+ZxSPuSMrKqtKGDY0z
Ri83RsOgeiJsGY8Eio+DWN6NDtXFeH4c7gvoVJpOa1VcwKZnqghP6AtOTSLK0WGR
Nc9/9P+GeHBRDpMkS+LjfxoPGDca2nb1GFK5zlIBzirtDrE9jc0PqWgGbekPx7jH
HhWMpjIcLO4B4IiVPLdKIHMWXRV9T2mD6whsBZ76EvWqpdBonkHAH+UYnVLkYt8J
y5jP3CFdWUhZptlCryWsuTgRVc7/qX1ztM72MeTn+MJ1a8WlFLE+1N51SEkyCvHU
0avmyLymn+WyLA60aJ/V+HbGRJoQkSKHLY/JyCnApom4XB129M8/jIOxrc3K6UAo
JbdDHonOaVt7mJxu1Pc93WZoqt0ELz+qV4ew08OIkDgWdT6zXO6k1x+bvRk8MEAU
PUN88Eh8zg/gp7YXi1854WOTMBNp7EnUh5ez74y2Et5qkvp5LM1TyWDUGrNif9u6
IG+npTe46vFv4NcDVz4nIFrJ7WRwJGPky0rjxcSfICAccNDUUzSEqQe+cbhSUw1c
jzlChUPqtdVaJRiyZvt2qzhNEEq3KgIMJMFNCwQfzft1kdLzAYptIJOz9q6Xu0oA
gfIlMw/I2PoIuuxK9RPdVEvQWsnuIecmbZmdMP1QBPO4+x2/65UaxlRQS5mK0B4L
nZ+ThG3DdXHeMeJ2QO29iyFAELMx8TOQ/2lpqfm8q+4TSUMZkv9GMR2bYlDX/LrL
o5fr46zEO2teKwFVcd5cCUfycZ6RgTNDuTRl2bMK7TlJiHbWzwbOJqiubXfN4gxj
2s/cNGbc1KfxsmY2U2Zch9Xad1TtlXhYvQy2w5xN1PUPQYcpuHCgDuRbwMZR4Vvh
0Dtn6Bye7UMLrk5SpPVQIXdgO4k8Bl+Cah2G+U5YX7S9iYw1a0+c5JH5L/FcsT4M
8T67iKq5C28hq8fL3xuUMhohhCWdUJ1BgKtJmAWlWKMKyfBOwrQYrwdVR245T95I
lhPmHM9gv6+18JdJVNqKaGN/7i60Cka+YVH2J2748h10flF+8FeRbLmMnv3cVxdX
M4dHzhhTIQJGvQ3kBuxil/t9QddZt0r6FR8ClnzzeJoZ4gG7N05rX73JZaInvge+
G6fkd4K4RrKpE37gkeHG+X9Uakto9PYCDPZ/onUhrOPBKJLLxBrqgkwjoSWILEgX
GixrLEY3r/mIWVB9HQ+5tVDrJZmkge5kPVslI5Tfa/oo83PjIrTv1ETIMs2Q/xWp
9z4FhjO0lJLD0b+ZMG4xBNL65gULocpC+1y6zsBjKzs5Y51K5pLqc+nNtv5xHBEl
nbXtgnp86fPE5HLinrYqH9SgDZCntB6AZ4bEDwQTaIRenllzuNjEAABFna7niR3U
6vb4x8OzzE1MOfZyHaKNjdQjC2sbDR65ZdFbYK4dXowJmJsrX4IyUvsIy+LCfqkJ
PywgSoYyHBk77s5YAER+0t60v2pguqOTaS49Ix5uw7kIWxKl1RLfvGxibg61UlID
OnwGpsNJ4FlEQimdLXVfGP4my61+CSJCIBBCTbxCqrBubJlMzdzrh2MdJY4hO+tl
3aRguhOsHv4lH+y+i4G1uzvS400AAE1awGzl6IqcJEJzFqamq/wtCmDPoHBrJf4I
CyVa/hgxNrQ/p4DQO3naU27m/k0hPZ0gnt01226ysvsXPRYrPXsiWgr0AFf11wqd
VeHIADPQlkZMt+qM8ntu6jlb0L9lJfb77QODDQmg4AtThq+BGCDlisghFGbh+nDB
UPEYOHnGZqqWFamQzacjhiu9ThldMP/OBw9cystPdPsocVyHlu1R6harJqMAsb44
4k0r0/UzhN9bRi1QaQhkHTz7jHvnrzu8hcqBQmeRDvWD/7VJruXqwIhUqK+Ndlgd
/a0sUVVce3JwgJXHVJiGSw1njr6L3nsAOMQ+8lfCuOveGkiyyUCmHVlIS+5N/E3A
UN7XaYMMq6nIMlXSvbSJXrF1bhVEsz2Hou7qQhTfbtCLtkRf771KW+3xl++n6/yk
hCUa2S2Lc27w+XEVcF9S7qEK9/HnUORIWv0N47LOhEPipJnxPUfFL0w/SqJ2adff
vzhHLi8qI6/wMvMLLGe15N2QtT+ot1j4CI4vT92pChyIDdfK4Oft9EEdiEMXMGKZ
sz3m2hn70kHNm6BOiwiehMKpUpHT+bIKUmDULdTKBR4rrlvmxLtwtY1ISoPQohQ4
FDOo02O719kPzCRHDoLwraz330NLXMWlqw82H2bRx3S11IO5iBh5JeLx6u2keU9N
Wa5IvPC5e0GUHZZwdzUKllLrpLniM5LDykgBY7SaSLn/64YKfgI7U66J5FQw9Cg0
TZhtFvmZyYVNlVdPduqSFVbsMhDYfIRn8LDBJbIaJhRtJ0NjjOUNWtxO8ts9Yfe9
bqI1+/nKVNGeo1b5QcUUnbo0h0soDiN87yuhBAHOki73hhcojJVfEV0CZ8iAZcvD
MXFCJ/Axs8Gqj4zJRfm/+lDVMyYk9rX+4ih66woo6di0kvqg45vy0nP/PI9NXjvP
mc5NkYTTDYXZY9mjHlv1G63T2jQpiXqmgmNu+MY0o9IQFXKkIkGmzuZ3gDIqoFzl
OS1w3uWPw5e8jU29ygt7LNKM2wUkFCZD/R10sG57X87mVn80JChKTzraS+aX9D7P
YHjQp5QwHYrfcB0BUKyP5CN8XB3Wq21s2un8abYvMGGIhp/WObyCm/uSu/3usw3J
CUMO667IXRxb5KONjs+c9aH1cCutzWqIUKUzCPeDeN7Y/Sg4DHEc2wF7cfyECZlh
ndo6+57xVIK/THFa7xp+Pl7WIyjKAY+UZn2zCg4sfxCX29JKSlsqXOWX67P54rdt
jC3rwAfvXBqn/g7lrIb3Ngnn6/Hn/swTZi3a60x1rwisEP1wZrDZixuoo5dVjx98
0CU0dYR2IKPuSkGWDlWFgwU4CROXcdk7YBdm5c+0j7v5N+NuNJubDGxbOodC/hsL
xQXAUvYfMGu7lSZf2OAkMqfzLWcmk0+pf6GnUBGtab6S1tcHRCNR7quPgV6T/Wtg
OViwR0QaGvjeowTCrUPYHb407bZLsdib8aIBBEFIU/LhF1MwfeF+dgjG17beZ7kB
5EsdaXKTWAc0nEr8Xevr/5u6A1VAk9WXsfgkCBgNqw91suANZ27kPsUOR9e++XOQ
TiMdI+VLHcgcCxycTXeZO9+xNwK7FcgqRrDhN8RreRTGtxeXLxeRzK0Y5z3nQZLr
W49NK5QnRjuIIMbnpUAv+uIZuT17H6s1K5bF0B1OJJjEbWQhUDUIZ0aF/LuwUYW7
WfEE5F4kbGM1KIiy0CW08MoUvDP1ZCXo1DWNon6BWQc+0T+cx04JE4oIsk86mglI
XSNLqLIGITmX/wIhWF0/JsM3JZfmc2rPH5edICFPwGFyUbFBXPenPagxNA+aW6tX
jqVQId39NT3TkxndVLHVkhM/M7kCd1iP6X/ex6W5v2QyKS82s+xMiYhMUIpmCSei
RIwrYkLRSpQV8JmUieoDjzplZ6qs75mfVsIiG5m4C2dedKbJlBYwbgqowMe+ZDvG
KIuCL4Ac2FkS+FZ0Ot+62Oc9EahG+tce2Cu+W2CQbmbdyfpdI6KVNFvkTfPHT+Xb
NviVT+hJ6Pa67D85czRl0wGjpA2x3c/X2fzctQbQmfyLKMScHdpIknxnU1e5yBps
TY58H+GFj5/hmLMShEWYt6algIRSSj4Em4r9obZekXD+FJkfdNSFAgGt7cfif+qe
Q5XIXf9o+GXiEbq4w00WyJICUByeIBOFR/qaRnT7SVMLr0O5rBQjGWet8d8JcyqF
OtSTXYayjVbWoHPRXDHzyI2CLfS17w18ndqBiZxfvRd8isKxzkNKpeeS4ziMu1BD
j8oi9s3DXNpdP44UmH3f8LDxTxsb+rXkSuBF1Fm7XTiJk6DW7C/u2j7mCLvJIcCX
Pkreliy8n22VmuWzz3+0L/HYVyqwcQQmrpvDJ/WADrxswF0lu2UeLZDU9rqwuh/T
WEqmywai/6yd6a0s3ngjI+QdCslFgtpd1C/OvplZjOo8XlNkcHWdpRgOEddanW8x
mM2fETlDvpRyGGX0UTyVoi0WlMOCPVjXuj9sUd+LppL99W2jfAYe+oxY7gNTJ+5h
zLcMQQKXSRw13Q9Pe0F2RMUSbHce+0dtUpF+yu9nbE8igSXNcf4ajcpu+SHXJJus
3353/aQMSnuuuobaZ7buHndSxNmXd56z7krpYMwp1ZHll96hl+/hUsuu7wZ8pp8P
y6YjRzV0Zt2MdoQlADFVGHmuIRnieNVMeO/QYu/BKslQJ65lWwBsG1yCYkqRY/YN
p7Yt04DvKJiGHLX8Omts1n5BIL4OY+YYc2bQRu5yPho+bzs/ejmEtNYABNoMsbNf
CFJ2I8gDjtwLrTcF+0Rt3aBoLxwyrw3zOnrwI3zy1/AYrZApCHFOxphq41qn3RKr
+XNUhVUqFUDn+1RWIDqIphmn3uXvGlva3A4hlQW44r79Xk4H1NLrOVrD0HER5/H+
8q81lg+hAEjB9FECRf4uRKkYC5clU2Jr0iAf0qYypmWG7+dsXk8AKjPNa1tbKGzU
OSFirs+pKWRiR6OLVrPWGX2byklJ4QsaFd4gqqpW58KcHilsrHAzron3YpxrCuy0
wXB9dysHjn1ehILVVP28jpEJNRARjrR2WH6gQ2Tb3kKYlXNGBriaHCZ1P6N1yY6n
aaS5dn4TI2ctNatcMS3Bzm6o8W2OYEuBikbGmX1ZS0ThNkA/2aAHXKIZu4NKQV/q
LZVJo2DW5I096vE1ZU9IGgWRvAIEqIoCyp6ontCCGthQLLGPnIMvSuq0xPJCiArr
uAkGcBef9whqrXfu4HMv9bnv8d2Xz+M4P/bPCenAixlVww6M+ZOjhIeh7izX0TCU
ehz/UV3bSyXYEbtzQ13o1xOiUoIWr6/lqgtLkwz3gvxxlHWJIbXl5eRmubBU9eCh
M0MLym8BLBhRAulSRs/KZVmJosxH+YPdHmiQ2XQfVYraaes5Vh06cwHL5Khti5P6
SLLVIxl5V878CIdl7VK9fCj9yCGgL7FJIbxgi6CIge4XEHc1JF+LYqd0JHDFQbBL
zZADKQyj3MYtRdEBp86i/m3QsOjV1wm4aN7HEw11j1WU+MqbvQTGodNUwtaM4K8E
fu7gbFUH8W4bxy8w4cp9mwxxVxlQc3C0msnhR3TQRIPxF0vv+Qqf1KHXc6bZ6h5l
8jJPaFyoA6GikeiID/p8+68GraorkYUYKNX0PBDqhE9egSDeBCBNB/9CCQWDCJQE
t36lQHsZFwC8HPia0USgskjyzmJ1M5Nv9g0ZKpebU6NlY1XPfVXwCmW7cE3u1OmU
HwEOMxeZLy97+KWQaaSHOVWDBXU18Fs3x+Zyc5uEB0b/AlqGPSSkkb5HhUmcn7+d
lTMx+47Va+3jrNkajoI8myzYMxeZ5gHMSde+751ZQWg8nNcnxfU3nSKxhq+xt+Xe
B0dKW127SZyeVuOjkuPoFN1/aziV+n45t/q7KNbwGLz5O1DeGySLWvs0odoXoboO
cEvPMA5wzMKyfSl09MRKM9514bpYVvIdiPRYB+3McIl/whee+RdnkF+gANI6dvhr
xV+jzKYg3AhWqW1cP96SLForzmBtx3ii2t6CdeL/1VUxmxLXRiAJftJKxR9bcRWP
7oboJrmbRN0CZAky5e9YbQNCedlRg3k6o2xo/sj5nO1Q7yUSZzS6nXsBFJwVYTmJ
Y5Q2cQwEcv1gCioMZHlSQEPP9Ra6vkgwdapHazOmHj0f2lbo+hZJvtRax9LbqAGE
WJRVU1H1YIlfdxuDFHLFWTOGL4YlLd9aiyinVHjpK+HAk09in1vDv21QeFq7n6KN
M2pjg4QrOGzp9d6w6bZukpAHh0mAOmPP6HbcMR8Xsk16eNQYcAZIGsZ9KFvCJ1Yh
gHElRmNc9azz99vxWvzlR/Z8PryOtk3xbv+eZ0GyFWOel7a279JdUwRyF2rIqg18
/0++DR2AH74aceK9e9DPQcj2eqEv7+2bbxnHiD5uUqnYYbot/AUM8v3Ri91hEySL
BFIEYHwiA4GXZymFAZaRT0VycTO/ZBLVwqBYKqNYYswnUDx2uVaHIeuUhm/4rvdB
8MSxQ3m5X0M+9r3vBkRa+s7T0GIP5EdWparoQrU5b65eY+uYiM3WeH3MTEm0N/Ya
o/DQ+WrxuWf2lMru6UQf8ygzmEhv/S07pOKS3IgzNvxGuIssm+2FG0xg76dHSsNq
VnkBnQ9NZBXAUunCpJ0syMHfBYl+HFHUUXQAxzXPb7wYfVzig8z5cb6haY5fvdtA
oCVzWrLBsgMBUSHY5TrhdDlRznfyk6w5m4aRqnAhv/Qk1Zk76dal3RPW/4Cr8pxx
DS9DilfuvYkuliKAWLx+sMdi/fw9aWsrEeG1gnLdLomzWKevpd6e+xU7kWgxVF4O
LzsFSslUUUxhXPC4Cuog9UlHED9cmiYNhDLE1hHJkLQoH2buAtrJSe0tPkS/Z/q1
/gT3g9jRqvZGqLuoKV1GnuM0zEy5FQw4yYgI6Evx6FWNVex5D/2x+TjbdwSusjnd
bt7Y4QwYjHhfEQV4qyNNCiR3VIwAxTJIDzwGn6/X3FAukyLAZ6J4ven5odB6t7sk
PT2z9GxszO0f4PfqEg8V360FAzDjVBiZ+6+UK7p2J+3A9TA4yy3UMhtvBXiTNbcB
ZEBSfgna519Re6apAW6OyH+YrSPGPJ4aW1CsqDx0BKjzH2QuCWR9MwBKGq+che47
yOOGIoa/2nZpXhc+EqXpc2MXqS4MAzkn6k4bYRyDZTGKakZjqAHE9oshGW+ce5d3
tZA56WZyXF0Nipmgny3ncyNpFPJI5K2NKCDJn94j9C+jzuRFXCzAg1QTDtRxTIMp
pvREQUs0SWo9ZKPjAG3sOVMukTntEcI0NgdNfIREva8qqsQzEXPrVGiFgcK/K5cD
yjU6ryqB0ssdoj6k+kLm8+yz8cP9dQ5U8rnNU399RjSI2do7d0rUhuJm8sHwF2JX
Wy1thVflOnZ3D+hKThTTk4pIRUxQdGWNQ2RGQn479jYoCjj1oAJWrPiGyGGzWuKl
jXJGyHYYc+nP9mn/Acann1Fbfz6PRaKZ4OI5++JVl+FWJgu8p2vK1bLAUv2B7wuZ
+gE2jW6rAyt62zPasfgSrxOf+jm1MDBZST3ZegXcixPPdFBM/v+8ZnkKg/Yc+wOH
IvnkxMHv0+EMYcX+eOsz+rLCtrGlMsu2+buYonPrepkSVJCfvEtH9AfinZrzvHiX
OTxXoPMf4FXNZakqqQystiBpFkdk4Z2AnRNKWUt8xY7thcbmKuWxLwAcbZoAW7Ny
vwSpAKqoyh8unPJs1eFPmdI1IAG7crI0sNvplScn8D3Adyb5+EOXTGU9RQg+3PY0
2pMwb22cCLBFpnYENiTk/9BNVCKi1h3aFF4atWO4SkOvJwsONoitT0Gb7M59ROyL
WYl3/z3Qbw2FNzo/0zUltG2+jI1b58c2HCZ1niinpbto/Dfvnk2QD2D1OOza9OcV
G409qHa9bA9amrs3OBREtuV3EsiLf7b85sFJHA7wO7vy2GWLxoKULaUNW8E78o3q
LFhPxnv1XR0Q8FLNJrUZdTA+qVThu5C4kOXE51ACMgTpLsWAHLXtEiLne+LTvmcu
6p/ta24a89H0GIy02AotVB9V4EfUOvdKoAi2LjNOuV8G3FceAFkx5hkmPnjyWJ0Z
jpQrL2eKmNQnU9rTfMwKFBq9ZCcQZ0UWG/nZ/+E9Qa3XutC/uNS5ptGYkTE29VEx
ZwQosKBFFE2Pc3ppof5oNJx2pquvBVIebCFEKjR8WZUnEQ/5Jg6edJirwWiXBpQi
1oyw2DRn3Y79PyBd/lJvpSYS4d8Y8S4E+2VyxzqQxgG1xFwEsKaasaKOb6Np8LR4
x3QcDAxsz2pqTSjT60BQPG1gn0Q6X6MvBQnq5tW/HTbgc9mcAftrrWZW8NXM1moD
worTtzcb4YptjBbcXw4kdf/FtkQSmcUAZVk5qI342qBCj6tVXMlOQcg9moyhyqBe
1X51tzdPSFq0Vx6K+mVKydN2eHXI0LahKlr8CTat9NwQAM7417YoLkf4K3wP88Ik
I4OKK3UIsVubm2Yud//BL31Z1ajje4Ob/363ZvpQKpQcsJ4VPZ2qJinMymwsI7Iy
xgU/m+XGp1u7N+c1lAVLzZJghrNJKB8H2SumKG0VbFd5elnqxMa3XMocQ1SSdHmi
f8tZmR1PjkPEFn2BV82ZoR9fr2vo2KwoB4iEBgiU7cLXNdNi9aPrgJadzwCQNm9H
rQA6CXx3qbKLcgS8Wpx3ia/joF+WRED36aM12ACEXdpkDtQNyCsDHmq9Cq/TlOts
qJXMMVBdKeLpidBGpBgO3IZCgpPS3wNg7xDxILk+ViCJROaDG8GgOKF/YTLCEr18
kVcL9F9En+iw54oXb82mzZokb6BTc2synVrV1qo9jUSmzeTE+43SeLnBZcKuk3Pl
Db99q3/8WgYb1W5vLYgo4sP1EhZQuLV8wJKDGDK2zwVL3SWOLKOz8WQ8OSiO8cIa
c7IJ1gwefBqvxF8wbda0xyKKDe9GVHV4uRi0rkXyfbT2W/17AFvMouXBhvVQZ1pY
jY9GdgfjUpiNxDKi4zSSds3r3NgJxkbbL1X0oa6qMEtdSg2cQ84/IXe1myB+P5eL
nqCc53SF5Gm3pzNlizZSfC23WgpOItZQf+Q3u3q76Yj72L2fGb6H+bu1l6mHLvtw
NYLi6xyHKGQbqvZ2LVaDuNYw5Xz39FRndQEjgxs49vFi5sKY2Vb8dbeymiwjYQcy
P834I3vIeMspDMumIS+V3yKlpq5hqN2Hq7Zz7p2WLtXTK092eaPtqoIv0A+I5Q3w
XMb+5HqeidR4JjqJA4k+qkugBiunUtaOOvQPx+IL+5lN8ivU3Bqo3HNekK1vw1Ya
ED4gcUXrLbyppf3w7Pp3H/FIzRjhrXXgLFIE24Zrm5iOd4UhgoMEVmmLYwvdsFQ9
nNFLxY9Loe8JEfTljo5m/5NhpBrqJi4pIiyLn2jxfKl5vWJOs48Ot3iY4d54bapt
taLxCCzzPhNBH8pQnoynQnOY5vVMuHBKFSUD2K9JLqzLxJFYAR+Z2yxxqcZQtgoR
prHOaIbjF3qXrCrtvXy9tl4h/C8GeH+T8lD1FSt6fdGnuxWro4deF2y1LZfQW5H5
N99ixzqC+LzoE1x7Cd5FP5B6hrgnShXUXpv3R7M2qQeNe1e0TyNXXorl3qQK6eO2
2eBOJ1p6WP7n0frAw2I9CVewB2WIFyKqn4RKLYfZuRRtyL0r4uAooe+qSgX+vw4+
PUPina5jgN/+HDyHg+GEVg03D3gLubsvJ5s88lSh69uUPVR8TP8jGhgXFZXa4seQ
X35rMIt5DphTTVKSjIEufgb0ShbDK8y92Bg83AY9qJEjn2zBiS8Gn7wp06MIfuHr
Be5e902Kh60OQja44OEl+RnVbj85Z1s9vaesDsfsZD3uK82NE3aQV0zqUi7j7R5o
apQKyeL0iZkeDeL4Pav1XC5MybpmkK5QuP87FpCvQuj7daPk++iV7OsuRwm4t8zS
YzbyTPKvOWB24mZj4bOAqsw4zmd2M/54MbAm+6l860WDU6HlpOVrYIgbN5XLXYo/
oAlGNAFNmnD2uxHXEr3APFFxk3BQp4KKaPzTDSUA5T4nWpU88OuD3+fuXkxCjBh/
gVUPjWLo/qdWlZHGKHxCGNWT0LzNPbbbqlkYcCWH68/5jKOJ/0w5cRKuG3WGBogF
1oIpDtOAK+KNXCHMRRiudKnsBbnWvveT3ETAA6ye2WGgcoWYHuZJFxMMQn/2JvqM
SnllEojpy2RCGgKj7qvswmqZMiN2mpRWDRteY2TkehPT8scIZRXGLA23HhR7Dhvp
+BTfBhIkVn87eWcG12QM8Iv4ap7nhxiTI5+hIpF58CE/FI32+6N6CN6kMhxvXUpX
jLR9tBNDsxoE7K77VVpBjfbbnqMk+pXZhKAU+S19ZAryUMz+sDmMmKLlr+MyCi0y
GsetZwYvRZZN9NDJnsmwREAnb47ptEkGNLFB+OVOnnFtuxJ83838YlhIERVzZsJQ
dSXva9E6BKSeoGB7sMTHLnzYhKJK4v4hwV+yhl4XWcLcLatwv5rO25WzXzPi+oFY
JN2AEuuu/gzRAkUCbB0+K9Zqn4TH6s8zRU7b7kyrSG/NAE7Il4P2qkxQ1pPm2XNP
EX3G6N/B35mkBIF72Kwn214WiIJ1spyWMcSDxxdp1vbw6PN9XX4qqws7e03WU7LW
p0M2HCH9SXRGBNxwSdZGnOaP6fsF1X49GMlwa1oq+sThCXx8WK3HGKbp76ULTOs9
YX+94gDC69yDvml3LE1l07qTl0V7ehmnM4T7wgc5lfXpFQWfcPCGE0vPPp74SW4q
v1jnwtP5Z3LG6kAX7uEiBL/fwqp4IVthA0lmF2PRsbQ++paqIPHR2QXJ9v/BVaIe
BxGRaZVkzvcVHDo6QrKpnrXW+u+eMWeQqszDVAE+zeiXGk2QcEdq3WHFnSdDNIcu
QiLrpb9OtubK/a4ncNFIWFExmUuGjK9Ni+jJ+QfmH5VQtNF57dzZbdLGd7mJLcQu
uL1FCdCxZMTy/imVCFv9jU7rcmLWclTo9YFm2h+vlir9yZBpomTMtT0Plsi+lI+6
cp0mubgv/DZUZ5UJ2xf/ghjCBf/qNDWlQqAw5rVtkZofVXzKM+kzRnyDqiFICX47
y4elOe2qW00RSvP/aI1dKhP0of752CPSP68BYB+xs8gs8G2YowQikWZ4ag09W9LC
eZx0s2ombU3FysuZaNGJcFm2cm/vYorijdCWcXEziQO5nSLGbjJsTsDwh/F1J5yQ
Fk8vdC7dgUbP8jPl/druIlwXdW5TRfUTG3dOfSveTn7rBP+FCpk+GuLzPVeenAR8
S8At9RmF0rPf9sP4G5dsg0049d8yBlcCBeknmCFfbbNG7jJrn0H0D8zxde0du1t5
ZnDjjBia7HgN6pHIAViUn1is7Zner1p0hBxrnpUc0xnBtMOVLfs+e9+rToyStlf9
/KGfW2CgmyGmGjh9Qr+Z/HXtqN8U9QDcCiNQexmGFwKUU9WVpRinJ+KjuvYMr2m2
82ZeaEHJ07eFo2+upZ/j38HGDK9fwTxi3xgOMZ+5bCaScJo/6yrrHYD4KCbRKJGm
7cPi5wuGDpPxfbdCwoNgw69LDHes5z9p6B/IvGjrXnF2+PmdWoJRIVh68LhddDB5
ChLgyTuuAfMw/3IDwAJLkoZK4k7jeWmy288R/BSRrc+lj9vRGKrPEx3CX6YvOLu0
WxV/veAAQv73jbiTjDzcm5rbU90wSX6vmtAoVNnal6Z3DdYK4PUrsngl9Msbldz6
E5PKxULwM9UPFhidgnoI4aGLbk7mdS1ELBWtlkk3kPr059w4qpaKH3NHYYfY/Gpj
YGdZ8fQfbl5g5ODlFVzyHE0t+VC1tGXK0tTW9hCMPfdSF063QVgLDb3BeBUObV4y
WxKtIKE6YdPOJGGbHdGHNevv7SbgLTN8c+GUx4mzOpx8GujV8VPFU1gS5cH47SrJ
p2NS5BCSOGh9mMsC4KiHmDSaI5oILceP7IdqafWOVp22foLBaBFUGB9McP25MlW+
kMFizIp8Wtqr2KN2uwkAwdIBndyzzidn0bjUOGQlDzxEI0nMpXD/DTDkQWuktsKv
NeywlRkK89sbAMXWfjHrWYqypBUoeo7seK6nRtOtShkwwFujsET63CPLmA4lSXyz
a3QH6koUJLJ3X60Fa+A3upwAH3lrCP1GgK0WadRj6bDxRAutWIuio8G9Ko1eTNYk
adtZ9mzvXyb+f3ltuqz5VdDt7qX/av4L2ew6DR72W2XcBt9/6mBY0NtC75xxzfgW
zV31eSiny0Ja7ecSN/axiIgtTTEb/ffsGvSUmJtx4XmhMohxbvsvRX3QXgjBm+qB
k761FRYouvn2/YOOxX0GoroUla4af5Bbo7ZHS/qEfTD26LoVZyudo8pF/0iP4ns3
I2NFxzEijK8uJFYXB7ZLWFs+iYvGXtkiNhXsVPiUqMxsc57JzHN2UDFJhUzIJOOF
Za9vAog/tHxmDV07KQ/Ox+bi7ysrd4bo6jzC/tFsqaXh91QC+D6gvnrOkI+TyOCh
0nzBBbXzBF8GgNsydQR+Rcve9JYd8ZDRvJ8BrxvI+pvVZx3yU8s4aFQ7P1/kuIBz
TMLs3ToA7M6K9QOdCkbGSTFaFkvW1U/XPCWaZ4StewDg/2/vKKB/ixdnlHZjwL0h
1uF+H5NX4f4kHQQrQ9Rh4eAHb4JEJrUE0t9yZC987WsK6GgfxuM9Ss0/ZnmiTxKJ
anYJOLt0LKseCHohFEhTuBvjsUMikGq3JzGLrki8fxSuYd5MGdQuvVkZZjxz6ulN
Z5GyeeJF9ssuF754J5N6Cxjv3ernfPW5v06RNYlq0zBrcx8paKucrE2oD4AcnZiU
MXkCt+K97koRkoOD2RMocxnFo7TFIlQWWjUopY8FZg+uUUzXscEkw8/Z5MQTNb/l
NO74AvCnBkw/JcbC5UHptYp50IJxsMpVkYyYw/EpKz7DYF0kVnor6WLj1UTVOsXS
0NMRPSngl6E01M4nsgxWncYQV1HopLxYB0ttXYBQNGlBvIDJIbleNw3rzlFmbi9Y
d2ma+oYsXZGqAAD0GALIs/P6yuXgPrToRs+/cGqWgaXAufkF75xFZsiNbrIkCi0J
bTzEUFscmtIWUI4VJIwRBb5ZYqVqjcnGrEu9LNtynfx6jBc5Y/pvzCzFei0NRGm3
Utcy4peNXHlgsftAPjPyrCJQSuO1RszIeMUW4vBxDrSecKfsPv/gZ6hDu/QdW7uQ
YW0cwDZirmINGYJ5SMRw3LuxjP0ddx4V1A/Rr/TUZh+9Hj0I+zHAqEpcqgintJzf
JoZr35mZZwo3XuCl957gWCLnqyGHxyXF4H8VRWSKncAivToUMNJ5CeEB9IpJbDP9
d1blAKyaP1/sO3vlB905hfsaAYd76xYHglftUhFB5PhQHiJQxYB3jZ8wGeEW2kpx
21BWZ5jheGiPLRCQp8uYXhno2aCnaWkMKnjH3gdQs4tl4dQQ9W6xLkOU3ZTVs61p
nSUFjCKocVHF41zKT4VbR5lMet9rMV2PQSXMxdBvx9shXnKYjxzlPWhaqmRJUPh/
7gyld8lxD8f7GG1+DdpsLTMvX0Fv9vuVwUBF6nAQn2UwtIdJv31bMnQxY8GGpzgw
4/UyN40C5AzGvihFs8JSxD75k1GMIdzlKijDdrqlaolY7S3G4bk/C+1ixQCS4rw3
Vg/PHH2/FL/BTeS2ehKfHpx2fzaj3H/yMTezl5evCITrnWgIabVwt+2JC1xNJPCV
w8I8jZRswXbb3RgFsHJQ2gDqcuwf35DLbhe4nFLMsmwI4ArnHMOj4x68NRaa0GiL
aqAkc0Vp6ZPuusth3VZVobQr6TBsflmT9J5Ewn7tuejcduKxlBsNL87N1dWW4HaY
yJAA7BzVBTu7Zb1aKpinOU+Co0CtfdVsAkH4EEnXgcutv5VlNcvRjqsGAryOphhX
uVghBXeZaZv2RuQbxj82I6NtSXBcno69Iw6iwHh+e7iS/Hd2pTMTRvk1l+HsAvmT
RtEDK2jDezPYPQ96yJYxMHR4Q+NjXI2IIWthZJEKmUKH14SIJTmZPwx3isc1oQ2h
fYe7ozbd8963szz6pf775clE55LT/BYS/JnM4HGzNfOIr2snxPprvjji9OshFaao
NrjsyG9BU2tH8MKfQsaZOdac9iqCmfaiVCpSDudx+PEWOb6ONTAM6xHsyhM+drWe
txvLelLI5+ppy1TFhGh0A6x4psErSgxwKWrTmlfugU2GQdrZeZSJUy4QE7zCG0sP
nLlovnJRN5W2COt3R6fu/ehWz7VVCS7JGyl/RhrmoSmlZDj8RCRRGFj4+Q5Klry3
ZT51xRwxkNR7t4+cLPw4GcokOKv2BMVs6gQVz/n60cwjkOrV80J8+CNZEc5p2Tbp
NNM7OwAETEZnXHjlA1TS6p+hGML3U9hPe0tMgy8ltCG/NVYy4bd1gfm5YlwmBQP9
E8yh+nImVXfeJx1NpdoXeXg7g4wQ9veXFArwQyOsXTSD0m2aX1EyKwYWI4x0ZxWy
rYT4z1Wc9AFPxWprySCupQlXrrI17lsVNpn1s7H1DOFubl6z8UYiqe2TCYs931dq
4n1Kgz9kWKlN31EtW78wSZIhI1C1+4XlfBEAXn2AjMT2Z/BshRpDa6n/7aCatup/
nmZkn6NA8xBxqXxP4fkIT+nY3HFEib9h2xoB6DMYcXkkJU3k1KU7b9ZuiSo6B9ja
2m3MhtXCWKaTDwRJRqHXJ/7+NfTzUkR146l0WC2MYRlh4G+9u1mlXQOr7gWmajS0
uiOi+NAx3Z4Y5v2FBRgBTJi22Tw1QcGTKImPYYhHiaOuSH+S3K047mqWgd3gUGsK
4b8aN7w2xBjXt5m/Fup/iU9TBoVv5plXH/LIiwil3exu8dwZrVBE+mArAPY1H1Q3
/7fgOWlBTOfPrwthVZKtxKsX/nCgJggQMM1pQkxpd13wgHKoMKpwx7B/EU9ClERW
NZf0GSWUIgTwHpg2KZiPspMIJ0TJ3rHmeovhrEboX6Eivdhmz93AvQS5V05sbuIY
zeKp+lOPpVHO2tFRFs1MviTOu5+JR1DU9m3S6lwN05Vu8YhPYMLH1ZR7UU9kyetF
CN4yO21cHfeQzEKQT2BroYORutApAup65ThgAyXzdArcIOL7Vz4bAMqrAjOoX6zL
GUQGWdVhWSctYYUlMNZ3rR4Ou5tWwZD3q0IooWfcr/Cv+ThdsiKdzwZVY8xUByFm
TySrAjWak+u0PxpwwlfQIaO1WV6Y3FRDO+ZzIOAG3YVLNqfQlQnGcXg4Ajw0xDmg
xOpYnJqsnrgkf5uze4KrngpS1V0jxoKnzN55dJqhy2BCGeX3kdKe7YWPwdIib4C7
D5l6t8gFGp/djRzouT2cP/KWHzv6HS0wCZbhS6QwTMJ5HXBAl3ktlR0OmocYvbAO
SAvTjnwaS1yL3FFBlj9iJthjVCAnPkQjW5LsHsW+a7gI4ijg1KYSdSHcDWxYgceC
GhA3lK8WQn+oKLvzc+K/sWEjBOO9ZBUEGeBIw3sYwGM+cMyaw5J6QJUcLppygGwx
a/ibNw8NiT5+mvtwMfTPUKsZ79rGjXN+RB/qXup9vdFQdWyeXVTdkiztklzPyYXW
MERPWebac1V8ED4blIxY0fBR2VQxMwETOMiio2mBIBVjJD6ytKl6Siwz2P82fbeb
Jue4WyoTPX56RYWrKG6JShMKWS6m7M0ZosGP+pzIk3fw96iY0SRz+6Jj1dKFUeHX
7A8xK0U53PTUj4A2ORHMJfVLO6rBRbpLczDP46+Ai9WwChVYbqdYadfWfRFWWDfI
7teb4uJyToi18owvAKGrNAihI4hgClTl1OaoSxTapn+PoMwKAZfCAVap0OY243x8
WX4XLV1Pk/kGyjJ8dNRHk+1124XET15tBvvVhxujxIAXLTdZyh2MXVAQ1/Ue79Su
RhsDOwz8ifkPH5A7dC9ohbUdyPSDlWZgrwsto7pVTPmafaCPpVoWq9Q7njIvBDlX
SYIjBAM05rLSRGc2+Zg37AWWJKoUvgT0/MTWbsLi/ZDjQWE5Ndg791U1GJBHGSCp
OH5sov+noEc/koXl+R8lWFF4Sq/kqMnavzxmL2jCRnGlbtoNZRtwSHBWvAJmsz3/
UBffu0HfhJedBkTjmzBljVXoUB3Ywuyck7z/BjPMUzv6dJAqS0FM93SXwoAE8liv
eVOSVFOIvgXZ68xSO2mwqbxjDz5aPBSmqYwdmVauMPF7vTvAqMa7n8MMLyTOYFi4
ebKVAE/Tv2Ko2PDSrj0AvP7/G0nWq/vDt5lMF0WzTBPI3QXggfa9itDymJ/gb1wj
AFS8vfNWyurKWIJ8jB+TlFg18RLJ5oKGW6hKMWa8uyP+ovakk2uyQKkShO3vVX5C
Fc2naKW/x7E4aWdjLpnAH5TOKYhSMB5hbm8AC9h6aH3tjcssjaEhoFFpn8uooSav
lq8/Cm4j3WsEyR9kq9MppryyPudXNLBdHB2Jpy8PpREXQ0rpx/bNC6tDGCMPw5A8
hIwXoo5+ptZnBqzyfNC7iIkTZ/5o9Ffoo7fHr9OYtiqbXIJKhe3iiGKaO7wckxPa
lJ9yeoFz3wRnFT02OsGScIeVKmiDlndKEArYdNNMqZGddjYVl6dYYWXheerznBgu
kOJJFw6gmU3NwZlEBseUhmyj9lNM+Wr98KZGfJL5GQ0h6aF7DW/etZk31AD+19ul
5uoNHqUhGo+Q2Jc41F5x0k3i4KkFxb+YAX3Sr6P2WDbuyxsNF/WnWOdUmYiZwOal
4ovu7XIbq7r01cJki0snQeaxOUEI5D9QF7rjz/bDxbNEyRv7ztepNqZzMaT+not3
B0oPMUcMqRazKWdWQ/RMPhjEc+sYh6qpdQvBR6R5+nnTQOEaGx6eb31MwsnfB6Dy
7WdsX67KLpwI6qD6VgXtmmB9z1l251qYD9Jfh6d9Enjgut14Db9k8kDrN+y/KJUI
dsIyNkfZByk2wHNs/0c4taU6GxdPRyv+THBKsaPYTknFatXPaiiRVpR7ytzbLPW3
V77saEd02OcN7YsMlZKailfNWpBInKav5ESyCW7UWCIa5woySgAuzl0aP7UaiHpX
nZftKQLVILwnGEaJIy6UyOfL3PeOr+d6Bx0YGSBJf9RLZoSmf8KhZuLL52Ourx5L
mycq3FSkUmh9oi1P4KLvUptXEX0+dU7pkmAfavLIFeAYJV3k+OY1OYqnf8ZaypaF
ImRDwfp6KnSRb7iJLO7tR/oASTrIZSjkNwnhlnypFOWUE+ZiP+SvMmNfi8fhJaB2
soN8WasoXQ/mR/VHws7WYN2Y0fAgY+pDxe8qb9HYj9xwyzMcPCbY+SrMQMLQIG/7
5S1HHki8dohFEx7ICdsk38nGSEK2TTmcxM9gFvofe/cEuRBe5z7MFaP7k9AoSfs9
Hcyj0aJWXWuaIq3QlFdt1aNincnD+8yXtuxtKfnzBxHQQPo1h+kqGo9AKiEjjIV/
ha6sMXbueE/Qj7OygzyG1xI47m6Qq2cP96FF0qHqTi8rfbe52tBCdJE8zd7p4B7R
4nTMHF7sSIN3/9IUHSULHcqehx7VQVDDovEXQ/dSoq+Iv1JdoHUiO1CEqsPWIwG1
tyoAUKeiDTf9tA0xD43NDvu3XuGT/qkIbvEkvCKDDp/H0H4cpVrup1AyAOw+o6wz
enawTKTQ3ZyACG+NtWFn9nfxw5EzaKw9IeJhhWoy7p1Ao8WJRHtbOvAXvPGnAZNK
RaTKM3STpES3KUtc9vXcb0jhAJM/ZtPe8M4q5ffw4PIO6k/XhWF0+9dpKOmclVwX
b2hmUewgPqFzamPUsgAzwQvA9FRl5E4IpI2ip0IVD63tbm1KaP9YNy/L7uGcCKfV
vKRUVLeoVNDig/o24OqNolYkpOfsKJ6zrsiWdRiB+U9wP5UqxjkYkGRhCufTRwTm
zS7cgPjg03JjdEkxJIc37sQ43d/rfcDIWzR20iB1genf1zgz/RPvgZL3HHaDmY0w
AmUY0hrRo3g2ESouMIb4AGEuArYKjsGqElAASrsLth2++23oNgIt+wy+eHfGGZE4
E1wdq8mdWQi6Q9IJ5Mn+pYlKlXaOofqgvT+5aVUBH8BDb9lYHS2ntjvG5fxNfsBz
60g2RXFTqefYmF/6wQIlxSZOVrkp017sAiLOOaV9ZLW9EmmZLsUMFsvFNdtxIgYo
iXtg9WMxEfnttNqFODII+NpBzQ2oBZpP6snqZvbqZLz+KDwpDAL9TIjXmUmZPOIW
kdnuPqnqQ4DvEsyJk8isVLlHTO6uhyj8icIv9NJkrSVV+N0DWp57RMsKbx5Vbmuo
6UqgCqAflxdfiDZhRoU0+EVhPvxhXipZzZdBjOUI3S9GKw6laPPIGkBHcfMGi2em
iUS8wlB9W2oGaRZOv0lDBAHC9lB/to6AyOB5jVU2KxAbQcUhJBah6Gr4Mo30pmpw
r5KaK4exw5Xd1MVKvjMLXTCnhZeL6MT59UZpldMCxhg6BeXsOPBdJkdL0aqy4P1i
vELNCww3Ia2o83JdCZ6MP7AAyzIhHrAXip8vNUi18kLEjY0liP6hDo3ifnDGiBl7
1pzIBvM8zmFqacdgxgJKQSLg5jFfQrMNFq7zwdjtkcAmwwa/6avWlPvx7Rvaconn
5oVBQKGhuzmQuWIv43KHFs3BVVlhr3M64lhRKlm/mhIItd2emwMv/+q+cIR6mLKg
I7CHkzWN7MeWhuhkS0bSMcXmOsjudpjDS1QsLjoWybK5uZGsr7mNvoZSuLi6FEIh
1nbnDIs8bkaxNnmWTllS/G5VAEpA8pCyq3qrah0yVUv9LzQsmz0BpDWVb5FfWDp3
p3n1LmfHNsEwakwBDnTJl7new9wPaZ98uGpOdao6Dne8JEF0sBkEqIv8hw4KaK+J
s5vCTDFTM0/e4IPQ4mtSIbyq1ieFMimsfOxi2iLt6qHD+fvpKAoQ8rGoM3tAUvMi
FTCG/tsHTybIMV84yXnALhTstOcKLG7egpmutFWGZsQRqdLubVYsTC3ItjvZt+sP
oWaGi/E3tezqqX1ioR9W7M+G3O4vB31vmTTau/Jr2St5Yro4E6kr7nezSf318/LW
c9LY4VzAK8U2qA4NgoLLKpuGJbYfoIMEixYZtzDxAIr8e3Y6MOzAotXOdxuZsAOf
H1uM7JJPmuLy8iBRnZma60nx3Or3x0z+r6iVeLJ5/xU65tfBFdce90/tfvT55MIe
GoJPqzQiDvUyykpjO9b7LvzSwStl9Wo6M32PUfqsgw8RrBimDQxQGt6/uqG+rRsj
kX+Ng3KDLvx5lCd5ZMyHcfK6nnOUM8QbGqcAhGAmz5x18swfrhRuLwE3Eeo1C5Ev
B3PbILVfGgBUy/ed0/i91kcI5wLKG0G67iv7XwHLD6l0+Ocm+4gEgbIiKVzrhpGR
teG0cqhIgz+bM9TqGOkFtQ10oa8f0KdBABROb6tuTpa5lsoD6QQu/ee5cwDikcis
YVhWAdLwr+n+XcGL9TnDMqsx3yYuym1Z9NI1F2A2hXzQGWvt2n2vi0q1w0+AVpHo
P39olXmDSuYwCd9kEI0EHbdflnA8tC9xeFNtZ/ja+ezNry7O1bZ71D5YpnAxo/Mo
9m6GIX4Qs1ECQg1BGQrkS/BDzvzNGTq4rKRw+J3t9sM/uO03eJ+BoMmhgG59qjeR
w4cQkET6qqt2l77/0DzRXfPBVXw0Cx6+KSFn9Z2OTq48al8i+6rjbMKovb1gCSn2
zSklqDuS9TeM3bJiWSZmPF3UFSAyGqDtCJJT/fe+ADpNyHkH2FZTwrQTp3mYcRKU
u5Ec5oalrYFy1dWHN9eUwjvy8HMsf4spySXgmlqVKWiVcqB+YKN/hgKCivxv/asT
6MLglgJBsCtO14iV3ijWXZQaSYDuCpPk53A9ByOWuW6Oq1PrlTcr5AxPYjrt2zt9
TWPxaLINVO7UayTx0S23i53ZCounSLlz20ALTrOKuqPk9wG8HQClk1GiwPlBmr8S
ooVjrTY3iqGsGW9vrauLyx9Unvbw7KauGztDTYdaAy/fVByMDoHr+mDm4tsUbjy6
vBsqYvitSgGk0Pm6JfehGXAvU1cXpeh/8pf/akSyLqJKQMO2iEvCWSLDGWUojJL7
ORB/tpUxQW4VBJ05WDhS1eqmVeZyN4Dg6V/BH+8VuyUgaSP+FDbmZ4ifgjCex3NF
Eb2+I1uL0DSwAW0VIor1DFmyvlViubX1Y3XPWsg5anwIyLV2y8UbdVlzOan0Jn+F
R5S7H5dkTqTOHxhNhn2uZpCzYY43/+04t0Mtx0DeEBXtdhZtcY3bkmAW8Atcaucw
WRm0mMofLspZ1mVQh+0IptCw8D34gbz5KMk1fsLROf6mAGaKQeTTMxlcqJfiKaxH
DKFVRaf3xEHuR46B5z8ieLdKxKbWUME+EJMPFmlMUpQizrGTTqOYJxJ8khoeQXlL
i7sIp5J2p+b1t65x+MjOJ/Gj63jysksqmI2AoxfFMfkoE9X6+9QxzYJ+Jfk+U6T0
iVpEMCJMNyaa71FXhntgCyHmreoterHPibZQ/sfFa4qslM+H0YcXmvUbBjrUamfM
je2rRs7NlFbqW8HRWKTBPLsaxDH/9Vweg+gImkkS2HP8jrNn+02IuGIqFkpVGISs
c3RRp1J3fy4a+ArfZbFmDcplPpt54aI+hWYMlVo7kGdkJktcvcHWeE5r3VGnxVnF
N9v07a2VZe4/kczYOxNl3WXT4c4mFwksPYOf6reSNk41pdZk1TvaYNB064m8YDCd
kZmmFV75Wqn4yX4iwfWRc2jRZ7hMsFZ1QTS9Oze2t/mm9SlS6/McGb5yKUW0hifK
ea0A0mdLU57c2qKRXx0Kc3HQY72FMV3eRxzBa7ViSvqy7QCyMZNqEPkEUAqHTgBk
ptiTKENHUfrF3jVKgNLEjZ7J5aU8pSHHSqMevvXHplvibJhLw67k5MqkxaeHF3Zo
iNSGo0YszkuKjv0fv4i1FPyrmdkEboBHNc3WRt1ZLntETHdTTcpLZfER1wKz5LWi
zZkJHuCBu7TtQzywRPynC6ZyIxyyTqPUzJ1Q1RNt71pdHKvMIxpaa0SRoLWmGrkK
7zRSpbQfoAYWUKaFA9BZddF/Z4iPmGX+sQX14tHGXTa1ZxGIIUOMwjC3rze4VFQz
rtnRxGLPKgrTmCRV8nSnlXND8FZt/dM4liHJUTJWymeMWoumQS4/ROVRg0tQGtro
nLM+theClJaHUet4J4I5rrXpVQ1LY8MyqwZBkYsyXs1rLLNONVVP4mDIsGb9wX0q
B/vrm8mqlBhRjq9p8sUgUiYAuMGCpV+lOiz1pR3ayii9J5cRuP/j+1/TFXwl8rqj
2fEuA7Rj9yx50vO+SUCj+1n3ZL0RMyCOzUJmk3DIEAlQ2EHM6ySoFxEB6t/kay56
QrD/4ETbgD4Upo6kxu0UzLgLyyBnLluLOIaJafsc8l6v84ZIlu+xqwsRxqeOE4oc
m1fHdoLM2ST6ewAiYHN/vBEirGCc30f98mYW8kv3xwUWWK8+7F5p1oD/NT5fedMP
IS5y1kOXTDGynSpHQ7PrauZ5esb9CPQuBiaEhtJESGXIRVRCAZHpP0Vh6SRfXEim
PGZuMQ5wBVnTPd+cKTuNEgbnw11kTi2n3F3ebCpZ8tleWgbAFcKkUpL4NDeK0Xrh
ZwTawF4Z6FGOUZZn1t4qobc1FaBvAf4w7Hi1BkKNYd6H1Rn9BBsByJK57eL58Ond
+oCDd5pDzU3y6Y+/uiwc3muP3FDenfN2qZjk3/oQW/Jw3fJlLJECKjMKvo8HS3kG
KCheWPiJqiuiuJ+5nFJSrmmhUtNhIa6Q/pLKQBEp1MgN211ikYsf9Ml7qbHqaT5a
JK6o9lyJDN/k1Kpy8ITdJ5GYe4HQONsZDDbJEKFLGJalscQHEb5zOP7FWD78Ad92
ndhFUZ9VnTMU+CA5nho+EI+OtOe7uSp7RyvejjavTBdpW5Qs12W1OehiV4UR51He
U6Q3hGcE8JM3hzlWVp089c2r6Eb/0VoeM3D/HJvIUToeTjmlkDz4HCOmVqOOE8FL
14G+2Nuq9b/qVBLFKai2lLDxIVGf52unvkgtuHNF/tRti/4BIw1mz3QCSnaV/Z3o
j51mFiyPNnCOIwGzAehkK5DdVNI2xPlQoXrNF+Xs8bgoC5bej9j2MvSfR9YUe7MX
LRjZgLkohk5r+4eTR1EZ6Bth4SWln3Oqei7mK5JcASef8Rc70+ZPGeOqpvVz9ql4
uFe8ca2+H2WAcg7P6r0yLfg0piekkvLRnJdHeY2RqJEUZP+dAhLD3JX4jZdDFkuz
Knj3Hsh012fMOEmihyj/KNJOgCvTycrA4guuuEgze5j/8CYPh8hOWrcyMw5v7cxd
DyYqTeyOBxSwgEDY37zV9cRz+9gz2OFXCYC7xWdIuVvOsq0biCYaBOMlWuwBAcqB
OhS71+mWUO/aaM+FatSvo81Y00Nl3QxtDa3qFI8+Ulnu21w0E1qHlWT6F+6dBOrw
S57AimYziOIH9WT6JFpDHmzeocoW0jBz4Bt/pAc907zt5QLkiGVjkB+65JwU1Ok3
tWg2TbO0pVMLKjmfVER/4tUQwG1q0lbfkIT/hz6EwocG/bw6oXxPUjoddQKdDR2N
3S1BJ2RljIcDAQZqGZr1EsKYX44rIEaQqbofgDFKTJn7KzcAD9+S2sEkmte4IWcV
JFd+rLNrTnaflH+HiL7rq+qxHpwMR0ygbWT0iIlp80PLN72GDma9P8nxT6vy/WJC
WtXYLyd9GeNbH3GRTSf7Kh/W0qPxtBcoKxPa/ZfZvtto0UC1Ln7tdTYjN4yfalAz
yQ1kdny4bHBlkaSXfd7A100GW2eCvXzTPoHOPuNQLv6esqW6AREfcNOsxqfhIboN
M30sFI5z750wl5m8RV0Qauh9zo970I8QfplCDnYLf4voa+n2qJqpj/HeNz/lz3W2
piSFQjy/MbAuoU9R0V2TUoqJuK07zUNevja7bBpzo4cw0oKQp/qHTTH9SE4hwveX
o1P9TsjzLDhvPcJ9LdlUBvnMOT1KRMN1qfJfTTJuJsvJEI+zBQvdyjbMtxdS2ExA
x5sF1z2YDZFQXmcJj5ihxMI6nERMDgXqSBDynS55qyPoivCkvVwtFghbEMoLHA84
llhBXbNoyiF/PvyPK4HSHiwKuVswEH03fjwEcechElXuvaoGcQz05WS8BDAnuhTl
pT01MW5Hh4fytskhtWp8ugrFeltcDATHT/yJZnzPTt0U44LIczeaIMS953tfMtOD
stFUSAphQ1KX7SARf/EmOR+TlWcGIezDiH2mRcfy3zzkXZSNzlxz46JHmj2rAQrt
306jcPS2Sd6NHyrK6Z4bG5N5IhHej/1z47Un5ZulMa62UEJ7xlcL354hHTsZzbgv
Q2Ely4o2qWIjVoQ4QDCCFcZDso7Jr7ojL1lQxpSc4Cl2S+rx6jJGy05wuByJLC0j
pIuvl7A1QNrYTttWqMpYtR+/Ml7DgsYVY0x7d3kcqfMy3/P7JucM5kCz2E1UOmz8
TWYt7xRXLQ7/5OFEzZUKdvk5ACxGKny6BZbG0D9qiD44/VvniF2sqn1MMew9JqIB
LTX+RN44qlT3gaWbuAJ9Ha76Tr5K7Zqhi75ySxFHHXyfAwOCkI2unqzJDmLBqbQc
2SRr2BukHbxSKOviWkhzb2BAlec+KRHdAwAIXfFtmIE3L9XwhUEcdDsdnmRzvQu2
KegyZJceJu5z4fqmjCc0TAZNPz6Rzp1usE1CFIvQzlu6/WxU39X0DcJMU5SULE0O
mS3L9+ZKdglFUFH5eeuX6cwIpZ8h8UgcvHiOm6hb/NN/YsN3y6m0f6C8N/UCLxQF
1M4BPFC5nkJJLdb5Bu1WDr93YVVM1ECwV1SaD79G6vzu0r/bfiPkl80EZCUIB0xR
GIxWTWEBaqWnJU+fTrN6nurZ1SVVXcwSTDY37sSxBgjF6T3/NeLiXkLumFt1A2EN
Dp0eskX84cUKbWeJmDmB4dewPqaFt8NF1ojrxsyQb86lbEAbsgxnwGAdlvguf4/L
Zijvm76ZLcW03dNA/8JhnJLmuJhbXu/oGZUfEpUYwQeJdrqy/7ZJcVRQX/HBZT7Z
6hhXHtWipssEnAHCx3NxEvibGhk2TdkCw26Efog3hOp7PDp+Y6eyZfmihfXF7M+P
dwtg5Pka4XyyWNJuOX1C+rXhmT1XnY3KJaBbjyRD2iC9zRWbdYCGT7QrXf3sKlSS
/LZxDKoxm3ox4ktgxvfkOLM0HKcTylINWb41ipwIB3FN5hLfW1qWrwmE27CVqFVD
rvTH4FtMcOoBvA2mfZkLIZwCIXgopV37fHKujXHQeLHLDKY3JevySiLci0UKc6yx
ZMY82yCci1JBip82JqGtEGnrD6o0PbjGHqlO9wEJ1cAeco3U6Yv/DVdEkLWylDcy
V3I3yDpCKUOTUasfSbstmAQ8a8+WqPi1kYPF8Y5WxStOIHPRXau66yz/veHk8Vh+
xvDG71IMOTDf45WXTZH1Nkce5h0KjffALFqxzjtFi6SICU1N5AoYDfKa61IYZzhy
CA76Y4w1ZEkh5kqj5CBL/EFfszc+PUVv0IlPPi7wCiCRgZMjuVeBmdDDhZsRHxaE
4mqcQlknjfb28Jtq3rLZYxYxEcPYi9BfxjCQaTqiMGxA8Qo2siNv6JRw6cdyfb4H
kxAO/VEx2Kx+z2jeXdROUareJIepu8+31tnGYYP0Ot6/WVDw7uEAkN90iCNIROCj
zXHoR0CLa7fSC9YdZjTU/cXx6qloWA6zDnrqbr0NYc3C2e1MmDPv3nIE6J/IPcjY
Hkbkk2spL4GXVQzhqjDi0PbxKxXB13aPPUhRqPE9V4f+b9kUzBkPcenIsZIBy9GR
u6p0g5SwcAh2RIWACv2G5xDo8R0A9eXt58SfqwroYOqUIXpQxvc2dn7BOv8+Ok9E
BiTjKEaGmOOLKU6b16je7Xkw0/7RMJp4UOFsWC9H/cs7Sh6H2C/DfoCRPI0BfYEA
ADSj7OIt+LSYPFZew59L5xIg7uq7uOxN4psaECXeHo1Cd1KE26+i9NKyisEn3XWM
/aABAxfEZsbuYMVut6TRnfsI7m4ZHC9+DmFtYglHsrMGC+9TS5sOjtsUVcUlU4mu
F2TFt7jsZg5K2Ff8wfjlDuwhvUBZIXBw4WKBlwpokKZDNXAEDIzOlY5unjXbrjtb
jKz6RgUCX4aIK/e8Uw3lURbdNjxa6pR1SUlwXsaduHEgoB1j9NY7qskMMhOSEyPj
djDdWMdtCUYFTRLXdFmg19VHl58/rolAreN7TAmzGPuRty9S9wcmlsmItvlx2Jke
TDKkWna1prpJo80MGXx0LzbW3OHtHeSN8nEbw3F59nhNevj+BovQW3E5fNiNpsBa
hTDjWMkbIKxH7AiJ3Z6SByFX4hL5X5SeBeP5fGKJ6s6d2tETID1pdPJXoNYiDTWE
fRFm08TY4ZRM1SRWSBOk+CIiRvtNHTNja6f6g8gG3vmuoUtrvQ33uO2btifCycUD
3krgdkpwjFRB/98uMX++gBJI5eIfsbc8ekSP/PHoT3vo8qsGMxWkbsYgP/iDuULJ
V1La8cTTqaz0O2TcgCccUdOSJrmahqqQ699Pouksth8nblY5KOtFCmaNhuPSU9bH
l5TXlfdCyL40cFq+dzr90uwHBDpmtx3OWVoR7x3aqjRrwhdh95nVds0mRVxwYGKq
+qBI+GJRqZLAbi5vq2Dg3dxhdmdYn7VlPHOcqTZoAonmT5nZ0CT3BSHr1dAj6k1u
W1CUndC45K5O86sB/Vy7NLUM7YDAgGJ6gg1DMLzgLroXLRdWTY90fwlSRD/CtN7t
l9SnbuU6AxSryxb+m2/HK+27A6DyENwp35uQvYr97bzgo2n5ABmy3m6Sv5zrM7aD
floSMT8zYdr4vau8B9N4N++74We80v1y5FxP0lWgO9up2jsZkcdmgz0kKDTq4S8G
ULFZKbGW5GarxSzH+uukDHNpu5U8BdP21YSKEIPR8PaZHln6w/XamW7xe+PJiQLZ
QnZKONjtKtk0qq6AYdbp9TBYdb1wi5KmpEpkbE/ykUFmPwUcIen/JJz+J0c7RqyO
NkWI9MXdhpVwwqro8Zru0p2v5YZUbfDhm5LygivlnzBD1q0Pv7AEM7caeW9XoPIL
JFyYFZzw2LUBIqoTl9eupGiktYZfxgA+gAv2twvMqoVUaU5WEKRngMpyKE9MSnQb
GzUcGxaZSExTF+sGLYNJOgTjdQqqlQ17LWyzoavKqIHhPJlswNz7JHqRQNwNi6Ow
U6qXKycQAkBFPSOvxeglPFoq2Cw5xMGkjtHVpEuNWu3n+r9MHVUVYo3b306b9auK
sswOVAe3t3d8ALzjQID03A9v+UhwyyXC6oTyoL3eBBvlV/cCN7LiNbGuvwXHxdyV
kuVnNCkftw3xgUp/FRjbzyP57vAOJNC8SXFVlPtlJKCCO2FRdoNl8Tb0kMxhv6z/
zGVRc2O5uIRWGgA6xXxDgBxEftnYmDmmU4Xk5X1mJHWGC75AR9TUsPRUJbnxqJ0z
RpS6mT7tZX1WHwvrzVRuTf7DWdTkf7rJn4+/V2PLtAS8AYza4knYMYDiHJoO462i
shmv01VDR+8qu9ExFX+NpYXmDzEUFU2Xx0MFWOt3geQjxKfnDYgsn5LU6uH+NGBO
xiBShW8f3VtS6beaFewGpIaLW8aRgLb04pYgc0p2qnSOvDiNAaeCe21IuN4bW4Ej
kbb5PSziU9P7CXdcvK71DgiDdF8tmUekA/1l7mbJ2vR9Uw+4vEt40MMBSTvHMorQ
0yhoUaYA4ArcoNrZUmBQJODb2Awi59StxNttaJpSC2CvDdKJAN6xC1OMHhe9Ap2y
MklqAeEXm8XxIBsiWvAS/g9gFrWLwYj1IVgJnw2Byv4sc7qLNsF3g5QjbZPNFpd2
uEra3HWcnnb1hOq6kqsSUXjxz7VN75SJ3tjM+y7M82u3akBUyaHzR/XqFiDnvVKP
jUYKTmBOFMcRw1PA9TPnI7vVBvzeDRVjRurTp7z8LlQ9PxaMNXRiafDzHJGh9QZ4
tpExUKv6NhvSraYe0FTf7Hub9vlBqkeEZpu58ZK0MAIFje4Qmf8F/kMysDGpiMNm
8iH1cYkKtD1xx9y8wFgEWbnx2wt66FD7i1q8eqFulDSBsxnEFLbQSSVLDtmISFpq
EUWjHF1NyY9b16jL2QGxvy5/PCjrzuWbpi518Lo11ORq8PKjf+GtJXb6k6paGrkn
9HXa9WPZplfBB1LcdNasKyeK5Wg6Dl3n/x0mdtBa2t2ixb8p+JXI2ddAq9xjZzR+
+SBZKy7JyMIAKnxpHGdsUPEL1TrGnDFXUMslHfWFscvAC28Zd7EqkH/VlNv9s6Iy
Gp8lPr2GUBpQoHTGcJ8jyPiVFcDAwvbEzlS380ADGcGJXIhSXxeeAURTXyf2z0ez
zkA2ru4Pta1snPd4FID0XcTQaeLmXLfEcpN+BHnrT87hzH4xKrrj9uk5KnBcOLr1
JyXrEOFE9OU23JwfMSIwfhj8VS0Jt7PtEIewJZugXPcjAMCgNrcyujjebV9bXRLm
l4RC7Tv1wx1jrdBJrl6P0jo9Oz/ESndvKSyckg04sFgNI8sOE7CVE2ZRuKI9eu/v
A1YewqJWxKMZ7PjasFxKs1wUgW6nwCqHA60PaNcWVcEfckXfH7opTE4b5q7wwBgn
N4y5k9hF+SyrYYKIfAcRlg7m6hEQGAVVTcWrModo9TJSQm/3Uja7pKvCII/ag8bp
TT161CpF+yOB9XWrfMf/p0Al8ApnrwAHwPCW3JHdFczJnZLI7L2rn6FFmHwux5Bt
zE61i/M/G5RGFGaHZAxixQvcq16tlqVZfqgaClWQWT9AX/8wbEE21j5w3cyvyyHK
+NJiA10zISfliZAs/Aup6NMUDvo+pTZUZAAxJcta9sTPV875H8xrTmgcuQgeWnhz
P2AHnYCn6iyy0DCnauvscGfXPtyt/Lds9JsW2UninCvlDh8DJBrTlO8WIGDaOTPP
/oVm9pO/yi8WamGwgLVrKUTjspJbUrHBFOsnyjjFgHM6x+/gX3j9+sX0Dnz2v+Op
JTy9YxVC0kWU0bz1/X1NGkf35gPPm9XCaOFTMNvp/K/A0CR4vaOPayI2IvA9+ZIk
eWHqJ287pApMwPe66VfIM/HW218WwyOxqRo4SXEmc/bTFO/Pd1Pxe4N9oxofthXp
dxzUXkqW5QVNRxjYmTgSmjR65agxnc+VolBew52289tXVU+ye9My9FEbmyGWp/v6
uL8q6hAFo50OrRO4YbG9hKrQTfSQ9EYdmJCDAzjic4znZVpk/jQ9gieN4fKYCaFu
0Mwkn9gW0J4eUU7leskLbLPrnqaVEyTWeNsfT0V4epwSbh5n8PY2TzIPhUbbEksp
8Nk1+JiB1EE6+ZBlUDO7sz5qpd12rmvuGSCmfeIOnBK9VuBnZhFH6lNh/4WUEaMH
/SlZa8NlW2QsgV8YHoKkjgs+CLefFLa3lsBH1uw7aH8Jb/dClg8eO+bVFaoAdY1N
1WYISsJfx1lCobP2O0WNJKJA4Dly+aaEI/0rOO0Rbhb/cxrSyOjssQNhbzuXTIqA
KsRtloZwaOXjLU6cabAxWtwUA9QI0UptEqTCSilFwPbVQkJGsd7vRQCPvXciUkLo
W3V6JstQLIr7xu+LaHMkmyvmmXS/x+AoMe0zc7zXsrM4CRJ4GFxZ8NlZx7LEMHZ7
QEQ6CZlywPqOBmR+oeu7P2WSKYFXAC5FZHTAnAwAH/d4xCG8+yXcQv+jUDLUR/K4
asPVasdggvuFiDyKp40SIwq2mUv5du7PT17jE6BYgTGwKLPjHwF2hmXgV5XHW+3M
+eSO/xyJWMQrweSL85Kg8twZTPBE0jRAf+Zgp5TC8AjrnujUWAfWTHL3wz5zYbzi
Yq3glkM/2HQ3GPkj6w0L0lDNpzwIY655Sq4Yz4iTE97eCaq4ERejUOKoVwlpRn1B
FebqsbPKONmns9DoLdW4nVZlXoTCmkSyTgDY/Cdx1fpNWNlh+BsZpgAerYITAw7j
jokeaY1l68YlAE4fxztoY1LLPv2cN7VjEY9AeeNRl5FMqb4Gs0sdQrGS6wQ5xLJk
jAdmlWpo0CeH10M479IAWgLcYHc3oeuKzjGXY34nMqxO47Ia8Fe7A6ML7T7XNlyE
Tfmp1OF7mF8bASA+P/NaP47KRtMDVaqrPjNaYbANnUHCAe9oEv/YLaKyCtQFzKPO
ZLQyablvj2r+TKhnp6DZ3ApzJ4fAEv7DxHK1NMWodt4T5YCzX9/W0Ocap+g+8aU/
0+OEMDjYiC9pxdDiRd4Gra3GIhfx0syubVZj03KhFnsSak44vAhBV2b9Ab9TDil7
NQOFro3FII1qvpub/oS6H1F3VR44EQRF4aG8RZY6+7RhWkXLNoJnaHJsKufXYLON
qMTbwhBk1DnWADwipw7LmcvBuGEV3yVBgKgjUdOsT6zIeBCgOLKHG43jRkS2QtcF
7IEkVTPQqI3ip7ZzmwywofYVBVhjVVH/zaemFax399P89D4k5LDTeawPbEZWvhB2
UDQshveLK4Xyi+fsf9g90oXuOk2qh+1ET5nQCZlhRTfExUoLRb6Dd8FqWsfptoWk
oO3j1IqObUuGgdaIUP+LwT93eCCP/mJ1flvQGZ3g0Ti7W5YKS9LP4N/gwmw7PXok
trVAAJnEZcNoq1DTTNwpYeIXJ2fQuRSYi0u/sBuDCAG+H/KXoFhttMjOcIlgU0AO
qS3u1Ky96GDvQMq5zw+HBeVgvQXAOdKArtZr2UlO1eUByUWPSSVYK2C61Gp0bx16
FxKDQs0gbFj6YQ6vbWoqYlgsDyIFIE1YygWSUfSnm8jXxpg9J22LWhNgFUQyapYp
iJbpWmPBkEgkczwAqSW8UZ9YD5r2UPpcaM+wQYS7YjU0B+DbDp4STUfS8ptTR+dS
0ByXN73ea88E2PtrNrUKyzKbKrz29kDJ/yvt3HgwLKrY+2g3IJ0jr/uAdt9wU6Cq
uq+P4hDP5XiTIojmCkQLkARsH30zZAqyFgpzAVRS+2ZMMXZLpyBdFVvBXWufaixL
NSHiUaQt7IahjI84PBoE6wIy/M3N3KXVh3p4WP2mspELSkfNrl0z++KizXf0me/d
9gl3nsQpiVlYem54IsfDM4ERm6oJZay7bl06gNX62aurwjpNi8WXOI3r/L8mtSpH
hkd1HF1e+OeRj70kSLAD4ZUgWiWsRPT9wWAgn7y+/Nan3jsCT7jOTrIm5SMJCwH3
Tw4eJmh6qd/Ag+Q2ijm7YxpCEprPmli510M9DiFcDBAJ2XpyP71+Hq8SpwBuhNwB
JjMj6iAzrmWVayRGeRSXsp8oLzpvqYY6jZrZ0dxWNh3aHG4wG7dokU5BWmGnf3AM
RvRmOc2abx6+HbafV2awjmEYCfyR4MtLdRe3leM7b5AXQ8Eg1S6MJM2GJAmCkPsa
EnKOjcMufnQnbo+zpy0D3q2SfntzHylCRZ1Ro270jgyKECickTihVFghEOv4YcpV
0ghPy1s98HrZHbOBJ6Ov7ERODA7imQSLy2XrmddLmBwwc0H2tSJcDcvo59gIeTzt
AyKpX9NlBjMa+W1OPGViaTMzeE4Jtxvbd6i8dAl8+hlCEjwRHUOBSQgTlv8kahGY
cDhhxZ/tFyoUd3cbazABzPpzlZr3mE6Kzh905+jE+cDGs4jLgyFy1RSCfZSgdGzD
VElHV7QiWGJtuRaFOgELxduQalhbcXljbwtmkuUT67zkVlsBQhreyXOEstC6UvDa
xBOMQW34cxuak25+jUM/vEjB96bi4FxO4bYwgk1Pgc/6RbYLz9+qtfV/NdGcZujg
apoEt9PzRIhSJp9gKU0He0+Kp35ZyeT3E1kVU4ldR3hPVDjA2XBZr+jQRTp0djwn
AAWQJHbnJ+KGEm9/Ses/lnHrubJLQ1MmlW8G8J8UvAbbhe3UMbqJDNBC/9xF0MHF
+MadVx2kxCudHdU1YT+f6bAWbuoqFzKsCwWgovvY1yaTUnz6gJR8f6H+Y0CGAKWK
fVqDAJVtlkryVRiQ1OGSMP4YzNGsV/ZXWKjM6VFWctNnfPj2V5gSBtb3R3wcZb0p
usp2tElXESwKphfwWpwYGNZDmTvQBaPzyrrQSkEU3wZqqVEM9PronI4AGQ42t+lC
tq53n1QL412SpPXc01a9GCM6mf5kmxvwPaegekN3ui9MGZZ1JcBdNdmVoc7zXa0i
VNh3GPFuOgpoPXDdA+G/pYEyyD217onK93Ndgx2k1Zmgb2i1OmeuD27hQKf9660s
ozUERB0av4yIMcS0qspZpBGIQ0xKpPryxAzup1Vge3U55j+XOeKFpzPkYQOGGEtI
ztuPulHF3Z4SGr5F72MKVlkXtGmvN+GzYFTZ8PvvxUSOkikmYWz+cprJz9fzuxUD
JSYnLyVjP8BrT5RfVMqW8kZWv1CIHY6nTwABLzWh6ocwHI4tfwPToYNWpg/u2WAr
As14P9Q1+YFfMzMfOEsSeSUb0BqUVoJjX6SophSLbOHKId2xL5GCgceV6oj58wed
SMkxutlLVKqELsLWuKkEDrMNEqMaBrcZdqtCFCJoH724BnbCln2qWQ7BXnYrtVfn
YmZEm1ELDnwXsBCcqjIoWo5yHKYQ0tf9FY4GX2akhSBgGim6lzAoy8JSEXvn9JrF
s6ZiOfqk2p8Gxl+bSdHD/TpBpBUXmgsofu0FNkUsUnJ+T5s+HijkxZKr+xJHVAHT
7LK2o8br3XKgwVsh1p9sr7nPi+ty8VKN5IvtfuU0xouRs1x3Tem34wSSMzKAJWWF
o+H3EFQ0GVOWo7G2u+UaqtpSiFhFVvkllbuVeq0oeDWDhFGRUKbMvRas6hbK1Xn6
M3qcmUnyqt+3t6gpHBi6BtH4sH2GVfvdLrFwSTcCj2KeVztK243M95Q1fb1nxaCE
W+R7DDhJWk8AAQPfRNUNQF9v3RrZquPwzFyTJd5U31x+TjIbH2Q11XuM0qKYu6L7
AiC5cKd0XwDcEqfdas6XTGDHZiYisMOafMH0KMFuNnkY+xd6KAb1NNk1+H+FzkiW
lrAPIX3Kh243MIoz+03NQkt5ms7XKeK195/ccvpODd8kzVVQ5H44NW1FuImYUE3J
ECwurQ/Rq00+l3nGp0p7nB7AbTxwtnCLr7/0LzVvPYznsm1oD88XgyYoph1t6s8z
3mwWC0Rwubq2+hVUI0VgLKEiKC3Nprqz/eVROTtjeFsa9cMSb/Snq6xu+vQL88I9
bP2xf2WlXpD4JeOofxPspA9nnB6njjmKtQsgJ3RP2ferQYKF1g8KuUpq9UcBDmmw
+eybV1es0ytHXEYRGGQ8u7RoInQ5lD7JxyFsUCrMfaPcGKsyImHS5egSUezfIRRH
uPawvsDWIDowCumgU+HFDZPRbeH1ZQ0mmoO/6kjgpn2jcic7us4YADOOJQCkatbj
HB5uMZ+6l8Y4j3S2HgnbP0uDJQLgeTo+rmU4olAidsI/A8RDT5YF8oK+nZJ9dKWV
8kQm8QRgwQ68hlJBHp800aY4CrY0vGr1hra7K9os/su12dmc+EhAmy+wLC5Gv7cC
Jns5LIMF+ExN9HHnKdyeLqUvj27Vg/fbI4NxE7avz29VqmenzgubaKD0CaOpUE11
KXimtg/ZRrJJ29fwAJ4z2WX3WhkdJR3WJ5Cncxz8XKnrEdz/zRoDRxF985O+iW6o
oVluo0DlKMDrsa9cUSvs+PxQ2GYL3Y/Eyj9DwLwk/qNw5HV48A4olk+hcz/EHesp
KXLHFYRw3FTYaWW4F8ZP6UdSAkyuRishyNdppXIGpJno32LR6lyftElolZCb4IYO
qVSxYboPpAHMTQZA2Iuwg58XyQql1rIWoI5Q3F0uqNAbp1wzCkEcAXaMao6PYCG1
4L/1lbX3ZQhev6gGvHBgkBUZlOKgvN7Q3pIqNiPsgF2NDJ/hKoDbfyXPwhFSxPQr
iJWdGlWLkHWO/rPvuCcqPihcRhWvST5SIbe6mIrB5LUCXD+yuq/blCxKEWEDxxUE
ZT+5lrHp04q2+wnFKvG0s+ogHBWwPKnu4AwJNH0PRYLHBZZOjOFw87R+40INL2/X
J2pCLbXpNFWniZxu1TxC+R4v1cuTNrzBG5KEoDHV8FcNFN8i39EuoPf7Y5hvIVah
CcbaaZDJKrGUSxN7QvVLcuC7RWFYZiEgvTbh8Wvf/GDD8VV+ttyChwFfpuyq3DKF
VqlF8USaDWShvAhXuHklo+oiKKt5j6oQrQc/9LARLNpoyafBtg2Epzi3RZBrja8u
UQUW4tuC9w6/FV8BbXwyyDvqeLxI8WH9ZfEC1JT+CIgxqPr+rZrRYvKlx7I2+vLL
MGJLCUJR4oDmYcrFq58UXKRaLzr0oA3/ASBVEVC6IaNcgmS90GGl3XlZk1L93QC7
wFLHpIf0m+mBkLJH5E4FJAFNc/kB+uQSTkY2utHkFNRlG4blD1d9rcYrqsJESfvB
itYlD6BmLp6Sg2ikK+iKygMdJ3XhRC4xVIK7KRFH51pUScZJy03VWQtsKPMO9kc9
cKZfJ5yGX5w0DxftsWhk/QybxaIWGDp4/MELzuVrlcxt8CukFKvMgxXZ+FFAJ9EP
ir+Fo+zLDIX4wTG8X5mf8wZ/O3hB8zdtSFwcZn2gpls3sIf8C9wr7iiNdUy8cMPM
Zb1tpEYKAvZWR+OCkteI6mcBs/5hDxnCNY3JzLfVEZMRu39hUv5jkZowTm2h7vwP
CnoS/Z1cIW+a06LKSxY3KtcB5pbOtvPBkykEcSUg0gF/O35mRhgg4uFyr6if1BrE
dtzGURNIMbmd7732gxY2YoI2RMV9wX8PKUQoYd61dwgyOSmN9yCw8hOjZOVEjxhy
Y9lWBND786Vzk7biBIR/Z2VgAFsSNuOITArRjtd2xgw0TzE8eUZChJohi2+p0raV
6OdfUsqqG1JX8eyfqCc8VcWuafRrsKDzMrHeCJ6op8GR22HEsDl6S0NIjRUBKfFI
NkSCP/GM+FssOLt3ydQF/HDHCO9HSWnbxWEp5WyrHhgCH8uLGkgbnFuTPmAFWd6p
WTLhUKvDIb2h7TgF2LnPIbh35bOPxnpqraLv582gUq6IRmlh+Rg2+qFmv0vkxv4F
zt3d0CvrL4Xd/x5pQJZZhdmoLez0izs5l7tojUuiwCEy4O0BQvLWQixKcdzVZ+Zq
dx1HnwcvROBwmiWJ+HBAnZ5mlPBMw1NVd5sKUnlVMN1GPjZIhR6qsFemnZpy7775
2GFhHjN9rlb0tlv63jwUAdB/wr6/b0pRy8m1A6LpuJdy6ajdvH8tdzmwcMUpwV1o
OFlG71+s8EdTqW6M4eevujfUTrK3lJH7lGqJo2TOBHkSDuHo0kD+swnkH1p6a5Fc
4nJ+knRCHUJjG+zHEPJDqgtGmZnnnXPGHdRL0uGG7r4+8Zyn2uR58cHpmsHY3uiS
uXyFCRyzGmW+0G8Il8lyD7FG+yzUrHeT5yYULff/tp6/tvujfgmXW0sX7pTXWs/v
XO1rkgVuKWIUpV3q8XTuGpk6bGai9PEHY/8SPbRt5NoREmKw3yvdyJwW2hV0hXJl
5AwzKH5Vh1AWPATOq46+Q5FP3i029W4pzk4Q9dNbPJg0wyiI+rXxXVNsnCrk+DRz
nGfkNFGGqcSjGw3LhgWLTEajoXcGzur34lPt/VsfRl84p9bJm9tH0+rc3Lmyegmo
43IqQ/4Wa/6yRXChcqPHjN5bdvCqx85soSaMXOcTEnAeFauyt/ozUQE1I19q6w0b
V/ZrcbG7hQ3ad28xPjMr1YukUMSi92vf3MkQKXww5IU1sIAbkz6g12dQqbm+0AGO
FQwLNC9CD6CCyJ1i76dvmgwjIQv6U0kgbQIqeTZDMET9PREPh1FhYky1wpD16juA
iusaYPpBkf+hkQ53QqLqwZv2e1/YVdWtULwDnTmmaJM9NjLVhsZbAKg1KENub1Ba
PzFJElldnGZAfubVimVfYExsz4SYCy/zP8HBU2tsUuoQ6EW572tUkn/8QTfrK1/g
nasfU+qhVc8b5AALGaRzq+dugpcq6mTMc/6ZNZKKzQdzZGzBk/LAH8xB4Wb56/Pg
EGHoDDJfyr7f13hwvVzFPy4BtmNQuG+M1hnbEyZRBX/6AdMDdyUjJ6Q7zmip5Z4O
lMMGeKlrQJd6FEDBLW5kT74N+5KBePrkQPZTp6A74NRVUaooYfOQvZEQ53fbzn7J
WTr051eeF9LBS/EqgCfpW+ve9c7lLNMW28PbbzM6T0GKwg5Bv6XH6KvoFMaaT9OK
c60gS7KOWY5fZ2u062IX8PCS6IJ5qsYBSKTAJK9K1ufAwjhxSCUCxSOFtkG5wj0W
M9ISs/vGrAwx/dlY8oklojKVPxvg0eKyLiRDDHuOQVeckQiaTZyKXvgb4YNVYsm6
XZ7cG2NfbGnmiCTgjsKoKK5OUMUF9qzbA2+HED0FkODVs+/s+MMCKp6Y3tVlCPSY
JTu6t4mSv0bcdAGqXeq7423M0Lf7rFXbdImWg/Z6ISI73sxGmI4yscnw39NWHweU
Z28WAbuEP1TTfN72kVLiyiVkHbZEz+O3CN0RHKh+h/LGULOIO4g7R0oxetCk+LLb
rh1UL365oUwc6YsMYEIS6JSoHUO1KYVdG1CXvyCgv4uH727EJVei352Ltv8CpVy9
hKKOwxHU2DJ3N9YoxV2GVHXrbC26dTrLeePHkRv6XkWcqIy8uuZ9zO3wuBrl27jE
eSF9O95tticJzGULRuHBsaZ4LYjZcY8ZaOxCsHYpvUoCOKTWWgBsdwDcTcyEyefv
cnjnytYjcW9PUN+SANglWDVnW5+2B7HbxAsHFtCICSjvq4isbZ75F5rmg4dHEl0s
iqxnJkibyv6wmpje2kheSsyIhWjkeuLd2CdrCMxJvLSC3aEQXLFJeGBxTdXAhQdN
mIVDS4d8ygD7dfgHtIjCKz8rj/L7V72IijSxReVNdfNLAwiUP8yFwYx0KGR6NLrU
V501/Hw5pATxGVtZ8x3rY2HQttBK/dPzRGIXkWGfj4xCrS1YqIH8iedIyFC02U7N
L/Ya2n/uD0DGzUSda80xes0h5D7dUfm+3AzuK9am7XUWRcIPXEVyeLlTVCW638zt
ESHIcXA2RlOYctoZ8F3/uL2RLK9V1TAvalxKkoy21aY+dhDAUD+Kg37teNW6u7hY
5y/BUECHzYOQdysth2HkLz6jW1P7NpIwXpko9DRWOAGHsuU5EORhHNlWoP5svqWH
deFS6BFiw2JF2XCajmMjduXj+/bk7QyvKq3CN5doJTzssYr8qR2OlNXlHA2DDhnq
aXK3VQNaKI/tHDjeFRT1S2aPo2pK9471u2sjnMAawvQVQ5tZKyuY9HB/FlU2pSlt
RkKTr7c1XSsyxNilE/XXgwWG8J0OpEAlxZSr4pjgLvNuYDFyTpCl7D8yWHdZkCR8
TKmBhzzhA6lsKTF8SJPOI1kdUzM00MtbwXfHllXJ04obdVDRchvQ9wmK+vUnPoxT
QgWr49H3TxGEzHnfz24HsYTiGYG+OJQS/ekpZlAaXb8aBm6LRC1JzwW9FgKcPcvP
XeQeyKnm4XlaimMsz0AQAKWnirMPXPUnjGQ1EWZo5/NCD6l1Of/ocS+Vcu//10X+
/2pJru+3rTa4MF8TnycGkOYQ9yt7B9CK4GlszIWKRgyl2S3myp0e9UtseMc1QP8o
4QIXk77tnu3rWEQe1HoMGuiEYDpUV7hftnIXQARGaHdvuBAXwOhiJ+LtwWN6PVeS
Uklw0X5OyH7xYMa0mB8Sn7pEvi5p+eexZ+u4m5WJAcCbgDj/lqR0Q9TbqO6ozzvO
nODW3j9dJdj1dO7gMYflo/I/NLCyIaDJy24+kTXy3g3rTepP9F0/TZ5TyGAkbxiE
caoNLWWdDjXUTvj8yCaZ8QzZeYV7PP0EKZw7akl+utnCUHAc2Ugf0sB7UA4jl0Kf
iYRoFCzX/uRj2hfw6Ig9D0JlzW9HByD3NRKXu7j0txFmBxcdlaXd0+aRNrMrYPI2
8gbm4/u7NDGU1s7+cdwx0eJTfu2yWnj/iQVPuBgFHkemLchVVfz8GRpIKgKMDSjo
qVEy2NM9q6YvNyw4WfjXS46iYBW0whY2G8jIQaidLoLtxKQqMmbW8QNk+baYRk5x
fA7yUCdVYXH62FAuBqmb+kuNsaJe/mAJZOAwxI7OldPBNdGKXUZ38bzGKNQDTI9X
Z5vd2uShVNRfEnv5lEXRYDqo2zLe9+4c9vhYrDgC7Cg/VLe60vywk6S5Pb4lWwTG
tvtcJccMDg1jo9p2jkQa+yBhbQw4ZgZ0vF7ucVtlm/lu+vmmA6Z7fMHWcfFlpU4n
t7g7Ow8YbK6gue4VG71sSIz2UoIjPAb0h1+xgTkltPekVkKTPQuGtW9xOg/aGxWb
cE24DByV+2tJYW+djJn0xr3JXIBrwkZ2aDLVPl8qLfwNLJA1ERTcpFQXijXbymyO
3ae2QW3+aWnrs/FrNpvl9u5VoM9I4zjv6pLOmw9H30daHeqgeaWrLCIvZkkbVcUs
QKgEjWRPpldb/x9C5oMB/uugD5Q2y9tlIZ9EubOhVbzZJ3bp197sq4jXnFah7sfF
I4Ic+AgpDheMN/5JHU1JGNfaWzfOiSO6rjeAY+igtvo/pfBxistrj1MUokGKkBcZ
0d5zgtfKTmkAPW+0xYqYdk0K5fPwVfdj3S348IUvGmtyGuowSt4X2YoKDka3uuap
6vodSsIed73bBcNWclwwFdOqb2eZRI1rvW0zxQz0R6/oKevj/9w4PWL3R3HKjye+
6Xl/P21zmj70ACvmAwyxoApzV4i41n5t5fq4efnSOJ9Uw7T/UDoVLB5Qz9Cd9qCy
jegs7jONZwggHZL3ouuaPb1pkSQdwfTo7bRvxF5dqsH9BQxV9DbOew2yOZZze8vx
7+KrTWoDkmqL+JXav5dum3EU5PgcOVzXY4N77y6rD6UENV692I7fuA1XhgbE34Vy
OmNf518vPpQbcRNVyGaieCAAVvdlHNUvkQFQPJXGfMA7Sl8IzQThHXgr6E46e0mf
2ivf35iJZUltzid7z22Iwk2h2GTXItIewEnGXdTaxsyq77HpHZOKhlFUzjioLMR7
3aaoCTJHwPkd7OVB9rXxxJnfUGi95SsdDJciAFPTmjX7K+gJ5HB9st1fMMqdvj90
1FvkJvuyx9BlF5ocapwprRVH2mDtqt543CpBhRn9zCyfNpGsR5MPje3p/K4DYzni
Ky41ZEARXavUw9NvUGC26IuxBERBNnAOp8f7bENOH5sFvUz+pWGMo181HuauX1oE
GKnU5if6J2A/bdDvufMyqZvywjpqTTxhj3gmFvBN21zd8gHBffG5IZCUvG0a7ga7
p1bzSAiYG3QWYmbZU8jEAokNnoG1ggCNBpAmr6nFJFvXKhN/iHHbrFp9u+S8H2OA
APiJwtbwO2taAa1Pm4mliZp115ubQvCEyDsxZ3UqlTb3yt+GP5ANtJ+hEH/XScxN
qYZEsMxc0yxvlMI2mBI2Y7PRD0uST+u55uOIHHsAvXrhuXRZDLw7+nSq5Ip70+9Y
l0mvDeQ+DI0NlsXLi4HGBO1Ll3Rm1hLEZk0ofhN2ksBoGzL7sbZrBNHg36AKzP7T
zv//Wqa1z5p93u3lSqUqNbfVpfJCUkZaZZQ1sThOZLu+IfVpnCUREgHcIWSH4TRp
zu70+0iTi1RUqyhdk9fFrxqk22/LivgiHcI42AWpQ/sy+OPCxUOKHikR4MxvAtY0
B7ZKmOfiSr4Q7DYjvVJz1psUHX3l5g9VSq/uFDLl5vIoPogQWkdB5+rRWqm1f1jg
SeQjb2/IaB3yPFV46zSrI8w8pSDXJ56/u9e2oEHVxufNHhC6+Uo/VBufS1QTEckI
h2eUQLdvoQPn7igF1KSULVplP1ZjZYUhr+l7VChNXQzS+jFYgLk2KSL5GXfXtjoK
pbz+K4OhgEiYHXpQfRd9XSkzsm8sX44VeKKFFql/gNNdcx2guH0JgN+ikpWRQLRG
jKD4aYqcijMYMNLsXm6Ck51BAQP5aJsHmtZtgH+jgU+C9KDBBFVbLEoDQW9hpOl2
yWjRqAlqcHLC0PVSIpzA5quVGEwl5EgjbsJstlyYJiRVYdzbawDkm9VsQBoonGSe
Xq7aVQex6lRuSdHkCdUM7uPi22RlxXXr2JFILwuKw/+qnUmry/OOF75zjsuPTf8Y
ewmFb2KH5aBSx+S+ail9Tuprk4AnhsApjPV/H4DhGawYujJ7eNYd9Xj9KYx5hyV/
JaUHMWkZXN2nAfj8v+TnTxD+ZyEjnW9eEg/wJ6pQxFuDfb0uVgfzfsjA2oDKBXYu
1W9/feW0VCHGLwf13HiQvBfWYivBOIMpDAQoMxxK6AL/AmCBFaT3LpyMNFXsvy5B
p1DERwGtrg3vg1l5SP1mfeBdGjcorbgu0ieFxWYuxAErJPG1Cs2gtHIyxiRpBQOD
An8u8bUn0A5OwNEZzvAMHMiANhQNLCSuS484KrJX5zTi821KffBOLMEQcEuBOveK
jxTdG/a2Z57/5IM27Q5+HXBVxDwEjqZF4/0BscfmMPq7TJS3bKWuLVwpneU/gacK
PGsAF0rPwvevVkWs2OuTts7w01bRbdp+8uokg15Fpg4a2gtwLij/E3e6AEwpsW4O
JKkPpDhf6DWIMcwi/g46lWgu0xmt7ZZbvWSZ1XYXCfZMOnAbByZdKB4FP59GKq/z
CQqW0Pf8ho6rR3BpI1r9UgkAusF7xRDylWhkl7qautLkieuindHiAN6nHAbOx0bd
DSAIRZsimMu8Pvg6H4cpXwY3aIZX81yVGZb2KRemBkP74CWUoVWduwcFHYkE1Aca
YbhIrBnXiaa0a13FaMW8JCI3bSrrj13K/3yyFuMdWTdeR1Q+De6o5FKYYlGo+1WQ
lXZyui0Cs0j49H/RrWonDr8OVMvCXKn5l2JkD3Jh9MQ1Hczg9ZSrAq6lmB4Sp+YR
FvxH4oJtEfaIHnN/YacqneW9TB/kwuc+YCUNelKsIxCFNdyW/vJXCFYXWx5IrlCU
Ruo4FvPLx2AG76gLCVk00mr+1CJ5Ze9jRSdjw2A+t1dq1bkzXxwM5gOWarSP7b/x
o3a4i44hhLH+J3lyrowO9ShqJb6B8oOd8iVCuJw+eIxtkGPrBBXZKGewRyZTfetG
9ikWURrbkX/k4XeWQ1v+WWxzRJUi1lS2bbNgkf/eDLnCgd4O6z6VLKHMKd9yzb6w
yqXDCLruXwxX2OnoGPhdIx/iPAaG7SUfwPK2AUKW59Z9Dqq6YBsW5YjiQp+szd2t
NdhqzFqvtUVtvt23uExc8cw+xS9Lvi6XdoJxWHMHcTnHCg4c/UJrvO63X9ANuQLT
4AOGNA6N1ofWyZcP1CIsUtEdMWl/3veb1aqLlCLbYBKZqlzaZvtvCmRJ0Kygtbzh
oJ1Q0R1bXEP7ZobZJzPNDNSUZmh1poG/OY3UmNQT8BpbEFnHlHa4ae1KP4FXhsIT
58DnBrL/ACMwBibDBBvpLDjB36JLDbYnQJ6MmMCUC5WuBw8nNtv8dgfw6NI0fS1f
IyW1mnesktvu+5X8LmDIn6KyF9wLrSpfV9cbqEBnqQAan5E7BoZHmrnMM+qGpNyT
0lyQasjKwSlMet/b/tG3R8AlhPLJaGPlrj+wXmoUfn6+mgE9DR+Jia4NjMAvtjAu
/Lrh73EU910mqMOJNPiAJ02g4fRm6hddTonn8TX+JZoJt4zmLyRn8ktYercRlmMN
HBuvpXSJJ9kN+lq8zmOuS9Tkytlv3Qxq/B0TpGr6QbmDWio9xlXgfaIQ+EKsuEOs
mOxNSG3aQsA/YZaBlxc/uyJpSmekVT4a4GmEtOuXkzKHeJvC3ZT5oNe56mooFNHg
RUZf9IbGTmGuTtFQmhEX7rUMHufkI+AS0ZgO9aY9EqGthlOyUuw1aFVh4dqLAa/X
8IF8vGtNxcQflkKvOUBBfZTSymUX19e8iKnDMNtM1Q92xI4N2Auf7oGM1TPcSor0
gxmz+NhlEk8kzdXyw/RH7Nn5uFGbJH1gPw2mjFYpm3leRC0kaHAJf3cVKqaOPuFm
smfAhFfoThXGOjxAJpkJmd5LSLizyBys5djqQuVXGECbzUOA6MXw2rdTFH9IwGiu
yvjKtW64/gnqnxOrYDZHjosJlbD/9HWvq4wZyTVqdftJBP1Ob17y1iSe1WMk15j/
k0tpBunl+Pmf4UI9LqqM2v+rHuxPsHff2HvYcEFz5YfQ8wBoRDH/7+FyGwP6e4rC
LHp5iJzDv2sR6ZjbKQ7zc1xSU21eZ4rm3S2eD14VRff5LIQbWAoSGt938IAxW3Bp
n0GA2t9uzyGXUI1JCZDSSjyw//rZKhV3J4jMggtPt1WlAwDZFxeucUkaH7CKk63C
vy1+qYUcmEOObtL7dQ3VJZA3iBlwBF1VsyfD00BqLciDJDzms1MzCVKMWG5A9uNz
6sfjqjBPxj1EexZU8+ptyUt99RaAJ4fpheWdpDCtoLzAAcZzRiR7qmGcKyC16xMq
UQuAT6OTJxZdzcrgH2I+BR3qtFLZHWAU5EnP9EjIpysBzeuAt/9V/LvKZ9YFxdPN
XKgW9ZdtXz6dwFy8IiIveKidJlkEOIBthcdiqraycbnembs9uzC7dCgOqBJLi0LD
+371hqGbwzG672y/hwRH9hR/6DA/Y1ROezU5YBrpylyzjrETIA/lz6XfyO7+oPUL
hiVHa/ZV9kgbWZ+p3YK2CZlx7c0IQ7GJfZQGJ7HiToO38tQhltbgz0pa5v7xX393
qrquQcHKEI53+y14XoTi3k8+dOXKd8ofo/yEFtC7shzm7bYoBZsZOyA6ne+LkxL5
NesnvX0f4ci/uL66IYanrxLRZ9FlIpF9Xwuo5+WhxurxHHy2VQo5vf0lyDHkByIj
r9yJqpd7J15Q3PuDHry7W0ZPx/8uPTgEiN+BT4UYqiV/oBrcUrtaYFjAOFj3OOxm
Pvp2nrulBdj6SJVoAE+wBU5aOjPHhRNIt3MVMa5CLWh6Q2oVBs0vR9YZVelrCaJi
FovMs4pOJfvJGLkijQmK7f3j7+JoOFDGf5xfBDNnXWjYtIRqP07Sn8sSWtSm3nv0
W6sJYbMQT1f+RLtx3TPa1wzKcRHHu9HLJqo6x0z0DPL60TVDo6/cVxtIOjllPS/y
SQpELAkGu/o6ANU33SCnJ9px++2JbEZMq/Cu6zhFfMH4LWDPbQF5MJbBrx7NXjNA
G5toy6JP4hdu4x+vEWVoatn/Q489jILMeDXEG5k1NYgsClIdAioBa1DLIwMzDuMN
V53Me6/yppzt00KJIA86934f+vTMDWybXCdqg4KnovOjlY8msZJe9VewzXJlQOhy
g11sA6N8InTq7tDudHkdiOadSMKwN9bRN6Hko7fx7CdJ3/HKTGjD76337C9Cko3S
v23TrPkrxNsJN1qMl+RcmmdkLWlTyQNQF4NCPUAKDWPOdxAbhlHsQ/0XCylxBR3Q
RqvEWARomXbcSpL6CZfbFSSYmseXYxoBoIXtsTt0ngp4W648+ph4ogSXOLZ5Qkc0
45cdt6SdK5emPIA9RkYdc/Ibs4hlQXHqVIUZvp9w0sM8N2lMUF2lDoBu7h2bCJNd
jtSuTyZw9SJcklKVlu884S4tUsaWzs64Gy556Q9xtoVPAozg2VP6AlcFtUcuywv4
qMyJmhxvqhrYDeqYm2yoHzzrL6wojJXI9SBEFV88RCaJq8LqDxOTsMoMzsL5TGju
cBJbFj4AuBeOj/cboy5Qe69dSC5AHtn3K7NeGVFGPhyvVNn/fqH4YVbYOF6T7WTq
wg/iBbr22IrVr6DneMM5LDYQ+gToQwIL96dO4DWjCE/u43GAYDTM+cG4PT+IG087
QkyCbsTU3/lSEiZ9wxQ2wA2UPRrv1BJPVcDD8tzlcWRm83sdpHbdvnlokd/FMQv6
iOXzUQPBFwbGnF3aCeC2DgLPeld6Nc+M8X7x8riejxb63mnocrED6PB6ClwOeahQ
lvvpMKlKeUmNdIGJjSKY++jsHJx1HcvIITUEaeIcjBH6Nf5AMIX27Zk0OnFfTp+D
ZWoyN3JcQZTjr/OK2y8pR9ZpkWWaBHbPPhAnL7igw0VMAhnThYcHNtP0CH6zoLQh
n8itM5VsrSbyaKx+vUcEpPCS+jopXYduvPvqxoa94yHyp3x/4cN8oUto0P5ImTz7
z0zvE0nZLedggfItNuOnn4GcdL+4Zh4LOmkjwJCdOCWstNEpCtWzDXvYo8cvLiCc
2hBWvaGyGM58bbiYKy732oZW2k9+UmNNlOxNMlPD/CICDC6pHAt4aqlTBFuHTXRs
Yza3AYi7wpsHlyHPLKiwMsKBlYi5o8GWjV4tEGIvId4YAYdcZh9Oy4zD5dtsuFje
9VArZ2/9zjyHneeQjRgL1d+XYdGNE52ah3OMNplDR2gZOLz4FOOPYGN84x0sNOmX
/NwiJKgUEw8Meam58Chr8vvHoizDqTLml6MuprkRX9kME37aKsKdjekQPhlxwgW8
OhArdSTYpmYXRuw5V2o6eOequkGNPNRuYrrtbfGAsy8hXfO7jqsk5TuYIG/59yvP
4I9F9EFDCyw7pNlyM4Y5WvbKVY+LyvwAxq0fbjonr2lvZRF/huXyfE4npyqYBPHv
0/nQv3h/M2/EwK4y3iv66asCLbnhmZ/Wq4PLzC32kD93OLpOYKJ8Ua7kxxTW8EMz
nB7nys3JO7h5OyrM+aOscbgx4bzIJEbK9qG4OGGC2HOhddMsBKecOF9leaz9RXI2
dWGwbhpCfHQQ5j/8Zvrhy3VCgkrRJVykE8dth2N6ZPVPClZA63bv8+/qQtR28Mry
UDokB+xS9lLcXPtFtAPCPA/Tw4TcsKzHsoOQYGyMSk7BgkJnjZa7us1GxvPM4mS4
M4sxxnWW9UrZdsJxeANZij0P7UjKHp6kosexb2VvCqEFyQFWHIhkChzVuBJvV4oX
6ZwWt7nQmC0EvRugOkdduYXWYCPP0azg1kpEin1f0itzJgzTZkuCPmy2YGGhy6nh
B99NIFGXRIg988L0twmDRfuVlu5rfs9ny0fkTFRY4izDIk0ibrWNQ0OisbU32FDa
GcyRJGXocXfdk5aiL3PjPV4DqPn6OztktQQQxvCqKlcCW1bOM2sPnQ2ZB5H8saU5
SvN286uu0BOYLJ3NHRdkpNKQfjXY45NFiL6IhD7RCqipgIYQykIWqJGvVQ1T4qEQ
tzSGjdIexoVh05byuqwMHCWZ4SRST1vJCIOEcLReT2XIlUG6ILWiZSAUJp2cOKdZ
53mrEnhDfWwok/ecO5pmWz4/F3YMw+Su4x8/NzJpFLV3IUoYvbqNzPm1hZmKzY51
A9R9txRQIOAJzIbmlcQZ/rmzw6NnPzTe1GJYac3MDBcy+5kBcvxhRXx93bkBrgVZ
83k0w47Wo85dEYbHyumr1xmZ622ddqaFj/a4uLvNgGDPxXxfwKFI+HtMC0chDdR/
Zy8zicENc3d1re1FY9skW6P6YAUcWtqq7vfmS4SJxjoH5MdNRBoD13vjz2zxerhd
9AjnE4BfBsOehM+qcvVmztE8/Z6GklvuzLw7CLEdY18QTcB/IijAV5QsTx2X/JMe
CzEGBECzH4GpH7ESqYjygqWWmmyMS5K3Dwgy6wRaBaRqGtUfl/xXVUmqjr6BIV39
Z3ISmQJLev51//2FlDQ/w6DlZHMtIg3yPMoY3eu/iyxOLcrDvR72FFwzg08jigi5
Yj0iH+mHWTh1uNmPCrdPuomecis3/TO8aV9LQdK2iQKtIm4Ted4kd4Mhk0GZ3k3T
3Ra0YKVjIn0ob2x2wx/VvSrLzYabbKzoxygsr0ALY39tHk3gCyMzk5VF4IiOHRzK
qRPTHe6/BZa+aE+s7VLtJEzvqVmWDFcOxLRFiEAZi7oq2RnhVy5NEqgBQtQeq8J5
x7DDhAPcQ41bkoT6Bh0yyvHWgjsx9er+mOG18EWmDwgiyCnjkBQb1orIKDwSbZU2
AGv0gQ5WNgtRfMJv4A1WItS9+5H6u6IqlH410keHu3qxvwsDq+9YppRw/sn6EDNl
wKbVdfldl54vKqi7XsmNpMZuFrVP9Wb1ZwfYSn0AbMYoPaUdcMdqn9H9KgUsYSog
3PEONxTluMnAuqsoegZ9dp91XtrHGZ8Jlf8CEvmrYVUAsdmwJZ+vFjKUH2nrOFi+
uMTV3aMS+TJqlciP6+rSNkJ4dZgStnQvlhEZyl5sHUYl4A3lqyRm/bhGQHZ/nimk
1FMdu+R1HNTycg3Ye2YMaAdP37uQajzK+GIGqMk+1P1Lq+GgeHtus8YMQ+hZFU93
pKIfjYKpOCTmu9yBbVcWJpDbWtAbmAt/a7V3xaz9nWISWqpGuZqsErr1SqK3oiIp
BWPQcOFzkkCllxFO5Ae3dbt0ddZCZs2/hRCXtlh2raaBZOue19uqoyAjcXYwnwMb
CEhfGSYZhPOEMWdWw2Y4ln5pD60Ni0lCB916YzfKWGQ7jn1ZDFFt89U9sNL2QS1R
rj3bkDR7O4OQAL6W9XWOeXDx6JVyKwhhWXitO28/vDbZdKqzZnbihb56O3DoIamn
qdKOQcZdB1wNMJCtipy0srHb3biVc9YmdHhOdGel4k9iwQneg2si5O8gaMnUasxE
rjh/PKqoqkR5a72xK9/sQ2kQlk1Lw10YodaU8QmI6617P6Fx3S2LeL/bP5NN70T4
ycl8Tg6hKiXGx5IWzY1+RYhi6RidriQ2r7m6jJobg1nrIr/xyoFr6wbAtVc73b5x
U+hdUxK69qu/PimjnobTDITQ2WvvA5Gi/Ghxu65jY9TSyodjJfnxXCJyKm3wMqrt
kVO0vehBdDvuf7D69kMBQo0De56+afghJjWUZDQqe7u6KdeqrI0VR243aJq/Ta5M
X4MEBTcqQgCRwOiOK6l4DVzXJRnQQU7KJbkXWaISahGdmFxuCCnF/Z2d/yo1PIWD
ls+pAvsm33srOPz5iioYxMBTlXpPJzaHXdvVkQjxy1tArgdMg4bg3RZyga35btHk
nyMEGGPM83XU2KEqlnAutNyThI+79Iat/KVgBhpkgrKYRvEeo5giXQjQfPI21d01
iD1VLoFqoGYVjD/AwZStJI3xZWsx5gsgXYQb7QP2GG4NtlAFwYApl8bVymdPHJOc
qmmJQps1r5CEBRnxhEp+J49AI0wCv4kuIq4x7B2Ig8RxR7VOMTGwjxmbR41ZlS28
ioC+U/qg26vSU+E4vr0r5g66oh4My+dmbCURAV4Jun8Cb2+Qy7Svj6oilz9jMhpX
P5MF6YgvwnOX/qKkuW0g3ctchpAnHp9L5ZOXVST7Ent+MvC2Rybq5l8K08XySsae
w/kutgnCl2TfA7dTosojRUhE0923Hkfoo/bA2zPLw1E1tEhwmQ6zChwc0oim3/r+
fRbs9qhq4DXMrTf87KdAJw+BRxdHCQrs+Q9ekD7dnmrSJKsijkGPCYCnsFeU5ok8
3fnmNXjp4XYLJIpiilWzZSgiLcNjVVJsKrNXvVS4Thneft+3kn+SJDIFYoHzLPUJ
amPBYebIG+FG6K9TD1WPxbfWbs81xXqegKD+xrZ1HFxKmtUg4+0X4rUCQXxdcFog
3I0Ljs1AwL9E1YZrnintE4/a/vCEJ93kw63LCndiHOY5zoKpejoNFld+vADxzTRT
ZQpidziRx+1eYLX2KL/Y24rgEPBk+U75wPUviNRNj9fCMLFKSgsmyguxDncZWtti
v2Bt/sWpIURDrPCCMqbiePngT1AkrDhMitxlY79W/4yFbn9X10LMB/zP7rg+HZcD
WR+onppIg5jtg8CxX/reuHNsuROm2QhK9HFjL2Mz5SlEad/nAZYsejyDeOWCclY1
6uBrM+InX8KZlDEALxBPxK+90qFeT+Dpz73owg44WLfZuMR4hw5lBFeY1Ledis+0
+/Wj/XWrO+E6ZJJbUuGG7P2NGSGDhUOHTWRDb/9qO7lTKcexM6G6u+3S1AVphoz5
6c9kKEe0+drAEM5wg4BxWjXscQLxDaEjM5hsXdzRKb1hVCye9wFr4o9NCiTWqV6v
RlGgMv+4+2sIgARUrYnL5nTyM4N9gEULpJ3im60LIBN5DGhG0UhAJsbleuoH2Mus
bHAAiNpN24vV1iaB9/73F1HaqgHIHfZ7tManpL+2j8PbQeNEA/CrWvmoK53CsRbP
WmWoeNOPczN7/cmZj5r/jcqrbeNGSq2u95TM2pdnHheUHP8BsP9vomtECYKXcZqz
fw/4uau/xZKFaFkq/WuiGGcTtpew7gj6U26vAPiH2cPcQ1xy0m/VxfZ9OxlgrOvP
jonOI2zBtkejH2r9Y3/9TOwGQCeODvr1STjofhP7gEqBEa51D9W+3ubk9MnwWfej
BnVz868OzCVAK7dHm6oG9RKJ6E87bGUiHLYgVdLuIYRGtWiJ+qkgBSNDizO0DghX
J+dubK31PAqOjiZ3qGPyBmh7jcFl+YfKFnJRxSngZUbpKCwwx69/DxpaKoRYFJcq
kY804jWbynVKtIGVzpR4s3q0tqoUh1jS94nDJm9Ahp5fGaa844kuT312jyUV9mgD
W+STJSfGSbTrBABdhPXPm1LFpfPU5BY+DupX9DINhue0tTWdAe4NVgrLzeWsQavV
XiYbleyoptNB13VHOtK33ghFGwZJeGeeEQ4TB30+f6L0tHYKlTdgVh5+BHOCwyt6
eJHNfwmpKwJOv7lbcZm8+hte+/kh8+ZLU5+TLiJMBdakYGxcmxdKqigteeyMKZ4I
6gZ2mCpZr1lOPwoEcaBdT/5+R+u3BaPtSFOBdIcspZ3GTAIwuQmEplf77CX7RMRt
GF26Q5WUh3ejHvoiDzMwxicwKrk8eBrTvRubb6MriD/QAjYAz2uOs4kOlI4d9SNW
7jIyMUoflqpGDSTR3r61DZu3IEvyrQozotN9zZyx/bVKNDX+MkCvpTN2LBQ6sPzh
LKZo1Je5GqaXLhG7hBqnuVj/xu0v2Q5IKCKE3XIJ30S+Z6NwXmMYN5uyGK8Q/2U8
hyJx0zTbPuodXqXabWQCqVZVEmnOoZvt0SmkQ1/0iwYDsHZtf+v+oq+x8EJiqOeH
J1ofl1W06ZtMia+jMPMe8yKLdF5Pi9jZxSejUetPzdFNFjgh7T4q9QnMoySYX8RK
+XySj8crXU3NftlUwB1QDJ+qgesMastBkRpxevm2sFzMwbALKCcyujjiJCPz9LVN
KR5SoNwAP2m7otfdO6GnLHvaZqNlqx3hfNkfqui0SzkwhnoJ1z5pQTbuKGrq3bHi
fUulLSWIwMsFa21mTYwI3FUhPFn9jjNe5WH847N9q+sD++XO7gTHoVgL89Bgszgd
nQ5cySlYgM6V7iJvVspMtJ3utiXC35L+FplnUe7Sb3b3okAoF/gIqKRbFRqeAm1H
pCLJoStXcQ7OALq5WIxYP5enjmf1tZtof/wPff2CrLavH6mdGakv43IIBkcFWIpB
UJfmDQsOpZK+NYZ+OMlYquAKARqLeN+gxqyctG7Ph4pXsN7ICrWmHLoQ0wAazTre
oAupp7r37Tt4JxgPlDN9gtg/Zx+NbVtMuNH9Wh7RbMrY+NNgtC7ywrLwCcKblu2z
Yv3+BBu9s8LXnVPZTyYaSOozOyRWRJGvmj5Cm2QwFnIxN+emCRNdf+IpOhG4cESs
6UGP07dFFkm4WV++//3vBIEVQV0iK1LKToKwOUZDWWrhEqNv77k1A6Vohvcb6YzN
gDAeDpahPBmTOStdz+SK3wXO4bW5DY4rNLo+WYUw+YUj00s5GdgRi2raQJdX8JiR
W8D1JVXLmbF2KTYr3lFJDDC3m+Mi5TBWCA7VjRXgO720qoyc59K0g7nsadG/dJwo
37EGFl6NAVN4JXBYnIIHfagw7TrX/krNNWrxITi8VCkeKs4NvmtXXqY16GduYkxc
0MsH7nyRpb83gkzVYSE7tjLq2dWTKRtF6SVVKJwpkSHtaWd0/BvwSJQRqI1+dcoc
+A7XkeElP97BbIw6O9B9OcjIx00ZipXgi+dTmsefIHfYvqjJX4bXKB5Ra4x1r6f1
T03XpWHIaaC1g4F9zP9IEWGBbP0K66ezCYTjb2n7665RxAluAi8HPE9tThVIhg1p
Q0fX/pprMUH1W8Asb5PBjD6H1K8zn6qS5HB22ND52h6pbNT1KsMki4ewNVa+XKZr
FGpw0hknqoxVrzdEcN1uISDFlYZuiIuC162KwoktDUwPiSuqe6xHwyVyuICJjlDR
shSdZicZz3etxhlIMomHCCWe1/OExMs/OLU1kT2w9127rEBtHUx5clL+2XIZzwWX
T6VDZpLJA6jEBr+3hzKXSbhrI8gQKtoEgdFbLp0OF2JOwqWxzjasE9fwvYn8piF1
2OhqdEvYxrtixYoK2qp44NCE9K829zdVX8mqOIhhPGH+hx80j/RGj6BLOya1gx/o
Lk2DIV2U1ZBgjZcNo8jvzJ9ItT+ZFXgyYsMHxbeSuaVqHSEULauLyefFHoKBQbUM
wRdkW4JYrlcPzdJRf1zC06DkC0G23SAy977jAPPsJeLH/1qCF1x87VXqBcKzJ+8N
VVboGrXtfwX4BqakCeeejbpvzHcOa/pTqkocaldI4s/NUoUBp+zP7+EPNhzHAg9m
1Fnyzo4yHLwxf1ePbqA2kyPdxFzts1ZDqyf4+erHvwYAPY0pmlTAnRWAMuVAhV3O
Ivjw+FukM5J5QjQbB9zzYihOm8i3sPrZy/INwFZokYQWEXfu4csWRs6xjulqcRwT
jO4tv+WKEK1uB6LRXr4eFDOrUyUMc59e9WLZ2ubFnpDVDxaFxaOPuc2vtedHBidN
cPvQnKHdNYnDPUMSiV5Wa+a4VzNo/kpnvzJQRry/h+f7DTYAK/8T9wX8MDSaljY+
dQZgVXVth6iK3nBxtFotWKf+7GF64cRMPd7QA42D6+MAMzPwn54QpMXT3M3c3V8T
1i9H8SCigB3RaqEdg2ZOgHiGXzb7k0H5lG8+hGXZS69qdvfOfRPIitnG7dEEzBxV
+XV3E2suLIWdVw2lGKaAAytVx1JZxs1ZP3Fx0VGZAOuORaeOCrpTt7k3ok9Aqdhx
8iY1qQVUgyedIyoMhEvkkWqUaZJjA5H4FY359ueVEc1Z02kaKjE3k+wwyr1U5zbE
ACjViagFNNUNEkth6VlYKwXfHsnvfWVFUhKjquIu6I3EY8GKgejxckb0jYh6wvvv
5OmNtxU0x80DAOEGUvI0ODEykioe6UeO+jHKtRepGoJllBs0pomj8sJHkpAzQfbG
Bv10ftFK6k+/umJsfH/Wq5D+n6GpFMUYM+4EQbfgY4ehrhoYaDfdc5u0zdiHvw02
89vH2N3E4kxL9NxO6ZzYlkoZk2YZDPf668CLbzbTuvShOarcnajLhRugSWY9YOLC
IJ0XJ1AIr/0J8QWgrZ8FCz/0LlMPFC29BviGlYZMyp1glmzpxOr/CeRgNYyuXsXB
dQSoPId5upOnOjJI6lxU22jVMSw7su40bpx+dwAgC8igCd2uKI1QIMtYgD2REQT/
o1IpBuORXnzVy4KG9C8gHC1MLzxXi+PCmr+N4ICax7QGcOUujf4b5yiVM6i7ghCU
1Hi2fhBwAhswt2mxwR3mUhnENF0ZLKc0L1u6n2W3n241LNqp7y/SU3z9VKzQwnBt
AfCCWo/YkTAkZHTGa6elHaNOE9GULV7Ivhk7ku2b5aFg51H35kmyIXprXEL2csv7
FGLd+gOaX8rgRLRUf/owc6PHZyNauQtYiaryPCoc3FZ4/c6Y3s7cnyIhIhldccA/
r+3GGhjRZg1VNXPogoGh/mqFnysVKe4h7v2wrFIWQXhVF5r7vF8LmU6mZdi+jJdV
gtZ8PAZcUEOLG4NZxDbz0D/C5Jva2a7yjB89j7Ux8DdPXIM3BdUuvzrNMhWCZcJr
EkG0XFKxVOjgrb9YoizJ0bHWJU7zFMRi6qk0vJZvUO3514WEc3jYlOT1uZXqb3WX
LaM0ofMd4w6Cev3y7nF2ZYQgTyspxmRXD31pTU2yLD99GP6mHVCJrnq9nksd6CeY
VdMauQckyZAtfyHJSWAR+eijUuwSh4VjFVzcGUBMtGC/RqHs3+Nb84i8A+C9nJoa
gJuGk8vbvxww7Ra1kPArU2sm7XaL3cNsFJrXast84a0lFxYFZUZzjWKYiOJ3wB/j
/OLC+Lt+naM8DFIJiPAkqHnFVQg5oUqt0gs80PpSfKPaYUEyHIvPfpbqxLOOTrBt
bVPIIC0Fre+XLjFQVHpaYe1NFuwcLXOlPydLe7KRsKgpX/mRUWFD8A9WRThsFoRT
HvI2tnDtf25zoECA/9rTOuW13+f0W3vd0WV28c6NUGaFTPJd4+JjQjTHsuGHuAh1
DmlgQXBsHYMmAbi839RMfwr4hVGGhSHQgFu+fbiZAsF6aRnaCyIW+cQRcxJjItBv
5aNgEcEiKu/5kMuJOTdDPv6uTEH/MlXSlqdB0/jc3rH4ki/HMd14kaH8qSrcxBF/
mNZOYt0+gf7lTUGh5ykliU5uft7/MFAaMATbG3zqEiytsNnVo3XplmVLLys12oFS
uZYYE0OA9l4j3gZ/9WHYVvIPfpj3+1FEFiPnoF7g+rSnJvYmshdd3vh/KQPvngFD
eIzShVgfCET9d+t9fjRSx8aN0JBNnNJSMqVKW06Zvy5ZT7D1P1DxJOvvi5SvMHyz
r9jX1GRmo9kcR+fcBaaKBLMSvtOnKbljVsf8ohYKrhITiD+auVZ6vxjpVNTZZJRw
f8uqKyu2QeqR/fNUU6dzoEeZLlLZfgznyRudSQOoJDr9Q0lJ5sOWa0VjRKBQM3ar
8386xlAKcj+mT3Ku4wfMqP9Dh1rvkmAtf0kiSKM7Orr7K4UUNCu0bks/DZLpNDEz
ZWRWr9bChyQbkYopGJIsdqEfsn2VDgMpGJUgGQlWzbhSueTrZSNSFh8zRTIYucBY
US0KF03A8fAJfvC8HhJIQoRXD/8gjMWs/4Tz//wxWZwTRUAtu1lqcbZspxSvwsrs
K2qStZZ/2KsU9MrWYJygrEdlyd2ADgYMHujQwD07+SLQYakM4IQSAWFthZcsQPtS
j4VcbvO2+LoHaXpKPfnRP8tQ9mcH0JX08Wj8ys4lG2Y8qrU25K6gruMD/6rZ/ho1
zyAAsj4oxHVkD08CXrJXxLOoqY3jx0QjLEfC5w7eUfwE7jZ7wEpEDu47dYm4Q2ii
OcEr9PRecJsaF+Rbu2dhzaCP1sAZ4xmvqN/lbEp6pNK87KZ2OIdJ5vVftObOdRz8
ghiWp/X89WJMdqwXB9XZqgL/SKzGA6bGJGVTxh8KKTFv7rRBiWnFHj5Ecnrjm/NR
JOevYKA2sdKlG77CL0+frjrEHMtuiJn/gcQm2p6HSRERNoTAjO3Xwlj46wLanw8d
lgSMnXrL6BNxEr9MqrGyksrQSfjtw/ugOpxG032m8KkYvE1Ik1D+bEBna4O1vaql
2Y95kzZ7OhCoGKeWm8jhw4SLRy1FQyR5epvciFFmKpv9qawoBsbWihySggHolDU0
e8VjOvaoz/gJ6HBg9B7mB8YufkFQd8rzK4jzk7SF0PR/tziLXpgn7d56z5ltlXZA
Zm01dSm2Xwmg8La1Ozw0Alh0FPlseCb4HQwtjPwJRt4CGptSc5wC8wLZVJ/fXSM4
U6TIvWd7EVc1pBxF1aE2BEz3ksWnolMzxv2rXnJ5SzZtEPFXpMXG0Kms9xY/B9Ht
J8tGt8hGuG8bHumbL/leu9dL44htexA4XM0T/SAq+7Ezxu8a52AM/kJtdeqXHdFG
nHnkybYCHo7a0L2l9rJg6GUoOtHKmKSopKB/eW3g9np9Jn6iqi26xy2Lp4zz/uhh
//JR6HK37MXZ+yIoKnSTmlz+mr2VXBesdHaTuBGQt2bVL9UsGd4dhwGGpHjjIpn9
3h1VvHMVvIm/781RSvrHomZUtkAlIw7+1XvpY6YJ0TWPyBkG5+w/5QVA+FFMiILN
Y0xQOfzVbfPqFTbe9qpamBeLCh9HXlw+3dC5hNu0opiOoyDUzdnw9CMMPerqi/Ah
vlZbM7HTdAV8R5M3VT2U1Z8FCTgnZhcGK2kNHo00/xMv+woJRolno8wK85c7nVec
YkDP4oRWotWHS5fFEJ6Xv3ua5VTPyMsVA+zsOytHcf3l+gRh+j8gNIe5552Uodlf
uSa2Vljvb6kgZiE0lfQcZcm0bVngLAZBfdgDM3+a/1udke/y7QbaISIQx2m0kaEV
fhm2yGaVPeWzICOM0/O4yXvoKmOpo+SDuuJykMo0Fe1llHywBbjWcgA59sJ5nwle
RpCConUzVVaUeMBLqR4zWHCxwGpwKaZRGdCnvHkRam8h3YES+k3eUjzxuVkNqwPM
34jyJf7KVXSVsRY1czGiFIW/sPj/b+/CYEBBBhJNyDSrxFUE0RfAumoTvlqLkPC7
ORVR9474rj8pPA+7//okClK2Va8GjQtUOAkuW1gIp4SXJLEW+QS0+ZhQBZ34GFkb
/iWP1yRO3jgQhNisHsw+zMHmDWJLEn0smyTkPhx1zANOXW/0oBdWnQNqGqj94oRE
oZ9P04bK51RFAYd+qgpsPtzekYzt9UxJ+gHmPVv0LXGPvQgsNfms4xtGuOHZvH2p
RY7sLbwbICJg1cz4Fyn4coHJcw3alOOx1iOlSQUwdj5hINBmFGuTqsdNh1GEfU6z
N9tgaAan2QA7TLSg0EZv4w4oZhSy0aQz1ZF0hKNFAP1bLeEYHxNu0D7sWxYCCmCi
+AQ4wcXqa4+aVV6XPKEhH8rOKLqruZZP5R6lwdH+XBvjALdNW1+4jk2FdnOWvwjP
Ib1LezuSsYr5rv2j+DCEw/GB1ljjGvn+deU8OmPN+Amt5/MAmYmVvMFa4K5aTP88
uSsVg8lLz8v3tZOXm5smrg0GI21Js0/2LCY9RXxU9HG/nztpCXhFB7hdf4JgfIaf
GQ+0jfHNdMegVDO5N6CudbNmlHZ+T+Xnp0FzIY4OIkweL4hcQ7VkttkjLxSRikx4
sY2Ou3MCyjpTNIzAbsRLXRSoRxhpeRUyc2qEmI3dvOxp48SNWsbjV0kk6fCZ0Fc4
h3mAAQjWk4w+GexyFZ6ookizZD1O+pn4gurecHGAmdMXeZBg+1dk3UJb7Hx3nmYl
CDI0gbM3tsSR0+1qkvmZ8H4pQsZRE6637ZwWa9eDwmOrknp+5/NR2GDqsciUUvEr
UpAv0eYEpPDHFoLON4rRfUm4XCaiqPPPZ/CRRnm06JnUo8OJlmTZQw32dDm+a1Wj
hB5XptABz8LTC/qWpkfGG4zow6oZgs2/8/5unZ2LzuErKCiftVkWTLnlB7zAu5Po
JBfqfAox/Anuu3pXammJ7Z0Se3STUY6q5wQi6h0NWTSlzb6wi7V13nu+oxX09HFW
uGgMwCVMhkjtZCSjyPp49JvabqbMRBoIS/ZR/IKO71A+EcV5ZGhNcrx5DQreSxGq
B+w904o6JSSW/I80wwJkijgWnIxPb69l7N8gWNorXQKvtHPeyf50M68avlePm9DH
njCEa5Y0cX87fcGylw05PglDEq61NFwZPRqdAqZk7oIvY+uu//zLGppCcvFFP80v
wdsUi5tvo334oZqmHKsZVcejlB8+gtkm3VAb+4zUO02sXVe5bovECSKkpJLrXa1K
cFwaep8/wBN1+9yAS+EMT4RNv+4qz03bJrA3pZTTi6er9sb1bq3PfG6Whs2WmTpK
oS5gABVEDM7AHpu8dOkHL0hCLxoINp83BckfFiwTlOwEhVysz6C071bP/OcqxR92
ao4Co+/AN4K+9rbUiajwDWfs60EgpIilCzkFy40X+EekPqy6m+J/J8429Lx8EJPC
xY3Boc4Ba0SJs4XeCMq1RUn17Tu6Lck6gPVQBTAMLRHRdCfCPJG93hBMftbfEMe5
DJHdqCTU2eXSeyW9nd0p9KveCtX9Jo8hj1NGbv1Fa9/vjC6uuBpd0C6fHFz74xYf
iFa96otaKsWMwqvD0a63iIz7EamRMefx2D8eVa5z8RNxdfYBCoJbl4mBjGoc5oeK
skzjzus1gwQZeniT6W/kLQI2UHzhcv139DHBDyN/VDOs8Bp3YFKcBq1O+znAYnAD
/nifD6J13jbY5kyif/XTFMhe3wQIvnJXaw8EGXy400oXDVQll7vjlydk3fh8pPtc
Hz+0P3Ikje5I8hFXnMg7zX50Ew3+DWGEYihWMgdsP0XixqR3KTLYJbcZk8l86dld
FFOVOAeauslCtxSeOC6OQH4It5qj5giB0zxADt7PJQWGBUhhuhmXZY4Ys3aKrhaq
M+EulmgxKmA1u9GbH6syayRCGByA1Wc9VqtvXqBUz28AdUfZk+LkddRa8RDrC0DD
/ZFfnuHTTC5Dumk9rsAYOVXCE5uPDI5ovchQpCpOZ3CklJihW5K7oNXyfhSMvwJ5
DDpClhGkezL5wwyH4OtYQBVo0TV3jri3CE8GDAKhK0ARbQULN0JGGo7A3okXiA5J
ZCEySFXtjtvlfqmf3KG7t4UibxuUM8dFndVczfyDXXrWAYXF5hsDV/lPMPib/44F
4kMmUiygTukNRTBFQvHrV/CVrc+ehS6fCGOom8mCkdVrOl2J1MdP7UYEEO+g0Dsl
P6L18O4llgbpxTHT9Nm1XOkTVdpqgADiUI77v2CYR0Ug9HUaB+XORma1bZBTy35W
ruc/NIImBT/eDEi+KJJ+ODoy1Sf1zeguMdbwICndvbcU7bHdJKlL3HV5PyW2lHff
A86YZ0bRi7eeaZ8xagok/lzxcykQRPrCXPViP9ukKg7iim+FhYj7st/5X6qt/Zgk
rib1Jc0sMB7RJvEL8y5UoY38yeKTWzUKJcGJmL7zAws22K0vqfrcOa/zuNu1Q663
DM2DzDqINOMUypf67M4dFm82HulTgn5BPNjNQgSBhdHwfTVyDOhsi/4LVnI8kiXU
3++KqUZM2QwQiXZ9B13whEynb/i4sxLlcWoc+7ADsrzzTC8mHssq4uSvgQmzXpeT
4QzgjQwjB6CESMXL3BxJhsjL4UvOL+KtWDpVlF0YPdgMhjLmJGSkafEp6AgcELF9
fKUK+lhw23hdvdLs2RF5KhijzBjHXy/sJfCyShOIan+rciwnnoZ7cStVUN6MGAb7
iQ/hi4EE0p7oGQAWw0J6y4Tu6so4bqtp0HVEHhHnGOvNKauaSeV2ZEd8R58RXEwq
zMXxm+Sbazs00NIZc+CIdIQCQeCCbD+y7mhPNNamAz08kceuAcqD6cCd6xnnSf4S
ooo3eZ/EwHzPKtxD6YTmL3WRNfEXP3OyXLxaLz8p2n1ruWNV4A9U7BP67jnV7Yze
iHbawrKBMPA7jRW910R9NLNFbTG8vCRqY3HssBSC9kioSU6eDK/ni0+pr2ltj4Y4
x/kYzedL4uPMuSmcGBwY6jEljqhcEbNXlZCvPq4zxyfefNiq3zEtCrhe9khKrXdK
gymDgDCKFrIuDBshW0i693dfoGa7pu1Qm+hlUgPuAjj4PVL5b2heKJb/hFjW8ed1
beFw77w+/5tlz9yxdvcaW5OHouubzGZICU3DpQejHcaMPd/7d06UUGct1lMdKYrh
2TiEg8kJ0UGJhNJ+Gj0iBJmqlsB5LYZb4F9Kgden6SlwuCMHXYQXrckHvP3wW5SS
lNFiFtawCn5AkqhUhb3sZkIlj1lW1VPbyVbBLSFn1SeCBh6dVc+TlWy7llYlOWz3
WYVvuZ2KkCJiHNoRDXkpUpZIFLfiMByFs4bF32rQu29oHoElG4BeP9R6PT+Rah8P
J7tsDPrcrUr66buIhOtaTYk6PFn/1B0Hcm3zDMGq2tKfMrZ5yTyUKYjlnNJwkqIv
YsOsz+2fGlOrs93utPAhJQmRHoqyeGW1LUp8N2xsOU8njbIo1F7+NE7/98X27S3z
UTOzDFgxwOIKZ6RrNSM9VB713EFXMGZXtFWK0GUKXoZVXq+Qq5NtNVO70I+NgSVO
2qh59+SWawJPp85EVBDpvYlgk1uiDlPvbeI9BldvCpx2IB7jkxlJajo3kLh+HM84
DBl1oZBQxiodgjt2Ym62rABi+nZ5zKN09FzcuiajxDHQdCi7O7eJO0OYpGkYJBaB
BVpupuCObvk6NyUvQ5vfKTufw74oMFctjC2p27pL09CaoW1js9AH6idQB3w2Gjsj
0Hy9fAJZmXmo4BCyPIKOcK36Fz5Ezl9xlM6L3AaAgnIYE9IYaCT6uYzVQZSb2bTl
zT6CUB/QoawIH6C39EewwezAxYrNaRz2lh8RSRJYju5EBrwL1iHgAYLz3cgMRluT
txCzN8Y0f3CmtTTy8LBzeX3CDCbpM7J7L9/a4m5dhFqyG5M9dKT3AQ06GPeZ8HAU
hNdRrqY15MEOwtsmNUmMPZBQE6gjLcmfcjFvNCBTFnnKhEGQV0N1Fc3F6HT4Cr+e
S/ErjH6FfoMwa4VDh2143owVCfJ78CnZeGUPDAsWTYqwBo2iIRsPh5HWoNXoeQQg
XTS81cOuDTYLxcsX7Ka7JTRl7je7uYOVpNvpEq6xDtNxZuHfjYtaPzUYV4PXkGLk
cURnCi0ZCKWAAlT1pn2UVgA6L9ds5J/3E0M/+JSNvTY6Hg/k3HLvz6levY7oIi9E
cZgBojN/coBbeFgdef93pUjQM2u6HspfzXYIs3p59eA2yYJo81JM5jaiBhVXYMyn
5gVgIthRCklHQgHwFcmGK8dXVWH45lo68WQ3DU1hPauFGU3eEtXh8kYxTaRELKpK
IURLnSpkkcB73Gj7YY843F7RMq7qoyoc1PptUsBm+8RJta6ewXCAcFPFACNqzUxP
/bnCnWzXg/tBUF7HDHNZNUoGmnfSa3WsTcjL9pTJO5lzZuVMttH5xO+ehS2Pc11x
S9xe5goLhZuU+imyuPprF/ke8f9H00z4zZE+atcIYqMQ7wiFWzCbRcQi/0ugmQ+g
LMp51dkWafNfDTn+Jv3oXADhQI+ZnY4UT/U07QvaQCtRt2qbaH5yPjTiu/YaPCEN
FQEulygAnyX+39PIPXn9WAWF9+gAXPuzPMAxh41kMjBswRLrazy1nOQKKFHgmLyS
W3BZEO/te+dnvsoI9XpoN87074lKWzmMfYRfxL/Zq+XIgxvW+eDlqxCadxQs50L+
SDqCbibh2NrfN8AKfxfN4DTgsEOTieiTwq4utXMOiDC2rXmVfc+8JsqMrYAmIRza
H/8fRgjQIm7wH39Nyuq3dd8GG4dniD4S6348joVt7SGUKeKnSQP5/TFcwldjPHkj
qLz4DrFyqJq2Cj8U9zb5O40ysmJIbZkkY4j+9quayv5UC0q+KMeHL/ZXU8ecAxSn
o1ju1jqlZRqPfMxPt20P4/9az6BZDh4rLkV9nf3kHmrS4d03kyP+CebmIhV942Jo
GzL6+igWrTlcTLpTpWyHy6DBFD3i1N+aSePdlvRNbwpkCzmz88RwyWyIi7f1t8MD
OmqBZuZ61GtPBOpYa+aVJgbboLUcOiZL4dhdNQiaPgUYZLfjP6D3T3U5BDPp3ZNM
k17y/01ss/JbyiTEjeGAP+QiJ7lD75CIRhivSA3CXC6GDV8eKALDB8JoogUfhC2Z
Fv2paZRB0zb3Fa5aDQup0zjgpK8NhsLA8fp64x3MNM0tBidZ5qIF3lsYTkco2JLS
e3f4B6e9Qqm5NjOQtqQubAVtqM4FS13yATW0TiDI13kbdxBcKdaHwXO1QCNSWgyP
RoO9BIg8ws3niGTiXYt+/6KuEx+BK4GC7FAcnZ85hQRi9+BR09ve+xsq4tNbLlsK
tAb11iyVzY9P6+VU+O+/2/6lz141N+Khb/Ztp5K0ui+CQA7pWyVuOakSDi6v9KBE
SXZfbnyTd4xm/mrVx6CLVyxZV3uyURsoEz5xuoPHsgvzsoOWHUrjDL2EKkWoCMxd
pUn8Jpql67T4WI2yi9lLB+/3guOdpgE8SUcn9Jln2QfH1dOARYHTKUlvoE/Uacgx
wOWDHLRvLDInlHYK+A4bgQ98SKxaK4OBtN/ibPZADRkqjfcE2gTfGLBHWvGblVKo
k6jd2OgMaUOg/8803vBIEJT1p1IbW6AVUNeTBnyAc4mI42gSqSuj1drdE7FKh0tZ
1xHGUIxoubhQPEkLqszcMlWCstUbCDJE7VGFh3yWqsRPz+RKY1RLEHqLveQ+7MU4
qqo14JKUlT2Yzl1Voq+URsJyqrWH01tTecIvA58DAbllgAnJ+Bb+JzKdOlTkN9Hd
vADZyE3enXYMlpZ98RHRBGy18IezSh3Q0NMkw5XrL1f88TyTfqzsok0EY1KJ4aB6
QoZ6LBbf9UO0mbg78WtIWqKh39h/5rSEvCBUlG7hwiTfaUEg13tTk+/Rq3HIN2ct
efgPNwri9vduZ55bFvoTLQWyK2yGuCRfQfHnliENRsrLefCFnyd1CesslHZ7byjZ
g8ZjEPjzEyIaZUfd0ilG/7Gl7Z0LXQaEQWa2eOnkEP9VnS3v1gZUERLlfUZEoKJn
iHzjGGRSI8NxV8d4SfJNE1dJKo5LIdp+NnJct4PsWIyLIRF8nJ0X1Nw3p+SxaU6Q
ofAFKdeoCVEJCHHq8MkwMTgAwpA06QhxrSr95wI+IWjomlsT1Z6NT2HV752jzuGI
h3pFskBEyt17fTO6syexWJ6vNfJ39YQlEo1deHpP7t/x4TXvPARKdFhsgamwI2e6
djbar0ZhLcoUOrOAPgayJtZx4pHDXrhW2fbmacdzBGnt5Voi1JHVM7hi99+f3yBf
mWwKLqazzlZKIRQEIGnZ4+ojXS4nscer+Y0YmAbQjxIKn9w2nN0g143w2UmdlfQ5
dvp5LYdbV6btqx3hmggKBfnemCRGoHOgA7QOWLX8ZQVIF2HiKitDsutXZcIg8z4t
8eGYQo7gfzGwdxFXQnqJluh/8fefPA2b9lcBKIV6dy/Kh+5rUS1ombkaKHWw2WM9
qoyzCo2bE5FJXc0VwnWZWn5S+/Pd6o7cc7KeDEU22GW1I8/ls/OKRRL51V+b8PCH
vfxWEi4+JPvlmoZeu8V9V4i6oTeGwUcr1zITTSi2IfRo2eHjokqONu6i3kjabRmE
UCpfw9pquh+yNFooaKKLDZnNaTUeLDmKWw41QaV4KosvliOE+dM+Pyuo500P9Rjn
y5LgMIw6LZ+0wd99t504wFB4nsIPROH7jKwQ6pN8VyP1kPdrqKuEtHxzSHyuZTfm
MlqZT1Pox4thDXmq3TVC3HA0VK9XXXeVCjfiEBxVg0ugeYpoTJn16lS3ptT8ar1M
cfrscUl4hRd8ExB8Dnbnhm5AjQ7l7eLlrSQutxgHDiCdOArNiXExT+lb4cvTqvCT
uBYZFtwJ0SXRS20V7xT48MACLqc/VylC12tcd44HbvSX4qkzzFRnT1ogxUqIrep8
lvpHL5dcWVS7cR74nfY6A3LVpr821LoWYKRUVdTLS0AhGPASuiprkmjRVNh0s59m
uyfWQQ3m5afUkjroKUuFLSXLtPBzMPn9NV+8dRBFaUQwh4xjO2XQe94Oq8P6C36t
hSXSKBT5rJqRC5pr/6Ph3WZuQ/iBflR4Dl1dp5KnMoMQn0KS6TzDdCd8VD6YMeHG
vIkyHBFbf+/v/GYBW2sV5TfdDKxoaaUhBdIGsg09khLuoPX7rcF73Ce3aKWnzjw3
Ma6Yy9xuucbqMUdNE2PdLXZ9eoFdqWyHlyqCowQ05yUujvPHqWAGMqF/8eJwcGRm
s+34218UtMySyPzT8rgu9eRT938N+6LF+JKMDal3PjObLPK3xqJuBupie+iMzcIU
0/npob0rCVt3KzX3CRysL9VVGowJS6xddDVxlj5RiVwIzBw9GuGhYf/hSBdN3UOw
EVzRDy4PUZH14xBdyTkt2srdKm7nurAshzdWmO2jlWtbmY45Kojo4NUzaLyC7Cqr
dnjwhPOe11p7TQymwhYHMTWxHr/8MkNIsL1h7uJxTLYPMnwFy73PXspPRnGB5Jxh
kmnCTL+E+rvBoom7GaCNS7UBHLytUj1jpGnoUp91iK0MsGni7CRfbacyEXytPAbJ
dDqRN3a4WdNNa9ZegrVtw4/2Nvgq5+uYIULZNhcEj8hARtdRqS5+DbIyLs9S+mqL
wNwqxYnLH+G2MrCl+ywJYgxFUEQ7urZqX+AgOMwd2TlDnvHoNdGon8Wa2JOZUM/8
xACIb5GZUPFp8qx5dLFsvM4llnp+cTuoOxY1syMBddTEmOlSjDsDWdQoF29K82Q6
rphB6Xtaffn+62IoyBjP66g1hb7AkOCG/VkaUti+7IThcqHw3temqWRG0rc5J7pD
6J9GWYBu8BcbkxWed1Qkl95nhIF/wCcds7puPVNPcYPdIUNzqPtV58Cf6Z/yg1bD
gR8gyw0FlWFNN/DcFzTSeP9XaZg1hxEioF/Nt3Enaivti6pwbVV996CPWmMw4wf3
YqAFqU1a10dtTQYkHjtL5esEGaHJlbR9J2Eb/OmT2l5NsBoQdfnMBGtn6UEBw2cr
878dqmmQevsl9X5MoIyPJRwxf6KeJTQ+ivMl+fblpcneHDk8qQ4Y5hokdtwcwofm
IoFGqANVfD1M7H+4rg92/v9Dz1A8F6j5GkvfvUWRKGrYAey1oxjpW0EJCsqhwnCH
xOC0L4FcfdDW9akxClMEI9p3kOA6YCiH3JexUD4EleteWQ7EQPNjWc1YRr7YIjCf
r2J+1e9DEsS4+VaHuoHgaslKsl9Z6+DS+BF/xCOy2WYQ7XNWy/PBh0QPKhlkIw+s
wivJR2KH2JZz8a3ZEUZgfU+Lc9hVrfa6Vrrn7dj2h/jIKfHJFZA/SeqypA37pXzs
hpWYppWmGzC/AXrc4/IAQuauRaflMXitRty9ZTfCoVE9PWl1ZQn/j8/OkC9di4K3
1kgQDlvrH6VPuDn3DtX1c4bm8jOMNWXVhzONnk3mccm+1Ju4mfkymQqe9aL8y+tm
VFG/Iw5LyCxDNpdRiVFzz/8pbGOuXl1oAy6/ymXzl6A8Ni3Bpmd0yqsIozAbUA4T
R/xv9Z1/YfNN9WjjqDqNtLgwLWiCt0g7hw1XnK/pCkOFuH1rn4pGvHOQ04mwmjnJ
V9eH+V63n5fgObBgaTIRJwbzkMasqGmTnH3N/lHXwJu4ylRXa7g2laG6RIQ9q2Im
pMOCRLwAbz5Asox3dhXD5cDm0hkgbhsJFN/V6TDKL5t58tpE9HDmD/xVh64ejqUI
Q7pqU948SHzLEvNgCns6yOtB6viUtz4/AEZZo2hGnf9Jz8pTkRe/CUpNJf+1TolW
pwJNBk9ms6h9nmGS7JRjtmrDNw+VHvgVpiplXkBHVhccK3OjyWpNpHugLNz+huLX
L4poSGZL7LZkRN0yWRit/cn03r54tA0F5+ayrp89G3gislHqdnsRUSxc2gXwuOsa
ZWUqShbHDcnT7J5O3BWN/KFgFeJf4wEq6dIk/3zgBJFyNQ+zAemLYF5jozMqIbiB
z4PfUYZWKV8LSdh1L40jLwXCz5ihN1kszzAQQu+/2jDvXD2sh29r6irE9bO7SYqH
oWpiEaLAd0nEB6vNxTuW00O4SXEDRSNqnIxbVkJRhjAIvOXioMnR+2hhbSqRRyQs
kyZBqATFnuKJSLuX6RPL0BjCD4/RKTJuX9U+9mlTYR9UYTD++BBP/iHzTWlx2D0m
CLd3Q1AjpnUwpUsT+hOBLpZL8XvuGJTH+fvWKrw2P/gWzxbjsncNeUBzTuAnA46+
lOebdlnYK4xMOm/oob7H+VNn7VPVmrmLQq9PDzdTd84zKLJ6U77CkpvCx0kx2p4R
LsPgxmoo/plqWeRMEv/irXms00r6RG83rTCXdXMWm4cBmzIQtI6M85iKsJ0/1NoP
ESMpkhDK/YugATojgqldlH8JcGXmKAkPsf2mGPfinfWLB4RL1vOxqUE3gBWf/wG6
yPAErei4IJsllNmtIoZKHEc8Q7pqK2fylsz66eIIZngfZ5U4aY0L0rbHW/Zd8oD5
fIO67rgF93lzac+dobAOkOPGgCV3JEPQ74+F+6jHsgL6B/9jxYC0U3uJYafHM0uE
MHg+LMTFXTm+ULPdZKj1HIEtshopr61e96zQ/kQY/832mvQLgyuHtJF0X/dN/aJo
Q1CQMl3BHBBh7uAY7UCl0kU2ionbOB6cav1RyCWwN8IZv959oZ0Aj0cf3fxZTgh3
eLE9ZdOc4oGbijpqecpadfMo3Vl69tUFedtLlpM+z4pVugE/9H0eG/JVzQdfd9Hu
+d6Cr+nActA854+qjrNm4Rj2VS1nnbxAwVs2qhJXffEqeKoTad5r/TCr9uVKRKZT
/FacGMaK2s/iY4Pbp9oKy4SrH7hfAufI8jh0I/2r6kzjVSuhFlvi6iaSDHza/rNK
zS+Pda7zqmHxAccTZ0oH1LdvM/ynHGVBci5ljQPzhFo2ZJ3gYVKsDvOJBxZFbB4F
Y9o9+ckaTjoBABZm5SFHukcUKEuLTAawgQAD4Ee1C5F5hlhCqLFH2byQ1I5/YguO
jdfnfXd4PZ+eesujNfxYmya29BCvoor4FcHHPvVR76PzsH6S3MByAU8QcIwKwBya
dlFUbfHLfiLwiG2ENuOAHcFvqA9+xCQzvMBm36jpJDVYCpcaVgJOJsHCmk93CDXu
ddi0CTIMHZ83MWhxVHpRG2gmylX+9z3FTks6CKDRHJ8y+810mRWMHaZYIgHtRUo+
5hq+YiBaFrgiKhjaWHp3yR46wf6BlhDgKp8K2sRDUEhBcNL8muEnJv1aFpa2Rv9u
7XtXRfcDPcKqA7rkfvzgk46hCSNrpdraz+ojcWcBE90Pqr410jFDSf25VU9ziq5r
8w9YlxmngFG8Hb1P464M83PBx2fkYqYJSbLvfUVy7mXGjHdXD7J6bsgpOplC6Ary
Avduotq2EQTyDdBdbbne/HEXSc3PiXdsh8f0AzLvp9iJRGfi6F0QrsTuqz6ZGnIr
hTXfCnALRIpY23p7pfp5/05cAY8DbLXYcoPaCxXmFcMcVlDd7IlBxyQYsRNDE5++
joN5hslioc3xqMXupbGlgfKemC6nBfMC3g5+dDS8alwUFORhPgG4amc1cGN8a7LA
7Oltb/bf0PcQzyTg/jU3JoKOQW40pt/+wmAjLYYqM6hkLAx5/nnhiYdeoXOfbuTd
8aBJA/z5gInCe1DpjSjEECn5Y6Gk75cKsdQ7CewwlapfQaFYk2J18G6j5nAc7wem
yNWCSmHZbPhVtS+ZoBSCuxCOBbh6DnwscvkpbOxsbDLUJNYewL3j2c6/U7ah8JDk
AwPOgAdGYedtQf7O++H+dB4hWc/D2lSLuiKSJP8jQ6fce9DERPnKmGBmr0ZVIESQ
tM/1dGP5ASRbhncMNiPk2+68MoD94Yw6u5j3vC+H4YVH7+bICXy6/yTaUBLyE7RN
MXzBfpYKjaRz30R0l/YcY/4f8NatuAY1BhERRT/k6YscS2LvQfzZkruWV4c294EM
Td+uwEARyPuxqo82oLyBmBUmKVh/aikMrUzaMOiJ4ArApv4BpGqBYeRs6jDIv6YZ
vjzsea1pdDImD5OJ400bQo11+D+fy5nv7Wtj3WKrXjJiEVSAZV1isocmUxkdIFXl
tj3yhHHBKR7brDS5txz9TJfFKn8V2wKuL1YSHbNfpt3kXhyqMvE0O8lnULagbSrL
1uWXQcQiqIDG3M0+Qb68mxluj0QkrcAPjTxiAw9phiM/f+mLLykUv735iKmth0Aq
IqVvzWDYIW1JiQCD1sm+pnnuQJ6+ZCb8Bn3DrDhq2+OIHBIyi8bb/TKZT7cD2kAa
uL7IovMD9rmMmCwOe208o42vbUsgWlIgFbozxC5/Tj+mG4OvQX1TxYaGnz/NJkOF
aw2/ybHBE+UFaM3YHJZN6SSbJQvtPPL/F4xJs29TwdD6fyQTWi6jEdbSPETaIG+S
SygbnXqqwDNqIRWJ78vS/DZuFKPjyfXoHvVAGphiMBc3M/6+ngcPulzCd/Qp4lka
wQbggOkCOhsYyNlJw4HK0lB3F1aiZgOtN4+6MzV28xKjKSF6J90dMWL4reL34gz1
SLvLeGBzaKnqtJJsxckW6ZtEPVdG+KNvaD4ruTpeGJRe+WlyNZ+F88VH5bTlXA2l
kDkEe6Al6lgBDvX8easIRC+Wg3ozqxrJtCpSMjpGe34JvepRhK1v6+6d3JoHjOBx
RmYLXmenT8TIp33pTIwLl7GXQhdqrrYnLqLOSmX8ycn8BfV1e5Pr6ctUBxZl+Oq/
G36L/j0w75PIu22iAEed/5P0lRQ+1tj54SjMoX5j+rzekVc5VAOpIf5MrViMvY08
CQ8sfUYD+uI1Mn/HD8eaWwdvq+E+0KCpMOBQFTn3YEWWoSc0Yk+nNz102k2rEhw7
i8K1MSEfMCpgfM2sJqi55SSwqc8sFTxAlVEreOscEHvcxyLDz2cYJi45Nqai+AX4
Zda2tlLhaTH3pLMcikRQQ50nNzPUtN4KIGI+8sEsXXd0mOMWwVZVbYDmAMGAInnm
JR8EynVV0zGKPkZfdZ3+z76SxbQIWgjItDu+zKYXHtvVkT++bMCwweeau7gkr6CK
uNZYQNCMef8kOdR0XHJ2QhBn/XkEidBZ93pI3h2dmi2LetFhKpecl3sSDxX6xk6s
80OXvBbN0i1UQwR69LvANJoKAkOiv1kTzspuHwUD7QkjFx9VbvjYk1GgSgk4nORq
1HOB9FoKMwvKA2VH44hwCV24SO9CZjTgDDZzg0gFPNXzbZs5lIPYm6FuWjZ6rLd0
9arC8rS4vGke4KwD1Q08gJ2fgvmWhLldBQWXFvBxOo6WUHuaph6nl2sfYgSUu1J8
SJPpw+kmQdcDEhlftv3U8wYQ2nkQn2uM2txtwHGq3qi1YVeL9qUCAQ+HatWqUZ76
AcGIKJpmLoGIzfBU9DCGdFDUQVcCl8sB7VsmwTItThhk2Y2xdu7A0JDHocbxbHnK
/CnAkmIRTITnHqMg9E0Zj9oPW4UjCuimfHxClQkUgOsPDQDKmBA0A5r9xAY+k4UO
ugEiNej15sVGBHg9OLbcR2QtUQcobPUPTLSVyWGTwK6pjZDvoYU+DFB1i+vFq9kK
GkyHHs4eUwwsm3i+HoaQ7ZdJrniIFSBB9acVTKWk33sGgrXUiYiCi0O4veuFp6Pz
rQw9E2hzuXYDtHyMrHVF0NR2KbBEabiKLzE/oWXUq9KZFG73J7dWxY6V+9CyKXOi
J5gOx/CX/fDdf8Rf9byVH14f5KWpoS1OJtMgVBBbPjE5MpZQkb6IZt3I+x3dbFuP
nMiTohA5wvWXdP0r+qYjOfMybwbHsxa6igziGydvMX4LAMhtvmyVzp656q9fSjcW
dFXS38J4RO6xmGuvVmZC6Ju4ySoxTFwY4ZhOFpewB+eJUWIlh1RY9WVvwBN2h91I
Mam9iE9yz5+/2IBCRLBsUh3yJbh/ec9Fd3DAa36wPmISPogtuKUe2hLIDczuKg1B
Ozzhpj4Ued0FA3MJlzNb9CXcxHHY2KkaTDqBGtPW0u/rXgQ7TU4K1iRRq8frgkqu
t1CeeYSb/Y/+rXownr+zO7QBzNLXTjSHxF2VYbsaaFe0YxcYblytqbOCwQWi2SY8
ohVP2EamkSlyVgqACeHadnjxnUqDA5OwJJuawMeORVWUogKJZgFyVrDhumVm5Imo
x6gh/vTIpwAd4Yi3/QR1XbIbiQg+r+vg4CC2ynQgNnEcAumyhKmjbtK6iAoavHad
ztJLxnDZGk/2F83OTq5k2JFfbdlqI0CLoZS5V4rfYKDoQ93YlcF/i29VSdtms+89
kah2gTNkIy+oSvX2uQ2mI+rLlTP02dEBTAatFcMvWE8+4ovdKMdANylaK6JCyGqJ
OQZlYt39BiTSTimRn8CL0qO5DhB50pJeaoPaE26ZbP1r2DPVDHMaqe5krePwd10o
051xUpxkI2DRFi2KPP5LBL1+nq7/OTjEgAvYzZBMUWF/g27jW4ik47t4pABKLnXg
IhBIeIadvp7g6bBY4Y9EIQlfF65/NxmpL5PTY5ODsU6ZdVV1xH4d8rWzUSPESSeV
nYjvWWKoJjaxtU+sbxZDrhos9oXmHeEFTesxFObIepDdah674QVkgYLTIqFxSg9b
U4TN/U+Lx2ZI7op7x8VHHlB51QnAgZDiBRJk97uN4Fc3OGl9lxMkwAEvuLjkndF/
cMhGkR9dBj3KaeesAQscVNXHYGheZoTFUT7kULmhLOPYYKKgrpe6Bhu6zItfCflN
ZBDQMQYS1uNg7kf0hIr46swE4v2gjU8UKXtglkmKc6Cn06XMQOaVwWw5QW8QeGXU
eazqtxQBbA43FU4fPaPgH3R9Gx2oneWEshtt3m/fIRXXuXHE8bhpYENmNE90PY8+
CzWH/MZEF7KZe7MbO+K1RQBgZ4rqm+sFWhH4U0p3wCeJEHUDa7oV/PMTQMQ8GlnP
+noPDcau6bOmPeNh+GdGjQmhh2VYHvSR/WuEIceM6FB4LE8WKSHeR9JaZ94QrXu/
FAd03/JNt8mcp8wvAN4pE1HWYovpM7NAZ+H1yclj9tq0B63wfOGdW0ESNfPG/1Vd
5n/sIVZBpNXp95luvtpyZWwp5s0egyPFasgL2gcM3G0XPSRQIwUpa7vE8TzTyml2
4r1OzqdM1Gx0YbYUOm77+Q0CS/hMQUX0qbYFhyP5nGj64nb4fD1iM1e7dLhqrQGR
KVgclqAdKlg7GVfW3x8gVokVvnYLbUiN2Mx7Y6ju3A6GfHVoMTZUVFmdiBehvWoy
lC7UBTNmDgy+v1ZyGUzMEJnuytKh5mzwNPbPhcjBb7vKoqYCyjlSO0cgyinRlfc1
lDx/4a0DzzlRhZAD/Tr1iIX1yZ8AP/k8yrM8AbCI+ssDhfhASNTKqmt8ECYCzmRs
0eu654KQnUmGqKw0OWnTHipqXMj95ljw6OXTtF1uspaAPwbBAdSya/Y5gb9f2nmV
bo0m2OJjOLW27n+YkBDtL7h8r1pmIR68aOGbHrwAOrjZP3yjjTVKyLW+uNZS+Hio
t1I1QKGvXP16GRqXTJf/yoJdMiJ93zcYWDkMe4IWLgeCm5gmLg53sw5LENQKOPsj
ZL8zclBLPiU3CB+umQtRtbd3CGoB0ylC9tmRPGhAwOxZ1MIhhguu7UQRKMybHVC6
GV9le+mXhKZitHLNWXLjTvtmWqK/ZaL1UtSSJT8yQ6SH4y/XmzztfOoLd+kKbYeu
A0rbu+4EhZ6R5vGgu4tEDK22CTdibStMiHt3rZn5uxnANvgzjL/mxOH346+WsA99
Q6RekAhInOT5bp3Hyr+h0pHd78AGjU2E5jEkXHO8GFGsH/MyIkn4zM78JGi2FTPt
MgHSIVKhfyL+Y3fxN95PSqSapP+qTPGblno39l8Xn9cKana0z8QJN3W7UuNrmy5J
ufHgY6y3QFmXt22QzgJWpdL/rBUfGf4UXKbBiEOcEOepmq+7iF2dS9dak8qRIwxi
aynQlbmP3rus1Dh/U1rqioq1F6a5tAwqpoKme0biHUr0ir3goVDdGz9JR3+L9/ic
27B73RcW368iWPjK7SxTT5cUPmsr/LCumldogSDMb7uXmyMqR5eOcqwnOYrWoGub
26/GLAAzxiQDdwlW+NVJQN0IM5m85fRNN4rHttwaN3TfG8DKTfcKJJ8SrvzIbiX8
fKbvmuwitx+6IJZCIu4Y9s58ul7OVcXP0gdxwos3b7wdLLXSAG5FL6n7RIsRm60X
FxB1yRqh4fzGUv3qj6XIvlyYvJwuEXyJCdi55ig075vt60qdX3s3Tkoszg0CsMmb
LrtRbGTtqOG3SbCvPe7/1cmjwJZtgsD8TpvhtuYYc1MwkgmzhdoSiPdZtxDN1Oac
/skfmQ1yG/DLvIzhr7vd2QV3D2LEeZSH8QinRxu3/88d/sZDJPEOLCA47UBrjgd6
Ys70Vw0hIGaR14kFvV+QkhT85ZwBszvt72RagocYj9nqsOHmH4ZukIfwtROVy4oh
xVostK9lGe5LU3/jF5QG0HimaT0RJgTm6cTG/IGhGxQMjPCU0OwgEqIQZQG1evlQ
Z5kS1hTOREqCOIbRfAEfbZsPsvjoM1FkN/Mj+8FNsnzZ17KuaFNV7adsLuP14sbx
ZxLr+1toeNvqVCsWQZT0FBchCOO64fu/RRxa2ywKFquncxC+v5AJKzlB8c2eZ8ul
v3PXrJkwiRdC8p0TkWqSliOO7H/Kzn18hZxXf64c6h9vxl+COMCRLRHqoY4LXwgz
EfSjMajVcwaU9DYc7jOfmr+VgVyOGSeW72cFipRNe56qxDkWWTJ4X3tM9MxWzL9c
osOc51BaZqvOtAuZi5FlzE97pVmED2doOWYrL+GW2+vBLHi4OI0XrCICf9kRgrFd
RrtnCsj7p5x1T4+3753MoK1O0yR2TRnzYaZG37xySU49x34FLGMJFr9YOhY7Kcpg
Gea4dRCH1qJsentbSoZPLcmrQ7iXgLcMQJpKGOUQlFh5Wpms4Tq73TUydnpEbjpj
ngr+2on0hxe5W7j1hVkDOBxoZmHAEffWk797iVoona21UcFBv1mnKS6IZ1JKy1RX
/FfBlGNu0Noy2a+yW5Tav2Tm7deFzIgVNfmwJzQhnnciwfajSNmllZqtGDbvHdZH
cx8zYU7DqYFLBz2T5rttriKleFauRKkHZQNyYRLzfsOpAbXFVpaz0Kuf9vJS6oze
wiCkZrOQ14LrmmZTYDjXX6tDajxyDVWgOAXN59JKPceYxWayYy4QXC/RS+qZt1/E
MYg0bssU2Z7Fmxx6q0qRr7QEQnHSVOKs3NHMBUxIMx42W9qBV8Kt+9E3yuLe7fQB
lqsVg55Ve813KLUwQ95rjM3NR/aNGpT/vH/UF+0FgyvGRfFA6UPiMK8I9+57MmH3
tAoIEe9nEigEWzoBmVhFmnVWUJameX2LdH8DSpze6p9nJt05ZMCoJ9j8HxZZWcGV
PMTsp5Qfp0t/XgnJa9VLpCMaxBI081uT0TaDZR4YQ4oH2CzKUD5FY7qf6lKKFTiH
SNS1UdBcAdCeTYfRz7/8KDxtDD0gPy6Fdj2ZIEHRrS1I9WRF7q33SnDS5rZvcsKz
agRSBgvOOPSB2AcNcrE+BHzc9WRT8nqYeidJ8Kd8rWMl5OY/gmU+IwjCkxY4JXNV
lJkg+HfHXhNqhMHcIM3KO8fLVzH8EbX6fyTjFVtJg3mhnMfUwqOAoRzwjUQre+OJ
x73dzecDvaaVVy3ELvYGpRxvozV8hQJY3vClFMMfpNWgfGvvOQ/6gcw97BIDNjwD
OPYAsl47Vsy1FW3cXdwtkaEdlAN4PRNqOC9WJ95Ge0DvkwE3GSTemDJu7MO171TE
Xg/5KcGZ9OvGrGXkUkhc8bt8jQGXNH5f7cUPRBc5dADVpwg7lDR31tj6DyxdADmU
C2KlEs9CWb83R5WB7OeXygY3V6EjhzTjjYXej5bK1xDWroL0pXwDQcZ7eiXXRxSK
nW4z/kLVZfXSN0h0AbSNC3XzWR1UsB0+Nz3364q1hcVGrHnXzCqe59l/RzlKoPai
xzPwK+vjU96aB+Bvgp7DDrXCNTZQCIW3EqorEDrQHcDh6Az41AbFOoDnKwI1qXuK
E/lukV/pJlDh39x0t6ngNqhek9r1PCtGSaEfgK/t2qzMa21LAX9h8GmRyx5iqh/E
tu/ORdu+IKEBCty+sI8TUFVxIgYKzOCQk+27qWrFCsnCi23w5nkoPUvXgRiVlaNZ
p4I9hjgdZOqJWtA8t7milF6OD+MKdQtrj73lZApFQsFX0aMWRYSbCk9yT5/iVIWR
zdhO51IrkwAw6Oj1rftnl6q0AQxEdPScms1Oxcv+V5BOgtLzdDlH/7Hin/Xxb1kU
a231grFauPRH8iWJnVu1UO+ldjn4ok1Nzs3JU+WK48lahL4RO80XjoJr3seBEaJB
+UHXIamfPQZ3jOMQ037qqj1Zm2wL6R6BSk7pksvy0jMZ7bYLG4Sw+Q9emoh8kjae
dAdZIk6Ck0iDZxZYIf+Oo6MCpw+3YNoxaq5cXehGW09+sGDRbv3X/QuQd7Neu1oK
8vyPKPZpnYLDBYQTr9N5ztjrwFVa7AMmpS/Weub+EQyL4ZAcDmEZ0wVeNKK6k8XK
Yj0UaCUfimBjOlVTloAS4RhQvDSY2xRu9gvSRDXEiDsejEGwekhAXBacHtEasIBk
ulyWMh5tGVySDhxJhQWVPlfpNIHYxLoFaPt5IETzGsDz191GYNyFQrdXqtkPu9W8
z21B1NpquoaRL7iZN3bFuPs5RFGg2qEJCDsWJKQGfqKlSuYOVsvICoKrLUl8XWTX
V/8D8bn4HwLX0rqADVZXSxFJSZWTjqS3rCed9SVfoxAqDvkAepZ5f18NEPCFQaWQ
QZ1fxJfIMA9cCUNOB1ThdYB1LyJqOXHcXg+T739ph6Xr2yntV2x6QxYy0zUjabmn
jq3Qk4oaVHOWt2JFMJam2kYG3HlXO9M2Bt2+GEHIblcnRYVAnOYK5qRv73YFo4c1
rZdvDItDEXerI42nRVA1D6AJc8K3NAKbVYUaF5nrR84B9XZhD95U/9qV+mKJnwyS
pW26HvLK+J4D70iWiSXU2F7HzmuBHVNk4Tv4/dfC77mzxOq67kGvlTDrt5AVkjMc
uzpLsYPezaPDQktTi8u8T9EDjb9OwnS3QsSXEcVoWVhfhpJ7CFVRMQBVWyACWINX
ONZZ5VzxBoqF36Z9ITzvipyVwZAjIOjizvDzaeLRkmCk6+PSTVdlXPNAo/uBu5Eb
aSYfzN8e1Kr//PcMve8oIZhwei+bOvbTg5bwSTbk2spT8KGNrD/d0a0uuCa9Opb8
6zQLKcFn5Y+//3jlQ9tLowKfyYjI8NhU78FXzeJvcKMLW/O8A7qNWd4ZCIQGxETC
dFnpZ1mV7XOGxaHujZxPWsfg9u1s5mM4h5jx3+VTIyLaoWKlwoQkNoxOOB+t8hzA
PVJ834M2MD5p6kM3GSZiWbVCd/f6Mh+nk0IsXtbRXjgJJMLNWwp0V5X61mcPlGFZ
v3Tj8BJ8lUP8MttmyoIQhCExHCMCg18BoDry0cE5MvuNnmpqresbFTjvRzire2vx
HnmerbRrf770V8eBV5Lwk5FZbIN96g8kFJzINfInJDjtajEaFUZVZ5ISGIQS2ZgO
rPVwLFCG3mcvqkAgHh5fSBLglcKQ5KKAnQxe6mlSjkU/+j91T73IiRnw2zFJBFwG
9udGuVpTw3zIIYmTpFppUfz6tP4rDZBJiAMa8y5swVRo+HrKXaQuGf6InsbaeUBX
58c01QXyJCSPNO0dbB0GXwA7WX66ZG+P/pLTMsJVi3bytkqD6irB6M1j0wnxxai6
PRibQ9kimSQvvCSoBFbPxqyD76Bb91yBIStsi/lZ1J3Q8Nw1XpgUtWRYFsjHGmo4
1AquosyuJSViDR+LvtUc5lC2tVJ6l7gQpgaUGqJlgrZkEilEHGXR0N/pp3JwgztL
GocUMsQAqvyPX6HIaRcTUS9E7VEVfkkgS4mPw8yO6KVomgiM5pLx6I6BLkF2MITp
XWxFu/57tT6vWUN7my2/SXDFyC0bKVOwXH3RubBPo7qPLQV/suQyB3LmnNf2+3L0
kaj3O2WocKqKgmLnvAXlM5pSeTkr01cVg8nq8Xwq4051a0QhzrZ959IXETvTOKkU
ElhlGuZH15ZDRWQHPjRz9ZZ9wxydUQT7nx3FLcdkouBzKAP/+wcAsh+v0zfTY9wA
kXHWpY0tqDmj07zk1QstrkXpaKX5CSA3Jr8PjPrKteNk7ybw8kshQvsnBQpqhRIb
tVBKNMjnprzzZQ3Tuw/EtcDdDP3lDhJ0/UtOUtBpTx3ZjmJ8Lf9PcMxzKu7JSEEm
7GknTMK9dUSfjs9ca5zbAJBGiFPKFDzSG3Lh6b7xxJjj8XHyQB883W7incpWFfID
2sVcddJbBm426/Q3i/q81hayav2CwlN4/TKuwbhr0JWZg36G6O7RhuaSbaKMzH2N
1CD3tbsx/62+1Wni1NBpAMtfDGE/+/m1gF9AzV+OVtQTSaghZwdxuWy9iveEpJ9J
QZWEtaQ08UIyXupt45eDgJOP2inpKiODXOsbaz/RHB0qYthA51m5f0rwKLcxoqRx
W8Z/06IAfxbOrNnk7NGZ3cBlDnyafArq6UIWIxb6LXD2W1aCuymKs0X85nP+U37m
kgosYFhp8yx7anUgRHCEzv8Gj65+DeJ+KhsJhEb19BAk2bxpBL9TyG/PRGxmdQ4Q
VRlzLD+IdN3TcdtrgBCMLsv8/x2a+yaosGvxe2REWKohDRMDl6/Hvp5BS/2i51Oh
iYx8DyRWL7Q63bl2A0vud3Zi4QQUcq9OLkPE//AU8FO309ekGLg7XeNol3U3ZmNX
FhTKGU/0NRj5+URK7sZ6EhICDc6qhQhlu++6CnhBKEBVrXVD3pNHDuPJlXkkQjyD
GiHK7LAzb+fFzIy/gqdjDIXsvuETTbPuG6wOV3Fl+v3BbHNiijJ8aJ1JyHUUgmg0
YEDUVhbX80omXLgXd4UmtyAzcYCs6nEn1oQNUA2eGXssNOsTvYaLkvgbp5tEe+Ce
qZc0UcFurduvl5KSn1M5pa4md+2iug1eBnml4punnSmttqIhy+vN47/eTOMjnl9/
Ss2bnM1dRuGf5qDUWwrfLILqbj2F5jJrCAh5I6uiW25dD4U7WPL61v6mLd/dZxkh
Q3VJuvO2VHy4iY6mcaKUL7jQLEwPEa02sbDtzMuGRVFvXpSqjFGm6SNAu+oKd28c
U1uBURaIpfp6NjmEwRfwQRK0/v2mUYobKo3NLWh+GYIZlcjc0yd/RzDA2BYa72fK
UOdbXhOgm2KEzH+2G505xe6T1JKeREBebxFovV+gtAdnut5CTJb/kkxpOEvY+CHq
lSXK9cOvYiU1Qiq3RxJEKSIH7Bxq389+rn1GcU12se40HT9VdAtjxwU5wSJWTigj
zpJOehoS+QqjG2Tv2vxWQeiOBu24G4kF5o3vgwlbmMZDXn0P04KpLGFAlNLTYL3D
LxEs/+oWvWITlkGLzAnp13odzzSwtO25kdinNwWcgv2Ypy4DTBH0tlaXEIXCunBk
qcmtDOaEkS1ZzPoOVxehcnhhJnJ8bKnVRp0OlB8OWc/ysogX1lEyd7eUl44XgTig
IqJ8CM5XbRzuGa+xRFBlgKeHY+o+3KrMMw4azqFBucCHKnVUKfSJ8q6t6krAPUiy
3GTrYokzw1fVl95G78rmvzqYb6k+baYKJTMgStoQ4VrkQtmtHRRFhYRuULbtkZYQ
2vc0OBV7AWWfqRcwy6hovLpv/QuoRufOFEgLKy45hzq29UsvE54vNBBpGtP9WyL/
X3D52ys+rgWXNLwRwkaueAGDjQ1XuNRaKp16BLsqMWxbh+aBKT6llTVGXhbYinn/
kaWKaPH7mZfXfPuUs1tHl6Fg1Lu8eWkyTYq8M/ite3q2go27ff7SIjS5WCnEK7k1
kOneqTjUN6VO4JTIPn0a/jrMC4K936Q1aJaGPk/2djEixI01/qm41xGJ5tqTamUF
72LcJr0eFYAUhYqy0oaydKZW4tsnH2nlJY2N8h6mUpudOIx2IJEgsdoMBqm9UMVD
MZ+mN+Emx0393EiQeQzN4GIUt7wLLRfz3lugu60bFdpEVZuQLCChG1sjhHJeS/6l
OliYzGfBMgBH9kHJw2+q0MYMlRN4QRpkprMYvL6mN1TCIbjqBZX9c/x22GFZjDE3
uSxoxyPJFuUlSW3Z2E+l+gC54KdiF87oPS+2FHvalkciwMJYmmr2R1/R/WZAFYgr
XlqXk9uwRXXIlyxzzHY/bsh+ejFpwW6u27htUux69llxl8X0f3WdkQqIX3t59zLP
mOnVv+YIJjIDAzYym3sq5YTspJiOFQf7Y/diWrNO4t4VbuxK6+SzPRooo+VoIYBp
/18hgki/u8sph41ERorZ0+r9EKMjLNr7VwPCEaeaJS1/ZE9L/MN1lRGJ4JIPjb55
ZBLk4n0941A29abLWKhVFruERzN+aoXpXTDZWmF20RLZV69oH4oU6PU5GfE6TJF0
i0zuo053ZauwY7NJ5nqSBMzAY0t/g/NI03lEAGwIZbKyd2d0y0aMoC4255kmZZJS
AZ5eA+2njgDxOxjE1TGNvVsVzx01+5sBO1vqKxv+3XcCNYueUhtP67JttjmbiAB7
cNgzyKywYuoAB8gcCLAwf+w+/m2GqZ9YgYxzV1GqWZMBFZzChFabWiRw1eU34anN
sPQEHUYqf49QLaa8/fS4gH1cOkE7v+r9Z6b5DrTH2KB1G7wPMlR/LoHhEpnEtKg7
2HtVx4hVcbffpmBJTYwk5HKQzR2BurT2I9haC0iV49KNQ5mIpAW+C0AJnUMucFI1
dD28gYc1FPOXWa1un0FJvrBSh3jIp0kbVu646ehgT3sBGpPcyZ5axtH6Oh6Vm24q
6+f+sgTq759zHUOjd+DtNpuFGpuXrH6nF4fY+jL8XzFO2qE29xJhRH5rHxW658se
xiH/DpUcpqioeoi4tRw3v8qEveFlFUgw8zqxtXJTCOhwvegmg41KGIUYS4er6vi+
s5ZYfGLkgRYeRVn/MuLop/YQ1FRK6d5HkqzMVQCrY7ZP5sy0VZ7pXTsKUZfubebx
ZW/465dedVuSFSvtfskIiJBDbeqnZV1Q+dsQKeVOodehbcvKwirQP7DrEi/KfKLC
D4QTRdr22C8xPGrWsBHMgzdKA70jJVZkU8fYObhIhn9mphybNUyYa1F5DR3kYP4y
eJlGtcBYdwUCy6nYGE907gsIFTW7m88NtkddnFrIb2rSZ//FeerTYj68CCRBlkXi
nh4R16OGrQ6hRj3/XSaH41SdLOFxh+O9E3Zxe8Td/spUObIHLsxdLF0DkRaMGKyK
r+hBj1X1KEIf5pWeN2MhRxMsUTVYmLQQ5r0fHfEHfsiWiOEdW0L9VC2nNokKHArq
quDswCVAt3Vq2Z6xpP7rRrkpKkxs8vctVtDoJxy982XD2cKw0MWl1b9al7D28SVp
TipXnWFK0g8/eNa6QE6CBxSikHJ8ZiMfVcp5ZudVBgTKiNHoGX5yfcsBvifK0zV6
vDOw2UE+6OnLKHXKW5ewH5IBcNolh03CI7dhk3zaN1Uxqx8QbIAdYmPVk0dNi/2l
djDgvQADuJ2uNJ0PvR1zhynR/abnX5zKjgkdm/zXafKGzUhaj23U/RaiIv+5B7Nj
ARvnylJN8l3Nel9Jg9xw0F7KZSBFcal9Liuw9W/SfI/KhFmhduhyyS6uh61rh+/x
Y/r6Hmb9cie7znGiWZW5F9j3DlZ9nFXk3nhw1DVEiUzl3NaimbVX8AIZMSIqlvmg
bWjz0PAyD1BSmzN00omeHIwzZ0mNfqMRt+TIAs5/I+886swr2R0xLdaKYN627YXI
sa8xcupsmnYz/WLfvbDZhI4Nk/Un5keFHb2H2dLSP98CnsldXkwyWr3G+ZfjDKLf
ZK2qwTkSeb97BJ76ha/s1/Be2+tHWRJ6NnMUNiu1DQfg1oBPWmS0i9dBESxSkHHh
zZHULkvlw9/ZnyaiVqf5OVdGmYS+H+GglRGgfSURaPt0wb8tAc0EeolDZ6cFMdX9
m0LUELWNr3tEJvyw4hQLiK4VOAW0ZFSvIs/hsOJzu8guClQjzquzCrzNZKIC3Ajb
9WNeaV3/XKAF9NewoL3NDVJhoD1/sVb5qhEdyuHXNewTw3GGHWAJkadVay7CoLnv
bCnfVTTzKwDwOjgIsvZj5CZkcfBGBbRgkHeM2Tc77OIUk4T7RDCEVLfTnaHIoMPL
aIQZINvMmgk6yCipoNYo3IYWOiE+kfNOa+84WAGLjISrjGWjCzOQkIR1BCU2APgc
da7HK4+aZgIBJ8he1pB1vNW+Hby6lkIHiOn8JskOD1NcuAIA7AJl0SXADsYwFf0B
NspwMvzACx75MuJ0jMfiGH54C4DC42PTsc7AnJQUrowHLOaaj8c//5JY1KTqEUs1
qoNQIknxGEODTdW4+0RSAGoBYEQAWrQrGz6mmZZ/LTtVRwSbnwbJ5MZTv420UJnT
FgEVCA5PO22zmLgzQo3d0wEZdOMZVDTODkNFuhdwQedFewxjk4iYYVIFZEVOCRCz
Hzm2hNLHuz93TL8siVWLkidAOC9+01CNKPN/D5SztKko1B28jd9Aek/tCloD/S7m
CETUTIXmG00tIxaXOdkl9pzQDAPykJ5DWsJ5S05wi8rG3N8eZIWWoh7jWGdOTr9q
1IjklKCoRhIgtv+gERaMewafj25VqYiScW3C5NHsPvzWWRHhTa7tIqRgt4uXD4yK
f9torXia84Q7XJJHtt7QVMEGkXh/KwvZwj5TxAWyFhr2gURLk8Y0PKRC9N3VwC15
c6j7m68fv8ER2qTZ/3KHfh/bzhrfogfIE2kTYkleZdVWj2BdReUO26N2nKmsFwNK
gqjGOnPKs73U5PuHDmkft3uC1lQyIhYsjypH4bp5SjxZk5GD/YxEGb3zQWSMYFW7
ILWoMu5bee5N5ZRstQxbxC8ToC2As4VfMNI4ZUPTP8PSreaQc4UUMFqaJsCZcybS
N/foU8BFf/mWjXFu2kvsdYY6DvgvPFdb0Z6ukBwxhdWXlQ8W9WvN4b0Z5DucmgaT
Nn3/lDS2/8j139h7FrnbsD7Tx8B/k2OT++dwkxULViA+PY1LO8KghuPGAx26rBe4
jlafXTTnyPGhhN64C1rLRpb1W1kKbOpg58Bf4tbJeQi7SodcquDkBkDljo8TFgtC
fsLCLUAn5peL/TYGjYIGd3xnFfdWPOcxeVl9nkWLqPYKyua+hvM0z8yaym/q0shZ
1oHUFEuySxeTb4XOpTK7MHMx3ERkTvL9HU1SJg9ihfsjtiTZegWDP411HaRa0XWG
7fcXBDuMXN/Hp1fH/+pJ1zT/phdI3AUTFdGuxulw/sCgmPkWLwiE9+yyZGKUVNRT
dgzBCUDcm2BkyjqulqmzQiBK7DF2VWEA3dH/wbweHF3JvF7eBlJeyhZB8mbvs9QW
m6C740wnljsmBsi1bswmj4WSKGfCyoqLouCrZchhUizN0Gd2Tk0PZYkUoBv1/1zg
0F/HvPgtWEaFQ6KGVyboA5g0r+feZrMetXiVc+KeR4z5ui297QtVb/ZNp1VaclYS
FGMwCEcBsj8xuvo7d7sJXE56b2rlrjDKS34bdT/lodxNrFGbtPi8617sY9tg4uxS
tUlz/SvD2BiI/NwUQLoD00JRoq+TxcinYM4q+3iono/AUxKRQN62cPbHnHOlGCHW
bvC/Nodk+YIL1R2z+zx0hsXgT10NOT0hwAZszb2/wGEdhVPagP+X6vn6PnvRTWtv
x/sE0kFqvPyCMHsZgNWgank559fT5udLPIDUUlHewx6z8wG4eOVf0mlAGunQ5Zz1
oQIyHsJ+ywD6HO1d+WMliiX23MOEg9KAX7RlWg60abkG5rwg783lvESxnq9jIAct
py++64juYHx5tY56uJ05wSx6vJRRp/ZqasJWk8kb0dN/D22X1Bu6MwziSLjyLVmD
y2moFfFLdfRHQUopL5Bk6ul0cdUikaM/UWMWoogWm4c7ukFx3T/YknY+n+Y6NcHJ
1yFmwlZIqxp8Ch5R0zmZVhmWREa7UXZHUGzDjUPc7tN3hUKh4wZkI3LXkoy0QO49
B+jZ5nK/5M57oOzveujpGI8Hy77JDmXiBsAyypgXt299H2TbX/A5CxAqzE/cKmk2
ELOYre8+6+qqKl3EbE/1JpmmbZY0re4ywUxmY70Q/cXnm7ainfUXKyi5koXgRhC7
TqnutXmsH8G2ZRvQRYZTJENfw6IXimVh2QPmWgZyX7PKS15nuBXZf94Owt34psfm
9F/4+x17/+P4GxERX053yPis5AhZZ0tPOQPARDG8iXgmBvDOKQpwazvRkrLoh9cE
5lSzdGpsU/Y7nofciaT1r3FFUuwaDVPkrQyZsbm48hkZD2yAuUrT1jv6MDVzromi
uGii+aFGE2XME0jmEUyvxgOKvsBv2XLreolwTHxFoZuBcrMoYk6+AcOtzhI+KH7g
rMOiOTrMMM4k9AATQBlvBuozk3aI82AwgWBFLi5oxC1E2iBxGYsMgCO6KS9EotOK
MbPuacRCi/hQIikXurNtXn3wNSI6uonwSAsXCCHMvNSC7GbHNMeFWEgf62Zi5koG
UmGEfWj4ym8g8c0OoyU6ewkSOvV52CqjAOS4nd+i3fTpKaxlExlada1rWmVOSKfM
5DjWDwJJq8sg7HwWVbk0hbOwT7KwiuvAHyMniQVYcQCE4O2EJ1D4zZVoZoE1X0ru
CaL5jIiQfF3HOx7e4zIQSFSBvH86T2AxFz4FwEUk99+nChSAD8mKhckm5056nWMv
+9zDU8H34S8OFwLuIDW8CF3JdQCNeJgKuuOw0MDUmiAljo/GNOfjOL31GuzAluEJ
AGzm8LaTQ1JxHZ84SkHOkusxG/1QK0Mla+rBntfLDAFAyB4yI35FL3GznByb0l0X
Hpg8FwLNQFXWxSXaZ6v+mn4z6mxTxZNfcrfWwV6+25/REr74nIZkuuRWsb3ElFEu
zYgYZv8Md2uUUnQPJl3FL1hqAaAS285gJb8JHIPlpkRLpaUabVBwipgpj3dk/o4m
3PjTwpPLyc9yuu0rNExdI5BAHJTOBZSXCD1qojbYgckOWBBKeGM4twZD/zGn3epD
rQLfuMRDQDhfcJzs0b7G6fAZqJNh0ArfVsMsW4lp8N39ayp5sSxWZga1Iy8OjjeO
ufXNCwErv83ueLOtrKsL+4QZ00ty08CsOLJbKKfu33pR7SqRIcxi34/Uf5EfhF9g
ertWehH1OaPe9bQbLG/FlRdwcAqrzyCE196Huq+RLKQu7U8AJRkTX8dpz0z4LAaA
Wkw73VE4+ZN8L5uFa6m2+7zg1S0zb2QjWpQwA6bAOqOKalgFCa0ylxzmw4KNCayT
0SzuPLdbmJksKJUKzczItqXuVAK9ygOZpUy2ee8YWLtgtnoiysTv1XLw+hwk0yA5
VcTiTaJtLhI40vWkNNqAecvdYCjNiuuwWIUkHonOIWrjjstIq3u6JZRczbqJ8GI+
SIeA5EZsE+UzHPAvi+6tiIRiwmYcAlDFioI1WnWzlQxu/fmw6o7p1IKDLe3FKPh+
+eVEvg4vqkWNFC19IfRYZ5Ao2fwV9URiFSdV/gv5bfaqN/XT5FMFROamdvheFNi/
iM188pDvXVdwU7vcOADbVyQcJ49+p/Pt5EyrEzWqE1uQp7PbDcVEThtJmmRtKgmH
iGKOBsICr7SjO+r9UpJQH15W7TBi6p1dkTzbI1uqb5W6mtwFvOYRdDeZlWOF+hoL
dkfohM25nyzwxRKOV+/hHtOWAxW5Fy6mGM9hU0KR50eO1bgxefrRpBPHuMHBrBkH
eAnAgXw58u+WBFeqBNypxvfaKCcPpaHLGRlMf7agu8XmgOkBAtiKJrgUjsIOLtTJ
AJIcPjYCPYzCD18HNvOSCcO1QUHanQn7KGgjBJPvuBPg2FHruwoMahsRLv5mXwHc
puY5balvEGUg2CCl6w7KDuV1cJGvpCY7slgYAMufHcq5xnfIR8qCh0gjHN6pW8oF
yuoE1hcCfTz3RbDHnrxHUXb7KmAmAdfeo4Okxf1c2pneD5n5Ameuga8o8UYAZNFt
lvLsJD0grYP1cimqCIRXsVrnqKjKEEJt/8M285SkOjBXvQIJ8Mu+2ZyLkHgXcFV1
M0BzYkgV2Guv1Ah8xxvV9Q03lW0YVYwCdROtcf8ssB8Huh18Imy/uMLrcW4CAgC+
v3+urmiQ/JIXmILb9EGi4h//M90pLT8kp+ZZZnWItJ3eUWNPsOjUy9sE8BXYMRtD
fz5FtJ1Q/Tqqs8qp1SP0u/oEMSSM/53A5rTJfbRn1z437gji2mtkUXNInBvxqOZP
Wsv57tTsGA6cK66KXUFn1kjNR9vugEO1ZrifVrftX7qD6sTLjK/aekhAhrohIrsJ
tZE5/iIOAgAG9JRywPaarukqCu3xRXNK74eFGAVjVLfqYN9kUIufpVZ2VJKCa1hZ
ojJXL8Ifvuh7cgdJvyouyfh4dnz7HhGbwqWTxyderAk3Ln2Yky+GNqyZa61g4eGK
HM9SNm87zG5YZud1g+WYC7IfP9M8eZdbRwOgk08QyiAHT/BEJOr3yZRGM/K1acJF
krcC0Sqsc5oXAjKuVWgdbXWlHFvUBZcxdfQKVI6LRodJnLhOwzAvNnrZOC4+BINE
7Kntd54Ea431KtvHWBd69f4jYFzpRAhaGxjW+qdBvW9AdiUQM50PpdfJK+4kFTpa
4Jr8ggQcr+03zkcIr88CRN8HvVL/x1+z5l5QwH4nK9G6uiqQOq5AksB7BoL7icXR
U+LErff2gNACktO2rIyq+vaDea1jEe7kp3sRBx03zPvLzwy64FfBjkg9t1pm8C7O
4KZ3H+sE64rbVzfzlMAndWEYOW/rf0ul9kLOMgTgGXMg7Ez2gIqiw3dzboAjai6K
9B37YOvF9RWj9c6URoEP7v+O0AZRHm1b5+zSURn6bXFZ1nF/3C43vYZ6SmN1mnCA
shLtNDKgAWwQWd2NZY5xCJhhDoEyKpWG9K949y8U4byv5giZ8r34T0hnn6j7j+SI
52uoIoDkJcqr7sM7iQka6RObB2khn4saoJ3d5QaudUIKt3vEcIFW27WA+5aNssov
iOh799CVMTm4jLbiO+mL99NVLfz9Gru+eQO0VWg7gG4HRTQSENLXEHaQ3H0cl2Ml
e9OQni4WdCJe5Ss51dp2WDdiIsdLDvWoKrWv3utdjM656wte4ZpJbCN2wpBVswsE
QDlfYtEKVlzP3s3k0WEPUIBNQZj9BEViGvv14zQUrkkD9Lpk8+sz6yA3a8oywFRh
i8ajms6eZVMLz1CCuZPzRd6eU9/JxRAhMUXFywfVKyMC6qiw9yRB15U91158y4N2
95yEILkSNCwYNACSIlTPkO8BwNT2V9i+JhLbPCtE4kzkv/ycauJ1Kp0RB8sGpAyl
KzjngHz+K0PkT/kOWbYrFT7nifiBoAyQiEvrbAEt44C7XnPS5uQEsFPo3YiXCN99
l3+wFD6QxaVfZ+dKgz4RWHnnL1yYgBO/H/jrsaAkYNsfbxsmdtD8htA7oyrBZJ9+
9w/DaCD7lbU85c4V5mEGJBvLU9xhuzNwsQIM4b5Nwmtc94vvTLpjjEiBWLQJncNr
aL9SzhKaGnaeNADamiwqRNZU01S4wiJ5/cWYfhn1i6/lOJgfch1CQRMIE+5yHnnB
x3rnTB7T8ZOwbbAym+9G3inw2Dpuyx2Xj4J1IyDNOmSDnsNnK3XL9JtqajZs5k3k
MaEjSxMmSb0AFt+NVJZLKaP8ycx1eL8t1K9AS00KzcotNyO4zvQLlgNnzYCm/gfU
a2SrfVleYx2s68bYTyn33GF5ba6TkoOGExJH7FYe4xHmd8pXHYF5s2siGabL++dI
SgW58WxAUmGw7VzwvEUQOOGKw6nDGs+lgoI7eV9UG6Njl+IhxBOkFPwyOD7srDTk
8TqiYPzmu2UCGzfotsSXo7QtkT3loF0OlLkrE/XoaWNqhv2EEc/RrAy2R5A8bvKM
S95e7k8Ri0jSl32fS1o5VxboeEQ55fJcQRyQks2B6mtZl8RZmn7G0JHi50IDXeRU
pmNIrWPxbWYn/3yCugFUZxHXKbpNJL9V+8K3pdmC0/t/9UcARm7xPbu95+vCrbSu
zwHGWGEBtZK1bgcVesKEyB8siTibkFmJZaHVlX4CX8ynYWJE+MV+9SRh2KlWimu+
ftdpCBA/LyKjKM5uyM9GkMw5ewFMW+fv1jnOKG0uzna0nW103rTqtrTHqtjloBk1
7ojzl8DLlk5Ys/XqplrRZwRL7B1qayk1ol6XmNDbdUHI1e5r3/8BEt/CL157mLHh
4MbuJjUHxO2vNmWBUALF0bRpc+2G5FGHFXNCnZmaEXVdv2+xaKlxqV5w/AOBxXOp
YQNQvdu1eZLR/LQZmmvwbb7VQO9xWXwZnGXH3P76V8Yu4cjp+Ijq4/kcvf/+3LU5
worhifzHfUOIvxu27d3BFzcWQtoySmkykv1QyDtSQ/S4Ueq2MXhvjkwtvITauhbu
VIgjXTK0ja+K4Ghuyh3lgEq1VI4K01zY+AoRn/9uzoIhTfOTMYPfQL3FS9NlPaRG
li/FkOmEv/SxS07CdhKcLByCFLpeMfqjI7q2whNZg9iUPFVztWOBmKcVDKiawAYE
VAzSsjjwgpbvssH75/DZePpktLY9yvjzJZ6Tp56l9/7Ddl5FiRCVykL7U56QaXHn
PQKLKmil1RKAp7AHlY3GQyrAS0XQm+ToliiFaEpWN6R1NLtYMnV5GMymuW2Fimm9
JE9woP+oCgfdKVaj5MUEvoFxnVkyQxgzyfRGv0LtSqgaYsU+Ftv16kU7A3autOgb
38JkVExXNVttCg7IxMoQG7VTLzbPs2Puch1h/4j/KQXreQDrZBLW6U1hqPCqTqmN
3/bO6JzAHxTZTwGzhXx6H71esYFgb00pfyx0ferPo06NaabY/eGp5oBIAQdgEWWH
ysYr72dYgfLJJa3IEfdPugyTqPmofwSZc66xVhExJPMqVH7F/RDP+bqYlnd5I83j
f0E+vnBpHfS4auPrDm4qagKSp/w3A42Gv0Yk9Pw9RmUs4YRyESf8+tuyR/Nkwnp5
nQTcWf1WQiKJYJYMD/sFTbkBzrtfUWgWiKjJ0o0IJG2J6k7fcJVFWnsce0/tCVsJ
Zn/YMVgJl+wAPZxkifc8kGxmNEFjkxAe4dwzX/Uzbym5ivbMdI/yZoP8LpTqyNKJ
iNp3VMYq7RU0nkbS71dEQvdqT3tBfeocPqoWNkpf1NXWHwgfykT9xNfv7cVbz00G
5u7awP8rOX6SgfSeQAIBix5JFl4u+teJdYt12/WEXywrnEaCzwrcSlDv8fqCnCKF
G/pcf11POOVKu2a2vt8baS9ktsLOBwEkQU+q0i0OpXsKsRQttz1DYTMXLb+VL086
4g4p6qXFO2bQaGFlFy3WCawMegPjcv8jflzv0RxGrYGllEz0EF2VaPgRic3Qu72d
XChFOknCi8mtLNVG/CF3fYwGOWiVZObP5YQ2gHS1vEpaCfzjkE4oOjFM0QsUkr8Y
m6fLm69k0ibEIilcJrltPVnqlZd5AHCTnoXCcgUm9n5tn8/KHoe+SUMVZhAoSmP9
Ar1Rq4JoBKZv+S2Pebzt4jaA09rMZkwPsGGqbtd5HWRXTQGJ9lBpZXXUvZhMSyo3
2SVlHSbuvOKdctDU4pF6JsKouORb8DgmUHzzdZn+PEQl9fLW01ziAajyZPeGIRJR
+1g2bIlaEWiiciztKSUafzh3X2gndw77XoIjhKFD+pwNDGgNBHqIcLma7LJlQlxb
g8tyfiiXX6veVQz+uLgvcaYEXK4/0ID9uK1GegOlFdBW+EoGtovvCLZJmHjRiffi
KLQBTuWgx93fk0oCwOA9BohNNRbrM4OA5N3hSV65T8bIbdtFOkPJSLXGNJnyRMJe
VRSB5iCeO7YfHppXBtrrJN5kcyZxPDCmEzEqQ2GnWj/qJIRErgSPlkQiDlm7ii2X
61ZcvVIIguvnJV2g7tAQd1eK/TaOKwoeDg6aCRF0MmMfQtoXJEEQD/9KwB3hliUL
cRSqm/cQICOoaqA06+eVfZ/PeaAdM8zuiQCtZHIExIrZVhzlsedstUOiCg3kSg7e
4h20c8Za+8thnah1kcwXRjUMkKyRpRdAppQPpxSxEXw4EnH74moPcir+/5ASjv6M
vnRXWN4SPFQ3Rem7y0VDgYzGEpYF0QzsMQHryxLZxVsIp8CWG3Ck5eLJ4BfKDt//
3WU0LE9SgpD/hCovz6RNZhgNHscl0D4tj41HI36kzfyzkRWc8fEOoSygBWsK683r
T0qcOUfTPkMQeldx4zRhhg==
`pragma protect end_protected
