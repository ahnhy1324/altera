// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
g0LJFtLsqJftcmwhG4jDNU9kWNvdBlGyhu0grhj3VsieR9XeGlBHIhNZ41U7r51j
mEkkJ/bXUurlT2Mq60HViimvwWcrpbTak9D0EkbwjpMBAPPGeNsfsHdkcQbQrYas
45G26Y5g53Lk1MGy+OSSSh2Bc6/w01GcK2V+6rMrOBg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24736)
u53pMrJuYmu/tWulxHjaoCpWw5QHyk3MFPeo/JKoO9x5GOpbuBeLkuFZGNdAg1ul
P07Hgk6uqy8mhKN90LUNfMBPKF0DQAoKQcTz1i3AFwUFb77y3uO7Za0+ehG4qVsz
XWQ9aZon0JuQtOodv3eruEJdNcTBoMCvXxYkQKMSmchaX6DMau14EjOJiTCa8T05
qf0lUC3s8jiXkoA8uojXtvsKFR14Xzmcrwns4wV9y6Cq70n8sEHD1gNGli0iFUQ3
B7QsUXlLDJQ7I/3Us3qBIfj9VBKO68cuTRFoCp9r5vsB4/h479zY/cLnykCL3vT0
a5oCAdNdIXavbit4yZXVwrheHCaIqNMMk2XDp7eginJKnGHH3d3sfQYH0iIMgwE6
YphT5Y2HmjS02udpGziltz5ymCg4a1exaSWdYdkHLywNkKgmN70ocWKFnWxNihpv
PZiKSogGqyKFEiUrXsc4Culoq66Z0dPsmMQ8rmhJKU+ITQ+YpXCVE1s8UKpl8MD9
4tJ1FV6TvGdpIoO5HB316O3CyIUAu7HpdAD0cS3LkPKJgr9Wb95uW50YQfKC1BGf
5yKwZD/fOV/XTGJ4axkj7AHb7JzuslJjZm49/OoDTGrAQ0an96ds94HFQJrNXhGI
UNB7640zz/rBrEF1rReUd3G8CxfIlZkLS+99T4WR2euZRC3nYlYHQ+UsKfMdb3Qz
1hnsOyCErn8Itwm5IUTFz0Isr7wlfGzPDEnMj2wAt8qkN3Mp2/Ua7HfdbzGnC4C+
9MtGj4XApg22vn/wXTEfblL1Gv2jdTqMedTEfIXSzFX2dQaPnbm4RsbjAHQNNjE+
1LvmLrpEVTqmvgXtbPqN9i3nRm9QDMMkCaQFyzHS3qr6GCThoyGCC8gLfqxITdn7
EIo8k1wZQ9Yy5obEqf5Kd186NDGcHTPA6D7y3Y5+kru9VqsbneRRB0NSOzjbvort
8wImVv8KydXZY4A9Y7WDEOcc7wVK83ALZhHFZZ6S/XYRkP29HD8G+pRuS7bwdRFj
gLivY5B+A4ECPC1oRMuFwlz6Pbw62hYoRZoHFDmAllKsp1YfcT/Udbq5ANwVRcG2
VfPUSQQ9jugc8YzKiPyP9eGixOlDc08wsLPG6Imz7gyRiCCC+soIhtVhRgC6ebBK
eAkB7OYUa9bHqUDceW0ZB8n8HyxZ5fJ5E4Ww2dH/atXD3cZDSUzmOlL1bjqhbANl
mT2ISouyWNJjMLT1GHaNEQEIJdprXRaStEdY6rgmXV+KZa+dE55TB5kWRe0uzNu7
TUJhZcyqKNW6TwQyCM/m1PLnO7As6ceRuJ8dDQUUd4V/D920VYnabewnpB15wM7D
HEp47zVQpkRhmbcI+gxxoYG2/1bgZXHxYrLd2EcSOSRWYIwZyeH1HeaDSjrJgrBb
58KceoiR0VRtjgZpwi0gh4ZCTC7GBsk73BZBrrUxK6WjxqCymd2sK0hU5xw12c4R
dcEEC7w//LGmTST0WtsbfbgHxwSDS97HAk5wRC9lh/h08SJ9bi2kwvvejP72GqT7
NqsHc1ulkSHyNN7vE0fqy21efd0ru1EV71BXx5/KE50dB/Jcq7YNjzFOI2t7UJjx
yCZL7v7sze3Mj9l/JYHCASX9mheuzIYnoPkXqe2qVZ0oUe+GsaHJTNYFrE5/nP0O
oklQ75QR3ZeSUvHpC+m66k7t0tmKyXNH09e/O39aa2fLkCQiFcjIhbsHGxRFEj7T
2IbFb+OKcokJsLI4ycYTnEIKUMw0Af7n+21wXBw1MZ4uv5+iCJR6OHAz8lLnzt2c
Mg61h58Iim83fAh6ccZUIHuD9MeYevQrRwIhHf4eiUuoy8vpn7uohd/9QxHhetJq
gPD0JDpOtg7SyWq6SGJbjro8mZAdAWDRG/HJnTJrU/0JAkH1zl0sY4Q7BuHciMVI
AGTpIy2PNk1785pN0BI2DzYrofAacF5tbMr5x1RuDibd+Se0OGxVf+zidNm6cISA
9DP+osvQOnfNB+mUdDFg4aQv90Tptks65wtYd+WyF1QD3dLK+FvhdhxSkgYhysF0
qOBgyQdQzzgfto/TM/SCyoVzgbwT/cpcbvnTNeyj0uVx7gKSGqDXAZ7iQTwT0Pe6
1tWm+FWj4kP1ykaW5PbNnRfpWnuxCvJ8tzO6k5kns+gcyHZ7lYDfqabWedoQrc3k
xJ/ybfhW0vMArP+xQYRBYUqYvO8f3UM+kHf7R/Hi3l+3/GhNNjRpCy5d6XF9bj51
CLqGS1CdELAu8jmihAii6YYxPBBp3JxuMqdyXvXyGDC8BFrwxK94T4BN/4TInlw7
2tzG+EPFseg5kFyJQBSd7vrVFB+d944TD4urtoxUvBhPVabild2VHtoMha5svyGb
CfXkIPVxii0/JVt9cBzHJGc5g0i0iJDTDNdl6XPSmRY+NV6uA3OoWLk2eOlDm+2e
Hexz234UUFivFmlYK5q/ps3V+zFqT2DHZs36HVifQcIT1va6HUPmBmzUeuZ+UTsB
AKLo+8wu5PYzLx4oZNVMXz6WV0AdPvTWpAHZSwfv6476LRp0MKVvHrY5+YsaiOr/
exkVVb5sTx+xjviOwRI/8o5EOZxHoafj0+7zW53ilmW2LxQZu1U1GYMTTRWbkWYl
/BvGWiEbm3DVAxXX1vHsDA3Ck9zKanaBoZxfC8srKGZMhQ0/hgMLsV1SKUYhBl1o
Mg7DlszBnSk85OWcaU+6UOcVbkyDdZ3OkcYBIY29XQahyzqeZmjnmAI5hLZgHNUq
Sm3TrTpUotTjowm5HC5oQNcSpt83QrCBNUHHZSWm+k5OqoCaFVhOWrXAmeuNzQ91
nTZ8nz7Zg7xVXiv8hPv2EsUPcHmuxmauiEzn2B/54NpnTPAjTdwC5/6uteHrFnSE
YITKtsQZvXA1VZE5dfVxjXGqwwjTKHsveQGe+hcKKquZzcAujvELJhCDrwc1HOf1
WbI7mL+x/sxhcQdMsbNYu33+fZAs1DUxFaIttqOGHMRCUvk2gL/1XE8xJm7iUdUz
ODNHUOJgiTjBBLNGYFXI5LUTEpWtLL8gneaU+cgw9gF2gyFQahSPaolletM4QlMC
zTlYibCMBG2L6+BnW6i8RfJyB1/um4jWSfreTYRLlgufL4hMxs+P33VLC7rzfL1B
QYwHcUMKU3olb3xgFy0+1XQuRoswJ35CmtNrHFJ3qN/tlv4NmOBfDJe7WkdiRh1o
/NeRj63e+zieM4lfS5luI2dqM9rMVLOfqnjdKM7+fFnxnVZ1vQuU+cIy5CeSjpMD
7BX3WCpK+dgUc9jqQ2XVDJERD2AY74ycgdlJ+QlVrjyNciyZ9VoB+pRYHXjhVR95
WvjdwQU5KNpVQFcmrorD2zznz2B+r4UZIMzx+FpM2Pkp11FUAuw3HY3vTDCd2vni
WsKh69l6RF0fTlUf8gNzRWH4dqkuKAGM5/D/jwEVyOjzRDjC/UtDLD43O/rdK4J2
S6WnjGAPjkNl4C5HpqnxjsFrLscXg600+byydjqXHYq3pgZgnJyqtyBYhxlKqdpw
1H3z4ITqA7pIKLGwrL0sAnbewvm10KE8e8J0JLLspGfKlUwxgqWTaZQLB9P5x6U7
lKw5/dQSdUQEt7oVaCUwsMbqh0U0v+nCZ0ETCgL2GpHAVe0IU1zdE255LpjL96f6
URVs6nfWq11kizVIi7lDP/pFR5/5vOKRIpEh+JlKPXufVPUQQAnGa/wAZjxS58Ld
Y5mS0ipECeqrog7kzDm0NMva9a9V1TYsB0b4Jv/yxe4pK21sR8GfzpRm6Jo3QLB4
E/liSl84+v3cpp94oXUtGrYWkGHOs6OespcoFKHq8XtU2gsKGTMvqH6wkR/fUyRS
ArfnUtT7q3y2Zzo1bQv6PDZQH88slczI9SnQOH1tkzKly/UY663CaW7/dpkxBENA
4LZZ3ZzaZ3nY4r5tQJ0x0I2J7cWt99oPJkGNCpgDXEEK6vu7UchUjm9Any9pf+8d
nr5yB27vJb/eIkk2tapMHMZCHDXvT1y8PTMFvMOEBXBVP3h954MIFrWdpkEPCsMr
5X2wJJF9zJ4Ub3UGlZe4rRNBXbUut4JOr0p4CbWnLW+j4jXffGsksBwDEaDSCMGc
F2cp0OVmhSeJCeGp0A31J7/F1DVOIYTwGs9G6Gjmli+qyUKlIvAByk2xEHpppKb9
LvP4+6Rs4qmCk7N0v5XHy4vLUV4/AfYdg4eO1xmFRDPbVwUnCT2w/GOlCG9u0BmH
JkdWRwuf+3T3/DVaR0IibbHIDhRfHdrhCepang68+sac9UQhidBgxTkSyTiK8ju0
E3bXThC6auaxN0IAuD2HEUwY7UI/0EjK3m1/BlC4NPK8GnF+/nfJfgjTxF2FuUQv
RIohramPBiXxIJsiyNZ+Q82efBYb4SjdRocKVjPuqYgzXHsWmq3mqVDv46q+grEC
8i8YZdyWK+/yZbC+MlwfWEG6P7KYw0VX2e8RZl1dRVFSFYrMMZqrLW+eB22V0oJN
0WMo8Z7zEX+ZyAw6+KiS0kLJpuT3RhGqWDj5rrzC2m5zAryZDM0N+esX956hs7Xj
X1kju9my0dN8Y1rmtMWU4LBn5jdsNn375dT8ufMjN3XNVr9NYQB468RQomaE9zVl
qLYUQJLbqRIk7TZvouHyqYYjSQvCPDBPDRZidgPBvQcniPnPSIai9dE85Jc5mE5e
Au+TEnTKwpyb1KBACZ98s1B4FBJ5s/iJpChA3IUX2ZlDRzHYHzv40skoMqEhV7EV
33cBbpNffcBfIHSmqZzIb7snzlPTDW5xLOZ1QiHwUEeGuZLkD/YpHrlknLe56XEi
wg66GgaFqpUHUcF+K9bPRW39ujPDkc1geaTgmuET8cDb21L4qyVooG4/1sW3NarP
IR542qu+oCS/XTvKav6jqMYbhjSoNz30GJYui/mpePy/evv19ALor7Iqm3wMz4o5
x7QLO2Js3HKBCA4boNvjDvxSy964cg9UnJlF/dtMh6iV9xt68JKKSZr72fYKpdpX
YdTyUp/fq3Sbz3C64I698voLWNqKfo4RvICnFEsbEgmk+H3IPoSAi4oup0EpXYG/
1MdRTqLsokSvTCjgdAro25Ji4//MFWFusB27JWhSqIPWenRdi9p3Ji0mBw5uIHQ8
5w6QIYBcCFEDHW4PP4IIuUR40jJGXO576rdsYH01Ih4pHI3QN0t1KeYE9xPOZ7xL
+rQDVNZx1Buui3m7UEHNEnKRFR3jvSvoRcR/TsFbuFS2bxtAkXddZPdL+s2Wne8j
AWcy0ypcThQ7ETWiPyJrDLjzz25HDX9X59d9br39dSVZ1RcO49C3AcdIVme0zqtN
81uLtNZl5a+xzIho50Jvt9WA+VKk/A+/gchdRE9Yks2O/XPxBo2MGdUCwPwlkjZw
ftJz1ITeFi6nUfY9DOiB1Q88H+xKr6YQrllWB+jCdq+X3ssvw8NcJhuCRns4xUO2
PRu3xsxUjqdXHMvXH2l5LfgyRs0Jk9kmARJWzkfEm+zG02E8eX92WMLn4D5cjBBw
qXMrA2RTw3cZs7OZcwfCrTomaTUqsDtu6Y8lb0xVq0A3X9MA0oomzGc1NhTo0/5Q
g9tiSPcVYpPalDPRnXew2mKceAcPbI+en+km8Dtu3vIlYFq5HaJmbGLjZxGqCYqs
y0hOSuKOr/eg7ASt+ohMIv9Jd/wwlCljD/smf244IxxTabOt+0NbKIluTwIGbmtV
ANwPv6CJfh8Ro4+X+AeYZQbLjYzH16o3D4hAawImOVV6+J/xqYagsigFpBUV5QvF
T+HpCkRhBUmTLB7Z/aWgYWHEp2Kkb1ruDNy46Qa0FqWsD8E0rWNnKkHStPG20YTV
Y+ees9FiGASppy9KCWJhdYx0/ew4IMAf7kd0pLL95+lzmk0+u1j/TH+h01YyfYQm
tTm0tRaC819Oe08xXM9hgCucfkhF0gTMN9qIVPrNENssnhvORZC7igS9Ocrc/xWB
Xk0lDs/Ff6JxfG26deW0EQfwAbqpepQV9qfUdoYu1VqPhB1OsYnLwwnFtOge0WLn
WzpxOX+xxFB4Nqv8CEXH4dB5SVVtHg2f++gbpaUzoJZWgbm8Ex3hLUGCioCWw/nS
8PGjw8Y7I9OOZRnL4pYxh59s9TRDO0ckQS+DtV+DQwjIOHe0ox+7Kd3ULxMXXvfg
2yftkyz4gwSQ4UCaIvmk3AvvCVcLWg0RBDdtMgpZIAGRosVRU8PaucYGTWFMuOCV
mzK0teL+e/6ZJDSi7VMIEHlEVJJs0PxnbniP36VLUZ9VZCYO/6a5zrLCIp+RIdDy
Sx2K9Ems9vzZiM4Y2wd5/N1xQV1tMrn6a680ZhGjZ+k/te/kHQiZwjt7b0Dqn7bK
ytf/FgCG7JDytIVqy8UnJljdoSerp08gwTLWdBY01E2TQfuVMdveLgdr9rcMPZn0
UceylU+rvLORhQHYAxx6xjoWhcii6l8ohPeIjj9YlDimEHTGfoB5GiljGn0xkIlh
/url/t59rNxHlOYnyyHhVepsEkGUTB+V1H2gPUtNHI0JCUMdiw/dvEgNyBmJ3qdI
53sj1tv//IJ5gcX7uYqvJmgWZ+5mKrPAvXiRV0DRCh0lNhTMTUDc3BRdaApz77BA
yCZZiaQz+FD3XQQVxOtcebgwCcdN39FmD16C8B6mnKa4Bl85KpCGQqQXbJtnifaL
tUxws/mwXUaf2Omg287TnAhI2Dxz1Y/HCz3nrGtYozcQaZtI478/KPbWkD0Jn5oL
iTI8uGYGhW28c7CLaOsGgEm5DnECjBpcbH2Zfcx9Pnx2Jo2yXY4p8gDNoKbIlB0r
nNXkXmA1aZNPJsPE/PlgbzPBKemLb9X00kmL7/odYMGFYp3x+d3KE6Jneefl0kPm
1TQ9JJNuWuIDm/JIJY6xF5SKX++NcsymIy6/DpsXGYO5xTfuVAsvtq2rIukw/aby
epBAOueRCOJ6WjyvUtugMvY60XVbirWXhWQxl04RJWUNNmBbK0XK01cMhKPXoJ+0
izSaDlzgS+euvOGbbogYMqAYYz4i320Q+qMrTQ2wq13iI3hFaeCeTHN+93YDuuAq
/47hb8lwpy/HxDMwaT4YmiefJJBHdQ7CR7XICPLT6VB0B9NDUHdtYcOf298aOFp7
dMgU7ZA0ATBIGTAqMpBspWqXM9zxlSfo47sNQV8IgF973FsyOK/xXkAtrcfeLzGk
9/EPCxiklwmRY5cvF5wCEucxe4i0A+ZPeQOQzucZhRbunenST/GgbCpgsJAqBxdz
pgt0raWfYoNgnflHeDc+jXRLjAqGO1bYLKyEw8Qb9rhhLxZ2qiJc8mM5l8xVtiLr
T8migBZ4QiqcmsrPWLg42RaeYrOQDdesL0rHk6gS4UqQuAx1QeqzaYERl68xoegW
evgfT7Z68maBs4A2mYlTH4BKSHS2ewbqFBv+3AgCju2+MFlQN03SnaZFJEsEj3Hw
1Z+J1EF3+SPigMJAJAC8QM2rjVRUX3aC1sdrUFjShsfeUW4xPH+yc5WB6yMxino8
RwyttiquW8t6gf4JLKifNpZHp78u4tIzBJKZbw1LzZl/i4p0H5S+4rPvisBF4x2B
9OSZMtOqm7NN4fXNuOaIEShukgMCNCwJMpBi+hjc3TjgkpUulp7fLEb2WHXRS/bD
+3LxNpFNnm9jf/qW6CD5Vy5syyKpFAaBNQ+E3xYbnPyiirGonOYPuoJFHdpiYDrG
ZokpR2G43I6B8+UWVL9Ru7KycunBPYuX6yG0MD63HeCsQWURflLcbvpMuRZq4bC3
u9TfAbPndC03dfMK4g/Y95grgVGh643MJ4eX5dg7e+qO2T85CawEYdzzyP6bgmmB
qMxFhQ1j94RvszIb2wSs/3rtJrcLDrbL+wMR4Dq+VJcU1EgJTiHNaRbUj5kaXIuG
J73uGpxV96jJR0x+4k06t597zOswLlOgYn0Mwv9sNTFTKj5hJ7pEaxEWdQuOnJau
BNKGMTWrGQoScx6SuRcumtUmJD1GXrFYie/SV284QzkAvk/ZJgl7IvcaUo1chcF0
8GvVVTsiW8/2naPRnQd2ylSpdb2gzWr59YjsswDGNy9WD4KBvLihUku1qOYW2bH4
G/gN7AOMbHFv3s2E7NGjm59vkWiDhv0Ys9OSkB46J5eXz80eYHPTIBK2Zxfcdlku
0IHC/tIvh+3iJj0khZmaqpLv9kR3VE0B+l2m2d/CvDRHvZOTF8asI4+nfkJ9kGdc
sQELJ04aDTt0wm1WuASZ+PED/jdBVS+ByRd8d4v8c9fiI1vbPKrJ6tpL6lMzc7bd
K+dwKpgb1oPPxthfnqi+7kAMvUzi5VeO4yq+FsX2Qds+A2xmiJGrmgq/OND/iIzI
1gd7eLwWv358UQ2tJkrWv0HzVuZMs9PqbZIFMfpPS6ldfQpFdIKrU2wIOdRuh6h2
EOojMGt0Qw6gHFFlz8GCvxFL0BnFSDN1OV/e4z/r4ObcmCXGFFRM5E9i7PlR/wqd
viRIMI5jHobJJf/Z148cOHznBDpfx1nHtqi0i1XbVNHOspzc5u+DWJVIupEWsXhu
6PLe8zoL86HOHil37c1nmQRii9B3pMO4pVGndFkXMKnXPID3xCgv3/dCL9L50JJZ
289pdr297gz9O4PPnYjgLmip2Unabt6xTQRtP+FVORCne7DVJxv8LV7/Wb7MzZJL
qi0Nli1XtrELDaaq/lzuxhaeXEuxfuX7lM6tQZg0vyOyT7SekSEqcPc7HFPr6M4T
1RKrL3NnORL7cLJtd07ddWGd5PltZsM8Fu37BD7p9XYeLr3ZEKoFeqKXmwrg5nY4
NMTILm7FGQuWWMZ6xheGgLP4VqQvqDdE+PulcG1vI2wANGmGBqMNNMK7yfvO6RSC
MG3YQ4jtA3muEf7xKRZaaqeEmc9Nqqe514S4SpnWh/febXfuMg6beLGr1EoPLZLu
ocmPr2Te1Z7zQTIcWB9/O5V9Qlpfeu4MoVKa2h1TSEGhoIlL3tlLUu8ziTbvcz7c
x+XRYCcAN5DzntCYcBiC7BsKpvCrouuOyW6zX/8udpmL6F5NfAg1AlC3Bu5rbxv/
tyglMd50X6XQ1bx2OlocU9V3j9Vou5v0MLtGpi0uww4E1nWcivbXyjhE39kApU1M
kml3DE+921uN/cW1XGYElpGX636FhdGQ5fvHfrGjEpbxuez/v2i/OFiETf6xVp4k
m1E3f5YUBoVPJVXag8RL/GXV3ZNnJ/DEn7MY5ymoHE7cZcN/e83t1a+MF7fJ2jAi
YjtODttXEMh4z1D3U7M9gGJ48K17u2ZXNjRwvz/Igu92+LcS8ue/x9A9Ac1u9cjr
5EZtBrnrgC9Xkc+57i78CGrGh02QC9Ew5PKeHapspZAvJemvzZU481tPsTIG0IhL
XBYfe0Pbm1TbLsQoVU1KFH+JSxu9sUqu14rjTxsXxOP1l3/F7E3n7zHemcbN2ExN
l3YAZlDN0ufQJo1yRTMSAB0vj/jzHtOscaxLvQR0f4kGSZe9HwCtMRWOIif/ACs0
hVNe+E9u4/us1z3AsBB0t2z928oRHMmwltdBEmXYg7sdvad/tzetl0OWeIeI1QGG
WIOpjWPjMY/ce7H1di7zaK/PKMZibIQgklT7FcqTBsrWW2LuOoihqNLGtUbz/+Ns
Ceiead+RSDB+HgdH5nB4dV7djEV7EDmr5TwoGmcacUu9hfZHTCZaVsw+qZusXXcN
uEezJWCZAGlVyXclfNgw9YTaTibGvmL4X1imqXZVL8dw5EE8+tr6ati2FTQnufw5
UGwaR9YMrJOIAkOYJXK2IpGccOnFmWv6Nb88ZtRNO4Dl2/ZFrOwAU9kqo+wXEfyl
0puWr0TRl3RHDjDgTBvXf4vftaBj4BWaztbHFI77NJEYvl9d5afXyvL9eEoBj5Ok
G/GCErbD/NMEMrWLDxTW/UAWgodGwycCOWHurPFgJa7B2mQYGIhnojZWuBZRl5p+
lCsXqn+Nc68Fp9NwM++UGoVsd7q8hpR1d7rJR4tNbYUwIcWv7qlmT5Xe5mc6CPha
L3zKLA/XpKylvJ+exikNGwhhL+XP3wdAY+1LNsR/SofxG0kRKlPFPZQqhzDqGqHl
pIIYrzNZWhhZUdHIgRI9FrlXzeEC8V76l8FTXEQwTmsyJZNZdO+WidW3nn6LjE9o
eog9AN1VJTEZBJgzdx/znAgB4stPrqUOO7Htu1toRPwK8capYAR467n94cAfjFBI
WNU393jzBxEKM7mpocxA12m9mubcJkOhg2/QZM7Za5P7g2SR0q+Uj9yahRUDUW/e
UUSicrFdbL/x484EGT9IcN2i4K33xiRlw7Q1MOfajazMq37qnS+dKXMIyChqd+KV
9id4/7Fcz2+whoClJ+RgIiEeUHZctgt84Zj4oTFEBXzuCDx9qD+lI8FSVsHd9B0w
BzqO9zyiqSe+nkiPmWWD6aCinctNNQVcdMGWqS1j1NM3DAr5eHsb+ndxBQrBOCyH
e7rhgkUdTJb7z8/VWre3/BTjb09GZgDrhkQRCqcXcn0dtXDJzP4472DRBGePPOQ2
SsT7doJApOrPP5EWMeaq1XV7hQD+MqaLQgSP1c3TSFyU4KuBHvfoUMKz4WnT9xox
c3cnspJpj6p05PoNoP2+DBDiSfRlOd3Sd/YATZjx3YO1xaGZH60Wev3ldT6ILn4W
8Wyo8COpp8LY/qdRbBVxVYUKohiwm4M1bYmy2Ip7nG6Uyi+wkbugnSv+5F1ad3l4
P1VEgHZeY6+vc62YaT6e3PaXTW3fuqi28Zm84rPj0l3e7ouoYTIWYhDjsOKc2dTO
686gEfxaX4HExAUSMwcSiKOhIz8OSMktbamlxqluggYH/i65tFkv54ZdQsZ1E00Q
zYZi5Ly456Khet2vLEZvjidEQrXA4Z+QjlaPHmgd+rM218IkZ8y6wHViD5uUy7TA
95LeCFUMGgS/AnCuksD89+yFwjsRzRtAd6afa+Rjr8GTH7YV+QcW/m++HcvVwGFk
KeNBsReLCCFvcN/sBxCfL5Db2pF63JK7L+F+D2kNXVDshaGIszt9fZFfFtApvGM1
rhYyMRsAYjGtCmMXhGSPItT0MWyOtOKNSmPZ7imYYYGHQYGlTk9zxfYj5LsNl4eD
VHH2U+iaqRtE3I1W1rPgcmr2OByZj3I7Vz5SmCXTBSHMIJe+SkCHVuYWmTBENj5g
3Mxt6for5O+LsDW573OjlfmcKNxYaw0bT2VtWVnwRYFEw4isJ/OC/WWA286qtJV3
EqiqetT8xgN/SmxsQ1/aR9yhWCftVfULVC/+cDsr+q0aynOS3oJMUafxc4zUzCaj
MNqOftWTVdO2jeuYqe4RNF/v87sbk0cdz81C1jI7ZfMYbS/q4l6KlfMp48GWGJsp
dMGM1+WRdOZseHGoB8L9F3UZUBZedxECV1OGRTiGi3uXZUmMUjMxHhhycMOsOt6u
u81hWwlk64n3C/XHKXvUC9T5Un1g7nd1NYuaIRNyKTI30eHoV3MFOPHUX6kiG5Ov
2S2fmGopZatFLloGmLZhIlB3PeRDEYlpaZ/szc0xI0gmFmh5auX/BpNwhGJx0dvq
sNcLYYU02ixG+FU/fXnhCRzP7GSXfIBelhZU+0OtbDebt6Us63WUX26gUOlndaaC
iMcVOH61q+p8+jravMMvQ3N5AOLubeaZRqf5cS4oVLFdjtCVR1oEy2Z2NFX2w8tK
Iwjw0+w/RN8nqw+GrrSKEFDtdUG1RGmcugJTbGT0Vm0S19egsTFiNNQc2d5yIPzO
FHKx3okAu5K1eMYzV+U70D0wZO+L8Yw40bIQ6c5sTL16/+gwSNwiIy/W2nvjeS4/
tk8X5RhlxKyKC/h/TtLJoaa4uXsGwHO/TF+qh9oWK7fVvpKPsMbQox/vicSXkdk7
XmluLMt6hM3Nl6LXJfuzwoF1tGlD4ggwuQN1rwFLfJQC1Kkzau3/40EG01gfGhOO
BVWxCHAxn1LThvmofklopYPq43R0TBEHAP7662DChoDkjRjLy+WGmsF/ZVGROR5k
7IDcIeC9xoueag5Y5buggxrn2QkSpjr1GdgvPSTBt7e0AWFREh6Y9QOVJ6ZlVblL
GkomOvNXgOQayde+Kbd+POKflOccJaBXrUexlBfr5YOeDRqT7Qho5ZC9KX0Cm+QQ
CuhUjqcbuLVe89YrmMFJh6lTDEAui8RouZuUcoq73PfwDU6fe0LtoTIoXtp35VrQ
8/PI31FZKLraZqk+UyADBr3Y6FOLuYIASYqsadTytiugBWxR+JbAafDAL/ilijH/
n9GRoo8Wq5/3lpGJmhpSyaueWGZKUajsXF+bbldrGWDW5gGKhudVzZR/epW4QQJ6
RDH69X6AiCappa+Z2OmMnI+gxSaumvUmZ4qSjlJv7Pjjo3FetoCUc73tHI6E5hGt
W/AXEe5RpUaeEjGLqsfnlIo172HWICrOUksDxUzdZ9xQqQ+nls/JST6C3NX859s2
ZuoGY4wShIZj6DatKJAR5bJXzV4r88eShQthQj9X3KL1EwAq4ewqITmsIXy3SjM+
H+yEeEBgbicgFkG+K58Kx21L313ShIFWVTA15NuvGgOcaBW37CjqKa3gfenn13Vo
heH0dVJGOeqJSkeIC8ozRDmeDplg5gtwyySI0gQMlb9YElq55DpSf4FbV8DPe2hI
/f14R8+I00IkdBUUJkZcLnbKBjH/bs+KhxrXlxFI19+tQj4cnBccDA3mj8IoL5wp
keeY23orx/1mwByUQbRwW7hXcxgLebxA3/qitIkFntagSbJIIXvNz5ew/OGWzqIY
7fC0SXJjlXszAUShVGOXEYXffApBNNW8nB4HCng+KnsubHh3iinnV0vYTHoXZSAA
+kth6tDhNmJApGX4GjxItZnjb4oDNJHhtmd7RqtyxI4KdKSWOGN1GGe2h5k4kw0m
sCZq249OYp1lsSdnRmP9+5HZoAuBQLWGUtcOCkrfjKLOQwsbsyhCc9Zn+ZSbwTSR
9+0c1C2bH2WwkL9+EXlcRhXUp1AvbTnd7b1keoN1IW0UzjC+Yyn8NENX6dXGlUAz
41LT3aPrZ3MiLdSdn0luFC+QDEkvYNnKGdQhAa+MNVnbDPDSaTEcZ76GMx9bvZSm
01urlc66EARBae9tcFbGJeC3VJZLdo+U/ZUTmAuXuatKO/FhTvHmrNw6Q11rbUaN
LAud7+KfMsefVSszphPmZ/wMWtniLWyMPEVohByTp2m3289HSVDgYbWKLY7Ktalm
hKYf42tUbDXZbYrigsy+DMvcggyBC01tnAE3poGf15ry1OVhQ74mK79VmIdhUv7J
rxFvx0BRA+B50Sz0plLx4Ud6wo2qKObzRNnK3h927/pE+jtQWylUyUcJNBnUrAr5
IIXUtct2KiQTxhUPeiXqr1flzXCzUYV/PHz0OcEw8As0KX04dZ6UQmaCZr2RZ5Zu
HxFOAHXjnII2L0vANN4K+dusMS2zofVwp/x5VeOXnBCN+OlItL5vXTLe0wpcURmp
OgKxEQVddFB0K5Xz570ECRzcWncL9z4ffchB2XTkSaeQ37Swq1wCPtZtj0Y7jowI
e+Hb2CC+KEdXciTaI7nWaF5PnqLYDo25UL9/ei3iSjFoZwOsvCGL2Tk7poZMlLKC
wM9y0a9De0osvqjXTxBI3t6l4XT19qNEfxLt4n6j3pTvYlnsdbPqd/Pb2sR+n+1/
wF0gTEQybu20LKv23aZWPp5RZ/3lcHVeurQPiKs1GoSKCmnAXXgLag1WFFOsQS0E
IQPYQRc++Y6ek+n+MMadt94I1Ps64AKiLJ4eNi8Wj5AluLlxjndxegu3h5h/T8I0
tUhE8+ydNAVJM9tpaJiSOtnjor9ZTq5JpDzCdYfTxKIF3Nc7fr6w7hcaaskGqYQ5
RRQUc2a42bPjWpktl1A+hOYrQZHiC1EyYseC4/OZI9PL8X7l943jh2ki9Ikbm2t4
OxRmo6eIfJ3IsFUYS/Q4IhYvHfNMd2xhORGM6C0OXgfs3fFvBNxZV0JY5LjgNWFM
R8TdmQzIiwK3DbqLOIYnPevDiQYy3bMd6OLSrK8zRO/e0A1I1sBClixSsb7Jn5If
qI9qcVUAHUwhuJR2gcgBwbU6hSUjhkUQYpMzY46YpMuziNoF+jTSAjqk1r7LBaHb
yJ9tviV+5dY9ubSRj+o3ox5cai7pQRDrXZe8a8MUSMY86b9nqiYG/wL8/2Mvrk0p
9y04Gp0wpV5/d/ZC3H9NSlivvaphPPpwik7h4OVjdagPZDvP4mPkrQGh6PIzbqNc
10NSLHYgv/bpzvNczGaaKsmdWNcPnoKFZDanjPLOI0zh1Z4ffpU0L+9i3X8UWAeX
WhTWPSUWYB2D9/cfHJnCt/bM2hpx5s1nmebQUbbQ6sQpquSlpTIwQPvgSX9sC70G
isVtuRZmyZrQ+av49lskG67vC7VjvUrAjrFI21iv30UwuASS2MxbxaIwOptWxUWs
wFst2wA2yOKdiPJIFEwNetvD2kNvAbtTYfck+bBMqOyOtJMVtL/Qd3sK4UjUDPty
aR/vFDOY5zDOTB51BB4XUAFI47tJ9/BWseIC6nt2ikuinpUea7WucNkBaY+luVne
zSuSFn20nV5J0eIx/zXu+gmsXE0m3mxGp7W8+U4PEjJ4GWSJXrm0kvNEuZ2cTFTC
YHWazLJtu2r+/+NyDmfUaSCXFgHCDIv6FErhfHnrQFM6vi2AEGn7H0PFPBiTJPaK
lWgGuGXZqMm7wMvIceRJjXVZJZ23nakX7IPqUVw6gnBdTSaAYmZCO0+KXzI+st5A
S3GnFHrj0ORcRpJC+QLpkwDurLbb+EfFx9Qu5OAS0OCdApKgJDJIv/WBP31UQltw
VJbmLi/SVxCJsnZhBq7ipp4YRSvv9ecH/fUZrXTOVos6RcZMiSIuODoRUwABVm+7
rQyqmp8NyIXLXesOgNzHrSPEcZ7QuPElmrgL4iJ6rYfzSMhaFjPcHuBRSjZqpOeL
MTWyAkqc0uxiw/m9cJnSWt3z3SfrSxOpZFx+K4ktELlHQVCltdUqkJDwgXFdZkqr
NQM7edOxZe8PyaY7x2M1mdDiTwxnvqB/WnTBvSc5MFU6lyu6VEPHovnL4HRPjmn7
35WpGxt1CKJDsF0ggsnMuPY3cUwp5gQIc94Mk/faphANAZHUdmIPFrr6QKjyizv5
dOCVD7vgVRfYJJcJvRdB5l/TUNqHtsZA0zPe15RNr43nfglLFsf5YQveuwSGWK2P
sjcKMHfie2CDUBi+21BnN0HoR21NjecopvkV58VBXvF8UFoRXRYeMiBBxfbwQdfq
yPTHxi7h5L7//ezqJyBcYIczLdQwgk3sTHjb+RnjrQtIP6Wo5axXEQSdjCk9L1Xr
ecTABHQ9+BgMPHo5BiSbAFvqS5DyvE6mzuG6mj5F5Egp4nHj+Bii63SsoIVmRsPa
pBXdsVqNgsnvdmKb7dm0//I6jjiS13VGP5LXSTyJ/3V8F+1uAjNTRSniKkxQoXCG
x/wj4n0Vu1b4L5gO9cBkihkUTesk1dq547ADgQ+TgjoXJSAldg90gue7LXIypyft
oux7uxyeIh85fN+Wf2pb5ajgHnMovPThsZGBkR5bIjBGx8xjsXrVTlhqjVZR7MJB
hPygYL55AYvotku/li1cWd5mZRhHjRxlxGF2Muu/4xTxDRyEiy6/YRh+AN00ithw
SMpoXwdFbf8t7spnuA1lmPeK6fyLTCJz+CkMTj3j+toxPSBjywyLIoB2ZrD0ijeN
frFh1hrp5ReRGfvEkfo7jkvgJHKNAozKW8cgFUBGcDtDRQtWVwmVbVNq43WmZ/hn
8UCffVe70fnw8ZztxbDESS1J8KDsuHv/HID8uHzOW8WZLWEzy0vuvtIlXyKkcxdN
C0FERmYLebQ05ODt3J3EWenLvsfmCPGDT+nvwdKjsQh+AMiula8mioD8jhDG80Z2
kwwkH5BjEhuqtCd3QseQ4lyuzlj+VAp1OK9hK14adBorb/Vwl/RYIIu3DwVkESXl
tzXcF4rrsc89+/ilB/6qU1Awz/6H/TJY1O87oS3r6hfGBD8UGsCFFLm80D5YZ7IJ
Z2i/+d+qHUmnleUoo3P3CnAFkOJX1POYoGlkfWTfuKVpOFxCAUv0ynlUAmQc9nRq
E8OuWIRlkH8UQjeiRF1ZURqvHBpiUJBaQBEnBPtipjxqVvbefGzw4uD5i+aZkyTG
o/5+SKA1xP+NJZQOkgAOh7/sP19lG+c2k7l7tCaiLp0IKWuJ0rS5pQMwf3Oi4OXZ
t/CJYdBPja3Ycg9nV+33bI0gxMJ1hNxZJpnw+33fS5ztegxSAFJ8VGHZiusqodcp
PxbSmDxzToUKfBfP0HBnuWWpZuIgkaC6H1cGaZNBserePJYf98Oy3POmHlGJ0B07
7OybRDxvZJjjHgUgP1D7zyt+hpwG8/sa97LfbQml4i1mzXutND3PdZQmH5UAvjhj
8WrEYyJurBGmCpQ23GbP9WNabHwqEpeauP6FGX7+4+lpwUiomAQTmI7pT+d/O105
A8qAc6UpaxDtQvCw2NCfm/iPEnEtud0u1gj8vI4p2SMjeFTRQko6EEE06krc+hPf
IrJO8Otoj0vuP7p0TOrqvwtvn/ZqDk5SzCyetim9fJ6ORpQZ6QM68KFGoQJ+QKF2
f7QXIr0mO0/1bTqC5UoE9rYL+XxvDqt1YnvzpdbBH+BzZNt4OdW/ao9RaUmnl9ui
Gss504X+MASCSbTQvz8JduKBq0skqexfox3iw/URfl3p7SLsnH+/U5gBGYLC6U1K
QwEF6B0qXDCIVbkcf0mV5UPnxyIrJCAVejzFHVvZLlZ6En7NpGiRMetEx0T3Wg6v
YMBHsE7RrTqQsXtYdNjdvb9CYqgtLZHjMFlqMc9nvBTD2iYfpysM7FEI9hnmTm+v
3F1OHp8kUPezkjZUmKorEdr3Z4xMiJ9HcqtAUNw7x8f4g6dVGoq7ZPiEUaL0HanU
eDH46qsrwN2NyYH22+y3QZlHlhaDzv9oHeZWn7QF2MhQkJEhm8slK0Nh+P9KhpbS
VbeTZ8FZrhycafLApIBGI6e/20JywLpxwlFvVWnbIpyj6sM6QJBEvB7Zh4GUJd9c
iSWyJ2JiAucTbU+O6hQokolwMW09iwzWd6LwvoLZcCjxtkFaFDGli2lS4FOm3h5f
84NjW0g9u6e8AcfU1MXfYLUuE9AxrssofBq8pdUZqDldLyKNDhipVufcLNYu1aSR
vZrdWT2xQX1CJw78Y3rvdXUPE8I1pmYceF0quw45Ifrq+5rQOoh1+Mda+BHqqh/9
ljWFeNzlVhFDD9U7/Zwtu/dWw2Kr32D8n9SKuncVzwXo/i3794RrGgYx5HIJzqcb
qfoxe2Y1d3KX4Otpcq7cmtWkKXp6Oqvfed+iBjFzlfRbMB+koGdu65wOrNdnI7EU
ENzN8g9JrcgdN9grwvYrp2TcGB5KRR5YIlJmGD9VpGWYboqc9/2Fzf6cVGZYXfqE
lA6xYOkNm16Gq1+Na2lmEh8Li3Bw3xtmnSLMZdtZ5m1pDz9GmVd1ns5vuJCbPYOY
9/oiB1L682fHkqHZU9T+juqWUfirHWlIwFL4zhUuzSNmP5tjYldYHMZ22SCfM0sL
NSBvn4yMaE7DDVtqFteDWpEZhNDBIEz8iyCnCETICIptNA7TwET0Yv7KWsiqCgWQ
RVQ+SZkoTet71T+3xwE4Xb+xEEa+oXriYUcGrhiy0miie9Yfjjk2kuunqAVk1qpg
ypP2r1c93vvGgTELgAberqBJS0415LsF8hrjptduwWIKFzxL5kJ4RCwpIeVnInJe
JpaWDxO5LK0x8F7TDVaFMKJnkvL4HRPUj0Ltb1EPiyC/oI10nTc7ukmAwJ7IbkMM
i5dVl+B5Mxb5ElhM2fVv4nX77ZqJFrtj2ujEELsy5kO/F7stJ/Src+iexzAAM4SR
YkxiQ1q/4VYjpuBjwoQcwB/FbPDIOW5HLMqG8YdQbvTeNMVdSRRLDsvdRtYfXTSA
WRI6VkRzdHdSOHm6OIY0FKYW4rnDlZFCZ8unlKCj50v7yYYzyjIvHgAYhvTmzS6K
sXmrHHMYoHbHux+VKhO8A7S+FWCDRP519MoG4dd1VBWnTFtjEdPT70jNBys6Mggw
QTXhCx/YWU0yGT/aiRF00aKTmgQFAlj36+W1u382Q6f1Gb9oE2MA1Pgwrmg4sJJQ
XMP/jTDh9dHteVvg7xdHIao6CCfCJredp/uqJ3XC29JA+U4deIS6AgOsAB3WeE2s
kQmIfdmcDntAbwJe4qnDi/22VYCNiUrbaee6CaeXJOZ2PAuTV5+2m7wfXnGZO+zc
Rs17att3KABT15fmuxE8V77U4AZ3Pfbar9RdrnV4gbY8T8UhwcF/RG34OxsZsMai
fvGY6jPYzlTW7bxJPvMELqtuygWbo0PTfC5bBLTSNnEbTfrhyHSN6P2SZTZ64YnV
TKWlvr9aiMNErcESPsRx57QU0cGrGFUuA+zCjY09ZkrH4qj07PQxeJErJVkpdMVT
u5Ukb5FOfSDYc/OxN2F2tQ3dq8z9PMtl0+4s7EO8hQRJMSuUhe6Ih1cXf8e8Md44
HpyGmCM1p4B8gDwhoSZIU31tYi4RnBtx6UPdixduX3inpHlVl9Udwx5ncua53JYN
qtehjC4EhASAxBwvI5V+X13PTqoMKXl3HeWOYxCVM36JHqDIH2iDATiM3b1JZhxV
AMiPftp1q0piIt2i0Mga4Rj51vMngkmppQNqutTa7Gy+50/wmKDk3Mbcu38FFhuQ
aY6I/AVjtqWi8MQLObq+C8ivWtGmMbJbMld19XCnXdu07o0SHeQRkwT1QgwdGr6+
0Fa5yGwYd2aF1qsYEwFoU2R71fPFIukfgiUTrv3JOCMQN098D/HHiLfpwW8d/JEi
0dVniPrsivM2hhD/ShVL7vDOYY3aBr+YkSoXbcXTJ56zjVFA3/nyvJJHnSNZJgJx
neyv6XLG9aZ0S7N6H94WQ9lbmOPqOBn0xwsESMjIqVnFzskLMLpPd/wUva/BJ1jn
sZZFYwUwX64uWctSQX5at0CKziNPFWiBTOm3DUiQWkpRwlA53+swsz2QCv2tGSNL
7eX4pZU5oZ+U6Qtqs1ymlKnGhbNwGp8glG64WRAefqGhbjRwhjmtHRP5xTMuMHNT
8YGXr+81u0jRE6IEsq+RyjnKx3hzCTQHiV9mGNnO6rnC5INUkZhG5p/gOAjkgMql
Msg3kS0aFW3+n+xaWExVlR9Rux9VBZixTWeMFL5GSzDysVn2aDmeyMEDFxSmi5ec
9YI8t6/87Joda5Rc47yK42e+IxFH169kKRq8zyjoniiY7S9nEzDvWdvcqfsRo2Ke
Ry9w6eoBHRJyrStBQUJ08LugTklFZVk1CvucaS1JV3CElMX1h8wCxTkqdcEHa1ab
mpy2KHk731gvokHhfa+UJWu3/yu2vkcJ+2GctMOpBSEw1ht9qy1s5j+5QMMBOKdE
1UuLZP6K1Bm6FpVcGrW+IQWKZkp+2A2BYTcv1AZwiElN/FUMQYtsfj25j13d3BDC
yzf4fEb2SjiZq4loyfxfdqBlEkommNWMHWmjAM2WzDHwUmb2vvNLCvXeISdLF/tv
UhNiKDaLgYHuqEo5h1TcVql9vSl4lzrpP0H3n1pDZCowes5CXjLJZbNCK6ggqOan
/zuCSLQJShrbuPe+EWetX0Xec4k32J+oVdwo1GB6lnMibrtjNVe5Jpzyw2MxYtKs
JCuqcFL3Wbfle3ZswidCtHNwCJATykJtjO340NUXSMoOrIo432oXMHtEObEp70ls
kPBdQoxRq4szBr9aV4FRFSQaSHNxGY+u2ioeREYPKSmQbEWtnEcUJxF2RV4sQ/GP
sFjy9XQ1NHlxiHFnM7WH/PAMW+0/JeXykscvc3i96lUI3jwutg1NbZi38JQdKwp/
GXelvmPcw8r6WTNwClHkG5gwRT/Pkk4rjzn+cWB1IvLdYzTvrj59kMuL5IHEiaUY
z9F83WyA7JpF2IbYvy1i9Mu7HTRNYTnMwNcfJNywaZ7qFUOY08/qloHP47Z5h6fl
tUEEIyOGdgJQkrsekIkFAzCzfUicv9nHA5MSQlk16apZFnfxP+eH5gQRpgUcEFoS
KHoGow1ee5rBhN/mGmdedwp+Tivt+t9Xcfa4+Aye/qzo2gafY1wLYWaWhDjzbvCX
MejIE4N8FHBILZrKSQhfvq7Ey/yT25guGEZ4e4uiQLEfWg5EPIB1ygRYJNCg+pu1
GE9NJcW5cQKDQ68fu1T2hi7GZSu6vqNE2uEyZOQ3ZU9lppQCbzASt/LMsz7aH9h1
TMwdNHslsxiFY1v9wl+u6TR3idii39UK34X8wqoRGp6LfZaFSnIluVzCIfqIAE4H
ZnygQzkrztiGP/U9bG/hWwBEX+D6Q5HDqcjxtL5hAHuVtHIwWfrp7OaByo6gKCoS
hU7r5/3WsLE+5DkOjUugBWDGtj/rHoIExJjRsn5trBZTRr7RwSNWhICEsPd1nU3/
cMOLAov7v/BM5xFsQRJMUD1lwvdSAcBpyyLLFD/3U1pjC08IeGbvOOBgksJajZXP
l/yCSjVwtETizCktR/NL/z0rYV8DFd74ZK7LaGGI3Tz50A5kd3iCEh1nmbMbnZmf
izSvk9wlaZX5ZVhphKDJkzrL3kIhfA4aOrAoJ/TjlRugBM5F6/q0pkt8VDsiGb5C
+rXO9zI2rkSFqbBg5xug32ploH7XQGdm3P6GQK1my0VH/xzHBD5RzLpEHOOweuNw
6BJdJZ+1DXXwLF+M5Pu0S9XbBZud+d5D+fqSrV740RFNnbLoft/7n2nBBzUCsYsW
WYvabSp3md/rdERugVhC3i/1sM/w9H6Qhn1QL0oKReY/0PAQytuBWhX6NZcabR9M
mzPT7MpCpQTVwdGWCMuOt0NnxclhBWoCkHRSaNjpymYEMkxeXKe0YhdC4S+nwuYs
Zb5TNzy0dhpdEgvogiXflsT0MdMNavvtjx7uuv6nqz4noIaPvWrh5gAo2JawhZ0L
7lkJl2tvXpS2mMgb2OHuNwNsomOuZErb9bs2W4/ooRrrHuPTvG98GkqehpzYYZSF
1EvVXiBBi8+/FWdDDtzdzJ+wO6nQCVyjWagF5hJT/xgjI2+LOgrYegZXCM3MLvDv
P7pn3emOCpL5HfzcrYlYcEH+p+0/oKA8XMQxWWdFzSmlrPAm8wU8HaHFTp39WsDj
hmthj23QTynmlGHNgzj9Bo8UMXD/i4df1KvN5qb3PSL7J32j+dC9Te/kPeB5sZuD
Hk/dWY01zMfygyuayse+dwQM2rSvRCyuNyJivpgByM56fjExaLrL+js0XSa9hnGt
ciNTBnubAfJfuk5jLoMgFGmJRuYQeL3EMz1mri3LvjrMR8sQyKdf6PjhVoYZdaXr
VW6B8j5gOd0LB7f+aE/uPE8/eIwjsZLV4NTRs57gQa/nWv2QaOqsIvVRdMEGacaL
Xmbha5p5lUYvolWjd2ljO5+a7ApcCitYX/3I05B/b0RKMg5WUSjAzd9HVn1R4ZK1
kp2j25Zo+hqSDMUeinnbUYw9gh5mhlvA1xk09pCpamnL/auWnTxy2o+wsGt4xulj
B7E5tWlSjylOwLJ8v1rKhjQAGNWX3JEULvihFZDa15HD/Sgjjwtj7i0qZUhCFBe1
Tybvwv+0PYvL+Z53VR6lx/sOBvRRvFGhiM8DGBZ2d0zAm6YU932k5dHTbyk1/b67
ObE1tOxLQm0cYO0cw98p097NFZFUUmhuCgsBQAKgFnNXyKKwWSqCCaoNjlgQ3I2T
24kJuLSg8Ahn24ghl+WNce7AfK8pdRGrTSlo5Te30lk+GcSYTAxTKZceUVqSzXcd
Aq5UL8aAprh57FsuujoKx7X0GK7CfoXP04T9j98+N5bMqdvAVym6XLONPnHorDek
ZCpEgsIkFLn9L9DyG69wl0xp40VBB8jPTdWl1SKmWHBbwoxoTdfOmQap8jVJfVNM
caMLv0wij/NNXzOigr0J9Jkazynq/JlhIQzaF99yAU7mjroCsvQd/8OB/1CYtKLn
82IZ1cgDOHp2YOBLeXp2SvkzZYFe/91hnAKbCAeSerP9ETPZPbg3YW78+LFu27pX
9icilKBjvkrUi8HVd3hfs0vrRWMJdx4VZ4Mq9Q1fzHr/qSqNDvN49b3ih6AEbjRO
ycfYEVJwxX72WahYZvO1kqO0f4JLX3JqzfbpZ28z70FmwSsNmDULKhRhzAfd515g
TDzbsMBZFhVh9/8zwPSSwCvBSC4FfHfpTBCplswhl40ubEKeRZ9O3zpkwhksX5Qx
xxQk+4WxygoIjouGJrn0CD8g88AAVKlvYbDW50mr2iTuiNjg6O4OHPj/aZ6CFHmJ
ShhOavRfWpI1YrsQBPPiHydaLxmVd6c9O0tM1ng02STm9e6V9nhc8P6gWaPmqH4Q
H4RfUel1pmd+CgzzpxjJW7o5dvN6mVKSgq9Lc/mbSiqYCuNmHKhQNO9YDUj4zPyd
JfpoZqoyCNGF2vcSy/xZfIREPPD3QBLFRq1lLtBP8OHwqXXyDEEtcEmm7R7WxEcq
zwJ2lRR1PZlbbtkeUAh0s+GomKHRXiIWNk1C+s2jb2onjJfPNNgVxlUO7SjUwXh/
iEx0jQsbVhl0t01R95DfF0iH6G/Xiju3JxYLK/S7baD0/cl8Qiscpnk/sIRSGdac
vY+zW5edlzKCnbkxk64WqNlfUfmapYvPkSNYYKcj5qAyfLV9BEWrg8hl0l/4Pt0O
22MJzHO9SJ+/Xu0xoykCZIC7MsIviJ3waAeIZoqwq+wb1cU11bsOsmkXEamcLFxR
+3kAgNQZw3L73LNAiHCTjIZrmC5THgh+fV0KBGFGE0CqP2R6EdbK2XtgoVho06Vb
F4r7uzqO46kr19mEX9DKTsLch00dXZzR2fLTuMUm8T1QG4dHusVt/0dyGqpc0yHp
X/KTUpZCQBgNqQJdlmwLSsF3LdxaOprUhegAGAl0gLEYBS/AJu4M/KKveJqFuXST
KqLQGhthLuhEYFzki6PIWFBTMvKDnrhHaI/7EE/SOGRhebAJss56nCeF3tYCsJ7Y
0a98kqmBUEOkzKeo+WmdlwRr4hTy+Ohn1g5sHmo4/6l2Ek6DOw7pgGk0MaedDh7q
TYnEbyRr3YIACzXKBR5Z+OsCkMb0ZgI60cVXAojrn5081Huud6NnyNe0YwuRjp4i
K0MB00rQErqCGDu1mjaeASM4Ll3RErK0GA2Zum7E6GtAchrgoBLeeV/jLcB1MoHs
cBz7xPE5xp9l+WxTFuXsLDDp0sTtemqv0cflrceZQzn8g5Vvu/c9WN9Lli3DDNCr
UEuZ1DCbsytIrns6Ft+TITuQjJsEpwmjr11meuDlaQ4gzuEULzRHQMbtzYmRnYhi
KPEDMt7LBe/yW6geqBMvxRkfrf1MnECsn9MovIKn9HvPf9/kRsnRtBtkKQ773E7F
3MEHMVQLaspM/TPoAKBSQdncZcfFtd1SywlCOYcxTOZHY7PfiquqYXciG8jyEvtO
zVZ6Kn9mk7vDSYqqW1eFzGzjCXVuekSyF7NctcUANJn2uNToiTOzSREdAU8WGmav
TjwdFzw7s7TtMi0Of6MeRLsocEQsB+hOoqmOo1ojiycEZORoUHt6MQaNeiItpSmh
5dQF0GIEb/JUvxvBIOdm+MyconfZQDYkYvRBWVT4HF3Qg1Ibk/FMx6zYWHyrbBG/
QKWkFbJmpCRtc5kMIzPEt/LC2NGBYOLPHuJcHLHJuYSfgqbuDtOkjaN7ENkN+LJT
SSKC/I6jXR0DI+X6O0yBY1AMtyMW3owDgpIWHYO8sgJCP2VpTA6M0FfBYWQNgZXW
YuQllk7OhE8D0Ldua27+D1RZTtTMbt4v8Y2NDjOujVKuDcSizeJbSEsesUB4Og+n
s9vDk3VGK8sG3xsLheTzqzOmhxyytgWryFH+xnT46XXfGN8HPg33oZk43l5YWo5v
NnUz1nS7e8pmC2ldpYxL+EBzTvAnwsuEuEIVi0II85HanfY27C4rOWYTaRoAq+Rk
wFlxdXBwFcOsH2gOfCwPGzd+8gHUIjtRtvJdnMUgHTvC6iU/QaeMjCWZm9BkmVm0
T6YV9Wr4a2JAyTwtKsowC80bGkhAvED92Yi8QghFn5nfLelxHKI1WYb0vHvfFG/l
myWahM0GBFmQlntoID9+VYJAs0FGwF8dcBsStZLFmJb69U4Ju04hpd3+3fCiL1bU
YwVDnIzTxzWET7uhsDKx3fOLAyfRqTJ/FcsR+hTnurcojOawEMS6o08XPXsuRc8w
1xn4x6J67lAQAibTqC1sTm3tYx8A1fHKkSAAMUBV2aOPh4b8XG/JkPnKFDbDNdlu
kxW3nViPf+ZKxkvTBG7Sr3raSI6BA8syFvBV3kIvfbVsmZwHJ1QqQQxy9J0780EL
rztRYsl1MOFqiOapRMV2BYAv2gVbXAP37wpMp/wYA+6aHO0CZHilfXyJf53c/Rbc
PdT2gmYshNA5+ae+ZIEJAASxwARZmX2umnsEm2JLatCqKLFF8YTZOpcaqxp7q7f7
j3KJm/SMdoO9UhaCUHT11mkZxMJ2OXk6J1unzQl8nlege1+61Ww7vFWMRDgdui0G
ZkAjUOLmG/OYFyOMB+hrcaqExxUbHc3Pk800tnP+9Y1PX0hEctMjptqLHVm/RIE8
qLQhnkiwqUOfTLb713Vr3Jf7+azoePmetYwmDSg19GZ2a8iRXE0ryHGPqCzC3rEE
j7wNoGJ7dJF/eAbzier+p+P1M9dH0gJKtg8CzMDaR8aayHg01OX3lLN0+LsnikhT
owqPWhQqHK4j3Et8Gz+nohSQzpPcPyIRIeeqDlImNOCiVSJXl8m9882oYBkYjiC/
bc3AWyNxzoiWQYmClU+VoPK2HsM9j+6keF22m7LFntjk5UZkrJtyQwZrjTjwqe0X
uWVOTitNIvjyaSacp2YJ5F+8IqCSZ0TXB9q8UuQz4iw41wxjDhtbFnJbUsasGdPN
OQ3RwtQKKJs2X/XBF2kz7yX22PisOnrGbkE2KP910bNvMwXMevditWI2nvKCZmrX
EWCrU91m+pZlOo3E8wwwHj6X98LXD0GKpagqWc0YMN26APr55NiirDaLJg2m2/P7
XBcgg5gJkBGcmh3qpa6ZMtNTWO52ToxDl+fGXF4cuQqA72yVdGWy2QcprSalmYef
g8PyNZ/9vXokOTjCGruiWGuuyPwvP2MTITrGFmotnQolr5T0BxP5M8JdaJbaHLvN
uOYtTL0Bvws6uEO9nuOFaRDpjX3v74K8DnfeRz3u81lrpkcD702KxFS4CaDVKXlI
9cfG3W1XHoL/rdDQ/Pof4E6VJGWY2NoEYKyODJT4wE+xb1/XOn8dusD4tQyDk01m
7JkGRO9i1YfQoIzenOtVkcs7oesJjv2r1sfKQyzxogSOQcdl3TOZRfO8sCD/By3b
TiJnQ6ky14z9vmznP2tGDFvrk+20nZVu7YN8rwEOYZAUbg1j2LdBYNkGFkEOC3x/
loSkaAKh8XYqrUF26WklV+SvsW/tbgULaJYjA08stuQOKb0X+f0OB0RYQOQN+lhF
saxpD4PNEzBrD2IhJf22h8RnjKHue9oXMpjXbMoEdJ0ifcp+a8kUXLsOnXhYCcr4
uWC43zZnfM5izSJv4xFpp7ezyDqV5RqeHAAiwvVTra6ovZBj6itzAO10m17LWA4b
x0aibzNG1sJ0MYydzfSipxMDnCp8cCZ8DxzdYtU+EnjudnrN6HveVUqAS+gEjjkr
0UWXMqf+T1YyVZqY9ILNY3DmYWbnY4plqqx8nDirr/rf0fbD0+Kui48N/GUNtQXV
nhTNrTAE4UT7KZxiRwPZVxZtdaSP/rw7/PH3zUnktbQ4qGVWZI7NrJbJjYsyLf85
VNLyLVVQDWOy/IGJiR14iqpMSwVgQdOe8Em09PE0050O3AQACEA7E/MxSxjGmsv3
TkRpsOjysAHk0CMa4tMPbVRHdGOSBzGM/70jdwQ977+XONtlUv3ZvLc8PwRIQAIk
wUJeOKfgMt+4ZFuAb3xIbOqxWph0TlkyvOBmz4f7Y/h6u8wXUqBzx3oTYpoOzD4S
g22PMIHmuK2RK5KYAE7M48EhyrQWWbLM7U6u5jj6wjL4S7s4eDugpRQp7TvXgotA
YOrc9kDfGM+ie7e+wqn41/wUg523YJ4WmjWPAab/D1Tp5fXaSdLzsVgAAeqgbHrL
0Wo2rYNO6vSsYNWr4QDJ+INJCCgApddXoLDbTV1Otm1Dexm38V2Vw/VK9jgC6nYV
JmB8dhua0EVpgnC+QdKJuogm6PAU6gYA5LUOtC/YGP9t5J/sRk4qE7pNGowpaWrz
ApPfPCsNpwsRxRQUzMRCIArZ/G+MWdSEafeKrLvijC1fkmw6R1mKD7pJlBOMUUWu
nWVBjAeqQih8L9SPV5GxwcfEmNyDpq/XL55XIkz1sHfM3W7ikE4y3EgQHAWkt0T3
1Na86PIj1PexzEIfZ5NqTSxR8rOzG7MxnCrbH0mdkOJdWwrbKSnaBacj/+2xwRjF
HA17r2UP2MC780HXGVJ6XT6RiVRyl91EVYTCI7J6ftJh0axnEBd+M49cO7S2g6ir
AMtD6fdMgqIkB7d0G3xK5TA/q/J/qao3nxWe6SUZnCQeyuiN+vppXm3NneV5VIE6
WRIItkcFQ4ChwkCN0EZVkKUW4RtJjWK49lKfeR82gaMzB6KJnh08YTeQ+IrJwWtw
SvWWiJIRyPHFjCifRYzhVBqnuEtIbVAenWte0/3+HVVb+aWtnwVicJKEsZtjH2EC
W4MU9rDN0U4agGwti0uviUCvWFG1UyEyr8AYMlg0JzYEg7ro/lcNbWNEokbUdz1m
fyJcppWaOeXBbpV/rhGj6fygE2iskwX9voEh27xHNV70Qywe1osKaaSqPqKi4uZ9
SEsA89Amlw6ElSyh0W88EtbYhP/6Cbj3fu2x0irBtwGZwL/oLmi8nS0WWrtMuell
B7rJeVRmRgLbOSqw0olADNKW908L5DzesUhPWTs2HMh5SaHpbDTJdozLSPg5WnPJ
66DcsV9T/sDB2X59PF+Na5cfIHAgcaDkkiVDUmCNpBsZT5usT0ACXV3RVnCpIk32
UtnyAmtzPVXvNN8Z/L0NhzVSsV8rj5uiK810376WzAWxgACT90seT8TU9dVZomLC
dX+MxLqJYGQM3ng7W5t5J7O6yLHb4PX/9Ww6qL+EsAJVXRI8ZHWN1Ci6sIYygZZB
TLRCshqGjlolQa46ypi0ir6s6XAljzattX1SDPOGkCzcHXEC7bwgR74r05ByH4ym
LuIPk/tMg/FvGH492H+NTMqcCsFNe3U23IeekCFclJpn8ZpJXp/bJQtdRLvE9kYS
iinp9o6p0hCNuMtDzl3s8XrX8m/nlS71SKe/fgfxqqmKcFAT4U00/E7lB3uYrfmA
x/dBZVSPqxcaHAOtTNUNX4NjG//VsQCAj5LcTTmrdFlBqR8VxwTcZd4IeZx8phIX
WZCXQ1DRiEwLJEpaHKjmQRZralxwra61Lj8lHtxdNAV56P9uUJGJiy7yJPLdNlBQ
4XwnmQv641TBheQmxU1KuIknYmHMFVTksvPrM8KUfwqjQekV8DEN3F0+oHknnM9s
PMQmG/+BMWzUqj/l8Gwtomqu1be9c1Rtss4IvLsVaQ4OapGugrPg3vBQuxe0/Ifj
fMb4SYbyIVvkrFARmMwn2/XHBH7HYDPFVmTJr/Q7mpH7m/4hyBtVKFA5lw9quuhV
6DJT3M+s1Sum0PlE9AGwQw2kNLuP6nsHETOIY9AF//t5eUcfhsi1i9ynEKExgpVp
eQwfngYz1uJaOeSASP7RcPnWJpWVa49TtAGUjKwqjlwpGuf1+Hcadf2rOppt+vK8
6t5GfJVIgAZf7K1Z6gqJPfgxCloOSbS+8M4asTWIlCyuPZD3YnZOMOeMMkWrMgv8
foGujHBzE6qB4WMxr7qjt3AQwoTHTv6WpFcBaeVCKEk20LmrXd/UlEqGzE4a1nmd
8YTqlHVBh/6qEolwpKRBKT0m5Ybx8UcoswDkLqeG6WmLrAYdDTMBd7RxeiXZazt/
g899fhU1mUKcDn4A41YQFr5g/4yE73WlWv3QeyOtZ6wjqZfPUbReW27alCjwW9oJ
/raipQ2EL0MKG0Pprm1RiUvdEalVM13GEcx53RZ9w2qk9weOckK5QDpcYeCNjy4V
YZB5puJGgRME/wbUPQyulAGIvgF7Wv00kBGBzOZXwHsCF3rrjhzfF23lr4uiauKq
GvD05s3IGkDSXxBiu7LZe2e53w3OROO91hv23r67SY87wj4AOewDya5P/Obmznw6
a8NICegEsIOVfHi4lzeFn6jVBfLoFukViAEzDPl/ak/SEQisf7KF3ym+4EtJDTZ6
lsl3W1mATa8jNNmpN280Yboh0QVZ4cHjTeA9d1NmPxLEYlJBWXVSefwPLEzVwzoe
UVJrMGssRyFNlEK36cKS+qd8I3a7Mk91P3XNQzHCf99vpokhi37smoIiGtDgOco1
U9NxXQa8t8Hk/ktjH9niBrHr3s8t/iOE8MlJMnIF5DlF6dJQ+02fmTP1SGCWdCiF
y2c7S+B/u/WGeCGgxKSy/D2+5P/ku5wUuilQhZSp7QFKCsy2nVN3UHmPftCY8SR7
yRcoQeNCppfYoehHf+4NyEVCyoD41Ta2fdO8hhJULvECykaexGaJAD5cAb2E6Q5W
xF8A4D7Plig06tB+HABClaDSg2XL2bhPRa38nIRopa3XC/vljuEvcWe+oG/ask8a
nbmJ37nsy/t7xKlfApGOSM6nFrAbgM/uc7eSqxkimpr0V2+lxQdkNb0O5ZWA4UlU
bJMPDnDPg484kx2G7dwUXONJaV1j4xmvq727cP0l8Ea9tWNPZvt50WEUpaxW2PNj
44lqNGm02KI09V8sNpuPp/R7ZI7zIqf+KiuRQPtNe0+ntx4LjUyveXFSYVSwcl77
pKX+eKlEZ8TAnVeXb9uoCWVpT/7n7bQdsj6spkS1Bq8QyJRUWZCFGULb3SwsqucS
j0JMSyJkNPxNJl+hPoKAAI/L2nyjCFn5L3sIUyiFBnn2C32P9Dug577mJ4YXv40G
haxyznXXvzMBaLiUNI8LU8CWTFxUpTTmdUN9ZOiv429htogLAemrM4kAqOT/qgzk
t+Fzb26BxNv82GH1krtNmQqoHi/ygFLdndY2dfzOWmWKmNJVI6oz0aIwNCaBSUuf
TUrUz9/Hj+n1ALkwHzr1qyMech6Sqo0t5exl2v2cNtW+mvjVqc/I2AyM9LefsWFf
AgvaTB/t43kEtlw3d7jNFGboAK7cLaIQnE/T2nmQE1BBh2T5VPAs4a0/HGOBQXpP
jONjGbYGHjwsRl9j+uFX3kMZhQX4JhOqwFTH4oQp7XIvG7VTINsV6GZP8Gz6vGdv
NqXbZ+38gUkV3el9HNjiPCvC3BShzd5u6B/p/smxuJdgytfS6sNPEOPlupwHnGMY
iwueZc8xft0kgke+To2MHUD4jpS6Ltj311iMLEXJR/mCee7GTJaq/slPXxcoS/MM
4o1OI3nqkgEJntTS8cHR230ajCiFwcKQ2k14ut9z9+0cR7ACxXn4v0HXRKqf0r8j
IwST+sES/mRcwnkSpfoBdX7YUna8ja3wFttzZkag7IHy0oZBkVXclCEL52MG/0Sg
8Nfvg9/56DczudiCSbzK/7TKXxdLVucEP7eyUYbhswhlCDyhR4uZRLgFkzl0BOzV
sHCRTXCrpp/4EezhOmjw91tp5XaqUzINB1SPmVL5ZXaqDIFvn5mEM6yy4sIXXDZV
FGNLe67tBOhZd4EJwm8ZdZPRORcOyDGhVuCKSCovhogG8+4C/wCsw5yKcJLXZElQ
ezJ4k6d20uDL607w0Rd4YlxsAM+FMKzBHN5FIp5fgOatvbVzlpy8JiVLuYO9tdkM
bgB0X9CfnOr66pb3xwMDeAr6Y6ILk4/9smNlr61iZZyyYCBLr8mhLVEWFj17CgA0
7OHLcoi71FoGn+0cJ34jPma0ET9ukbu1p6Yaa99eNIl5av83bLI7NPAcvbdZ+C5K
te7ZnZbt0e5lLjTNN/GCq2a2WwZWuapCDqO1MEygTC6JN99mIvGUe0khPyBMUfSW
aIxIINKCTmHpgex2roWnnY3rtkpmjd/yAuZe6Qm7WjwtxiCUz37LRLqHr4GLXG0T
259+51/F1R5k2mPtgP59QI7cGAT/5Y9oo49dMr4T3gQVclKboLFwNUiMhAaRuQUZ
k8NDXKu5dJY8I/KopaRx8KlTefuy+G7MVlzgwJrsv5Vv0GgEezYBWcA0ET/3PL3R
E9sSXxQoZ1RI5UYzNq4qIvvlINc9DSbMhr++j983zt3GL84iWvKjNBTA8isljj+I
kakTGVlNcBCpMhXcygoHr6qjLHoOwVEtuNw0ZJnO9FgnSTuolAFEzoZdMOryoVnT
iZPcek1/a7jcDqpF0nyBjfOcFVp7xX6h3ySj9YQxyvB3EYDfr3iAWOON/um/BBxl
YWcrF/JGtXUP6lhO3m+vl7Ji7eZctsBSyGyb9Gti6/I5gvUgemTHAuXLBeijH25z
55S35L2QZ3pw7tvOKl8Pn4hdLCO+davQIj+5IZqxmhDwN87K7zQDKeO6uX5Dys5J
bSbepnQIxyGjW2Yuzohixmn5rs90Fen9Vz2fPp7L8rqWnHtecx/zdRoBjgcAbMDy
VzeSLQCaSw446orUfYTdHh8+8AJu2QwNVJJloTjvkc9GyAsAKAdlrUHQ5pbRDD9f
dwb/FgDiJh7PhM1r4sC/XRq5KKqbw17ccKpihWPxyFKy7Vs1XJce5rj8HHl6VbEU
19pGekuTlxc+TSBqNJ+MYK52VJ+NqphSH/uIgfqu58ngSC50qd1tAlgtMdjbzv9Z
B0gvhVazPkdFYAO4ipe7dT1+hC1M062tJfhkkqnZCypuuKyaYaIk3DtYP4agvUMg
JhMYhx7JgLNwLdoK8vDKo7QN4sx/Bm1z3OTOZxWlIcfjJ5mZwy7PQvMDAS6Xz/gR
AeRFRBXsgeD9TwrCm+jNRcNsdPdLngDD/Ev+NAgPjDNh/UYtbee6EmWTET9Aro9e
5GWX/XJ2NwtbL3xnwBLeiiLfOOubzOmyrXDkWgQaS/El8q89ucrGTGNwa+B8gUVg
PUPyt+vEr3014MjsRP+xDcEhTCzDv6y+TPC1hWa+kkYnPhmCDo2MLZliG0iqHyNu
U3K0egAgjp8VMjGQmvFMv8fpQpT3BUhVv6y4PUmBLyAO9dWRj1hQJvDyZIyBlWJq
svGS2EOYtke37GqVeI8wzWgu103H1n3w5NzLq2yxgAF47pg2LJu0ZgoZ1ZHtoM3G
Ak+A/i70qo/dSOjzHzV5QQ6cf376lFsZ3JEIXQ7cWjYUHA5s2qXczRmcBlkPNToR
zkzWWn+6E7MZ/qsuys1vZB94nCK5n6K89PAKybBRWN6KHhN6VLl0Itab4od1OcYH
AF7k+Gdh+4cq5EoafwwkI5ZHBznS6MkznZ8kAWsDE+dvJCn+JZADjPxctrNtE9t7
fVlijsLxmGEae+j+Ks5rjkAoslPRbnvIa7hYw8sKztB/YPEtGmZDOYsypoKzIrim
2Ev7bTEDf8laCC6QpmV8Bz+tziMFxW24TlsifFjMRxAQmAKdj7BII6nSF60lwIDU
lvdl19sOnp96YfGm4M4vO8h8mfkGUhPxej8+LsNEBjiQzDJnTtYntdWNuz7p9Ah+
+uNZ3AfBICNEuyRd06O0nBDnyWDeSsoIF4y2HGOhkDaMCEIKjmDmsEUWytFVoYjn
f5IyieLu0P9cKHUkwav+mlxPGDEichyudkB5wBLyGQqSTjhi6uQKhe/8Ou3AaWsa
zjiCrkqbRghA3uA2ZkrAtZz1HQ9RK+oBZn4ChlPHUem4PZD1N1RonRbmh5c7M1HG
YYyB8Q3DYeJnnJqVnRqBYpYlxr2S12kox48eDbl20MZHrf7wNxhOmcnh5vhSzzbf
XnEhfP0sOYTlIxwgq5WZydpkbHCTvcKImZiAzD/6DWsmcF+dnzY50CgosEMbzsB5
/C4Eyi93NEBhcUMliQVAVPWOwMSOGi5iZxMANultlmHrNySb2ND75ewBqtrtaEGn
bbWCUM2jmYHyFXUM8wuUVi2KFnRrQer/kpf+DRSmvlNrxjc1uC6Hlr3pQJ1KEg5A
J2aG7yE0yvIB0AC2yHLvIMsZwKRp1Ev8sBeeTE6/nRlpcyMgPTLyaJajFVfhxPA+
0VINGcEJZcGwq8P+MXENoNjww2btqpyiDgDsPaRM0SQiNx7eEDera1KbBH9ZcDa9
F2MQSyrlL+XZO+qfFWmJLQWjD7zbnwk6AbRYLQ9pZzL+KOpoTExhIYDCtibc+GbR
iZSvuVacRe/B0C4DkbKEXYkTBq971+ZAG4Y5QmiLu82cUuT6/LUdiPmGszNiKU+/
CR8+8+28/ugbFGo5VMBIGWxrvGHdptmMez8U54IC1idD6SiKDc0L8n7dIR1xbIH+
RRXUEMV0eFBOUoFy1ccQtY6Tjfou9/JWSkT9GJjevcsTnu3bpC1IuYthi2SJtdUQ
bQJxyr0AMkrnC46gcNbEGxm+oqOhr4hZqqYywNpqpEGyLUuSQYV51ZETvwEAHAd4
Y9oUmSde1JNABMvFF1B1nf3f9S0JA8VLrK39zTGd+TBE36pNCO3vwSigHAY7Z40Z
oyDNXDqF4CbRcn9cob+dnLahp3f33FWf3/xUPR1OrcJczFXwkDljHESEiYnxN3wy
A/BD/Gg9Mb1FmqvrJVY/a0QJTDF378OVd0WWQRD3Hfbl5i3wKM52jU+fTnRMsiVY
3+cysEuf4ymgRl/MT1ibL4zyii6wKFfYWdQyD7ZViGlLWrV60mEmMLsGrsklhL2S
Y3tjh8be9GPNSaxrkQmMEzw4OLMji64DSEzYt76lcvKZjZ8EXAVescCIFMPIMkf/
XKuo9lsZsoePEmvksuytfC03dFmSptddwxiwyyaCfCKiUF80G1DnWrRNwGYi9p+b
drSxQjyWXZ3JgjrX697whj/LVSwduzzT23rrYn17H2pp9zbWmsJt6q+sC82W3Mlu
iT7rgB0h+Hpwj3oLXNVH1A==
`pragma protect end_protected
