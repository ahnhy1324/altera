// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
n6yUe0JorGRUO761N7qYRkCg+CisQo//MC7aXzU83CXkoW/uNaYPpWE57XsubFXS
oHkt4t2rQa97w1OXxD3nlFTQNdzBxHftWZikvSe8MEb232X8jvBrbpNHu8Vk+exY
ODpK+HnpNy/QYX1quCSw7GTGzh/Qqvp02/x39YfLE3g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 38656)
qR379lqAS+omDqGWr5q7cPKjWtWf/otKR/OmfF2Gj/HFHi4dSp4KTEAHep2ZvGAF
KW+kTjLY5Cg2A9aOZNHi/fGQRjj70PgdIzReVuDzUAQFC4THxiMnf2gXVanOAJDG
GavU7aOyxJxf/fdnls2lSP15Co3AQi3BvWPqVpqhBweMnFh9/tz4823wAv5t9+EC
wEaALHn9JENz2CbFAeHEVWQb/W+zBs0vWocjzafbcOylAI12MFa/5Qc/gzR3qJYy
99HgTK3voiENLcsPKPN8lK6UsoYPj0WweOQfwwxeziJuuoNx44Qw/USXiluTdWCI
kMN1JsjWeaI32MCpxxdqvNkyECN9TyJGBI5J6jKCbB6NCMzsVOXWf8xfdWU8PAmC
zCQoBJdgShrQoooQOX0tVem7lX9mq+MKlAYkLfcVKcQNcagkhJ7+zNRm3COJyMWD
D9NzlREGnT4Y7IIIjjC/SSssDl6moIGruQD7IKPGf6HdmFoFeRy9mIh+RL5l3QNW
TXpTNpavE2svJUIzZGZhmcmUKqAO1KMjXXM0Kxg0kgl963uTS8MK+8yKoNjJOvRp
HI2Ugf9ynUA5FghJHAsYPzp9N/L4GNUdK46g2UXj6reuTJa+lFo+llUr6ZpvS9AI
EYuswYvSdrF9DzdZaNtKjfPkm++YHVlc7N7ruZXrYIjUAv8mVhRrpoFlL3HRfDN6
wKzJhIcVplIn8hIZFZ/qcEfrqLo8grmmHlr8XlpGAyyhm9ueYbO71fJg1vS5NVk3
GqHXDlVnB/cBRCHTsFzFIx9/ad881mOirDQPmmHwS6n1YvkDoCQptz0r1r/Ls8i7
eHuwHYtmrT2MM9rMf1Wxoguq6MMt4slxH+fvDushE9LmxT6OWEVjosQ9ZU8Hto4Q
PSmyRzQQdK08QlS5Gc+IugURkNnlIXlCa76b9w6an2ZpBRTcH1W5v2iPdJG+WCwI
7x+yjdWe9bIYveU4b0SFhJ3p57MLLFl6hvb9m6uk1ELo/gib1jE7VcgN2k+3VL4h
D2UD1U/YvWgOXJCGwmViKsrowGQryW1dQ+DZyxkSru5SEglLAcQzBX05yMCtNdNh
14cuZ6yNfgYSPkvcvFbP8G3o0XFLIjZu5gTFgRC3oHx3XGhf7uC8TxgPkAE28KSE
VvPYsLcaorNWCZcxGUfmUPZhcGgIz/dO6nBjAavhxbrhaAGMKDar5/ldfLOoeU70
v5xQ5ViUgcnRCmhQLEbfxkuzYIUxp94fMuyhYxnKWHH7Mt0qsC7MhFuhxQXv9oJx
3CpfYMsnrSujkxW1om4qyh2d5WuD0yJJYK9P5JB4b3PAq42G6vNWsP1guLUqDRGG
ygBM3yKFsDB95lYL+ZYxBCs1AFyfZSEUmmwgw/sL9lqrE7fvjXEvOtWXW1xoINNw
nYstNt67eQIsZM0hWJ4cXnyhLbPHPoUTvE/Zm+IJj70/rEH4k1xysUqPsNDBmVYC
ZbLYI87AP2tHuVq5OuaVtH0HXFuBrZgHrLoGewX7ufACRR5C+Op0m4aP5HG3hou9
3Qnx7TayoVspeJuUxqjjtS/Sqd51PZ8E7caWEy4e6ct8F95dwaK78A/DXrMfXO3d
cUvCu9QuYnLMi+gFG6KxP+M5pSlpeCD18Uh6H41aOEG6JQLeAUvMUm6APN81aAgl
UuDdlLaeRwLOjSmlapasbWRLhhz/yQ2F4T0ljkSn8ob6Hlb2EBT5EvTvJcvaKGKN
bFtUVXmXUDaIi9H9YNHksRuAmcSe3JhE6aCW9GJvZ/Ec40Zq9IOQQAfu6z56uSIC
XNqNQNhiZ9He8Bs77MjifBxraMH+6VADi8n514BmxwiNXL1koFQGc+gK5GoEaDfC
RjE9erCTovLXMD7jzxEOj+WBjN8gZl4m5qz1udNSlDi1tFFSdLLYbMaVfYXZOxHo
O+h4pka1nPmY17q3TDqOvcvBmvdFkkewxWiHtfd+ntJLaP80xE9jqFHtHNkY3JXN
0Qunt7lbEiqzmg78znM9Z8Bd70X9ft2LlnlXPQEmv4hW0ofkhN3fDeOAbfgK/ahF
T2XJenWW3yCONHq0Gmt6UgBzB9lBjewrTkdSB09r7dfv65ScCuEq6TzGNHvsjOFv
TkjBQbipnoXh/lsEWskesHkDyuGDiSFr/UnF8+Swtvq5aaHb2A4bOj7rCe2ysC4E
wQ2/9GnnFgV2b6+3C1Czk8kG7nsWMh2xgIoQAwESH1DpYEZmZLKz1wIB/sVJQot2
3W8zFfYjUkYGdm2reY1aO1RjwzWb85S1G9ajaYDfBi2IM3hKoz166X3T6kgzPON0
pQ0hGGHZK/wGbA+cLpU712G4kIwpfOq5StHScsdRlIyG7nFkHYElJobJLWo00IWK
jwT5QldSufvxW1KlpAyF4Nt+dT1Xql9t9yCqtg8fMfisIUQMsv3i123mpiaG6k1W
Kb0vpitxLh1WdK45WuGqVJEqb+tph1g9Bw229EOwM+AaIB0cCtZakm+kw0sWIEap
Vmwbo8NKEUtBiRNdNxr9AMpVe0f7J0apGgoXvF0Ca086v9Z3Nff+oWpS1EZZ4oT2
KvvXwrjKYUIn9Rniq10RjNWKM29B38meUd75/JT1sFCZyZzaiZv97dn8Gz8E1aLx
y05JMaqb3ZsPR/52/fVZ+UjAIsIsSshaTh/H9+FQonN4qDuZ1YPguLxvryZ8bx+y
0MPTguEw28+eASmCEMl4imeUSD/mzWp6TjkFJfUoUlnVwsGshB9PcT3dIkYaMWlV
E4xfORf97KmRncodfi5ORFX90e7pGpYrzMdKVXod4qXeZh6x1Q4PH5b3Us+utbOz
7qjKC8pNJ0IjIivVxsCaP6ssFaVTDyBoShpQum0Z0EbPcoKwgoId0Op5pDGF8JaV
kUm5BUU+1cpVIA/Y+WvWnIskoBK+SRQU5LZR13PDcSTsUG1S1kg5VHuSZa4vaJNB
aTGafuxiwS0lo1Iw3W3HqDYTEm81RmvAi/L5MH4MQmC8TvYtrQqxAySnm3w6fSdu
AHkTdNOgKyqTRA+buWq7X83gaS6SdcpAXKJ41LG4MXHGHcb4CleKBgj1JO2sSK78
UXhBVAsdt4WT9fpQtHIa4i3Pr2hUs8Q3gvRi1Z8ed7U5oe9ArCiPybgRXKZi0eHa
1LCXtG3TbiyhFU6/S8iZRoE1pko/7SRsZDW3ezGC5ALZ5xhq1iAUYbCRXQn5/AeM
MzKYhwSPK1l+RFmzgMSbYQAEKq0DhblRwffjtXei+tRyFJnlWEG3G+hklhf00bzh
3/Oq7f0nuEVCdeMXCiDZKnIRZNftMBN9tywBlt87XVzRg6lL/M2NTzfOXnMrU1Ux
/Jii+QLPFjIUP+57HbHUrgMzqmTjEyggKe508065udw0D6F8Y4l1WOAg6WA5NH//
BSS07VCZQ6fIK63TC4ckch31v5S02zcFwASEsYOAtcFIhCJ2S86SZPDNQKHFgUst
H9uknRNrWsFYc/1Q1C1nFAEeIj/rjJfeKpoK1Xis2weZBP61G5B9i9gYldH4VO5K
3LhzkQfMjMxIhZ/Xqij4xA1fPPkCQTsC0h7AuWLscQq2AU3zBp7qNiEtQsITvnUv
BBjB5+ZauD83sOebElngYM3s07rKqhXilq6DHphHKSKykPteh4FB0kQUkbLrIMk1
Ot49IpvpOvXsFmxpisFABI0gEu9h/wnLQkW8ccnh21Ny0yPlFG5zxSSXT+AWYhW7
QFIXx+B/7NQqg7vV4Wi6dvEaUT/JPs4lC4clMU9/+pwY/RRG6kBh5JUfhIkNHeSE
IcYMpn2jJ9cMu2P5I6BCvd7ke4gYeCrsj9FYj7/7Ev4JeKZeNj9KbHygZISLJCvZ
rxkqpWrif8owj3868hqMIq1zs1BkMfEsYfVsFG3awke/mBtj1fGsLLpOCx/zLLyc
2OA2MZkskgcB3tSQRhf39A+0uRPDvirRu1EV/4rLI20P0jKqD+EhGR3DG8VSoMCn
+mp3RbUrl4cdmJKKs+CvZF//xtPP5WYas/laCQNw/HvMjcJNJaO/Aj+3iAVEjzqp
oSoYIWF0TTfwrcYMDpFB7NcyakWcmKbB6QECV7VepS7zKeAezKdjowhHFbK4HByi
2tC0S0k/oy9+d1naGcKC6kG31o9kp3Wo5yUvoWDPkvOumJhboxFG6Mqhd6+8cUqF
QdGDQNe0jJhL3SnwLgfyprYdm8H9zeDmoeNTbji1rcSzLr9v4w4N9yucCCmaaUbM
HidThhfpHj0mZYOsE09h2qmoLwrTsjJcdQQamVUMhxpXzxmhHO4xXg07dgJD08Kr
osEo7v+uqBbjD2lvh2zsjQWyyc1RWpFixEGI4woeHOiZeBUkPa5C1t1Kt58EZ9tA
reTsKkiYkQYPLnNRuDKhTKmQ2vKRLKqaPO7UwyUvkYiFilKiSLkMAh8RYnJWvSzf
YH7eB5Rl0Wz/pV7FRaxuMtYnaaLuztZvScPKZnMCf7BePncRexArrDtED/YaQdqB
jN7tiyYvUiHUhoqlWa1MlLY/OXFUkNcM2TXvxnaam74vs98XBaUqk+mPobbwQ9pc
OAtlohDYahmCmhKAFidn/gcqfIKvR3640abqsvSSmvRkhr0rqLsLxZ2VkOXPPo+4
SuwWtQzeFRH+A3IDmEFmOFNda3p1uahVrHwjXl4iVYUzZgUAe/OJ5H7JaOyLHBWV
BniI1gUPfumwFMBt6iksyWdL2rB94b496ozl2J7AV3vWC869R+NrCZ5E/xi+noAw
8/lc1Dx3geN/wW40+MBqU65ETqLwziU3SmDzrOZUOyTEcZiXhnrVfX8p0mV38qbK
9lEmEuwbYNZ7oDB8XFP+WTmszAHQ7WOlTpcD72OAc6Juq4gORlCpuGcu8SCpfgQE
mGY5Ocj2xKQKrwHFVzumRuSujcNguNYzmsKF22UA8L3pD/cUZFj8sUfw7eUdlnas
PR8M+HoC3tVL1fk52y7XuPUU2WTHF7KNwESJISIa6vgyZ+UD1OotlQBsPZP3fcHZ
SwJoSSq18FV6H4+dI2kAlFox5zm2KoytoIjIe1914fEUUb4+FWFNXFCuJkC3JkbX
TbGwZrY7n1/WFboMDY6FpLWt99dGWfyVr7S2Sb/ceV1WTubMbw7miMvYI/5V/qHp
KF4d8+ggeSxphXXO/eu32Iw2tHHjwB+yG8fqlwR1Xg83ubhtHpFLzGUbeRk2nU3i
t9lMGH0oTped2jJcfhDk9Ci1MoLYxa53id+sDyoym4dHYLT5bcT3zNljiQxfHK3B
iQR6wRYA0Jwf6+/YjarW1kGNQhf5MPIUaUWxSevcQ1t33WbI5S0SDB481yba40LB
TU4xOperVwrCaUm05m07RCtf/bRbEDyuM1VbOs8Qav/s98SkfX0IqM2GW2mxNRf1
n/dMTTszxPZZv7ZKly22RlnL3bjKG0Tw0VShpT/4dDsqNI1mZkTUOTIHixXrX8R7
oHMsH+9G7h47OOX3SWFtDnk5CgA2rDxGsur6ntWgRTjZxM9/MPhYpDLW5Qyc4IAR
KWz5TUn65/b8WFuAkPOShWQjR8DPv/vWFfxRBuY8s2gpkKOrfrqeNrfdUzrKS+k8
JmwYFewU3AGPqccGDMBW3S6X5U6iaJcksPldA8AfssOHenlp0KmdGO6rLXpMObby
Ar6PqEvGbg4vK/SAFSgocl9bYiSQY0GDwzNKYBvOi9NsaEXtyIzhEu5BFqplj522
1WF85p46q5EFnZ1l8iIKMTfS0G2A4C7hz8ZmcI5963b2L1IixYPW6MelCkUEBdvK
5wBEtf19L+d6p5AGsputSLEIu4vEzyv8R07SX5RiPKUzP3m7wAHJeozyM5U3iL9t
hy3H2C/KqHtFG3VERKmL5426HParZctz6nQAygKHG0SpFTqZj0ANaIv8tj5VX83C
IgeOYiWLcjVvrlfrxWShqgiBDvJyyl3gowDQaS8xaU/incJi/rCQUejC4JnB7JBH
x2pAWBNMUqWKRZf4A3I5Hml6+Jetd1R0lTGP/mWq5gJVPc0yz+QT3uwiEkSksQbQ
4Bhi9iDd651mSnbKW7k5m/eCGLcSyC0OI3J0e3PpirZMSkjNXBRkieC0en9h1dz8
bVTGubqDjvmw7kUcnBO0uH4ec4nV54cWpvzIWMz2ain7KAOSCoIlFXvpc5sNOz/8
sTcfcS4wjYOckbEsDnL/zDIwdzNHRC2U3oiPfwCIiAEij74wYnNL074CNEhBEAGG
G6MV/e2iGKdZ6WQjuO+G+8Id4BxTQ05IM/kCnP10wutzUw7/ZXE/+kdbJc60G1lA
6pTbxRT37NAb6Nb4epb7mnIIpw4xFoqis5RSHxbO2IF4yd2MWVL9JQxmT1oz3efl
HySacanCZouBQTX5oZDgeMQR9vRG9dQQOPQc5zaXbBcaWPWHFJNUdV1fHX+LRjJK
qwUFulU6mYmM2NDbSHc0LbTjRgv9TdS8sAsf5STsZQcuuboWS0aPFnmbrGqDqyjx
EI1Fa8z7qGFBBgW6egnsYO0+598fqbTjxuFIv357ENNhYAmHQCYXEOYI2kktDv2x
NymkCG1UYkX9u/0P52juoNUPHB4gN6Mrxf5k9zU1jrUft5MuFYPv1xr57kG1zDjP
zGTKtnBp45PySP0Sb7H11fVSDvgI7xXWz1zY/QUwcexxM4isbCvA8TqrjaFxRRYV
uorZRxIYkh4HtET4riF14PJMcJyRL9dFh5b+5atAtWavs7nJYLjmqvF7h9B309ja
QgUgXsnKOwdTB8c146MpyLc3kC2c15jrGu5RVi7EOegBZ7bT39LO56wip3zrxxTY
MQfq/y+gczqAAU1KP/RJkMJSpei3JpVfCzjqM/FHu9mOmVjxWBcDeJ0Iu3PLvEco
o7aLqZCEArxMZJuwXEk8v8Ap+WD2cB5N9Ljlz2TeO8XUWUgoCO3QR60PslwYFasC
96WtQcQsW+v54fjpn/OhGgvw1SM0R+xRGxWp66ny+snR4BxXp6hB6cYZfDpv1p0w
tulH/Prlko6p9FyA2L0Kp2rZ6zCMKeSsIWGEZRq+D93wdvvlwkl7GBW+aolrHcoc
pOIFkIL+6pea2Hlb0qn135L998dKxsgDvH681BQnvNqz6BHlLyMSZfHp0ltglxUu
DO/hiFBrVUyOV7IwXS0wa5XCyS3J01Gsy6v2DZPPDGoTVzovwsn6/8nKiiNzxQfy
yZcerygtyaIOezG7/fJgUIAOILUolOYTQJewkPvSZ0ZNt3C3TuwNSIzt0L2jhrUX
nhp2ZbLygqlMRqD9A21cIYJMVtaKjIEBEtJyn9+gxoE4B6SHpLbXRfpGvTl0QlB0
WjvIwf82Qnb32usZp7piNwCSde8w3FCn9wdiJvBJ3JXJgQ/yV6a9QLfjKJvKLqBz
jC+7LY/k2jazM4jsi1l/JXs569ZgOf7hgjZ6rBYaXo2rxe9Mq2rVywbtmlJduYzX
IzxIcNhOmEZ+a9uaXBCBcxuu1bAExQzGAQzBu3G75ZtnC6nKvQM8P8q6FPTFNPVr
+jD3e2vlzEeoLLn3f1Y/P88w/XgB04xRCwRYTl57eDjrqsZiqsdXPKVt8Wqj2YZJ
FUnKQ1NJoo3j2VvKMqT/ZCsZf1KNJP4OF9q07CaaW/XpahazmskXhUip949b7ENS
ljStFTjSyZ9W2AAikZU1idZLd6T8bGhZ+EAJOX2dIpEMCgw/be9S12RyoLpDkuDT
cGiRn8+pVpWpVXN61inOSdSrrOu8DB5azn245wgZUYJ/6E3o8IVBAhSQH5K7Up17
rQm496Wr8i2d74gQ62x+/1Ff+t/n9ypnn15kpIrOEjLyXzlEOcIBIZXaekBws2hY
mmG/xwsAAa1DyEW0sZUeyCRNpRKt36NrOIppb7Ybp0V8ZAB2/2chVCZW0hjWTr3/
FHhkTcXq3S5vp9iI0BxWNx+ODVFG/tyCWR3mnFGM0WPOyRetoj1AMtK159g/p64i
mgEIp9itng2VJ5w9zLdwfiMIZUKfk2FPywjLlpFMcFPAj2bH9aL8v9CLmrBQTJrg
U+x4n9TweeXPkzyteONEOful3YldqrU63lOouo3LMqRJl8s5UhNPJBHdzT04vO5Q
X4QO8XsFi99a8bFkyZLFGQXaItdsPhzA/EBWOQiC9T+HEPphWnRqX57cqMcZqNkC
j7qryKZBYpBRjggtuiBL7O+i62kg1X9/NlWgPGocFJvMc+fu64zIZe6WfFmYrXe6
SXCSg5oVGy8oCGdnJgyaHovnsVE1ZLMC9/hxVhOGWD7jL/z44cFJTO0j+bjMyy+w
pxCOiFPlwObFLt6nMg7aiKcoyci8oEXTtZoTs0pvKgL+W6jqOtIpCiQZfQu6YhSJ
5JzhG2lujqX4kbXBj3Pm3kG8cIr8l5hRJ3a4C808mvP8COzEHmOO7cGOc96teMQ/
9ndEfOb/ChfUVOBvM+fDzRGiVA5H0YKSBaW4txrydNAWeXhSnAoT+tvEZLsmfk+y
Q+SN2CKL3fS4iMY1imbItav1WNOLRT0TCdGSRM3yEO8qp0Cfw1f88gc8z8DMsNX0
SKyMCJa9HotIDphoY2nkDn3u7/jrBxT0Oz6+iSY39MwMPpY9g/4K8V5fm4sXpTxX
Z69suYxpZX46YRDVAkhK5Nk/S0+3Xwjj/oEWZTx1Fa1+2JNMtHeNZ2XkF03YpsLe
u9HW47XclGCPNTs9o7Mnx+agxDL+tHuInWzusxGq0z9GntWZE2WY0VOLvKMNrllW
SU88UTn/XIHGB0rFuIyEQp1zhOef1GCu0mfzPEF/7ea/PkfOH7PZvDL9rZib03e8
5q0kH+pIfgKxzYkMVUZhMF5fMNc97m1QOVpnKbaQDaXeBzCaA00zmskmC1L/STYY
/W0kxJ4NF7Ag2MYSvdRxzK5/u8pGrZmuBTnd5/Vc2Kqse07zidm2ARbWoVVNxS+I
L2mxgucKDyr1lDVlRn9V6uAGJQ7IblaNa6E6jwbVkxZQNhbOn8t2DZiD420Lwcgr
r5F8xMRpERv818yv6g5kwD8h2Qv2n2GAJ/Njb9WEmoNSoRO1BvpSzRPxNRNt7M56
eQmS05/cBPx3tMhaeA3a6JgbdEjTBs1AgAUDGjbXl4D6gzp2qZsoLMdZ7WlbGl1d
5OupiZ0gX5Vrkwca9+lfBVUIGU6C0flPqOOFnBhmW/unI8Mqe5QifWBZpKmdaSxR
SvpfggAtadNcvc1WCJmZakz/bWoYeSKQD0MdjZnjr7Wr2uM18cTUDOGq5eT2lc+o
As1wadg26Qj405/IgH/xvS3j0WKfL+l7pZ4ZyJlBwxfFWvl63uuXjW8KVqmS86OZ
g6s0QvmxcR2PrQ1qTOV1r63602IaqY0NqY6eikRSCLIo1AhpDSrAxjzBNi6h2h+6
+o93bC+Rc531mLYcQGFm5MxUzacwrU2Aj0hKhjmbWEMySZKtdAzM2xKPddA8KCVU
5HUSmE9FMzc0iOUL2D6JfjRqhzV1VooAFNvYzRoo88vjNN2lip+MSgv0uu2qJMFB
OwTJ3gBlV34apb4ZxNQfRrbnbIpqhjOhg40JRvjsdGUg/Tb7Yrdbbup6AWViNlGu
yfBkUU3Y8lGZH8xj/L3PJC+Wkj2fcHHhBJmp7LLDfaEPoEd1nDNdz/7ZT9EBghXI
7oTdkqnMcwWVx6LxjNR6lyRNSiy2lBNqbuUomiPlNR/iMw6ynauRLmdhxmGt9Hq1
Osr7A7T7x9g2dEwxupsLhwikV54UF5QSLzGCKcAmWa5m1Aue4YKkZjzJmYeyD0qR
GeJv12CwIuWBdqKSuVJrBojWnfP9m3zbZlUX1Z8bSADBF41vKRkTw/mzFH186ALJ
zKrtZn/Hbigv/j1e+lvIKA2YxvquAJY8ypErzeM3CsazVZCc0qQlD9a4s91KzWVr
WXvdZ41897tyZrrJHM0tBgyYxMEtS1KthCOKKjKBuRzs5Fix6PHqNKWIKNSwwceC
W9N/mHzzAVDJllTcXdq5OWG/VM2iac8tY/xZzyCWRcajzoXUQ96IPNrUkNAvvYDs
Hyy7Vh2vk8dQgeWocx2+pYhcraeIcmQNiMB9RaSarCj/XhSJPD4swO2oe0hMNHKo
3KHx0XRLCj2T4fbZEGABlmNgOKhkTfqR5tXqwKxjixacGT8/v7HY0BZBXMfOf8bg
nuOs72IwVMrmLBE1V9/FK52DNlbVNM483WDM9S3C3sOGtvllqbZrYOMgR+FXPjkg
jfguAHhasVg9t/f3rME74F8I8XZxrbpRPdkgtTcLb3TGKw+OmYhbB3MJh544HCeg
gqu286G26HaDC7yU58ZlOkm5knEUYGlhue7GOcmWf0sszilmA+mrxxNdmZLKPq2s
JTxl1bg4d470F5HpmPt8Wjy0XbnAG0Dv8yK4pY1z14B6u0QdTDluopgRf99ba1Pk
ZVq/47gkWM1bWb5Z3so385Bf4lc8WF2xTeKA59X0GccEjk4WoEwzOg8hqeqp9h9K
RQGL3QrOvKvFDuKcp0u0sZFaKJgV7L9tEM2Bdd7Jw/YL5lzBbUF5ENpc5aNc0Qoz
sJ2fbV6qFVr3pIv+P7dK//mK618UGsT046w7OogHEPcpv83vbVU0gBsrSuewW2OT
S3QIh2QoBY5SoxHsIJVfpnANpaF3a/1UPk0QrXGdqE/wH+01KiamtgyoPM4+I6aJ
vCj0AhtAkYjJoakxOsLuLRCEHC7HHUxxs9zWFWRy6aZ6c6BzL3hsyDrHiTitfJAW
gyRo3rgJm35JBKPIxfFSfklOC91CRliKzb+quq+IqxsniD6etJjVhNSmo9Pci+Gi
TDmKp767NGPcHFQ4c8P3eTEU4t7RdAtMBLZufa6coC6ZpVqiMfYesZGep77HRBbX
a51q7TfjIBYTHyOMG9Lpip5KoHaxSaDNS7ZAa/a/TEUEELcFk8Zg4TeYuNyzwWW2
RhHSN5ewGIL24V4hQzHtFqYyd96QAxUGKHFM01uUmy6fqF9dWzrYpjHlIooAOmMu
7UsOdBWjN1LKyZlkYRNa9ejS+6ey1d5ZjIqqWqRLmlhAcjq/mjPc1EOdeDrZTIPj
6sw2lZosPhr/E7MsGTCA8GZYB2zD//oBs1XTEIwRe59vdK9GM3jbeS+uvTaFFjFq
9GK2JZ7IjcCCtqBqXDIeP0gxFHb7PZq4aB7nFteX1F2kIn6sRcPDie6tvoAQhEi4
hFRhL58ZEvrIH7fJTwlfpMJooMCnNHoOLpxuKv6hninq95LQ0WB8HGwhslUm9lAM
2kRBoDOulhGtdw0CsPaEMsaA4z10ZR7roh80XqlIqi9n3nVfTNtMBUv+HhoyF/3s
qrKzZIjXOCfmZ10QWHnsfuxTKViTrPjdDNz3Gr2SgQRp6cve/NDZocMf5rFcKJyi
QyGP6JtxbJ2JcMxwQKjHp2s6Zj+6//LTCgFkPO7a8OtFvqzCz7Ui0Ye/Mt4jSmUY
U9WXYr/x8ROPWjWJ16GQxiSKrrZZdOoHvbJ1undPtiOCidltuH22x1IsvsdOSg4V
pOR49SUi548jVao6sZZ5EgRZP2IBGFQoSbQlrQaAfQo6ObNKd23GR7acv7M/eDbl
5Y67ks8DBH0TecTaK290I86kq95dspgNDMHb2q5/yo2JS6W/YwPG4dwvNDu+jIFF
H5dTxxdrqSoFN96xO6DJ8gFxwj3+A0BOYwHmjgBxg15IYfvdinG3dE3d8c4piN2K
LCwIIvWS11qKqsaEx1RoWTySw8usATPL8uLDdAQsyJWy4WHSz6/rCu4DCG9KMAB2
oOgN0RkcX0IJA7QsPvb3S0m76QtaJF3JJDKI7BAjtWsj+K8zhgT1ossu3U141o8F
kfaA6w5C/0xFpJUX5dfgBXm19wjoAWjpDEvBx9E96MfY6hjeXKZq/hlna527DFsE
dhs0w60MSWrwrr7yK5e96nRmB5L7uTWsi7IwgH7YGVz3YK7RSp5G6RbnqwSb/Okn
aJoMBeKI/JWaaJ+6uVF3h6ASv7hmMbvrwMd0CeXrqjKFAKvJLmkM4JM61ukxi/lp
ne9NC2dAfv0+T2yq6rwSP8wpMqBaTmuumAkihwks5HYm/PjqPgm6JLthWLo1s4Sk
XwhD2p1VP5DoI/auXYENgRz8BomevEFLhu84KcxrQWULrM+nZ29GSh0m61SgSHTy
sRpueb/+lRrZxARFPU7vAgurb++NiG/R90pHtf3xF6ZjuRw9uUMzRJwXjv7jxftV
/06fD3MgUySKRjdwZ3OXlD4qw13PS49KkQUfjSuKApTtvZZI9PNExUNM3O7cCxlw
5OsL5U+kFnPt1vGE/fQrLpbghJtiZSw4LE3HOCF9AKq9LYMlXw3kRq1Z9aukjIcu
Ap8BOh943hazRDO4rcrq5ljeo4hggo3jaamAXYE9g06CuT7GwtTHqXSOzN8wGUZ7
r5YwAAkNbEy0bIZ2BDXNxXc1x9ASdM9DQF5QzDjJMhMyP7/5YhFWA5KlmC9XGnNy
Ri5QppyBh6+UIc11Jf6AQpi+u1D0h4/p0+SZiISW82rLoONCGN6LQi+UJYmMJ49c
6DZiQ/0c4nWxN4sBAYxyaWKxnfVIUJmHppa0JjvkD2xkCOsa35MtpyZd0dRderu2
U3bwY2MJFWFCi9Kj9H4PvWDC4DN65geywp12eVBZWJcUoOIQxugZa8fHINDK7JK2
RidBbWvN/fwff5zZyXau0LhmrWFel00nN5W1pHvdngKkWbnaUOl5s8kA+YV/4TLo
NS34kdAieItMmuw3OR9/uNy5KF6najeD+XA/uJ1YnCl+yUQwKyigqAO1sNFI79S5
7U2KegfBkR/hn0im2RzLXqsOqf3zoP0o3D/HhN2DLiO4UvFlryjp1CiilukMhXxy
I8EnDeKfTF5J9N3zS3dLZ2deDr6SjcFNYMZqebRx17Kc+7S/+F+gzohqcyMMA3bT
DMcxx3YKYLoeaQZrauODz25HUWC+/HgVHcexBz30eB7TBypJ3TdxRJt1LQm5kIK5
jp92WLWJfN7g+ZRuTCk1N/8prGIa3oX/oMfoWx1B2kYUNGoxmmCEclPqmoWzes64
ZOH0L0KnLpXekMBQ0pCOnuzsjoxaUUGDLQk9yJmARFzd4aMAjQLuxNwQDTOqxy8u
ac0cfVlOEpd64peCXTrAicyVVW18rJRcYjg4oLxMrbjZ+t/sztICyPHqtSbaFaxl
skfNC5HQBlVUaX5Jlf3MQJOJ6Erfcxn+l6gH4VXaZiwWWbm7k/BwTSk4D/9pG5hD
9Ik3UmKJjDOzg5HTuHYLPx0tqyfgVw85gqMPyTbqQQ1Eu4En6tTSVBTwQUNWJ+3n
YAvDGk77kQqak+pj9mwt666/eaSeHosr+Kr4yd38EPF4u8TfhVqq0Rdv1sx1xKT8
yI7uCfttaKjVeJesQfldAzz2qswd/8W77bJdDDBs8GLRZxkVp37CU7opkhn/nboA
jX6PyzrJFcVbpfdKY2eLJ9hqOKV10Yr3DlebEtSfcTQEodMWM3zHbgDQWxYLIDda
39215fsbfkvhy+vIxaGbQ2myZnl0kp4wvkduThGSNN6KEfaEc10kOXwBgIOAIV1W
3I+uSBYp+mmB20631ggqK2e07JqWnRSKkhz+Qv/qp2LQ58uZtOegVePenxmtQSUd
cNkjB2cY9josvaJ7Ou2Qv2xHiHCazqOaooCv8Ei60R4zLDfHBvl0puYnVOP+Lfby
djmJLzUFFWp5LnaEAEqidvoUTfO0skUN68pmbtzYBU2bhB/ydntLwbPaE9mS1A2r
NjtdP4HZHLwoidWC4K1ShObEkIbhWVBrLgMkALkP89dDN5RIsiZqtxEnL6Dn94CW
fQGW6nOe07h3WMuvHg3WO1prr90g3QGF8cF8S8eDpl7LnMUBvyIMNe902aG8yRKi
J5fiKJcHt33isBdOsrr5b/s0NTcfoqaFoWmiWWiNhmHN1ByGMW47Zumv2pLUPwjZ
t3OE6nlsw3R++fp1IUMVO3BPNAuMf6YRgQqtZ0nb6d3BmWAueCqHAy2wuFI1v3ZR
IPJ2BMiwaioiiy/3Dxuf3l91hTHVQBgrf2YQq+jIRh02vdzdIwdCONcAsfNUt0kY
Fay+TyTsB31NP5A5lj0jTViKrGwwZZQXs/PFdZjV2rm/NQWoCQB0xT2jCfxUaSdP
YuUThqzANG8AGmboRa25e4sacrV/uSA/RofBTV0Fv6tPLN3SF65i7tAVgRg/lbqM
Q7ejDeSlatE/n0/OfPPInz4LahrAoOnpt5KRHNxCup3RSnnu1yMQNgGgV09VnNu0
zNiVFv3bp08WTqP+4dWbk5fPPtt3iYOBqopW1azsQr8BzPBv+ICfWc7SzsIdR1mq
0dEDMMtN2Q/UjnPH6Qurp3u4m3rcGQtpTSaB8HCeX13n6irqtLGQ8k5D2u6XoItQ
al6foziC1uGUdiilMa2F3r35zFUvyPi8SgPgBsZS8p+9sHLJ4M4Z+k0YY/VSFEZr
IVrH58HdZHjgrouBUtr7JjrNAYKDqGzS6gEqyIahCgAspfTBFbatRcTeCQMcV7pc
q2p3UDvf5MZMQccmSokMIsXASc+UdrGK94e0oN1VLofmcUN7viwb1tfWmKI3qYEo
+RKAUG1hIu5gTJd2fzXYtMTRhrJlxx9Sdqwg4CErYOqONM4YAyq2SQAk95jR82W/
bMTNYs3EvD66iEbmZJvwuGHSpwUuMikA5ydQ55Nu+K92YNFC/aLxvP9sFb02X2dC
hVKd4DuVceO8uYJziTnQpYZn9zKfjkJfU6rcdII2Kf/PAIuea0s1Sk0F3TIJYtDj
UPUVBfRtcS3JIhN1CKjEk7AgoG95Qs5CbEosG7+lL5amn8DIqU4b5AGYlQtOot98
UDqOmqoVypQeqTbhKb+8cmOd0hoyeswry5oQMdEyNgaCJ/FnVmKGIAUvQPiLolkL
ziMDHhzfvDBR35s5z9hBPtD7Rt45ftqBJB/pSfYU3FR1ONGWEjP/L9HP/su1bLSl
3imaKGSOd7dBtx+nNnKZHEDmBJnF1vG7UQkafolULz3Ci8nGaRnDL++pRJHcMJNP
ApysMOkEWe4rmqwL2PciH0hG6em4Me2cHz6Mj4O4JhKTxruH6r2DMyi7JEnaWv6U
2yb/PCWxvOIGd6t7KvFEHYG1kFo8EwQfVbaYIri8oWoIMlS/Kn44+Q5PCxhHcrzZ
33FK+Xlxr0Nn9Pss37JY6IqeLFG9cl13Aog7f/psm8dp8dn5pK/ak5p10bAxvOZ7
5G1ZKnRk8Q4AJL4ZL/7X7oW0pT6VkyJhyipZag5hG6Ii/7E0MpNQQDlSyTC27BhD
B66+CcS9YYxgQyhJunJD7rKVIXQ1W1+6HeVf/kfWJsq7Jcp3lRWgnAnWcKjLnoNr
CuqLJhIWfzMLXjutixRJEXZZHje1354wlaSNFB7PFjg5nSgQ2mVzW+F3X/lcDOA7
p8jsn3+8TmW/hqsjqt7E8dZHWhjXQLvnKaEzRoKzRxnZ/7nizwFe9yJj1kiuSOU0
z1bHYQ13LEBGgq/EFlDeeOBDx6IHyoSLLPO/PWlT7Che82IbbB3BXEVuJV4yToDf
0L02yuytspNaRye3iv6a0s2ir30jqO/RWU/Jd0AY7SN4RACbkRxbEYLGWa8sPFh0
+1hGAvNIbSCENzAca8YnydHRoVqVquXhiHavQTE6eNeuN+YSFa0bAatp7EsGd12o
9rxTj6xRtSnsJ6Nfh4rfNrmoRaAqu9fe4KPX3DihBt2KqO+s0IswmnTnSrreh8XM
JwpRF9aND7H2JmqCEx/BYRfg+2KjW3QECdZhUef9LfA8lUu6R4E/LUqH+AHvWYL2
sw4rP85c0FMHR+Eet9tn/Y4sGy/YMdJaSncfkIR2JKXETFhEY1+0cACchmxbPQ0b
yBaFPrRw2gYsR3hraY+0OF6fawomBbYzoCCbzFFQogySVwi2GFFp6jRepFWCs8x1
7eVvVo9zrLAYyE8EoHrAgQmIzjCsjKnwgh7m14/UHqMO4s/DUMqYN1Ce/jy5Bl3L
JuFWJjp69mTaPO+0+jjEo2gYH5Llu5Hm6BQKcLjeBHVbSBoB8P+jjMnRsM+BKXxw
V3yilmSgjMQClIf3rUULRRODOt1ZSZ0b/7KFlEKSQqoUrxAw5W2/wU6NHNDOGAkO
yjBBe9KO5J7oM/6Bhd4pXRerfxr16V+cAE03nPlyvC+C09e6rSGuLX57xlDcuSWB
k1fKEHzdTmDHnVP20mwaBjWJb81Qs6yZx7RjTTHBQ3N5ryUvaF1+rvAgjru05Qes
p9ItAdcR5QSFC8i1KX3ENAEWFNa3eHjU5aG8d1yIgazpaXCIy/hhp2Vk3RwMrL38
2zWdlU9XZfWCG6/RvsAZAyOdtp15JippN1FGJemUFDNC/tRxesLTCIm7lhYlprnH
St6ZWkiqpCBbLcTKxlMV/25LUoI83qvXyQF1lsCmTYf/jrIMC4ETh3+i6GWPo34M
srkqqLtDPm9Op6BsKyM17oOyO4fHyUJYyiB1DbvOVHag5/Iy2rdAzP4waJ/uxamn
dKKO8ozhFPoaDS45EBmVL7KhVBb03Ensl4ywWsx7Smu5HeiZAWCIJEndUHUcZ3T+
Fbk/DZTpHO5szJ7r084tZTIzjzJOxhvXwFAeVHC3pZmdxChdSCJBuQWiYSyRzePX
F/4pVNwlojfBWaoa+BEorjLc1JCsYwdgibhPEGR30cxHgCHo3GmrEoJSRQH7kQVz
FW9EDo0Qbk4J8xJngBIJWsfPxQJzg+281TcxJ2fCQ1Ad/+j6Rb9XBWSD2S0pMm0O
KYmNArt7bU3llsaWhmDFXGuLr56YAnJkiDEDT3gWdPUH7KUh0t6SSfa7SUrMobIZ
tq8GzDlN2DeIYRpLhgxVJ9CSoa5EA/haC8bVSOEsu3hbypAJ2tG0S2KwyopkN6MY
xSXyt0Jr3u/l321RFXQdtMVBt6LrxDe/JJtwHnR0FzFal4M+Zjzbp8Jdd9LGwWmX
rydQPUApMy6YKIIuFuX4WpWDCE+GWsCR0Zy+27SKafNB31Tg4WCY5gUVWxjH3u0W
TqjfB0NhyG7doh0TtgGKK2Vk7f+o85pV+ECpTgnigbm9idsitnH9YB1z76IIQmcD
HOfcru7RSy2VRRICrT3aiErC42LQyQ8BXKks7SO7aHAh4RrkzfaZx0bxc3iF0miZ
usEHJ3b4LoBUTZNBPHjfEVTvwDlT6IhKV4cD73jrWrDUQ4opv2FsM1umzmQu3rgk
+kleyiyZxdsVctTUtFv/xOXdOvJwDkDzo2jOFvG8m37JMSNdzgxEIIKLH83NEB0X
3tqwqj7Ds8b3cXi9s8ICZn3YVSXDt5tpM0UYR3K9N11c+8X+CIGwlodlLv9WfSXa
2fUQWValqDVNtLvydY6qJS8GBq7Nw3Bh4dy/9rmDyFsuIav5GQVCBvbRf4XAQWsU
AJJxh4KID7oyMXbcV9IwIooBM+rXWtpP/P8P+xTh2/Uv+42+z9QjjuVNQiZfs8wG
9w6rvylhWs8fjSd/8zsP6E7Ty14S1ZXG8ursOtV3VxleRYs3jg3JPdt3/nCnwbM2
UhQoSj1y8V7chsaUUkcCAypCVbQ/0H0jKGw6+K9XhEGk+aHc3s89B3JlslN/3NrZ
Z/LHpIGCyBxVEvDhp5QOKdNFv3u5shaZKBf9Dl107l2tqZ8hq3VY2xhG4vmrzM52
Gi8/WK0ADfz1f2jxFL4YckR80hiZeJAq6FLmQlm38ZnBCqHGY37Ci3rx99lL5UzF
KpX6fTEq6G4uzktQxNhhKJcW3Xr2Zu8qMG7Iy+JoDGKKx1dhrONPCINQo9/8TFFw
CzgxoU8Zhl0BBbZ443gIpAPbNH02pT2JfmyUhjhxmHoZUwNzU7K2In7vIW/f3QXg
ln6DzXggQ+yIcAThH7ULVfys298qZkMdLF7pXDEd0u1W85gI8VLKhnupxLEc9jdx
a5p03jNDssyBcdx/D9toMEVmuRxnCUCSTNjzy8d0zSvnAk4WRcHIybOT7zU38BPk
RpSNEOcv1i7Vdua5vsfrIK+qIMCsHWr+UEi4fCGFb1Q9DQVRQRWMJGTlbWlxN8F5
SC5eIesvlw+mYwM9JKbPnT0Af0EEOozYol9yR/Tj2+cLttXYnlLuqgnavxW8w9AA
npKj1SKAQiB+YRwwBbjH/NiqOFFPnq4xRjPvTxqYj0HmHRQ+mNSRpw4WVG9/G104
ig2BGVZyy0tLh49x2M092xcZT2cEG/y4bIJ7sApZGcFIHjVQXLrP8qzcpnZit8WW
jmQUYPNKhWs7qL8FIJjOdHpcK0gSki9z2ypksFGN3HKQRPyJ07/BiQ42Yv3JL0Gm
6Pic8RQxyegmqGA1Ti1SDep7w6Jjogw6Rmz0LeKstLaQlfgfuar/GozeRomnjyZQ
mDUP3IIadaEJocMJ4jQNrNlKGx9rtJyhRlcoEpIl3OSuvtRo7B+4jLJDt+k7TPHR
7AynX5+bID2PbyuW/oNdLjQ49j9vJWIbByrIoSy/MeLkjuHWNIGl+jW4iZoUEAUX
INNWE4CfgUujuozNUcmjXve+2JyPqg/2gsInf5vTlvHl8lhS2uU1P8cs1HhNwsW1
Ya+GN02bqJk4q+DTNP8Tbco+1Nt222sbCG9dv5Db7sc0fpde6LKrbzQ/1BZySiCR
rmzX23hWb256X0oQfAtwIbVPaJptO4xryOE23sZE5v4Wz4nYEx2q4lST8rd4ao4z
rxD0eahtAYITqH833kTBLOoSKxGpQvw/PA13qs3Ua9hs6ytjvs9YqxeW5IO37H7m
erzLoWoUM89DCxdDqrX8tPv6FY0f3pNZ4BI0/dgODCld98X6zmu4llk+DyJB3P1s
7hnZyKksyDNdVaEyQ7lgf6fCWs7GEFXFneWguQZ1DJwmTNkOknGbqkll54agVcbL
QjIhl/sDyonNk9r+EnUG21XbPsydG0bWBcUywUxHEv9J153ithbt9x2a5G71kgij
HPpYi55fnAZfsPC/flrGoqyJc2v9VOIIRENWSX9o0kiGaqJHWxTjacTJ8YN6sMiT
MpH89a4vsIiMLX8PCR96+z+3aMJU1sc7rdzsb3AMIsmsc1ArcRJf+MK7pOpTYtfb
HfczoRYg4vOoEM9i70Y54rbsK/dk2s5J37Uc/MQ9SLnrYfFgZJxtcfj+Uihf+Isi
6jPp6FnKeVtvmO5HvOE9sluhvTtDkH5U+Ki1CTbkqKffAebom4EGVKhnnGlp7IxC
EjIepkUQTcNyHM5uGbGGLRyc4sGFXVCnwoJBtL1m+eiMCeX12EQCHGI7OG/eZ24W
FoFMGks26DKogVGgQV2DQEqrohAu6sWNoit0vwEOU2yovB7hqRXls7Yf5gh5mROk
GcVi36NmmysPu1VL214SEZS+HlgcEb9iPaBNGKmBEfJVkLzuXYTWpbafmcVbfwBS
7f3q/xyKPvYp6KcGIEEXMBwusz4ZF7x27B7GDTlINtaq8P/n7AfXTbq4CdtNxLAD
9tnUf1CkvPD+n0KGxwE1hK6IWQFXsFZhtvR+bBxfNJPuBnPXTIRJ3Kc4pYzLbcQT
VUEa7Xg4kWh46XaYGbC/vVF4wQx8IYUSz1IARJ39/I5gFuIXQQFZ5etHj1W6pA2+
bKTBlWW+zQaKllGRm1FTde/3v3oLQNgTt9WddI47JX2cZb4pqxUXB4+BtSYirueF
hTlcIenmNIRSQaCdPp7FzVKa35vY5tu7IqrJLhr44uCTCpfk9fJC2Tgfa5r1N0IN
KFzW0uj4cwKrgU8MbMYIYgHBFOMFtajMPfe38N6/jNQ6UcDQpsJZxtrrUNS4aIms
qZ0lOnEdHHWo+R33o0gaSNPGZLBIPIjoAd17o8v1RkpAyCTxdC/rk1UegUJ6xHxD
VpiA0mCYc3sDR7xkxI0e/L4FeBVB7E8+y6MH3cPxw//rSFke+yhu1KhzEORd6lCZ
v/Qypt0AZg4vmPWgAP+7yvSIAfD/RY9a78Yy9Z3H93P5C6m4f8bRe8gu0K+TWFMi
xoPVUGBGvwfnssZdsBeAkZeeLYwFDxcSjkFFyYHUQHawqP7D3XQ05eMKxGpPV43K
SrHklvrraccBmUJIyZFLuDAK/NhIXqeStp838w7oUna+Qb29sq7oOs3uDG3USHgX
d1W/HTU20Ie+hVK2ovYCE1f/1vEyxFoQqvWGPqxzO+cr7JU+ydMuxNXXN2clVlfc
fvz/+mu1XfUOgYC+wWKh7d7Pkdy2J3hWwDQBVpfcGbv5+6MNWBgUp0vBiVR41qXv
6bUEeUTYeJcnkROTfI9iRDmGH9cmShGSfUECGk01ikRkvZ1IQHHjVlYjZ2jCaRir
wGAsh0Bk0zALXXHxucj+rZRPEZeK4tmc4V957ogewGe8d9OgF7vE2QjaIbBCr6Gq
EmjDo6D04Rq8QDuQLg55soHb3Adx5SczJPRxPvReSoKCTVWHmJ2AdnaGVUn+3hok
kKmtNljTgsMUsAR09xrZTxuDtS9TJFd0SIsul3Ehx62CUDLDeXGbEy5PAG6aCZ9w
UJAiu0BCY2SRL/pVqJ6us3vVw9jAxM5/1tZQI6ckbDEI/GrW/qey/bAEO417ZhMv
W4tossiD1nsKDYKmtHiSXMtIlSVSBBnCKojWLQd7I8JZFmlEiVH56NV3il0DPfsy
IpLZBQ6VdmOBepxE9ws+QuO3MNtQgc1PAV7mwurFzJ9fyy4Pwyv+S6kmZyTsHfw7
k8hpCsZyORykIbLLSz4fgyuQEoSgoPUlrquCEGUN3DlwzRsSp5BOJHvXhQxgJ3gY
6fYK5zyfzChYAq9eMmSPRBksgHswGL6/YcidloFlBpHUZjfDUjjvQfkjZitBW6xr
tf1I7FItwCyACytpromtEbm4J6ZWSpk19rqogbbNjIUfnbZbuU5tt7eNU3HJVMFP
IZaXQYqspAvWKGf4X0EWJozPF50yCZsFnj6fwjt/fRFKpk32S/RkqO7f0NGN94dP
tcWid48og3S27Mwe/PLdrSZJyU+dS3qZL6hbvrf7t9ZmcCSHIrzF3RU408y7Pxbg
05AJKiUYDRqQvBFVTzhJwj/HCEzJeVRukLHbEB4YBN1OxJK9ZdqMz7/vVjeDkNTV
ebaEKieTRHZijQBrnJtK8Hc5x8061FPkLV/FDoA8UJnKp6FldI5y/96cLUNT36qC
l3HTKsx/TCXB/OPUwpBUtJ3KCaf8tI6raF2gBu4Q5WzninCdpvArnWT3C96n6AxX
z9GdvZHtbYvy4h13BP/7BEQh5uLKHZnOLWmPwC5DhGYJ/oHjnDuRk5eKT1huw/Wm
MJJf2zSQmCB+Tik1+R2XwUMpGRV3+Y9TWZGi4Z8Jh5fVCHlZ4cFzp2v5GKdcpBFk
5/PzkTLLRw/wp5fiRJZSI7xcK/Vg348h87fSiKZ/OMAgmudUhyOTEqjJrmjvo5G/
5dTHNaH2VAWhOK6brwsmv84Lg0c0Viu/D1MGJYmCiu5kdgiGC+WHTHVTDT9AHLQ7
hwymJrZm8SGp9jUXju5R8b3pGtnGR0XGXNMS6T4XsJ5VYrC+4U1fjnYQPz5r9+TY
N2ZQnoUyQJHhrNkg9saz2p06oxMQGpcJ+5ZyB+nY8q3YcdDekF2q5g5CwsWz0EbS
WTY5C7pFtM5Vf6lf6WFCD+N7flbTwh183R07UwNHw5dnI7cr1qLZ/tMl0VgVJFum
QgyGMdkKuGCFEhmGRVddMGICrPQGk9McoOam6iI4T9zo2i++0K3zgLIZhg+SsU0G
mMjMGAjnxmOGQz637L8el3qmk5CcCdFlzdB90/pw81sCrIjEtxDcHsuFkMD7e2Kq
qq3gCoxIvzJGbhNcvw8tCJUyevcZb48BSPnqgo/iypjhwUrAkYEgZ5WfSU+F5Ci4
yVavZfgMo5Tf1d8J2JLrD65teZfgNXgyvwTM8M1gJPNw8hDJpI7G5tAKKm6WLg6U
KV5D3elTKBRhXkND1tXgiqYlcxLwDm6kBa+TmXcWsX8JNy+eXkFe2CI9Ai+7T4hB
+aQt76TcRdBCNmroiUajAmbWQesWSbEgh+i2PK24Ar82KjSatffLFtE/vqrPWIF7
1DVD4ZYm6+Tvm7dE2ioYO632bQHnB++yjv3PSUBHYhCAOqmGadjnUn7pXrQYHnVM
Ot5F1823s891MGpAP2wSrIdQx1id9C+PJHpA12SMoLawXsNhiJE0cWu87YTYX69d
FxP4RtUKj8zrupGPecwnLgFrY1/D8eU602vBTnVXaHrXBgKHmPScIFRRBEgiU/b+
T9haSwnG7xO2mqUM5UBWwte5GWSPRcf1ARDkK5fh3MxdKoPvwUxAUt8Yl02JSPN6
hQbjFeTqNX1xGhKG5EP+jxx7D9fRxOYr1A8RN0Ok9E+jwNF1lGjEJQ0hl/CjQ3+8
AdaNqG5r6Sy7zVi9Xn4yneirZbSRhreHil2gTlJ+cZyQnJpcrbcP7BDxUDcPXEUz
VES8coDrdHAFL7lBysWuKEBGjsSXmMm0AQ1oWz8YMHA8TPgdgeF6EZvcHR3XSp2S
eC5gkMrn5x3ndS03sDv+tO4yBijfO2yi0Nqvz+IFqRQcbLQd0DvO/RCI8qadNRui
mVfPXAszX5Qdyusd+86TSFZt9vQJPrqD3dzszVczO1FXBp/CtCLi4F3Go5F7h5il
HhPTTGGIbUuZsTAY7041XiyTCr09JKWPdDshtVjmnGQrkMhxrADAXYTtV+x6dkNz
ILs31BGFuXxoqr0k7XWbvOE1Css2EaXxwepLgWMbM+PGGpuyI5soWE0CIjcvLFDy
0tagDffHDfcLl2+7SoKRoektv9El/2TZz2zL8H5u1fSIEQaP/Ffd1zhyRkOHCWfx
eD4gRF2Lb/fKbegrKeW9LQXRAeBM6M4e/YRYkYkq447Ze/geJ+vNwO6bl8fBPvL5
yPMldydLM17ShldUAAfwbeJ6AgF4pRKBN2bbg7AkbgOFa5jce5jAlAyCSBmYTZe0
RBHaZHrY4raRHSdKgBsaiE13P9WOtPj1MNp4KousJ1fXsyGNJLzvMKwlVEoDgqun
PZplxhQnXjnKuYew/ukSx+hGLAtvWK7PYaQ4+QLnuv9ABBz5wV52db1z8T47C6N4
aZ0XvPExli/mY6HNU4Ew+xlZIEqO0MpyvkbEcazVoEQcprVqKOelQYll7lrSsCw+
PUezAxA7hrrnQFSRmhM1QrvHwsTtq8RVOXRwrF4dfVK8A4GyVrmQEEswdnI8OB1w
oGSrHon17/oZCzuSB6YJU/eMrQD9M4dsKBm1VLISDJXsiqcreHlRQOblYrH/O71V
WeW5fdPAfb7IHOuX265kasGi4jzL3dOZrA+/Nx8jB0aeBfKfU9QaLb2S4CkJ9R5h
/Y4sDzrCWlsljVP+Opzwznb+VZlscfW2/55SWp7NUopbbbXGeOZBtdYxHZLWP0uZ
oEh/e1rEFwb1M70dxrhj90E/22oGcbCrq//nbDNa7hu5kCx7fDtG9KHGak65u2Mc
1owv2KUueltfkVRePPSZrfrLjaYrSU5WgMkZs5gkHHSsm+M5S0pBqBrI6pcgfbhz
o4Zm/MXzhyk/lRtpqSunQCJ2NQRifX2VuFEwI+Vn6tGc5nBaZlUSBRuxY1RsPAH2
QKhHeiRQi9vSp1mQKaFJVrpIn92Il7b1KNrFUXkTYM6EShVhvmpL+HM/st29EtOw
DBssHZVnsoNHWBdJ3xY/p/QDIvFpBeep5d+IQ3W9D7JYmVYbEboxHkZYGpkx8p2N
St+mXLlNOHapgs6UAt2mm7GuFLq0Z4h6K4Hlon3aUyr2KjGdFivlDKBHlG+4J+fx
ywuujchD5G+Gpm/uuCS5D7oUL2BKxPFvjT/g18IqbmSlbitbczxyMKoSG5Z3ouAS
+qbnZb7CYFAvUoGYHr5mD8RptjH1N05PQnIrYf1d8dV8vTukYwHflAd9Y1dhr5JD
SexnZa3101z/ofYSwrM9idt3JMImyVt4Y9zrEmTzR+UuMxpWScHlgOuk8a9ll73w
CXJdN1c6rxauGYJ10/7Keh7MAZUZiRu/F7Mlz2oT68ppt+WpSs8fyoZpYZAOZFZn
/XbZAs76sdJnQkt2IJSQ0D8dA8bKxpiTgEYAqikZmslZAAbLPXtXwZw8n0VY5Km/
M5lBbsKwt+Qsn3MVuuoytaTNFU3LYn1gEJMFPUoqvOtVgTxY/cqsZjPti1NJTU3n
UhTJ6hA6edqe7k/fw6nqpLVQ3iqY04IyrGKHdWXjYgvHjs+b1faL3YlER4PqkBt+
s++IrKxV2RHiru6NjzWy/UuaR2TsYojfGyuWaYyn8RcV/HvIi+yo1oydC7gJAm6U
46xuMbKDcpyWF5+GT2Bi1vIvOe/1TK6dzOU7ow3dFJ7MafhJ+tJ8SXlhhUKXY0zF
nM89ePQRUJlVFVprxGXvKIh12KQEXApVTbODKtuvRI9T54gey7MYC1RcNGx5lrGm
zIJ0FwsSDKF38FPUwA4QhKKzE5m4qm/mwEjPcuDhq7Z74MFBoVyreobrGanle06v
nkVNS4j2oxJqCIz0XJQ1GZNvVElwFiZUVZSNUW+9WqyuxH7kWMS4e3/UUE/PnURJ
I3bcTnrC1YDT3HKDE8Xpb060ZUro/9Ld7faLTxFecjvF09IZwQBKIcezjW/Zyzwh
8fj3wpJTLMQMnQV/+UfED+qHySL5vT4w83MwCtZ8h+JHvW03thGb9K7YqSYeV6vL
ac4KUMCS6ZCWDsIYPpJvopdxWREmRnWC6C4DebY07fvGBT9nJbv12nb4CcrOiY/C
5nqvjWi9k8yZh2wzqL+r2l2utgCVfMcpuV3UKlZOMHS/HGi2GRWcmpSiZs0GHtSl
VT2aZE+sJ9pfIcSdhmYySZfQjxV2MIKL6d3DXVYfPNdWW06fbfjhS+2Csx4g9R1Y
GqKRjoxySvHmEh0RC8p07sz34N7wZfbCj+VWGrL+zsH1bfUAS5kjk2+UC31WX7x2
nvv7Qlrjhbw6N1IT/3o57Oqp7hYVFgLcAA6KJecXshRbB0MHdJuXMLXMnXHtuTQu
Ju+Ao9MMeXypUt8bxBDFIwqm7jPta3UUJ6kgpfV5tC2+jfeouljdlI27+nDNf2Tu
87071CoJoM98IkFl8U9iBe9s/ruU3pd+e/oOnbTD/gwUfD2YoeoICX49bel7LITK
AkZyGdt5Q97iGhDu3gRqKAuW7d/jGwl+IHVg+1A2EnvPWlNaebM5azDjkeDy5M/m
e6dbHDfQTEz6sc/fgbsXOyhAWivzOwa+AKWalAVFop8RvLXLN8qLmSzzVLBX8zBi
OZPx6uL+EHgbzCFBPbpL7hgYUN2mfiOtktGu2DIQS64dLsPog7CxigBij9Ja1htv
1TQhrCp9z4mZYVtEshS8CHLGwjKUGr62PJn6NkLyMIMgfi3QDSl0Lj0ViEhVxdqE
Xm6jacudoCEkOSUy7L1Jd9yDHO1daEUXLhoqdhaOM2GBZYWLhwHL/00ir4fzEajr
G4C2kLQRX5X2kvwb3Hi71AtRKr1RD1+rjKvUZ5nKm9W1PHxBtCq+WQUzypDIvy9S
DhLNZ+CcTW2zM5THtApiT88O1EpIjWcqupiQiWwRhgua+NamTQmaOlN6dodE6WEZ
31c41ibrlTpBefGklaIc9CREKmGcVaMtd1DG0p5ez5m4q2zUX+xigR8i3C0+eRXW
T4bM1Mxe1eigakXEIwMnuK7hApfTZNDObzLJ7ReWwCH1CFuMs/SWVyrOS26r5qSc
GRNEk9rYk6oKeU+9ypeAvn5V+/MX92urEWDMK2bWmpIZ7iHp92H39xY57k4zJ7p1
SbW3CAB1OTXcJ2tqMuDwSK1P8XxkmI9zQUE1cBN2F7nFMr631QWmHZ33iVWCGy41
B2/Y4eHihYppaH/X3Ts0R41Mk/Jl538cX+2OLM3od3RbYPBh2b+qTLrM6ipNCQCJ
vVseHiEjhx5BiT7SPcoQ1VHLEieiwT/KM7KsijzdtnHKx44yP+NH+5XQxWN45g/F
1Expw7ilVkuJ2NcTdZLRFxIXk5I+Q2mMQHdDhhCL6qmxsaVYuWJRbG93PCokqvpe
FnwlnucJH2Q495fc6dmUBePc5ove5fj3EyjZpqgM5S6lj59Nb7ZBZCQ9QnZAppS0
vpiCRLk4Ahih0lIa4UpHpu+sKQBcbzc/E7XoRKvBPwEbV3w3dy11pOMQ7yCh260d
NY0dRE8OKY0qaJDf9oo4tOyRHKvndVCz546ytdCkMwlbcMWJ9ghUef2pVIlsEABG
OTRcrFhmmyuxiby6sBRhhFYZ2bQsrLUanKEATEze0LhoNPdDoSBNOCylv/if1u9j
MkqT+One4IrowbUAAdqetPgYeWlmn84eds8E/SmAXKbWbT1M+MljMThI4zd58/8l
2Av1VG2QJl2saYlNCVusBKo2QKkgeqzVt07cjvO6lYXCmA58zs9VE/GaTFYMn4Zj
6OyQsu/ZItjymwU/EGpLioHxIA7VT94HKpbnfEGCk2gUKnmY0kt+IhL9/+jE4gBv
z79SvM2ivn+5BrDWFSN8yJrdq5Fyv9KxvWjvbsj4D0EXaACCqvpjoJTzmEF4FFVs
o0/km/6aZO/NgBN5LGj2LZ9xXbr1NZOf3dB7Ng+y817LCkkjSOaFr9nsobA8364V
B6l4IBOUqj2ubBowih5cD3IuKi5KzSmbnSvE2lCu4bBBUIIaxScmZDrbm74S9ojo
SjiXVlTFlIGILCeo+uzAs4Dbb8a70+ZUl2IVtIZdns0l5SDDBNlAXd1AV1HcpRc8
gmINCZaPRN4UeLmbZlWcqkIyJSsNXAwvpcrk3kubj8i6si/2jozwPUbR59ptHF2J
rsjc8vDGRjfFgYgrUcmaMZFJAtBBPhzfsgNsvk86sxh8EqYQXWbkT0GjB+2KInht
24lNBTW9dyiIP+KrQBFljxoeAp2YhglgYFC8RCLAmrlOsTpMBpJvwIlG3OPtRtbh
M8IK3s81mpmB10Ef5sJEsSdLuBR9vXk1qQR96wac1zgTs7Lyp7mzq6uSyZTFSfBu
dgu5TG7tUSNgaFCkJg2XrsBqc02ctqFHx6MWBAt3D78zL6I0NHGBaQG+d37AvSEX
5d1NSewzvCY3PAWwLIRkLVf9g2oHqch00bmtZDrbp7wNeDrq0g7pZ1EWLz/6CHmy
1lMkr6zx9f/nOFbzhyXmjBkm+prxlcZKjCt1U07XNd2AHwaCBlyiMVcL+Vk8M0x6
ssee/j+pwe2hQq9z2smAQ0pZ6Gx0/oqIIvFd9aUAaVhsgocTCiLJVqyKSInN8UXR
h1vmqrcDXj3bG+3pYjwtUlb4+3ivF0CpvtjHNuAQXpme+l5CBjLinNNawR/id+QJ
uynSajZHSDgRtYReyYGp4sTX+DV0KfqEpPSi1XeQ8bscOX2ZQtsBY7oXyklUjTYy
+FCPKL/lxwkXhOJmRJq7luIwo5RvgPit/bDYEHhzjo7sK8KZLBMayJozI3TDT6r3
dBPVNAub0wj/PeqUgIW6MbcGFiCihea09PTwXHElJuyjavLyEsecDE4Bh69SFIN3
MhtquipHoZONcRJmZVsTC4HkFCqR0s/UnJC7cjBuyn8n7u3ZL+yUl0PUkFF5xZW2
de+AWwoCKlg3KCEvgyjrhLvtcWixZhQF2Ca24xn78R/DqZmFlAXR3SaPjgNa41ss
H9k5ge0E5vATnZJJC732cMddH2EzRiLrz0n9hSEp9io8kGn6QLS3YdRwveYEnTjH
34x7euxs4Lt3d7NAlGdB4mRGDlNYP/INXJ31/hNTwATP4uqPyvrLDLEm03zV2M/h
17H4rFxtylGkeB1s8zG6JpOIOMv7pUGOVJtbzqTraPX2CN8wdYGsDoBVgjeq0vHN
L5B6Z2v6uBRrqMIvtrRZ4DzuZ05Uc4VoHRzMmlvgANUa2qufi7f5qL6FbZEwy7IL
UAGkHX4NtjqhqjNw4mt5rshci0tTudCxR8N21NFvhIC0VuKsBZ1Dl8R7dCxZr5es
vyyj++Z36jhdC1AdC+eC0Ef7DsWo6tWmG0l2WTQ33eo/jP25+tBW/nvytTl3zyUy
e2t3ZCrhMZ6VCoCOSYO6q0VXTMNPnxc8JAHEkFlBEGXQ2Ju4t2fhrR/V4QxUgkE5
Y9t7VJUYy2d6mGW0vIq9y4D+WHRiLWSnAlplBDb1lMFGZS0LnKssoH/eHVKIBZFH
C1LylQJeuCfP8uvpTg+A0j2h3et1ImYtngn/KU+uk1mflPnfmjAwC27ievGi/nGh
ojiWqVt96LChMYgDFhBtOo7QHftpDn6mDTooMoyrrR+f8BXIiDSAiUCPsZ0TEoCF
Q0LS/d7uBa9y3oLD1mMNFqMOHhk5TxpwexCDmbufvaYN6LMwYgeZq0Y4gey2N3gA
ei4iJYQ+HsgZeYhRNaDED9fYMrp85jBX2SB3+M2O8NiGFkgWzE9AU3DINAmU2uIu
Pi7ncCQuMDMJhcysjG4NRUmdPaGVKfFHyMH5gefHPF4t3WunyA/l42lpxBLEC0pK
6WGE3KXpMzcsyi/YMc0gUKx5IehmucC1lFhSw47cvKV99bjgc2OYexhQPHUadaFO
Q/kq7A7/31g3XtL0MAA2TefF8vZRFZgWXVs/WNXbHvmUG2Tzqn0Lhm4XxBX54mzs
sn8/AJH6YMcs/nOnMqS5R7etn4D53Mu9Z7CpaUemYl6ZimxrE3xifd34wM1E7iyO
EzA44hfuSBq66hrQeQCV0hwkEnU7S7db7Hef2uLiWmU0mzJEG+asUXo6gnSB21ul
sw4sz4pPMSvd3UwLHPd8WTardzGY7om0Pl9Q+LjQl7F0yMturB92rirdh1NgARKk
eEDIpb2dnJaayJBNAWOOKyUuvC2zcokun6K87EemUKZ8PtiMUFnjmYk1cqFc5mla
SFHyL+Z7FFM74v4HjxZTnRueZrbTXfDZfcgadCQgHtTWvddz62BA8lFIxb88TKv5
lj6zTdkYLLo7zuGyT/YcTL1AF94T2j8cRVtKk7mZN8lxKyXf9BZyMXbv5AlH3oXs
gX1hFjv11SICy6oXD+lkL1VXbk6Di1NMH2LhKvQpoCapns89ExRr8cDcrVFqQGwi
uAdIOWXWwIgdK7cJArK1gQttaXMMiSyiYTyTsBNZyqSEWoinUfqtHfua84HAPZsl
PepW9zCCLlrGhKHhN7/19NN0iac8O66wb21T0iPkFeFyWql/BXsQEstvV9RV2pKq
PweU/VM9HhAliRo8mxtRRPp6TCMwZR8uAicx5Vgm02rqo3arPvTw/oc5N26gJxA0
Zr51tEJbn6czUnCnfxTvyf0wpZnFgGSd3KRf6SGb57tKRC1ME+ViKi0DHzEdCUVw
LkFAtqnyy5ePIj8LL/3D2u0JN7Gza8OVfSKcm5Zl6GKueJUehRmpi9irrpFIihQw
DPzSoJ20j9fL1yBVJnaHQaNC7eK8bxiKgOMME1lYF0fp2uQxQDsyPKE9Z+q+mF03
qhv1ovtJNxu2KFpO9HonsYdtB9VcA2AQfafEBC9sC8h6/119IGWX5Xk8lZo48NmS
Y7gIXqcEeObtp/DAGzmezxTHxTXahYG0FdMvHjIjxVCMNdr3L0+2PDNpTuU+u8aC
uX0psM+v73Du7AMe0jD9z4R01pN4R7vUKHD6o6xizoNNtNtznrHFP8TFN7az4tTp
TtM2jijqj6qCHZSGDplN5kfcVmCoMM2h64zUF8bmdhlmrB9x3FCATRh8EVnZEJfl
9n4jLQLshpEDj1HfCqUf+9CdjOooNMmKn73clmpOhoomLK4N+kuftuFCLTnhS904
fPMtSAFSrwyWwtmXXsYbTy6MVmSF5zKADLpF7A3rkXor4EXbevQLtnJsvDznIVCE
Pn4M9kYr4eJ290MW44oav0NSMU5+oIwmTb37QubxuMsyGqM8GTBVPfhr40xmi4no
0r042RRbQkB3AplmEr+KZP5Le5333EWmziIwmTG7kWvNa7Tk5qLpvY//iPWbbI/x
N7BQYyOf/CN7aHjpj7lucfIynNOagLmfN5t3CGnSnQMVNgG793AEd6mbSQH4oksf
QlRTU1XdP82Ht7we8HS7UzGelpOUVNhunGEeoazzogy/vB6nlJquSIQ6oz7c5awN
MMxSBq+z2B3vLMfBt02tQrpnLZkAdFF6bQwkLvT93s+XTNtCn7f6AvyI6PiUkeJE
BRIU0f9rHoSrWQ8cxP1PzS5QEtw+79GDrqDp/yWqyj/vFme+kHKu6XIvj5yGVhcB
YXmO7YOK6C2ClH6+QrFH2y4DOCV3SWZaDQnfZ5b9KjhopeL9ArREH9xnOSQe95ri
aAb1etkYL5G4iFA/EytoF2JGUeS4YmMlkx1wmfreCfCoZwVeJQ/RPWEofpJ1p/He
zqMV88z0vp9Wyj+MscX+qxbEtHbjj7PTgMucSvrvYxlCl79jwJM1rodqNZAE0c5S
oyNdBnBGuNbCi9IaLYTgsWKvE6QrDvyNlhy6GpHU+xvmjLxCeQcVpUGnJwApMiDX
hKq4FNErTHRw/w/5EFzyOUoZtOrvx1QpvDZK+wt1o+djdCkRAfmVfdwKSi3Blfcz
LhHUtTuiHdCcVn1FrIBrCCPwKA7gZx1Fxh9wiz2B7cyznOYcVMxBqcNA3pgvxxh8
to8W8qlsqJmsqVi6YhRaY2bIpkWnoCEjyxn650CFwNH6cPt7GKEfjyY6bv5dFMp3
5wBHXBaz/+1cVTwFG4EzCmoHqmUTmTUPTJipYdglEJ9ebu9mVePGW/f6Lisid3fV
kSYSu8yls/lKlEZuLZ0uwoVHbe7M1oi26rMA29yhN8AClBluMPBrnw2JbwIJAwjQ
qGfmq/kbz5iNP24ZwJtEDghJDpgbBvQhOeOwpfZXYuDGThgO3ukRKR0uquf7yKr0
UrxKaaN0d3oUYsbU6EO+M8s+If+4wCrmI6pnvqUX2aOUJCCgHEMVavdn/ERjI+Dx
vXQlVSgQKSc4ubXRZxHr4pxyFs1QbGLyrYT/uC3Vd7FayQnDIu2rbdWdOjH4DV0N
uYImyrkCxlyoipabJBIY112fCYVBEwlTf27+tiUA6KxAM0Sm/cYqtN6VPwgM/LpJ
KyCFRcFZMQCJOPALTpXuUJfaLrQ4/ZP7a3Sn1cq7WdZUjR5ydDvYLIpIqVL0Bkrn
3Wg4IkZ3btJRjDxGE0auZ1lTY1Jewj0X5nZFFuLRfr4wMOczBMlt7dBI2FQrQqD+
LOF99eGWx3wY/9MJrTIVh3DteU0CdnzxhUoxmK01JwkJjQ0uJe/bahgIrmQnQZFw
TmWpr7LI+bpzTo9Zxn2o9LFHs0IPRKaLT8THNkFEmjkOmLizKMGB6wrCXeEy42Hs
9PNbzQTNJTOmEN8Ul4JiZpNH/UM51vC/ogwVhz0ZfGl83k+xqtJK8QErR57hNJLi
4oLgwnv9PiQFwI8b4bSkAvG0fzZBK+cR2TWAXr3Om+XpVGh3rL7W/acYT9P9L/+0
MOSqHhuV17gLyv0iBihWFTpyPZmYEIfOpnEKYPiWFPlrbRW/KJEgpsF5tXQdy7Du
uwgQ0IK7sUcI3qAS2R0hNSRHlIVhXmAc5zWVMVRXzA2SwbJV2cfiU+05+VrZLZxt
1pBRkpQNV4VVlL2pb+/Y4VGK2hDW82WV2t8BxKgwiVRYpKDLhZ2CD1UE9o3vdwHm
fewqtEV98FI/vOZNwJdLymqW7S5ziUFdwcQhwVhC2rnLmHv49Z7mN1IvasQCIkkf
7tnXBvCOypWSLVO0wrcHm6hXTvC5NjByq86qiMb9WSC2ZVfzseyD3yjsA6QajjgS
gOg06e3HKCvhNjt/g4wvWxYUbgmy5gQxNkUSsX2JESO7t7oKHeMdiVMnukX0mRQN
BsNCl47zGRlA0hLkCaCBF7KhcQhy56D+ozMCVfWngss+GhucvZMEsjeRrde+XKPb
ni5+wNrWgO7UYc1EZLboObWUwe0psdEbnUZb3MKp1bvRwToV2NPy9hJEUjHn2f3h
dbs0/PenNH0kB88aHmu/38wgUxGHSqJeXHT5zq/lV7jkiU+c1RMg6+a3DASAb7Gx
TnSBtqafEjJ0F23XKAjW3I/FWjvvedQluK87Mnaa1xo8B4WG3Y7YMg9/9Vz0QF9M
yelC5p/LZIf1iP9R1FlYiv1PIEmla3d4j/L6gq6Nfb90fsaul9iHev+mzMsIKUOa
FA0DGOxR4qU0VdYx2ltWSsEvnMg7hq79sFZh6ZX9dShCwSCmF4sTEbIp8UPSZRXN
Mc/ZI9MTORtPHnaSMVJzyEOwRWlffAIuqjUUAUykWxVM7utbdPIpO+SbLXPZQKxl
+UTJpsW6nxYVBiKTJr1MFEp/TQy2HBxHpP8THBSkWFR1fJYQ9sKnTfTpDln6/jug
Yo8YlZgxlt1methytX7pQQlL0XO6Y1f3efwPMxcBGpV7m4h6Mc1FVo0XakHipd9b
gd5FZDdWV9ECkFYqfDzMWi5zXoYw724CVafrkiooaTpHYIS69R5olvZLgHkVIIpt
UYPzfNraxqM90abc+eFO7tD1Acpovn3rsSF3CUsu2W5NnfFeDmquvjMaSK9e+Wug
yE09biA00pGRzKYLaboaaXYBLXJU44AXBSmGynZE9ZELYQ3CYC5jrRd7348SzdP2
4uaC0Y5YBtcpQeuoxrGeFnt4rE/BlTElmZoxDLPzoJvq0i5/9qlB8ajWyU99Nm7o
xvN+NgA8p1hW2sD3T09muFupxVquy/wR6g+yix/RoRx3w/SdFzRuH2c8KYKR7EE4
d10YskQLfJGbu5v2dGFnqtkFW4UmyJUF1a0Vx9XRJx6O7TNh7SHWdeHcgxYPFLnA
cYjtsq/2cEtQ+mAYt+NoV8FZa82Vpe/pnyNkXqRRCCZpf0o9NFe0GEMNWfroak5y
KVWBOACBpUsVA9gQKg1OxJGDucPwhyu+2PMrV905fyMEg3jrzgDAyUIY/inMvaAE
NKt1gMi0CQ5hsk/Z94GbQQEKkcZAWuMfLWpbe1SfDu7eUrwxevktB8AS/tL7MeCa
jWHSrJtq4EiYr3Fp/djzdU6fPsxIQY4f0rwQk9WhnNBUcFJ6TFKYNadGco627QPS
a05HFVgwDIg1rJ8CvLwrzcMOu6nG2qGXU8srpB4dHWIkf2uEDvbLvwON2KwnufRN
5wsY8arjEq+7v3ObeizsVepWm5uie9DBS3fxcjFlJ69wbL42r/pfhjaU9UOWVA5B
HpwsS1+gBqmlCedEeXVnvGG89RDD5COxRJjPpTc7bHYxpY/OnKEJPwMxY86yzRaQ
zLTcwt3Aj6rRlI/0ENjnl325IKLGFP80mvd6npdZZ/V7Fy+GKuz8UiYzSvDcfQ+n
kSqeW11kQWBC2SzGpvEBOKghlEPhW44S8sfDJVR/KvP5s+L1o7gPfnin+MT9wVsx
KcTVFnxwyWGqJu4Txz9IgswxhnLHG74SLIdb7YpUOq0RwZbBgKi8dmkVU6lO8baK
mw/8wVjyVUva5cUYuixXIJzPnTMmMXLu80PDnp1L2VVUz7eW/iT4PZ+fqk//m06S
PXm7ulOKrq6xzz7ckOS/d/VNeGK0Nrr1QAnIIJHbeZtvaBKNcDzoeYFfWkHTwx1u
x/ij1Yxl/yQGf20xFNfG+1iLTo14tQ6WE/WNfQX2Wf7Nh/ozXtAlP8PqguQFOcoK
spLzMnEVdfIAFqyvuzK1GOP2kwsHLBLpI1uawEP8g93czzoxUWQBUsCRJMneZ/mG
6dPmiN+OqJiFmz8xmjv0KqhbhHYVZ1FUflu8pPcTJbOCyliL/n7vdxEDEPRTGEQB
3Dgyrzq/P9K4VFz/LMra2TBmdBvdJtAVFfHeUwAQsv6FK6dH6KGvDfi348YNaT3G
7PQsfrtuXlsnWiAaZhp3e5y4SdLtxdOfjiio+0jdmt/SQz7pCO1w1MXK6bfVlsHf
J8F16LmuscFMvvXRGJXO6OXEtf6oc8IQ+oV5QrTyXAziKut3kUb/fIM2VUwBo8Wx
0yHVpUL6Aj9AnYLB2InM6sYZ/pRMcI7I+0hmDBea7NuIKfyFRK+EmC4rp1Zcu52W
VQJroyLkHKdv7stAb1E0Nzz/XmXtuux/IEi3yAgajW+G5q7gvGVwq4l/s2VMp+AZ
yAJmXiRQhlrqyDXNMTwLha4VJdNlH8IObp2wl9n7TYvsba/CxZJ/waitRky3E0e7
nzzU++DiDAD3wroY2fOuZapXPkRF3a7+XRrVK2W7K10AGTwTXcqN/dthL3OUEmM3
ZaMpVjGss1DwnBmmHr38lNph3JT3HPSDxJUVa0jVAUwANGH295alvRBBnU1/usiW
AzkgPvfOfrGd3j5q778zDK/xZuOJ2Gg822+rPQfxABTxbcKbW2h5sfqf7m12y2LX
xxywa8wkgYE6W57CJTL4BJJRb08pW2LdUmLWpde2GxAymhN8dmzPmgU/aphGFRG2
Br9mM9xmKNpsINQzPCPfIO4xEjm+LqDaBOmm1va7Mp+s/Cz04pQhqJluJrvxzpLo
qbybE6mD5r8LdajNQ4r94G+FCJhIpOOdsQWAOfpwSSPAC6K5dRFYvg9gZaxf3fg/
+jOWMTmjraQKGGUu/aqGqBtzl1lItwASiRNE0lRDytzl7PnHTgI5l8FaCIpnv7u/
e9azxP05KKNRC3raHHL4VD1SS8D50VlmeyK28b0eKoO+pls4srjs7xzUiXS/DdVc
Ezw+5rBVKIjtAaIFWTYPDjGCdW8uy8moW0vJ6KWmFrrtKx2bVxOhqfeXCMFm4mvV
deeTlv5htt3jV0oMik2lPU+zLzajfuDN5AFpcLvOTbA5UJmMxV7ME/xGnuetwd3P
KzaQ5eLYXuPgK0w2WN9ARCJ4dRLwpf8e6kaFI20RddJn94LRWPEWeo9h9DyzDIa3
oOy9q4JUBaGFnvvR6t+FUYAYkgoUlw47CKKiPV+4Ky1YcVrPBtdhK40oHFa23cEH
creoW4A0XfTjI6a5ZWZxfzedPl+EKSCUaWd4zjfIn8Q2yR+H2qr7GFLbG9SGE5Hi
0sXEeNfaDdpKsMvYlWTiErCICLEc3CPUG4fFiCHDmYmUll8fT7uJ5OTlzIjd+HZ0
mtILL0RA/skc8TSkXcMPVc7DU4M7X3fllG6JvXVTb2phOJm5+0AehzAVc0bnai+r
6046wCVGfVn8PyjL3gTrzKeyaaMtbtmieCFmsK2y4DZSrgfYFbhB2OznO6i75D9i
ibE8M3DzxRqQCdbEcEC8ALfdJ8CWodEYJ2HxKfT4AllRQuc7Jd+JLwiXonR2Xtmf
n1ZUeVjC/adCG3jBLQYfXOh2wwOQ3kZ39usiVEr5nIcmF2bkFOnarANswBz3A/Bl
m4dhMHjQv5oaohSLCIeHv/uLUfbXEz+A14QkLavw9csqDWCyuyUSgul9aPtruO1G
LgHeAeqWQUkh+XEWKfq2b8ZnrM+yR19gD0nrz3BVDQBsvGN3Y1CX62QuwAVrWDC7
nLlM4b13Cb9r+CfVb4FA9N7qcrMy5Q3UhofEID0Q3Z0Lg70Oo/XY3djWQS6DCCmS
FSDDB5ehqbk8IVjaOQm2z7Y0GHB9T5UF1Cv8aI1DPCGKoShY/O1UzFSPhCTXX1aN
hadVrUlDcnaxo2OQxSTa6qmRZ2h8f4d8aXTfXSXf5OzM+VLz7nuKEjEL5gm9OeQx
kM7kIfFYUPrz1uzCy8Mud5c8jX3FjKSt+CMmrEF2v6DgYJrY9ri4e0i1H4evuE8Z
GywAQ/IHVLbO3df9B1JP0OsO1ehohfZx/YVFUX0o1Ri1T9Xon6bT8gbNDwEW5KLf
ZHohvNkpMkDbyezQygis/z7IeU8cCa5Gbb7tKoyhOm9fMSawI3WyseowStw3xu4j
3ZXJYYUKxYe1pbLWQKAHXHPHQUREoYtNxvYSCa24mFh5vyERCqvxG7WHVfCfAkqo
TB8cj6Giw86h0LWnojzfGHTKz342msSnsDnca37ZfalM25G9VVDTwnF4uuhT1I7L
r3vXvAabRmywAkoaDwduvYseFDSsZp6eKi075ylc3QEIx1MA61k0mV7Jfe+J3NKu
gOFnzVyBAMGibhbCrm8pSTZswFoAiEV8PBw58eWVlMtfBSW7PQqxZUoOfLdvSElH
/RlttJY1cxbG8qdD+aYcLYoBtYq2c/NoR4DLa1KAbjuouTBsqJYKMFtg15spCSh9
JMU+hIbbV15P4xoeroQo9p5UTLnxYy5iumE2AQxWX0bSjkSIbnlTB2buQoH0Jcrm
y0bZcAGM1m4K8SWuIvOLu7us+Jho2sbLcScfOZkEQlKuU/BGUQ7VImgY2bibU6eC
tFCxdd5ch3QZEs9J28EWj9/cmUg1SygH3GihaJWa+ZBG8x3T549oaobQPd45IaIy
bVjroHGQdMMNCo+2u+56FIugAAtlPVjWL8M0C99PIPjuLA+YdBiYn5qWhGbR11/T
L9hDnYb9o+pOGaKDsvAArl6eOvaF7bMj4MYJkJtOYXVNBhs40WPBbXSi/1Owhfkn
UyQxAG8hm5UULIRJ8Iq3dkYAaI80AemwmMZPd7yhG38aAbsYWnpqmHRtNbfEwWD0
FwiceGBeEx2TFqCMgNRVPfELcFHeYEPGsNb/dBAE+a96FlF/euMOIzOjOf38x6BC
RJTqX7oXtfN6mg3YCAJCGi4VUXgSb5I48z899PJ93ZDEz4NnqgwLcP32aepslcJ7
55LF8vDvNQM+B9AEqcB9ywufg+sEpdW3120oHRn92A/ZfmgdGjeIFcGwqVLPgRPp
KTIUy8xc58CMn8uEiyk9uKCQmI1WJlEgYFjwcn4IhkcQecKCXhCbZnk/De4i1xpJ
eM4U2KS9EpzR0zub/NO7xz6RXj1zox4C4ryC7+e+w3WBZVFZ647AiCRl1m3X4OOH
AznEkifBd6gSdCuRQwgaJVFD89UEU8nFeO+rWQ/0QMH0ICEq6vFNVlmw9Tdi/voU
NDYzMPLcZW1xero0p3LaG8T/NRIKCxHvhkvtvFMqZsAlJdFiGwm7UjwOCGhMVrli
YFxkMOacAKGXHXgrMYv/lRx4TGwPCbDyIDkF34arkyYMVtVHhMSBht5KT+St1f1d
l0ZaS91gzm3TLkq2V9+yTOp9mG00Obqcv39pQzBOGdBDMT2Nl7U1pgVeOkajf3nt
MCL6m3BfsfDWMZ6hlTOjwNryjxFFtiqWOGcALPHq518e3h+JNg5wKykYRKvzJ7JU
eMiwYLPjaeDmUkTRT7fF34A/7TounwPrVtFHkho+mPGa15nEuMBFg3FDAjnzBHDs
sp6PDCp1ZSnHxIQNAjl8QRY1u1q39j97yYawjDEza2/csTLCLRPeqB7sm9vdX6UQ
FlHN89Wz41cXIdvYfCt5Cg0ZUqSlWNilI4u8xVB6BEishl0xqoRwN6FxHHf6Hv1z
li1CqfFT6/2mgKGh9i5E34I73pQc3Pp/jJVvuWsJkxGGNfp5i/0N8XBsYUfTV9vn
vHeEpj/2ctMfoAVGvCfV4WbaadLXd/dydybp0v0xFa8XvfdAKVaiaYkkpLvZfuR9
2S0AtQfugCpQCBFT+WWyemE0yo7yodMymK82Qb24cwBaTKD9PswflW9l+pBEzVS1
kw/hEiACpWE/ElutliKU0iPC7mNE79DlK4CCUaUJLBYeceEzfd7nX4QMI93Jhzkv
xjKgwHFw8mvNKWsTnbS5skBwTYktHhiqXk1eRYgUAVj74RuBoxTIHVEwyqtVC7ys
UxQy1nzhHeX8g0zU56DqKT5/CPWgR+bzpUdRH+UiuqgHkY+/ze3v+v/UldGYWxVc
w0sqttQAAexoAsboUZwS7fhiaaj1aD0jORgsTIO3OJXkaVmduTCTCf98bvU+UTRC
JE2Pyv1YvFqR9Pd5XKZ0WwU/Uu4FtG+cdBXxZhMGu1h1aWn6TF1l9Nwnujjl7hxq
HicSTdy2awowdnRUnkm+/gReHQXNid0jBReL93Ur5OMhaDuV6AmHbhJ3ct+wNvrL
YbS94Zhw/unV3L3GxeGSlhlv6KdXWWFlVrRgoHBhfNyrvnPtgV87RKNpNGNEkHMu
XI1SywH8akFqyfWjBJBq7WI4r49ZXXYHJCrXf31b1cUBUkOBA/xFLYhtTLnf6caY
XcUCCwKYfg5yByDBX9TLGcHNdvaIYicKKexNxgHvJNNvL9wuXqX8Mb8+7RbqrV6Y
WKg40AZmbGCtbIisnxYhu30P1p2rQLcIkkncRcb/KDmHkgsVX61D7+De0+ODzFEv
R0KpOAXtznotTkQTln1pQof8vckXmqFlfNsqXMU1gdhrBnZddwgeKzCC9W+uTheg
Uj4ubEapbm382Zi9AV5f8UdnaJQS5UeMMOFUPnre3RPxNhEs1wWyf9pL/oJHEYeA
IO1kJOj0IWKlvOY5p5ztZzqOfzsTf7eSgfO14nj6I5ggWVreJBG6xNq/4301Mf8n
6XietAcQKWtcCglBPJ7LqhCMIk4Rdc/yxBEUOLNRy1dFUJWxQmnac3y3mmIlbjAD
oFkh9IWK06O0hepz3dFrfE6RFNZGh/+sEYWORpZc2va/Fx9Biy8c8vAx49OXlw59
VzJA3IH6dATyvfTgibw+aM3ZzHFPDk79zmDc864+Z3waGDZ8M6xecJCKgYnF3IWY
cB+jAkw8TPX1Lbvr8uUezxU+Fi2gUOrADNpSFK0gqQxROmYYs1gp5ouYUcwwnkEW
RkglHkeYvmS9dvVGDzY36SOD4p7nNiRQo/hJyfvhY6cbuVrFJubYnMPBlcEcuh72
Q8xctSTxks+T1dkKjZpe/8rRXZXvPWbxv2k+hSf6FA0GA/3xaKcEOn0D5MYK/k4M
F+JK/sMtHVZcJTIEdFREzwMCh/ibEcqOaBTwP10B1xafcidD++eA4CIUtAQxErIN
g+DWf+qs1wXvSbH48D1HItP8vUpaDyievz14T/hL5Es85UFizlS0AEG9tEUB5304
+mRFHCJebbFnB37f8TuCpIk2esxchxmfVjubFlxO0N6Cib+QOHoMtr0wYLq4g5QI
RJwX4Og5wj/IcAkek7Kj/5A/+90CYeNaBG4jHf3wChixVfwNP9tTx3UIMa4G5JdD
Pv/m9xcG/0l5XI1/LtZNl1jyLRx3ZyRKqp62gqoDdo1btGrqKsFYFo1YW1rjUNBm
NyN2QIDAgw3X13+7EXRhq7MOgZ/xC+Puch8wqP+VeJUiYA/B3H7bVqJh4wudT2en
9wNK7PesslWmSkF6f5iWOocXkaNXJ6cKrU8R6za3rciRQnXIvhJHt96Tyr1Vch4B
flXNS1Zu6DmsElVYjOm71+YEs6jnWcqQyNYLpQtcfSgQ3LhY4K9L4FlnYZRd8JCg
+qslcti+Ud+eotMbjAAyxqCcLIi7eMMMgQ3cgJDQpRoJuQ+fYe8ijpWz6c1TAmxP
J1FAv0sBhdNg++4E/T+BRWzkej4KRu5tHXvITYcWf2zPm+TOS2w72Ii9evuR0Dc5
3+aWtLGRe81Ldv9ivJzpYeE3VrqIfMfHVb3XH6nC93+tcfSuIvU8TIF9OEsAlmE+
uJKIRRKkUnPYR21zbV+AF2pfq77Y8qpmqjZgF0hPJOlZs6EqThk33/0R5Pan+iHq
72yn93EWKK0FVx8yN3lLUYd2ALqd5mbRDMScXvTZcbXC/icM+SXFuYNLdpnPGrmM
DLp85dphtpGesqYzNRpj6cWTDkeES9lsYdhnuipnss6u3gBNHIVrdEjLiuv5zxQh
SGNO/4VQyRm5s5Rn2zyq/OnFw87gg+Ctrl8VqW216HXBw2axPEVUili/P/bQp94U
orG7D9YHqKe+Wq6FtywwKirGQgzq5pbBky3oWdwJcFowvcpynTtSXgsIGQInojkg
lvaVkTSW5TlKY3pdPFcH3h2/pmf0EscQHpFHItqQupj3wqPfIJwHsvKJF/E/kFHp
kMCDqCX/8Awtyaz8OKRDtN3hroKVkUCxrkxEJ9jW8ns2e7OIb/URjBrRshn8B2rA
VoAGxSITn/6GxP1PrrmilXuvtrnpy2oPLyskcl3e5b0ByqdPIhcrSwmkfYSUsf6j
MLeTr5JsDprv6S+CkOH1SM3p4w0UCtK2lJhuKXp+iq2GrcCvBCm9gxbMM3YjC7Sv
8pJ2dxMK1fJeEHdql81IanT+md5uhaE0zQ1jOGYFb6VgXmINPmhgRWjw4G0keS8i
raQmqMsmaoUe6VoJc1jXodbrf8IE47hQXJDWfb6EItBWEuDL7IjV9VU79ZVFHYWt
kvO1PKb9FtXm6+enRzBzlH6LlPpurX6qB96jl62OU8mvfqhf2IsixKer8hc0aF8Y
1aEfy8S/46zG8F3thQ8pSVlQffi/04rjDyrrQPiDJgLMOFOcAOfJJCyauP0LOLS8
KwsqvhtB/LPcrA1KDJxY0VYdsKOBWu2xJerNsMANsGKN/ncmdSYQ/bhYC1cDaL0t
JWTPzfMfoimPWRTuyb1JV7xQs2KKDYPy5ZboV1cbgXdAXWCIvmM13f2U5ikTvtYX
P1ijrzSnIJYlUba18smWsf0coazTv0I7vw8tFjkhADpiYqdNBZ8fD+dr+WIK7Ejf
c2rBOF+eTWkPEn1plo7JpZbulFucgFScavMrc1TtvAMFbz+GPviZz7uxy35OVWw8
/uFi81YGTiJipOlPNUx/CIQw1zAwIVK6s45tqAgUQlYf//+ITG4bo5JX7j1n7+Bu
fs7r5gW2DDTOt7H9158j5J68rlKE5V9G8osPSJZ4K9DHSZmKc+U2mjPHRKDpqzfZ
A6onig89SkyVzLUmGtrFDsHQYQIK/7zOO6/Vr0/IVNvzvKWFWVzyyBebVlGbHNHG
rQN3LfYsqWeIxOlum27duHidUMXu7pRzva+Zwy30ESq18NcUbqaOwizMoNFpYngN
GEHxqR0JOsf7B9j8u68Kb955OwlDuQrLUGV4hXhIO2yTSLhk0S+/tdGYh/+1FS1z
FJNcIO8RStNI1lSbb08s1SK2dvWptWupjoQJAB4N6nop8OPXRQOmSB6z6CNKZ2BS
ZPruObthdAoe0hM/0Lpy+jVJsJykpII6fmKTXufuNfzwqgSfc0oeM8SmYmVx17Vi
A7z+K1IDKtM5Jaz54DNPQ+Pp/dfy6M6d2Ujk+ZEp9fSznVY9GWLwwC3EUH/zAve3
z5bDzjOu3G3Clruh2hDl6MPNTs/RvPfhAgolHFzGy6eX9yEEWhxBnSQeat1VGe/1
GdJALfYjvZAdvTHEckl+wlog/6IpqZlAU6AdL8l/s+AB75HHNOV2HD/j3g6SEe1I
Kz5hlpSTJCAm6qOPWIBDjsA+FKHdnNatsZz0DR9LV5QU2HC9tZIHb/Fe4eUtoTzu
XeEHUtr47KIcjCZaeiUUPsvGQXxiiC60STN+3PNu24oyAIwBl5q0uICN1C4h5n10
5ZHys4nt4h7mMFUJKVPdjXBV0JGOA24tbvlDEgklSd0/IL/sr+KtnFheVLbiDf7z
W3MXIiyclRzBtJ2fZ3w/KBqyNEdyqjVwVAkt98rZJ+0X8A/XtMrw4soFwcWDP/3a
iTBb51QASMAdwvb9HUMlMwTNXqF/MgMxtX8dI0qSh+p30FE/RF6ab/FSFijraSer
D0LdVhdg48itPGZ8sHRok6NPGb4GLHxuinN6pYuX9/jLE5zDUfu56ptdl9uZ7JPm
tJwVQ4v+WQtSTA5nVkK7QwRKqYIdQgA4LdG5XheqITDuxHw+K3cxZW12z4PA4ECF
sz4OMzaDsCqqXFNJFCwS01XeUCg3DQlmnOc6ibky1Mzt6lJmGxIVZ/uel/DtVl+1
cSxqcLPQ/8PlhtskKiehMwDNQ7CL20TxCdhty26ASXO44nWHLnpZy+mm88NWSV1D
rSItKNTspueCSIbM4+TPgZYj0FNMFIffV+F885q4zlO1pAmJ/tE5YQcHfLpXgQOY
o3jQzxnMfe9Fnz0XDxeV6EiGGaS53ZmKcDLxR48rUIhKSs3HTHWE+5ZtlPQOGR4l
G9YikTcNR4MCZ+h7Jcfw42DOs3C/v7xVecvVy5F2XVetCYmVEhio6EMFUQJkqbgn
ABazV1HH8yfqSHbchEDHhP9nFd03hdTnvCZQv3b2jMq8PBTiiJGp1nqsNsnN0qLY
pEvQfV8KrUSN/M0GKWVyoiZlDwKfTRNeVGeObxg4282fhdlW3QBUjXr5YIijKTDc
HhoDxRHSmMW4subC6iy8uKoZQ8TP7Ei9VYvCW/zRm2YC2P4Mc/WyUOyzPmnwyfLh
LpFz37MeolEbwO9ZNahj4VW1lRosKru2EQQSst8h0quRQkSW+LZXYBSxgJtAyG4H
ELezFkSNr5wKgjdL5v8uEAqUCoTP9nWNUgzV/qJHZmb+f1PWG2bgpt4VQ209Dmdq
EbwCJW3hk5o6+G3QgjznvFMtinDHdK+BMRjA6ZdatGluwhu3ySJLnG9GJ4lCJT7t
4GZv8jQbb/a+C8jhfNM8c4P2lQlAcQK5sewah8LJUZUqG1u80SjRGA3iLUhlJjK+
er9GOvQnOqIxZF8K+enpZ4eAOCQjciRCImVHquhf5PqSFyFq928gYJLXlMedZFeK
1OcB6Zp9fMT3dsLSn+7Bw63XQsBrtp3Atub/i3oLQBDUfU4Vf42qO2BtXjpEK6n8
SrMfJ7O1EBviW6PJy0nW0W4wm+spNSzrrb2FFpXYpOTWgYxXyXE4er0SsBZtnEzZ
1kE21iAWhF0oqh5HcyGQ6RWcTkJ8MRyvSBpoTuKDbbLEb1KBQwk44SqxVp2wg9zQ
ViFs7plAc/U4ot8IfUIZbWB47IkWHjLL1+yyJ7Ru7RdZ1gTQ0wu7q8dLWvBBnwRK
aHqz0HZ83NHFn/GtJGtc+75FOpfpCbOzwCKmA6ijNQ+BwSbKFM5ARhNRnM+5H5Yu
KicmAcdTqhY3DrY2HNGdhPvmsQjsf9LjwLiYSHHX+CavQEgWjpxCuFC9hKGDs5SQ
ia+Mf2OxqpznzW23TrBpFr0JkK6lNOkKWCy6qIJop3yKsE4VFafJnA/oM+hwiQhH
nBiQf7FPN82gL3kGCoNi27nJgTrukJSlDtqLjpxd5UjSMf8zcmORgNcoNLPvVim+
BCTHhy587a1gVFGcdqzOlIQkb7X5Os8HEh4rcOxqMRFrPWa7Vj2uJVL8anKdcT9x
yiFs4CnIvj5fRVxy21h8cbBOrCVAcTh2OcBPc4NKYZWQ8vBlWugGokvwN3L73BGF
Y0U8X9rT8LQ37pljfo6UjIphJOgMStFYrJaiTzwzcmdKJgdQ6y/QwLOy+1gbspdI
TtSFBA801Sd6snLrXaMn9OaBK8t7JzmrXPStCl8jsfmRQx79OclMGQsVDC7z0FPm
QNA/1EvT2Yxmxzi2BLaFDd8idbLYyW/ErxLbcKA0BT77rTBwbjno3w66JKD2nD5m
nk32BSEiwiJ1RLFmmgQYDxXuUTPVwIrlx0X58XQW+CvWNhuqb5T75LdENy6PeGpA
5jCvf9b6c1iymKAr10kuthr5d9GwqZHEQQQ22d6GdTHuwEXpmw61ge6ryP2tNJhc
c/Vb4U7wVr3XZeI6Yg+B3jITag06dckUo9wDypZmQU8ycKFvCMidE5qqNUMyTO4j
okBsbXyfQPJ6jLZSfVLDDEOnAoPx6hoO8og4bHaWQv2JOmkCnrq2ghSBoJ+MaG7C
yUFDDVFdgPcWJB9QoyOzDEKyOUes1Ov+uKp0/3hpJ4s7CVcgg+Wkf7+MqjlN7Tl3
JuSuU3b9/nTydfhUxNmyyM2jvevdbsiTpC/3A4CPzONTvsAH7I/R4xybW96hEebn
5D0CzLuqBP2W0FYvgcaj8Sw8dVFKQC4VjEZZZj62D7tUKZ6tH7/jRTzuxuDmuUAa
j/PANr1MBdLnpBB3twe+r5VZrH9lR7Bu2BSGv9T24UhckSEneAqwvhNaR0E0ai2f
3+glGCi+E2Zv247fa3B6+tpdiKHP+G5XTGS+g3ukQ+R800VM01efaHbPszXpcQj7
rooc4mL+GBS/Smdhp3hRKw5kqlz9VdMhlNWXFbicj5Ouh2lwOMf4yC5sBq+LCcr3
sf4Gpt3PQnFg7HW2W1HiEq99v9MokSDkmQIWRdO/+NqJ5Ytx2IU6wsUc/SaCJ5bI
ds1vDBaqrUk5V/9iBjmsvfku6hkeC5dhxM+VHoJuODUXeq+MQG+WxHNoXRGHuEiP
/YF5BNjZI1ZUc0BQb7WR4H43ygu2ltqxJ48x8piTRuM3qJ5ejNgG5BdseP/c90s3
WvB9UugIwyQ7cwhWtP1grfmHLqWgIUmvkUdQWcq9+rirE9b0T7J+WdJnufs2hOh2
fFAHn+5X2bs8I7LSwRvRu6G4v3JdDsmdqAEVqE1mKeJOfHogYtoZaPOENokg8NzK
62wKis1KNW5LFzRLbrmBwEP8bWyVq+mqQcK8172lzzEVa2j/+RzOD2s3DKO8S8s1
b9jdXM4RURjzmXr3W1jiMNsGUw7kVDmF5h2qkKDTJ6rXbfKLPvIs2cfP4ZbWE5ff
gwcXTlTjFRngpMbGG6djtiEg1nvjztRP+zQnStAgYa8X2RE8XJHobYD9eCCVeCLK
5zZnVEZO8dY33RBrFsYELP5lDqCj28FgDMTvuuddYg9a0p+ue1/NjTYRL7Bjtddf
iW6Gn0OCeqv5iBpcgjy2aOhwzW+BbhQ7xHZihnpcG5iMsdb/AHGeVohJo4EwyQEX
LfPivXLz0Jb3cnatXmbrNq6f0ArHvcI2HfE9k9L/xAdLHaSkWiDSByUMy4khHjzj
pmJVFwvUfwzeadwITTg+DC2YMi+ygS5WR5eMetnoGpAlMykvZb89uu6Z9H4wQkIR
wCdpxbfL3ilnnX57F2aDsTvZYF+AdtrDKUr9Mrm6c4bCqDJGqnNcKreRxXsvgvNI
e5sGO4nqrN2qv6+NqyEyk07zU87gDPlaMPPXe7yXF163po2vmnvj90/T5EzYZWGs
/db2LQ23u4WtqvbIhS5wPjmnhh5f1eHAaLp2fcw4MUPpXCMwGNU4z6GqwLUgKMEw
Lvf+5WWCe+He3Dg0ENlLwb7tyoVEVh1BWy3vT6Ybsw8IDZ5yteSHn3QE+e+o8LYd
IFnBPyzGAE1iZOEYdbbYTn+gNUKb6nOpRKbCxdv89EMBqz5+Cxa7DMnBqa9gvOJz
Mh0G/p2jZmy4QVhGzWIj9OS9P8Ga0S2orAcw1z/HEdZS19Irq2ulw/ixliAFW9RU
pAkar1cCnzkyZ3iUQJUVbYp211UgXRHlj33ScPSGU2dylvHPfEaDuZPjlaNiSbUd
r0UoS4g6cFrskketyE95EK7M9/NoYJD9PGAI7HkddSXRilzyWhBY8emug/DS25eP
SBlIzJ2w6815PFZv+RHWe0yYYrYaKQaUrnQ0xJtCJPkBPlWwnKGjwnFV5I0hVeu4
cItuiHGYFu4k3iT6NMfxsFfA6kwfs593Pr8thwAxGcPqMuOwWtkaGMOUlrRY0+cl
j227krm2tLiPSv4ja8EBC3Gh+qhhAXXmBHtQaIdZPgG8flcHzIG248GWDvmQmaPT
eYeNMJ0uWLlVuU7clpnpsK2Z2Fq8co8rqWU1j68UFSJYgfV0arT07KXXWPXR/RrB
7PZv2+FYKIGbU/YhcylZg0NJQLRKtZL9TwszJVG5xPafRZ1moFunfSJgnQRaxaC7
TWfWNVkGE5fw4JvA3xF5uC6A9DYciU5CpJ8n6F/hPiSpFTT5pgHYKKMsPtgBKtqv
cI7sfzNQMukkA9otq7rew63rrbvBlqQzVc2TrOB7G/bqfpO23PhMRk1vC6BILzsz
BCrrVP503DQL6fPtziL5omFp5kumtTVPqbHef7Ake6T5WH7O4Qp60HCrJepWo4bz
wcmtQr3pHZ2+dZhQw0c3DEGIkRNca0w6v2oUwhoRdkqcEPLSVvjxBJWH6UDj3U+W
LqaznUU8W48Lxz1N3ShhCt3xymPumupjOdLAUuHvUyhkKauvAY9vCS6poa7BkuZR
w8+W/GG0JYTX/vqWLNAXD9PxTGBg0k8NoLFwXJGs7E2v/9WTLm6c/KpkjDFa9hMS
y2eWZ5hXhtnW3RPxLMZ9xqdCCf7Amx/qUqt9U0clU6wG07q12GLAVZ58WgHmORzv
/C+p1WEJvI5mVkr08tFxhXuxK8nxoChmlSTmulKXj58bnFZZ/OpRHEVlkUsdpPIq
/ZxiwRaxv+Pl7WhZ4bPx/mix+/0UwuSMef1iy/4XIIf7rbrp3km6ivERNYnydWBE
cEsLOrO1CIIK86SPMzcKPbCyj+tuoeErVPs6xup08KdlmmtNhTZCDC1wnNZNTgn/
wzqbDj4UadDFiijyjf1QNoeRk25hUtv/mAK9d/WJtjNYKjDMLPSEV5MIzKrmauYp
P8epNowIq1oihOU5JlyZfejgH0S4x5frFA98P7oT60LbvvqAVOk+3H4zNJx5W0QI
t/fS1Ijuy038agPFnOz9hSJH/6Q6TTqvt+bXZTVOH5M/o3tFfnP1xJI1xsTUdmpX
05RncWsD+90jYg4YBKycBEYob0pRxpRIxa9j0dxYqJLg7BE0eTSRDW7VY0bSMYPv
T1J3ti/pg6Th8NCA5+UdE+Q8J+mTZpx0ALsp2RLWemHLYBFU8zYd6lDUIsYTwhme
FYPS/IIvIJ1YfQhJ25ltB+qTOmEnSm2WlVDXfzdSDtgcFm/7QC9nm0EyST727qIq
dl9FUbojIgNEJi8i0H/lIaz2PImP1p/CasAs13xa98IXkYeJeDfw9ap06zR70/ik
t7ZXzr5SHVKU/Ejwijs6ilF1cAF6A8CxDOsgWyI/93oKcRRwQ5aJLX+TKDz0IEBd
XnwAi9NAq4cv5glV0yh4W4j1A5cvfEcMKWWgsfi3qnLcEZfyviW9lz2jl8vb3psl
4Yo7PZAhY7+cDAmsILy0uO8246VbM7M9UZBiWobuM/iA32vnrmLvTO1+yFncS046
MuvTYpkFEuclu/a7T6ihTu89tg9D3/8wRzY0Zzq4e+MjJS27TpKBpLJpybMTT/Ti
+UhzaYu0nPOjJyqrBC7kFxObobOoU20c+WAhscYNLghUPozcZqyJLgMRj6p3Tic1
ft71/xxIygKj5JpxQx2ff7THLn1D+9AzprL+FFidd6+b2Ow1vW5+RvzZb6NZWAoR
r9iZ/+QJhWhijhY65vF74unl5zhcLVq5li77WLyJzNAr2WsKLDUzHkJb/ZQtXz/l
5gJbmP2+Hve57nG1a73u03dah0vuutCTD0DS4EGS55oQIgCQCBXsuMOISofKcdGm
9HgwAGWzoUVO5iDHa9w8Ua6l4WzemMOmynU4Znoktc4aOH97tx02+IkX0rceCsSM
fPLJVEbgfaYUdtjH+HhcmxzJtKDu0vtA7xDSYdh8SyMmDreAt37oNz4e1Dk8a+vl
4esw04LwzWAzPz5dduy/PGAWzP93YPbdAe/nlrNqIRmJZHsjPWp4kQp/pf7ndNf/
VmmY2nZwWPSi1vQmi295KdMvYE9fgldy9Yj6LYZvGKofRg28fvYmteL2WHafLk4A
Bgf975oA8oNGHS/TYU+SNyTRvtsBP3ZfCtfIqj9OP1yaWaM90hsfz3Bc8gd6WBEp
ZP1S+3gnSPFBQAJFNAgGT1ZfS+WrUByWTJkN7AjZJJfjoLSrnH0O5LcqIlWr1PhL
xrizWsjw5f4A/3qB7refGgme0WMjuS3jo7JxoMiZjDjD9lFs2/guqQYr28ij/bP5
ECBud56dmWjrjS016bsuVpNjJBSfvx38zU071lnOw/47g76oklBygDCQxpMMnxic
S0YDAdAJzzfGFmCCK445eH1okRCy8+DCalg+vmX8qpyFjQ3l2MOh8Iou5+AI2js/
XZwfbAkJFkOufIdbe5q12p5XX7l3+ChblsueXta3LotM+/Di+fAIzsduVJZo7ZiU
lG4wwDRN0fqHlysNMksHbgziiCQPDOT9LCs8kc/LXNn1kc2OGXKKx8Jo5PxhWtNw
FD6XnO3dqU1r1+v9BDEV1e6TyZyE06qbKJTdkNFAGMMZcKAlYWFA7dlSzIpXy1A0
snDM0dEavQYyqzJWXzxg6cGLgjSM69Gw8x0DCQs7sJs0AWBLIPMFqGol/6faQ72+
p+u7YMQgkZTiXn+K21vIADls3PgZlY4JwEOrWRYCIELUdwc5QOGXK3cdWWQq6C1Z
WbWoKKUNLhJWYyH7JIXCG+TRHnkQLxBcWT6CdpCEMQ5sZV/5PMfPc+NUTM7knsPr
2FigZshQttIsGNHImjLmSAH1uUuCwQYwKiUcczsKDDKlcAIG2Z6N+2eaI9VMH7Hn
pf8o7RzGuD5IlHJwd9OMoD5PP9Sb94hvBP7euKKM/xOVZEskyD3OCFSKiPbA3oJI
TX449S22d9cQyiUSdP9kjygR1nEO44QKPkK9uAQc1tndDaWsdOv/lE+ILk1U0Lmn
CuRadQzeoVPWSBnic3l/mEI9p6EavNpVYXoAwmamlsmvG4QWC79MjKp+8gCfUNG6
F7YseXP/03CdzGdW/VYqpT8RTtycOa46ZFIXNYQbcifeckyuRDoMyjdZ20N8/C+5
UtNg0mHt1j3mC/G/whUB7Hjw+NCvbG0/of3AwlfCdyn4aZtbPjiUC+bEH3ATlqAx
7c9glUYWPbuLhItgSHRVvgp8OGIRsnobpSxYik2UbEHycVaaFbQZEiZIPh9hvHH4
7Qar5FJI4GUTSduEP8/Da2HaIHJoADYRK8gvVitczFE5f6XEXIP3TkL+4L03/gw3
5tjhL4IRgvkbIh1paSs7KWXYBS3ZFoahGB9PJlOyd6CSeh8w8boXb4ZlHGNeibgw
qPNxBstVOpkgeKHbq5zp5OZ0ydHEFMg8PWyQ8WaZXbi/6Z7583BL1OiyqXOAOr4S
YFEnaeXVX1E+zIVCkmchpAxabeebvqbG0oyI973gCE2EbThDYFw2gH66ESRmteXR
kss3PLwmbqff7Lyoj+fKIji3gfiC+xZx9AsmxKiEcMZcmiV7dMeoV92p03w03UMt
xJNg8xixm5xOYTFLv6xF2DWnzpKOHKcYawEWRg5dB9NdT5VmL+x/TRpQDk0KQdG0
ea7b7eff0kSiYBMWdnZ93U14uMkKnwWojadD4shwi6VaTfVp3tFDK/bm0sCqZOWL
jysDjJYbnPEuEpZCNiLBSS2u4FQ1c+XmETChWdsb6xfk1sMHFJ8DPSRQnP857NEz
V1Vh9QtRGoY+ArEX2lxPiCWDyPZsb6P2cCmh2Iu/qbR3+KICUM7KC7eJrNrNDKXE
h/hG7YNdUh29DsBXv+BXdoA0RGuUGWEMiR/JA60ut4JxSz3jIYHaalWrBTQrwX+I
PDrDQnK7JkfsiCdyD0lcUmqE4Gr+gNOITwJp/10cstCJx75LSQWhiPNZaha6qVgJ
DKdMZ/Fo5TKKMzFkK8CGpzc+kQb4oOa4q9LRk7Q0/CWLExHczyZHwozy9mHkxS6k
GlIek7cGV+hgzsBH0Lsrkcv9R9JqkuAEl693S8Eg4Qi4JAJjYlvjYVfP1XQXyeDY
UHUGl5T9d4nbj4xqlR7zqHPSjoXXECN1y2ca5dt6904Sg/kW4z8FjUH+WCjssFq/
QYjXcGLujBrw2Dh7vdzLBwLWApjNw/XSIR3MeH6mOoOGrNKC6cNB37rwg1VwV8wR
oISLbmELkU2PfelQTCJ4zCrZgBm9WFvQ+In6o1XE9IvPgSi3cDniule3jKPrBa34
0Quw1F1jBoDk51lnpcWHqwdvCfeI1QI/g6IgZ09+pb7KxhL53qrh1RMyn0l4qrAl
Mw/ir+ziqZeAnJ92PYPZU6l9VOYNKuFBHHpdSvH9OILG6frxtbWsuwv/4bOkm7Hr
KooC9FnYoVfR1TBr9S21Oqx6syzQhjw5856YV7fJO1CMjm6LRbznIwscBiIpJar5
7wA3rJpYAJ0wQLgTe2LY4+VNV6NQa9wlQlromF9JKRwobj8XwqzPVA9v5WZWXGOX
rY0yYBoko4zgVaYJuuCxr5f85/N+naNIFdpmOQlXn22i8jaZaXgDyvAnsdF0dATV
xyX4wjMLOqymFxKgn6JsvgqWKtyDWHKUYPxJSn/ZDJFbSst4XWG1ZNKkwkOI94Ha
Wzi/PdqmqSeXeizZlYxldQ/Q7sSfpk//12szaAq0MKFrrDiiE27vc2y65XgesvdF
riBRYNwBvfpzfFASP+s1+hIGsAx5Vj6z819srJj+qv110Fetgj6LZ9jh/SlNxs1w
7kfxYP66m3WYIy073j4BsoZoSuL2UwCJL3sSlx3A0i5dqu7D7GZeLonn68uiZTM8
kvzX+41OcKcjWsNfqUsT2saA64LpKcZuGirrZjn+A90e8P0C6isVFr9F5LgSxkrO
YTDc1YKOkK1hEB9ZrsGY/IuFWYyQijMSh/cw/ciaTF/VWde1sWRheE/ouuF+yP9/
WziYbk78wvHAY+VH4ANZHq6dNHmtxBNxCo7Ve0N2msvHlGPhdCD7QjpeOdUQvfdn
NF3mYwoLWxbWZIMNyOz+uHf5MuEVCFcMRyJ3Me9usB30dgJavu1+k9ss0Wn8skBF
aJaCj8F6cIHPaiOy4yYsQ+0GyoXiryYoKuPUMxMI5IIOMOwrIjXIbB4JuDaxgVmZ
o4hvI90QsneGhswzs2Cd3Aa6tG8GdDOkXEjTaO4t64UFbRq65EGORmRF8x6VjY23
F1JEIpHhjdpj7pe4PIA8pOLoGpZxj92+8FEYCL0l97pmXJMlmOcBbVnS7xilA1RV
wYNKWR77a7zXy36hTnXGWV9QAE46GrWlVPZqBgYChsjxE28qXa23lJSPkDJARDBl
36/MkxxuY/qH9+InkAkvr3FY87YWQ56NEUoh9dL24X23Ql5P24Iu9xLLtq38CCRx
lEgvJxqou9WlEKGqHjWUTgHIBuWHkkmOicIsKZybrlCcArV5DubBJmx4YsgRwCyv
0oPeXCf0hhYOtjtnezv2qAxBK1KzsQyejU/BFdH3Ub58CkPDaq6cHDPoBgkdo0sV
KevGeV9xJKvNggLUaob37qXxDRy1mz3FzaOVJoKB+vz7Sp74ggKkba1ZjWVBxvqL
NRxCI3GVN3lwS3ZI3fIe6LBF8KI26brbuRaSXiOvzz7r5f6eBHN/ivDCAJ3tHVeb
zA6VDV6u348JZLEe5Zo+dsSmJOw4rUATkTlT8OtO0jIWXCTYPHYMBPrclntqGW8a
9EQzgdJ6oNIoRzUuuuuBrdMEHa2V3J5Sz6RSk5Dqzl3qss/PXqMIhmvCVqlTkk/z
pJlHMAD7cXspMcRZhPLuSU4V1W6uE1VuuKsJyfjnlkM4izbTV2DdBngJLmLu6Cc6
IZVzfy6H6E0JhE6I/HWIB7u7tpP9ngmn+sv2FJB7//tjG45O1/8bS1aC2ouVi8Za
MuwZlqoSoDS+8Vwr31McMu7YkZyxVZ4r0HABrTsx9Xz3UD0/pReL54Ns9rvqOqXF
csWtux5vjNKJEl2vg7r3DXlCOXCCCucmldafKOASrXD+FrVu/TOkAx9AeDki3Eo4
I4yhzFiY2MKRyb9pBX9kLCq97Fh1BwlEtSJdJmrQGena2h8RDPbodVD5JVFdxUHJ
zgGKsCC8ETBJptrjFVKeBNBtrMQaRcbtYPV2bnLWNTsVfgsR/mscIkgmFerFBYkg
tlywv54NkjN/jDyxk8BFdh/owv3IwAICUrTFVCrJtqfNcs0ugRDgJSI/yBD0RFh2
28cWWoDRbc5owaUSMVFgnC0Y+85dQ3sFDpiNdd/M6LdXLhDUyWYyb6z0EodR5pln
cm5ZobjMBW8rf8lt4l1jD0vqS8M8uov/Htp5g9DnX5DH+S2GqAsqpAqGqwP9ELN0
nW+ugteW32NijIpFQA7BxQ==
`pragma protect end_protected
