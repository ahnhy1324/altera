// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ILuAxjxmp8PP2st3pGSl6epFliV/7be7EWZ5vZnfqCy0bQrKIjKZSr2Dl0Hbao1J
4byqiKdBWQceeddbG7aY6bg+zvfJH+NY0mP4IcYbv3HfmalyGpuOa4Lw4nMfI++4
IymLAzHFSuB3DDken7eiHryy/UiGcOPYitpSXXDZwXM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 62272)
0Zh2EMZJAvHIgwwsZ9h9mujOImR+dgA34SM9qAaiaRI/3vNJaqX5v7QMniOygpGy
CyJZpOi3Xl27FiRdjVx/1Y+sp4A7Kz7MlTdX7qFFXyl1QeEClYl20EMS3hq5d8Y0
U0NsW9SrCGRuisohp+8h8Zz7LjOTmpTO5Xie+Ki/709O5ZRolYFM1DnlS4cfgM9K
lFEdEgWWjhNAYRO9qHFx9ST9+AuQbRU8e2+0H+BMWWYRyicPPc9lOWpd+1EueVC+
lQ8EiYpM2G4X4cKyr+fBO57MXfpSFqkhsegiCFcUXra/wkj5HvnB5djWT5GOHy9l
z0O70DIHupwv9p3rVpEEWm42XPHEacgUqGTscGTwmPygOm5pvPJz640Fdfhakqe4
TnvGJYeLcS+rFcuvG0Djvn3tZQUbSdA98dB0D37bhC2R9tNdZgY7K9u9d7NivLko
W1r5S5c61/Piho3XBmvexgjlxX/XwHfWHWKKeJemSLSwlNH8x/cLp7E+WWm+UVgM
tNzliu6f/qaW1Tcg0QUAgy2YI8M/NJAyTYXkmAT4UIQSCnID27WanpmUr4X6jF5A
CWyXFjaYCG3ysPmUJJpoxdaxhkXn5hooza2qqWhTNZclNKlTln2H6ndG0wIMxcSy
Vvxf9IW87F/UJzGkwV7Opojf4BgiVOVtLEMhX4jD9GWBg1gVCq+Edtvt7+i9Ffdj
T20uQa7Dzdlaz+e7ohKIyr+MI7i1xFDpDwdx0LbgYA7Rd6xNKazcGmtPZBDx76u4
VVDwVpNNFyfAhnOd7f8/ymCisosbguMJEGbmGPXTFKGRQ7tv9MxyXYsXmvUGU7kH
4QxmFdohOv1Hg7MFYQ40xq0GaD3nZp5LZWQsEEnhiC9olnaVEqMN8f4N7rFegssG
FpceDhThZdLKkmOpqWyAv3poWM9VMFfdc7d91LagSPKYe3qufc2MtFrYSrmSug0L
K/I1fUjhwEU+hQ4Ld8JH90jSU5qYs1NNaQgXYE8ZEYQJWT3sxfB0GjdNk5itFjly
ybTBkHw0e+NghWfoGZvlbqk6dhmI3in2oj4eauq2FsQTf4ZY9WMRuQGjcvpeVwkr
8BoRIpKF3Py21rTYcFpgRSZpMMxBOvuEianeqC+NcNcfxw11XM/9kXghUhOoBxjM
pUnOt7TkrrjaeeG9n4aBWB1m1C+YfW/htUHCssKhKRrgvWpUqH1jBvYXUmfpypAk
IH0AB3dJk25L7EgyqqjujeyuaOFvux5qcBFCbZevES4ZHkbjZ/8kWBIJsu6uMq6d
JOpVQF10GiJIpQGPsg26LKxK6FIdqO6KL5VWhpisH8cf7M518gA0osINMMrZ52JQ
uCt23q+LkIOtW5KiS27zTV+PM/OBSqzoDny/9DwKbfuYpQiU3VuHMFmbBpr6Fu6s
XvuIC6ZhhtuEe/hKoXXLYTQ0QQ6VofoarDBU+ZNYWBiU3ZdU8CMiXVuHn6A6kRct
+kcj0RG7+nk/QjvjVZsuMOD6G+Q85V7LVxfWVZYAoeoQ6dIh24NBeYNziBN+zRzW
0mic0y6VhFn/j7S6dpYziU8pMJlRkVb4BsSDl4kjqz6nLXZZeyjOJ0r9mD3Nk0JB
1u+Y6oBLWlmQB+ngxCwbzXSNNXjAILDJL3rNTqDg75314vCXSqgr79xMzAIa7l0U
p3t15esVh04WC7iPaPyfgfTQmx2QK8gJqb2PzTg5aUgEMAdU9cesZnoX4VKv0oqI
LQveNluFH7SjnY4xjAO6UI7NRm4181n9CeWLxiDCl0u/WGzbnJrvkW8Jq210UceW
/5sL6t10rYpQPRFImGUmPeLqokmTCliKGUaT+qq27nMPXF/bLRSwwvWBI3CB8E6d
IlCik4IkPvupLbHklOHf/dXE2hf8UjCkyrj6ZAuf0Us0lVw5DQ6d+88nipTh6HKY
kVzUFlPNdB1IZMqGv0CIkrDfJ+3d08Gg1ewJGuYMZQVNnhRaA7XOaUEhCJmQlFMi
oWqAGeINYobR2jeKDjsPGk5ICxuYFwMKfmIKAzSNpQ8UrevH7VuNYYCxFwBlthPi
OVggVYIXiS4yVhOjAixhcjtvE+84P9N1KyPUr7CgKFJuGeRzUTOyGPOqmJX4EaR0
Gb6yZV3NABmicO6yVe8l9FTbVjEqLNRWxpd03LM7se2rgQ73S/vX9eVFYNCQW98B
8mmoCZguIV4Kw2+CqRHuCxQZoFM8YY2qITHHVXFb0cjI2cJL462XFFTRYuFSvFfO
/V9sPDf3vyvU1BEmgg9vyS3TcdIfdbbymDXTYJoyGjatWTP5xpc9Oc/wXqFgbj0W
R6tYL/p9V4+t9LOQz2WAsrHRAm2drgTRM+yqbWKrVrKFKV0xxW1aerz+5j8RapY1
35bYFDy7d5wSifnQAqV2q/PAvmfToBKPM8R4aH5Lg67Ky9wWxat23/MzBeLcnIS7
tQSIYBUb9bWUGUV5vjdAqKKwjcmFPd3IVXc+8iaAETqcvzCLbLxInf97Jgii664w
6NC4ZyKcueWcyUfaHM2m0IXehl2eq16oIwBqbwBp9XXyvSgstz3c3GB88mkjwHfY
NWmSursTz5Erx1tywmzQ66+vn6fmCxQONWxipB3m9DjFd5Xc3STvBC687i7g2wnE
vkkxSoLXsVjpotwoLH4ZFwtr6O3FNSncA0B15fXJHmKy/H895Fr7niQg5QxhjwUi
r+ev8PxvNwsH4z9uUdG9fBb42RcsyIujEAlubJFUzafJ6diMBp8i7XT3Bi4BEPV5
HMoYwUIeQiD0c4Z9ERa2lv3UVZcYjkq+L6jED0HDov7EpoOkEKaUME7l2436KV26
BdpnPZhitrcbo+m9GBCj8Qd7tI00VSdzBZF35kEefHZ0wp5i/cjGkkEMiIB0zd0U
W1kdQDTiXsFysE9Hyl9SwB3K6Wu6SFk/BXpry/evR9CqAX0JxA5Sypg7ooe15eyl
mo4ChJRqcB38SzeOkLXSkR0juzBoO0GBs7RekrLsG/7TcOS7oZacW8Bdy4NTwTsY
XKTmcNWvDcmpW16/SczLmkuNdRs5rQ9YocSxOc2788jQ6RVU4RNOkihhJv1MM6x8
hGkRAFbONx7LQE8Zq2SrdKboYHr2CYnxG5gRjyCGApnJQ2On3Gzhlzo3V6+ULXaZ
eIeVoKffUefE7a///OT3noK79wIHxEpfdsQ9fFrNrmtHrNMjd4cJ2XAoa4I3bhdl
w7HbeJF93pEIuD/3U9mzw+wVzVkQH80lmTOP3TyALnNhBheRYBms7hpv6SWZvDqa
esMjdQ/oVMOeTsUg9xStcoccd0UhlYYhhpmMYJRVftzfwqQWvYlRWw7ByEY+Hqjk
hsjg7M6Lr5UloTKdGnn+m0Kf6dhdhvgB1S6EQVw3kZANT3owTmZ0bqRPZ25OyVeg
Tpr0COKP1OYuJw8Yn6sDXxmp+qyqPc7CG2weW2P0Xi2rxBSLg+GmafxJuZc5giu8
WUb75EumZsmBb6LuoY2TnRTopINt1e3WpT7T4YmsGwV/QoICBfndmCyJ/AJOXFfv
aW8AKV5VWXccrtsEDgjxS21OiSyj3nxUDU6rU4CSnTq/QBD18SpWwDph2y8DvdF+
BQAEdY49WH99wQTwPmNmT16PZsTO4i4tuPfvUmu5fdbZ8xrOcwiKftWCBghfOey+
oDFRzF95OGwKkaNcK97sSf4aTFT7OwCFFPSQZ6mXVr555sbEiBNPdlZE6rD4zBRx
5jsOq8hV/s5PRO4BVRw9wFB8+y1+yNGDLc+Qjb9IQ5GdV5HbyGRxZ25G1gPHS/WH
WnH05o/IN0Nfb5EUXMy8AHWa4V1ylhFe7fO0K2EjXCp5KbBICOZaFUJYo/HfHhGI
pA21xEP5bFgcgBIUGZiLydr2Vj7cNwhORbFGc1kR2ISL22/CqFmORYtgQ84PNBzX
Nn4K37Dh3VpEdtR5IUDoQLDluiH08+X4Pp241h4qRBX1jKwi9QnqwIByetp2zHUr
KqICk8DotIUFYXVPFzRSos/gTM+16jwbfEqZ1y/rQODpFdrsQADQ6k55IKEY8yl0
mGHmsSFu5rd4oomPIZ0kb9IbWvn1NFpJhgSh+uwtjqWQp0vTYKyFHaXCSd6t4LFq
2DaBm7bwYdzQkgkPP+0y5xEs2VcDKgXyjRIoBmHcA4ZUMmkitmF+kdHBgoD8lwGZ
kEaDk4kBVwttqgzpvrLwacXeilJ4Wxj7M5ivWRWJAlJ/63HjzmhhdLlvm+oT3A+M
weWpTCvp06h6QpmQddR45J1NdyqWB4S2iNuKfxisISEhxGOXlYeVYuT3jW/z5bu9
oLeE/eeeqfTypmPwlXH5k2H6redDtQ6afEA5T7CegW8xHpp/isJxTcapmtPnXLH0
9nLXAb312q13s6u6tPK5GzwjKRrmaMvZgnMRc12ZeZ+O64FCd3e1QL40J5Du0aXR
cZkKfcGtoY5u39rjGe/VPN0a3N28kU9TBhYQxPgOI81EHmVUYrXWQqlTp+yddoa7
ywD1vywm0gLWNMErI1sXoBEQ9XLuy2r9QN4N0ksLSPT18lrYMNaUGG5mjgAzT5Mk
kzLV83v7xpMTroLTDYyLDT5Sl6gsgCtI3PtyseOBblEH/WwaCSGVB7hoai/qdH85
osgVduZvzq3OSd5cHUZFqMN8TNO7vSUzG6FpB/3wAe0eEp3KzDHPgsml7gpclGE3
P+oJ6qlu0Ycu1MhJ29Jpxdho70pEYWMjBuX8VD4kLu3TWzaCQ0nJB41N+QYCgVcE
EjWmwF8bFZDspHPG0oV+i1eWUZQg11F09H0q1p1errLa+x2L+MLgcLUG9Ly/e/Iu
52I1//HS0Fbh/6dZb1wY+YFiDwfN6Jw2wi1PTZwbxkqR/bQpvTV5xYfookCqh6xI
fHpXG8Qk5abLVQltspz6hRkA9imEzCmsVxyS4dpLklM7Bcu218/k4CQXdMrpbCRg
EZWrQMZ3ddm30RIFiKotUfWWc52kqvoVbJkbNPL6Y/ntBJkWWygi7F5SN1W2AI0G
yiWfOeYG3816NQFlZajwX5AqUmVqQuW6kgg5+nI5/wr1gO9atVmIfvXAOvZ5kEAw
vZlRgcfpRuPgtPaMHdLKLPdk1UCoMYIQiWjt5MrEPW9W8fryeD+TNeDQvLWus2VD
cs3xe+TKzW1R3cBuxE95o5e5JhRKvgTuN8fYb8GXwybYhhQDNVgBE2KLfSPNOJn+
tl3mYKW9K+H+16ROk20cbAJphoS1xR0fJwIJn7YB3q9K2/KYLthSIVcGXW+wUkBs
y9o5FhqY1DPsaAEDYDz5aN2xTIkG4zwESSHVw+nfizl+Mml6s/w3wSl6E/JsWmYT
eUthrEwu7qBQGRuyI1TBNQjFC7ksJ3ibCc5e7AKC2SZ2juKV6I+fSw0JXt7Aw+mM
GS4mcA0aCvEGTQaubDo70t7wORRY66Ykfr4UtKNr3soCmgn2rSEvVcJWqSQG6/yi
MDq+HBhzWAwJyXNOXVRiuMpxNAQL+QETXSy0TJx5kwfOZ4oiOonn3lodUU4DSHvU
bKzNgFXQBOPTriT6Xt4JATe8U/8ywUvRYAoviWF7J7jADNX53c4O2wGdIo69YfQH
+V39CvzFB8vnRPBLOtQOZYasur8NNzBQdwgwno/55QhcNzDCjEAL+pC+nXxt6fz3
NUVYFgMEbAQraBy/PRQuoZGCJly6Fekmbm7Y4zWTebv1DPz3uR5pHMt+5zqgdzsd
qTyEn7/o2HuQ0i+gElaq5/Axboy3cbyUIgd5vYJkb1+FMCVOhsy/1FGKTYg53W8q
KY+dpGjum89uD2tJ/aLrQacV95+Ejqfa3ohsA6BPjVBebW6M+sBt+h15x1PzHjYr
ksKu+dAksvjPBR31fLcTZncHR5OXSnzkeln1Nppyyjjm+CYNh0tttEez8BIYEx8s
68ZW6qrnknoQgSlRLC/Eowrx8y7JcHm1HJZJSKwWpYcrZJkyjifcYQzI4VlKTq6f
azYwXST1fvCKyxztuoWigwkngzKC+vWdR1Zz8U2bD2GgOUyOzVqLh6eEHL8HUXFL
lFpie9brLHUQfQxG5oDMfZWhU0EoG81CKp//DffoC21JFq32q8Z1z0ei3qlAT087
x0vgTEkLOzPDhBtdkaAF234x4J6EdaNRYKq492LaQZ+z2Yg0gIoeJt20/Xe/4qwr
H2cugUoNwVvaVTe5PKEQ9n+PR66K744e250iB0k6pNcMsW/ogYuOhGM5/Czd8a/j
LJDtTpah6qDDjSu0yE3ezroJnQxGMCD9BFR0Wesn3YpJInpjAGQLFnVkH7LW+HHR
J1g5FMAAtStg71jquT5/daZTLGzpEMprVpz+dgQpvDP8nasZnPoBBmJI1Rn7q9eT
NBV9nzsQTL6AqT1tNqwyqZQyN4l/D150swhYof4q6BjOQe7DKmlALd2rk+rCdpzP
JrsI0cW8D7dKm/+MNb3vBBLpwDE5KNr8MgMNO+oohVKgvf7Tq3OA2z8x8Yc6XOC4
GhtlKHVnTByd/bRBYbWA62sxtdG1WKYSMPBUYI1hU5Zq3fI7lh9/kliz+xyZM8lS
CbMn+nLSv8uIwUpHaLTAPRqWgH6YmLkipHK9jaulFMvmCw91hYj9XtUF0hE1Bq8D
VNJTcnxKIk/KsLY+GivJkpTsT3tAiP4dJURKUqqpPwhFrT+ncOY5MxApHikBoUGG
OuA/tDAU/IZAHF5K1XAetLWNdvJ7moGprehVJk/iSxAy/FOmmaOcPJOaIoiKNddG
4hHpSGRWqGO+5K1wzbA2OaVr5lDAO3RsjJmnArg/mzYE9rFSY513Lh7ycEHv167b
u3YzeLTXbsOQUUrxwiJBhFQhz3rLdzAEsG9TfEdHpjlUmIx2UYSLX3PJCzVoPhOh
VldgBwjU9ZhFNHaHT79Oc3uvQpQQh/qaOsGHLtlJ9bh8zK647Ebaoy6b2IyCUwlL
JUMzhUT7LrIuGoH+9DaB+Ibj3EsR06Lp1dt0coIfd+6cEWyb5p6YJ2N9m6aYJcQu
ajaB0f0FXt1JG1RDHlcKS1VMtSZsA76H5BRDSqQxjMuddEhLX6Nt/RYJvhPGJ3TI
Uj7HMlk2jFKLEwxoo912fE7m/pj/6vEq3xDQVkdC1Wfa+CdF9cdZkRA3EqCHvAje
0TTG+0HSGbn3UlK5qQmpUKMUXiNMSk9dxfSIxIdLOaVMlmw1zZBlWlMbdL4jF4x0
5eSAg5fIgLyVeqiE0n80LH5zXfTRRSmltAhnWgFRCjhIIALNNUev4CBu+ktwKd4h
/EiddLUZ2S7u1x4bVHXOGbOpm7rDWRZxfx1ZfIqR6tlFWBD4gn3Of39Cr5G8vJax
vK5+RfZoyPUCiDwfllRSLRcrkccJKQeqVCmPXo9hytiqmji7/bJYDnTj5FFRfPem
qSpcqRia787QKkJlxyVYqnI4DlrWlDZqtVg07D2Pt/kc3oUK0fpRJhIYua4lMfep
IGDj5Yp7hmfQfzeYGVj0cThF+4+kq5J8YoH3Woyn8ljsHtpZqMkf1MI4IMZnKsYh
vy+qcqFkpoN2rEDvTdNiyeYSdKaaFKKGCvhF8zmG03b3hD391sxRvhsasIGlI0dh
WJPqoV1JwqyKw1iHePMZk1ma0QXX79yzJYu4L8UAJUl1cSaVzj9D32ZJivx4Emjz
wcgWYH/ObnvmUh8qP2BXwqH6fn+2v2scwbu/sT+OXC+j9cNjIYNvPnXI9Xs6eBP5
fwk0nparWpnHFfWrQ+NYt8vo01VSL7i3j7AVNK0sIOwDdtgdUtVmSglEk03tMHml
LfBA4uCo9C66XQipGhkJN9YMehSUgvaXCo95FLljAnJkGNf8+5UONx3vo2b3C72q
L9SdsZJYHIJySX1hLWtw4vbLF58CU0agmM5O0kfv2cDhER5DPE1cXA7SnkVtgp4a
GghYVaC3i0N9X1OYmqOjx339XUzSx4dMTOBaDqdTLJJpnrjxbCrzol22O2BPdcTm
VdFldnYsxFomKc+CQPgCcadwyyEMfR1/eVkgvrYZUm/ms5KjzVc6j537H9byUHke
R9OF+AcKU/ghKTT6wx5LNAvwH1BXJ1YH2H1x8w3GNj58X4HuvJV16IflrvGt89IC
pWUgV2+Nlz85vOSCalDpra5lK/1RyithwfPr52kdCXYplTKXcdeBKS0R7LoQSxUM
ghnt78KPWm8i6SfnMtoT7H4cQruiRNXTaM+STtqXSWiPRslA+iesJdoluCgdzjCP
zh8d5zqXkhPpC7ivCqSOJhHD1tUVjJ4tXmjCFzACn79WolE2g0KoaDEkS08/+M5y
V4ICURhhejqLmA2lGHTw7V6K4onVtidYoOR/zjP83oYQHVvWwUthzeUhOK/khqky
kFS5blpqd2De+IuW2dWrRdQKs/mx3126Rxd82BhNZdNgBXHriAVI/D9PskKoWym+
pMKokOQ0JBdHXp1h83+vgbsxeui9KSazkJiA03rjQdlJPYLO9x95NLEmrsgoHfEQ
MuUNOHAAq9GMoIN8Uat0C7eM3QWxLJIuXfjOFH5XxTbe6hu9QmX4U4x7p8AHHo3J
983R6kR7XLTs/hT3VMjLtbb7E3OJYcN5YwOxheNfHAdBjwQ4mnH2WxQ2taTEBNx9
UT3pYzW3LPJKmbzhs8BhKOhnl0b2boacQ3tAh8ZhgH4XC/L1crFa0GKX2skqnRyN
pYhtEEfSNb/uBRG4IAqreNqaFEnR/w3uOOMowkAVuBd/YdlwBT7WdzMzTDcSXkBo
xcmlYEWzCpzMvFRGBIf3Qi9659akfyxtqdRbRmeyj3LnZVP+8tnSiZoLBaGUVeP8
pyQASSr8XmAWecwxl4sLn4Xkfh7sRFjTYq2ZPSujB/pLkkvD+aNAU2gYbR/lA5HT
lRRL8yZ1IsHBStohqtf5sUPwPa9sJtIzFonIJbBpPLOCrJ7A4MOarkw74Y/UH6QL
up9/b9uoNnc2cZp/y9ncgzw0JwwkyQfWdik1s/0HPvfu4L2drSjad3SBQFqCNNw0
Os9iNy7kv+42dcOaC7IujwzGulraZWEzgT7VjJRUYabG5hC61wsJplUakilHlj9r
wrHU75irxZg7LvP2GzjJfltQQeWj1rP7Aag+Ab7OdhQF9y9PhUzUiNhWAYpAovMd
yVyvCq6Rp5lQdgDBI3fGFqd/aOdQM2KvTfl8ra1WgybrxfPhyo/SbE1rEdWGo3WL
YNeAqA6IED2SG9sF48wn/xREHQ4UaGYkCXv1HmNw0PZLh+0usjdd0NMjh4G23TtD
dk0dZPA2pJo9frCgdu3lu0GCracDuHy/OzU5Cu+FSYWANlJOK/UEaDqsVEm5cWjI
Bs+rnMWiA36fo9k7D0TtsizmH92IM15ksdUGTB1gsEl5u3oSUDkafc1GFocsrha/
zM3+cRUAle0WXwxelyg5k2a9dwdtGBUumFgRF3P0TzI4swG/FPHXDcYk9/+p0iSD
tEYqWwpKEAA6SX8+c3BJbNwiR2T6qvsLUbaDJ683WOYWyv4qKQotolmGsKeqcLpX
oF6Yxt283ci2L0yx12WhVk04ZeqL/BIMoy46H3tJ3Y1jH4nxpospxoDBXcxHg86v
MrvcKmb7zfWvIIyVbVmvCvIJmS3AWitMdD8oqTDa7of2W0lGle+M/6bx0BWcwkIk
9i+By5LYUJ+5HiZLqQT1wNCQ5RV8tJTnIsfCM05LQlSX7tFF2QQTqaf+zYIVYYj7
AxLQzKT7qfMzQ64a7xRgk2J9/HZG7vg//qan/2f39dSloTtwZ0KuVmY0cCvLrq/u
CGY6Tn7i0XrKwSrNC5m7EQxmI+fhkb9i0pOvhwgFOMRjuKSVZxHgj/hOG2Z7dG29
P3fj60H+ZpfkP+l3qg8Ot4q8/3rttH9XmACeW5r7FfOmAbhbvyrx39QES32IcZEE
LNWpKYITXjSDfjxtiZC+jjNeRLubBuIIT4stH+WS/uhi71qttddkmMxhoMBVGpKC
0XXObhTpMpaiB73PuNyVcfBpRA81VnMUz5qj0WOxnq53wTNpzaC9w7zcUgkOOUTf
aUObk8aPSw6yZXEnDrMnX1JSOuWl9gnut+JYsN0GIJHokQCiDHGx929PI78L0ww1
cAvy+O7rnElgi+yYX6WJGI2/MLJ4OOE2vulx+GaNQX8BIBglkIt362CwTve1EaJk
T2c7Vjo+VTZi9Tm2G/DtJktVgq9rmzsYIv42uu/dSTW2dkPVudK2D9xbA+0UN0pF
+aDAiS6BQG8VdxX2M2oDgjyaM9jt+FbdDvTYeSDYtIYPQexwLcFo6d3n9P50YH2R
4MsL1L3Ck7oJVI3Ncg6LyTjqaR8ZqcarnfGhXACO71DsyTMK0aMhA56wB17MSNDc
R26mqQtYoVVlJVAju9e23WUCxAepjN8ivb4QGG3/flp0idIrvdNetkPVOe89YEPr
1HCxCjXBJZY5QcWRR7CUjDjWIktXGxIMbFir/bVDRlSf7M5tqXlXQY4aF9ecXVlM
MmIYDTunzA2sMsCP61VhAtnarNlpeLOc20vNZ7vNWZDkoaK417QkNShyEz5m1tnD
jRKNRH83mUBpc+LVvoSL1ZpoiBSKXbivQ9dXyQaBsBImc/Nh1c0SD4+WLw+uqjrY
w4gUPaKScZmqiL949877YFo6xgHNjY76ZVeWaIyE1vMYE/BiavD2Wahf6/yT5jpl
8LlOJVXjScczv7SbwQr3j7C9qKGxmDIJaJ2Hk2zgX+jPirRhyQgw1yV4EXi8k1wj
HcRwz/cmdG4rz+J8RZZzknaRaMBTNtNzjrgPS3tRdemXhOwO0pLu1nsCA+RjYj8n
207KFSs55Ht+tbeafCb/bEMdg8I2zQMacsJXfcJbbeQnxc2/50TC4V7AonMZP0GA
OMZXIb6MGz9dnR2IgMOzqKwONfRTwcdXy6TxK2xOmpGuRbuZDUvT6wWTRHBvpNCw
g5rInxHGKwqu+7dizwNNnSFmXxV6mGbOiJD7qZn8CH746iT41RzPuRwMxVWh+6XQ
IlUiqe02NtMlrCjmL1XHkvf+LATdpU4AOT5P2IBFsgBvKrplOnNSKV4EZeyBlCi+
al9y98pnUJZfWMt+UKWT8dfASGISvFIFIDfphmA0lsbUW54l9zG1gng5rkEc6YeJ
vatG4bonVXpgu2QP4uY+7PE302eYDGwTXD3rSKCCm6gJPY3A74c+5Z7E7beaWuqq
7bYxJyINkZI4A64zNNfSKgyJvAdqfRDaqs25N2zpqr3KXbUmstS0PnmxzKXhrKs0
AQ+MjyOJuQLGn1AbfhATW0l646omG1d6VgSSfCqy+g0Q8VhFz43cMnhfX6oplvIw
X07BUYFY6DkvSzKDxviJz9del/J0QpysNqkMFKVU7VoM9zpOVWXGht+l+OnR7kTm
435NXZuytuPYghrmnOKuhG5MC2zD6tVIXG0lYurj+zpT8kxcFcIMvSQCtqIYm7NA
68oiLA+jea9tmKyJgdBeJapTtUQvlwqJIxhKpS9sHOesV3AXgy17lUP5NYO57XYh
qFmHgseGt7Oo7+ATVnJVaHICtVVDd4HisdgC4dD7MTnL9lDx6EytY6LheYzq36fz
b3f7Fk3viMx876RaSb5t+aZZPGRBigSS5G+MDHsdLKDkH1kaTmv0GdZYHjkwMh//
Os5DMwbRR6V6tyzlJYyQihlRcVRab1dcyv+x+P1CAm3hySjnJ9W2MoX8Uwx3n0qg
i650rABR4wtzuwceoplgGPJEyaAq7Oo6SgjKebLgAtpbC/iUidecmg6aSnyiMeUL
0LCxGsHufam6ZM3patsOFRoiTQd79KftZ+nlKxDNeb3xyzMAo60uqvPmfrpNhvZH
5itpu4DnsXpzC+o45HMwrK/VVu+hRK+DhJvV7JyKuIdic/TPQ9iuRwxG94FfZ2cI
ufwhTktfELFs8XExLK6UIs82iLv7NRZ7AlJfaJOrAnC/4JiLuaByhmsHKTz+sgV6
psM/QLqUaz+2L1ff4TQjdhe62plecIhDsJYUhe2YUh+IXlnneWj8YNZ5CAVVCK7u
O33832e4WvOqeH93L7uPuIMWC5uqby50VGyxANM6X95DSFOVIZR/Gu9EENXxd5c6
5zqr/kt5kLHdT+DSHpS5qXo2M4fiVlFWW67ZnWcg9V27HtX8FOx0AiLtXWKIDO2r
gYaciTvrBlJByCjiE/Hfd38wV9JBMURQyerpShf+7OYoyoqVdanWiZINqFHdSQhD
dy/3O48mquUcJPCZwBibW5H/syNHTJsEvHvwnQpYdD4NSA3WaRF7a+LXwEOLC9Ca
4nfYwXoQUKckogi2KJztgAa/SZr8IcV7mpyIZllv5RoKWkqSsxiz/XojSy8Ij+It
Ox8JFAt5dS/oz8tQ5CKFMlBlMCmLeb27S/6zHqaEQrsTSbH/mPiGprF+oFaIrpg7
DXqgE8ALPWHLgUD5r3X8cOkaQ+ZeDEasD7WMwzoIxPozDivObruyLf30NvJnXxpU
G3X2CJq96jCqvH08a90Bbv2/nF17iVT0hFg1k56Mtzoo3hhB4vZ/wcSqhFI7smbr
38SsbN52dVPosp8PmU3kY+1u7UKeULcQJVX1wONfiHyZekKlZf99Kwo+JW127U0v
6mdz1JOKWyycDwTarB0tZvSJbi+0U1GjmdxLtwYmII1maoQWRw1IoSM85hZ/tzrE
P1n96L9yklaxsmTqgaJtKCvYfvOe1Vq87PsN6qELeEYKhE5TaM5srLRA53AoGIdI
+5gT+0xLyIUh7NZPWD26ookza3IIlYTKYXmxlZIBD61dnmeHrLwAMyeVkDXm6pto
XvLI+rLWSyL18Iq7NY6heHL2beDF1N/6DveM2QzT5gNLq8IRM891iSnCwizz1jOk
YtqKKE+LgXTMhP0ICL01B1mVPzan/9TmyvGNL12MxXtF4qzTCHd1grVMWCBRiPW+
z6Yj/0vYTyoUy3nUJTpDAoM59Ucl8nyhyQVe9Q2OoIuIPS0DD8bbz7IlFB7ZnXmf
1rX4QrTvUaOpLbT7+OndawYVQIXra1pJn+MYofK3+B1RbZ65F3fDw51Kl7IaVmVQ
3VNHKHlThQYq55jFRsXQq2ZZOZoDtCvoIdkPOUYqzLAxtzqAwihOL+cWaaAbpw99
v4Jz3u2awBBTaWLDNS6I9+kNLqZ60CVcAPvueXP618FrmMFT7CO08Coexkm12mRD
QmagvYCsoArm0vchnGyN/Wg92/BJIkIGAQ3oYYZOiLdZWGMfxR5V7zEwg51UpkQ7
HI5OvXT/BoqD8q1GROc1dZSj0YZLVthsnZ9dCd6+XAEohl6dtuZRzSZuB4u+rdq/
qAadgmy97QImAYOwFUPIlnqI628Tbyf3CmnVmwk27TE62tpDdAsMZ5iYYxuzAOib
KfKhQXoeVIZrdYc7k+ZlXndMgV6JTKWkcAbR9rgyVspMCu0GXCS7t5MkILfCiBms
tzykhFKcn4us6qKbJj//df17xUEAYMwYLTEc7XLLBDlQrZqHUcowzopxgKcV11Qq
+Ea4hG07JIdisb+Sj7O9yYJQizLHy2Y73x56aj0wl0d6fJ5sSXjSG/Jtsvh9D3mK
R9MiyJOPgmRWUa0ADjdO7uox++aWi3SGiVk3+Qjt4tireJUH+Lc7p5YprxREoHMA
3gio808OmqETv8w8AlhS6GBAHs5ECmoYc93LDxaYUlp6bV48N1jml7MksyN5pIJ5
zB0cCtNmz4XdcuUT8SWWkLStoQ3JenDwGLYi5cRdSQecS/HiYqbeZYPAJUD283ce
bxYEUIleGfayeNeDe9scs2nrrlw3dthP0ak8+Ckbfy4jjxADr6LCznTwrItgYu6c
Qph74jZX7ZOmaHjVlzsOblDgXRLnpBkc9WLTtiGTatOJ5cY0G55T3zpQZYMPiY53
DUNi28Gbt7wjeIpJCqBg3DJQnl2E07bRrev3CaI3KfTbJWZ5YgDkTb2uQggE/i2o
xua5FSrom//5PMzN4mDKLWk50vKWCFruxpS5tdc3JO/KzsCkJ3kLfTaytoqR4xm7
4k6A1SBU5vv9iZIBsMZak81ZHa8ThPIBmluczY0uzft3MAXcq+tAnkdwm4FQv7m9
CATpRQJy/CWBVyp0lJ2TmEqltx0SE4htzrVhj3xrzCGLsO2PHeVY1WAIic+sq3AK
k6qovlI1xLhCq1OxHCGnECVhkUqOVLBYOCfXUMC9BRmwhRTJrPpsB3IdlRUXp+f0
oStJl9nxLo71YHplLF3H0Swm+OXNhcmem7mkGwyJ+4HeLrdm6szooE7HyHHJZn48
1JAlo+DBw5GhX0WvValgbrxSVwAlj1H+IoQ79GI1MJZYuBkQ87R0om4xyHY2G17a
UFMdi+yH5akL3k8BGAFLhL1sR1/YSqrOeTJvOYacMO7nKzVzBBgMYDF1yrrsolMx
AWNLGg7Pzvql5z1s44pv7dRPGOe89aBOfM/gGG/r0lIKFoGuVMOKuionWVA4X6RC
tjdQ+Z7mB4JVEOoPnmEB47LThFrVVWsSm15IAC3YccYdym//JIr20vFVEUigbyU5
simKlxTijI396zp7mumN5cCryOzVmP4juhwqLo4ST36bt81prUaa55yVGkM9uk3Q
h4CYJj537fR+kOkFAkBzJ/twFj8rU5Q/ryo4485PnzNJOYM8wVclMwbjOIK9DGVh
9lMzt3lsuJitsM1RZIuVUP54+DIc1zSyfZewcrrs6lhSmsx9pz/US10Z5SNmVaed
/fSCEHQN3mQNJNkgHtvOdWYQxVNZxjeLDIb7LVo3f7Sk2MMptQkVDCjdsOgZq7RM
kg47e6C+OuyI1zdB0EXlFw9xmN5Ww3bU6BHFBw61+YavDdvrteiSTTcma0iuI+So
aetM59tU9cJYAiEHAhBqxlrycyp5wnsULUPQwEDq5SY2fMgNtAvbPLai5QO0bcJq
lBxHp1QSR9Bu27RxAqFnvpcuIMbVU2Wt2/i3pXoUUOXtzzj315RwoAtoO6IT+ath
/DANNW6KbMvPWi0QqM76ZNIpEsAfkT58cT/OtRAmosHq7l9sD42RUpgj0v9pYyER
/5/JnapnhAH+qcrQCeS6XMJabfpGZwuYkRWTvYdxzuwpLVtrz7VuOIb7KRQ7CD5F
+H/M4dQ310a9UgX0xpvmBDecnNLP/zlw6M3wDlYbJmDkRT5CP9rQUrui2LqCKlGI
oeMGAGD5yKb7l1HZfNq6/Z5yf6VfU2yKld7zpfRwzT8wYENsVlLlZ0+jb7aTFVCY
Ct84dWP3QCxGGbs6OMLdtvD4OE519vSmUN071CuX9bUu37qOsLzPOIT2MoAkSafb
79eM4s1nwG4ZfRZLkIeW7g8BHYrFXpSeHOwSo2rs/vo4EfDVGNovMEgZbecfM5vz
DXNz2xlr1rOhZNCxKuwEpU/Ff2eUHzg1IDDWBDhuxKH8fh7D6sHevX8cQq5QkCK7
okhS4SVOJ8wOKgzVCm0I+m3qn6xc/Zp31N17Tt9mjzc9jiFCmrdfP/0ScguUt+Yt
jiHGiil/55LfHqy6bnBP8WUlrY6NO3Oyn5cSQkz1iGcrfLfmpFEbbDacBcclEhdt
r+Z3ITxHBKmGZo9vd+qXRE44dNZ33wIUEz8U8tArBm94LtxdpiRFp04rPQVkXlPk
QGScHDuSxJyMcRCwsZ3oyux9Ex5mRQ+R0uRrzjXIJ763OEkHEJCM+CDbH92YqTl3
Tmoeh8eO240K7HGrzl1j4E4b8lgdCIaSrkR6th+A6ktWjqd1yrS4kLKVZyLLxPuu
7Ne70a+zLXEBGFZRuIIM9CeqQPOzYXEM5X5wyPQ2lv/162+Qzj1KgablSCk5kP7N
n9A1YVFHKLj0M3hP7iuI8b1F5BYX7bvehFuFHiK5J3PJSk2RI9nZo1R3t4DOhIuW
lXkeR8To4nG2FW83jSQwi88QVjiIN7SbQimjoa5hLaD6ZqRHj0BYRPP1bxrsO6he
G4eYuxdbX76e/HE3PNPdJ4XRsUxen94etJTqfQ3+0SVkT43rDzoUNsvrx7SGhajz
rwpNBquJUyGN8E66c7+4F9oeYw9AM5lNa3MHSfXRzzTWo+L2WJh4R/kCZJkGBEuT
EK/EEALP45SxZ0QB+i9pVeZ8EkTovDHlqpFd2gfg8hfxlsJROLeZbiIQCcs1X6UU
PcKoqZGAM8rUwI5Ph/50aG2LsE0S9Q2o0kmV2KK6eHKlezAvn7FxdCmWX/bwv0Gr
1Z7/3q360uSt5TA4thoGYoyM++9IvRe+uL/Om3Lq4NX8sfIKXa5RAyi289FUhbEJ
y/rPw2mX0MKclAgvUsS/aixJtaNcMTq8RJkueSlyyp0k2924VgRiqa4c2ZeoRl07
Q8X6v+pQ/LNso08G3rFubJ4IlmdUbzfYvOMvRrYod8PScSNmHlaYk+xjW09yvoFX
E2JYPt+pCqHwqLYxBqYzTLq7hrVaSmK5sqiPtetfkzqlQQhpO5uFWage2yYGSdRV
K4Mq8rW8hwpcm9rfqM/gCD6JBjmiDracqmT2RKbV9UNk6l2igP53WkNbBskyMYzK
8LNwAkuZeHhVmBcj/ZlXSCA2o+QueZ4um82URrHLxC2omHpgKpi5GwSW7m0jqN8K
b4+UcRIWWNopC+kuWPmaSDxLiyyqrcpq25fNZYUxOQTF8vgHajF198QRYSiJuv2S
l69spFpZFWoKW1bVIJO2aKm3YjLu1hh0wJSw977gw7OU8BrtH20ijDn407JWY/Wu
X9H3fbHlY+J34Si+2KBlu7RAZQwZuYLIHN3W5/85YKmqugEOvKVEWOAnsCsrGdZN
LifGdUdtgT7EhhVTLBnlymXTIHktTl4na7+ICavzn1kkpDNlmlqevnS0Kj0q93Ag
ZilGxnPDQ8+6IRhMrV1WUa/BWwvgtkvhrsPrbB7ed20bFdpf/Bpa33SH4q1G8GRF
IF270iQomNCNnkCiDFpBNGOs1NLUUV1oISmLCwPBP/KZpPb+i4hShWZyU2oNkpTG
pkoIRUG9mnnYKX5zraGRLNNZQqkYp/2WblH8CXKx7RQZexFqT69By6AIYmMIdZoZ
6Oq19V6tGuZ8SSSxiJyhsWTTNMtKXpYEDWE5I/Ame5SHSXeVi4LsFPnmDVPpdY4L
6VjWJkrxx0O1EauDCbKmpoWc1JJYx+DwfB4OcyjLYHDcTNApgOqHhWNa2+znqAdl
UZMNH2zGlLN2lpkMHp69sPrIp7Xal9RP9qt4Mf4YZ2O6U9aEOSGlMG8gGbl3zLWD
AFqaZPbMO/1xtm6eJqhB35ArnUvaiWbrs9wDPbKKrOpRknwtRkhUlSLIwUlnMAd8
/T/ZogJxscRSyGjsDP8S9iPVEn54K25AeQ2VNXlAXZ5LjY37HihqtQ+IvAakJkEV
X2htFbyVXytkm+R1CCyAAKVbetC321ie75wPnOYpl25DQQ9hLgJ20YQ/YdGVanPl
QSAAmc3EaKWfXT+003ZbzNt7OUCd5Uy7J81hld0NVfqqXSJezGARRWpHDgDNQTK7
Tb4MHSl8CW1LUipct6/f9ENHS3QAONguFOTPjaQ/0wvGxw+U7F6P0GTbiOYogkmu
lLdvne/PN8iVHwCyix64RyijqSiQSR3m60FCg7bZOjYU6VpQDyMUqlUC5odAIhUg
71Jm55T09Ur9tth0QC6VzXMJ18lNhNqr59Q8U/v9oQpZ5ZMRhsTD2TJz3i7T7FPp
2d84Q+hKyjI/qY+j6t3+CJKJKBoCGBrdvqGBeM2j5TQHau+8LQIZLjcbVcBQPZiU
bBgRtieChWFREjdSa5iXecayM9d+krohEDD9ddxRpUlDPi2Zb8s1sKbM5VvuTXE9
5uCgPKb9HU+3MkDz5ua8VNULxVhAkdRIcB+bsWtZq8FlfGVomAS2j8GtSa+8buu8
hj52IGQTLjjwjS2h/Py/q8LbasXaZdm/602BdP0ZfrkLIamWVnsgnsaYlj3l6XC1
zjhxEYYnjUYI2w3Clxa+S58PdVHEaCk940++QtrhesSdo+kpVXutbwCy4Alx6UpZ
76cu+NJxQKufHWF58jmy+lfSXUBz0kMts82LEI9JxZdd3mj19T8kTEM1rCfG6Gl8
Cxxm3echWYTf0E3zUdFkGy8UCPkazgsdmDxZpZdJw0VbqPbGVrI/7PFn1Vge4IOW
cFkiqyx4jNnO32GPeprJBr66PCXfmym5PrqWf3h8mNK8pWcR60OKhkosZmJuH4Sy
2QV0OGOt7Ajz5rYEKGOvb6n4zaZLBOWLT/fT4/CrNoVtf8/RdcMub7OWPbfSMy80
pYVhzbN0OTkri8TIhiNYTz6AEV8mjK++GDsuTtdeQFWiR14dOTfeIx+gR4I+OXeb
dcmGgGuoIU1SFGiXGhRapO51FXTnclE9NVAAI38s1XKQBukGT+TSfQ6BiwrVVZOJ
bET8MNt8fMnVfSaGKFwl6KddTySyM3jPCDYZ66L28uFXK+fvzxURJyMdwhPAaopb
h3+xqqJrOmDvejhfzLaNEPiy3OuDG8gys5g0E2btif3JDirfGS4tTplZbGpSjGBi
gx5P/xKCFHaxZsebBxk+y8MxxydEIadIl1HgWXBT9+g/10JwlawU7iKDKn+qcuHp
bl76oSj5l1/UR3htl07+bq/DRFDwrrGwDFwocz/UTt2V49zYB4bwVP+dEWoBbf7g
7IsTDMTLp0oLKF0w3T7NbmwcJ75p/2QKI2ovL9HcoBob9rYegiPqtN5KB22hpf6f
u8jtlTUIfWlCd6AUM4I1Yep/i5Yvv/UBc2V5nBt0B9lmJzHCm4/YEFXp4sUszXpl
FnNmZcmbo1dMWfNJscBPzdq6bt8jk2W/R8GglSLsiMUD7ZJMYEN+ZLtvrIPAu9N+
HhotQIw0YpTkb9SXaS/j1uX2JvLkpo6HzA4qjMtLRTRc27NlgCVDBbNDnqF/eoV2
rEyqM+v0/gzo61TsIu+KAxNNt/bR3+b1yQvnmTDWFz/SE5rNLmbbHFSEn1TOZ+SY
W42SJrDtfUeSMM6PUpLTlzQZb4r3TgRezbTB/nWb7XL3F/3lRWc9tBEfCsgsRlGH
rM4AT0lkjSJf85GFIGyMTW0efIelGhLUOSXyr/nK25uh6fqvIAbur7GvgSJt9qnv
hdHcKyO9KQ3KZjJyj6WD02yTgiYOHfGi3AK6r+zQsP0BHonlwiS5ELmjEOjSEcaA
Sb0FdYbv67zLjlwoyYTdopZBcowoCn3t+AASiQHHBlLZ0d2tlGSRBn7UcRolWTSp
GYFUP/emFibUa8LT8sCnRzE1oBD7uMO43qceyc4lvXd+xvNAeL+aE7BzgvgULr94
atqbb0+0TCSA19khkrlNzR8D9xilzvKlevjquMGUpAohLssq2v9M4/GCCs6cmIQr
x6Ndifx6+gbAxk0ehga27CaDi3CEXDhkqySu2Mw6ca+N1rkQyLaK0sdUcrD1dYrK
MYYYdT29rd470A81nFMZ744E9mHHnZ9jNbrDrOFqd5eD4q9/mt6Dkx2oZPHlf1UC
7sYx7vll6Y5Yc04FXXbD8P4qvq8YV0W/cOvlLhrW/ubvMrHHg6rKczo7uJ3HI/av
908WbY7fDo/Dx4qG8GITREqj+QU6GC2Nar1f0xrFs9sfPLfpwJUn/yRAXhXMUnlX
F/9Exmx2fZSud00PI/QaAvhJoXKRfSFx3JeO35UXUBX0frShhTD430U24IhsWBsa
s5EhephMEiKwlVi6mYNg3z3NDurr2WaK3jIr3Pk46u2Xa8Ly2vwIKsFz4gUKttEy
j/c8sVK1hphUtK+HGH/Ig+CUYruXWgMNqKlFOYH7H7BbotI0PmtSadh/tln2fth5
+zLjZZupZ3/QZ5yYqNAAxc5HL5fW3ewwYku4GrLEOGAfoHR2kxDtoMVNhBp8p8EV
E3q/PqacUXEOVR3vGcTGlmNnAPnb8pTgr/GeSys6g6Gj0RKOPZZAuCPAHpAA2KI1
nMBQYLtlxcg215xcWM6j02+6rZypXHF+ryFlTqBzB2fl+yu5KyJuEqqHZL29bwjR
md9MfeJWHWDugdEUPEOqedKb0+rkO/z+UQeveW+gAQeYoKUKleyMYDTSso31LXMm
hZPSoxtZMd8/d1MDS6HeM3jxMtPd30EMx35Pq4HltlEjZZ6Kj1RisBRmlGyhX6CO
3hY4+nTttR+JItgLewJZv/2kib5EcArIpC0fBvCaFa8uyRojxP+gjnVSbrehGSL0
hA6FkvQyb4xVogW/NuvEeYupprjbde36+ETEJu4MZSGbHB2Z+UNyBgSPOtlB0z64
CVoE3/CWmrCqHZct0rZFmcJS9bpRSLU1sKE3lhZD+7ctcJT6JSdZTcZDPFHrAy29
kTVvPT70zgCF1ngi1pFd03W2RBRil63b4mG4cQU7sNE5aQ4/sLGjH9Y5cIGhY0uj
FkorG2ghOxr9q5lmYZA1RQMSTY/mHN/tFPYBhAE36v2Uu87G063gMtXfR5f+s6s5
tr3tXtq1CSAB3abTlh4TNppL/NA4fRhejSv4kwHw8awKx3gsRm1xUdC2Dx2ke/EZ
GLQrncUoVkOsUCdlM6aBnwx8vE+jnypFnR7SgP2uqj4eODW7Lc7+4Jebd+McCDhw
X46oj/DPkkTAA+fJv/QodD+yBBjaFmoyLXQ+ixRSrMob0B1WwTRHMAlpCZTWCi3C
uATefqfu/yn0r5Y/rkNCy2wyNaebHK+DSd3+ZvVg5YC1oUAxvBi1F2pB9WnGADpy
5I4xvJjaraEdNfovzxmusTWHKXMPancx/t80k40t29R9PhkXQgqP/EFpPfi3SWjM
EUZhpaZe2ZNlPz7DkPSxSXZ0SFHCTq6/1XHI4vooYmC3ft5FS/7rx5sDv+absxYR
314X+Aq/JymjwvM1C+EjXEBtNtY7gHPHEaCl7vd15QhlszvynbISJh8ReMJ5oHkB
ZjGoaEGeg+Ueu3aCnxXnWoZ0BtXO2a8APolM+DORbEx7Mc1qEcKgl56ScuXuXO6M
wrRU0Nrn+4ax97Z1BvF5bRA0gPYuirao7OP/UFvihsC2Yy9AqvexOKIbG5P2TSZh
REuciJHcSM4d4czMnMU3fR56h1l3pav7ULsIe2nl468uhMObzjW95YmSI2HVcnRe
DMp+4hB49jQ07YwcpS9SDeSicyS8FMefi3ce5ey87sI5yfIz8Cgq645fkXCuDBjv
vyzrpMvgBtvWPrYgwPk7PFv17rgnx9EIlQsDryr0mL3uvEKrWG5oW3D/Nnw+VrHl
GLpgr0w8G7xoiNy1kNrDMyWGE7SlaGaA6++dnFIr8HkvaXOjnSRz1zYXsPgv3Jvt
c1HSjSmpfN8riSuiZS2bzsG72E3Re7xxPQZdQbDEbprZzaVa1kfY7u5V8u7MUz1d
3NQDgxnjQ1eNmjrDfX8z+Fkkhgq4v/60CS096SyAQxHPoGVpDyFYYcPacO55z2V5
qr54aZm5MgpfOf6EC2+bOJiDiO39eMdhsBdk2tt5rYaH6hnbA2rJ+5wGtQjJhjWu
vYZWdsBWATMclmDF4EWhZhX157WZfQykHGlO79iqEwIcio3N2pD6HpsAo5lPEzEB
HMDRCHpOkhzZlyejRTWHhmJXxUkHTs/mrdHWjTdVvpU1XIY07iU0bVfzai2w6YEZ
BHPSgiq0cz8RFnEardR3Vdb6rPEbZZ+MD4rErOhSl5udhwDUSiuJbIRQBfQuLnEf
Tp1PBhLTvN9Sk20103U7b/mc9SiCCBgcyNYXuwW8QVYxnYXk0LSGLUKvroL/RBKL
Tty/rDzycK8WOkbQvL0O4NicDJzNhq3URG8W8errK9CoEsAlRX7QkepXfM5Px3RC
8hnf19HZz2ddhLj0qDE8YrNwEnkR/8GGdERAJwlMCGhv4R6aXbl/n6xeiw5rZmiM
u/8CJ7dIoRCXcidVNH123JuYoNOGBZAJq7D0DD4Vk0cfQhGMf/0okAM/8QScK6BB
oYwIK3Ofrdskls6wYANfQsdWJLnK+n5d8zaQ/+wT3CNtJMpUIrqSsZ1wLGnpnoCc
G+WHn2T6G754jIL/bMmhqv1V8/Hp+DMJoR1ML+IdEuyVVwEn42rB2QA0WdkMZPUm
/kfR0doCfaGlgR+fdwyczNeB/fcYvwgvlpqquJ+jcDa8mFREGcb8p8SP3hWYbqfz
Pca3PvS26XIKD7j7bXUMUdJu6t4QOOjyvIm9qVBotidDo6UZuz1+K96E+T90uqTs
vEhmmVZQ44qc5z5MPApiP2ZlKmu3lOgfbgGoxUvJFlDosi6ZT5oeV3QG/mmk1xjw
7+iuchiW1aIooiu6XFAOXP4B0dPxVA3MFsqkGjZXOwk2wThG2Ucer2N9PIbVCSB3
Rko3JRP0AXrbG/Hkk97Y5aildzFCMQvxmzQzBEp9+IrVQCw1vatpVotGOlwVgkoS
sWFEELrWDrAFOjDuOmXtdqHIvZ4g6yXZDYLHW/wTllN4+yYMVpY7WlBIu+ErRLoy
WW8n5dHc3lrY0UH2XKQBwbWVKiEmqQaLjtgYu/f8cwCWIksZpKMCKziVbpwULEBM
18pOPh9XTFOc6eLd2uZnnYQJdSFPd6Tx8LoiriVrR8aI7hbcqnApmBmRtCpNC+nP
4B7A/yjmvskq21ZTONLJxx5oFNP2n6cLIjaLB5WLxRS76stq2595ONabVOHzHm10
w5Xbc8MMe058cBnyfGu3yGN0T9VPEubcDGT7OgAoEZDUGJM4UCWoLCNpNPikCBGb
t26R1p2htJmcc1rgMxakPKYPbehbTxC3sJ8WfMmLIvxRuFc73LMjx2Z+4msL+9Vo
Z7nZt5ic8HYk59t7AriYJ9I4MBErFH9b9xlEFfqf35T2v5/NmRtg+tj0ugODoijS
LLJK5I+YPbPSci7npVgZ4nCFnb2zMfx63avLAt87EDHeTDnWmRH/RtnN7Vt1EZoT
k6sgODHUCZU0MQ7r2uZ+q0c3Ikopkh4OksxRhQuED3QX1oYdmBjjVNki6NJXPFbn
ZOAmEuw8A58tWNOkkuLgA2kYg665z8BL6M1PjHOv7qlyt5z7AZoJVhvzbJhokOaZ
/5qtv9IueHyALopw5s7RtizMBSrUv+pL7yf8ngPtcEd1Leal4VqsPDHT/XnpC1JV
FZfjqI1MvfKnepAYc1MR09aHxREt+nHkQNBBJUN8GH0R+6Z759X+A/Ow43KfQLly
envkNWuLFOHSquGepvsAUa8GYa7lZtZr2tlHhCn/esCQhGfDn+ZGHksIdM2HsSkM
WbWVMzyGmGLCqyFjx15NbDpZxM9cFo8j9Io+ZXfzNbv6wieZHIOufFsgy0Lk5s6a
lc5KNaSfxVBYEkW65sZiDFWsE4pjCWcjmDbVkT/+Ls2ghuJ0VK9Q8B58aEko1CvG
29j7eIlLes+8C2rXfnozN47hN8QoN/JtXfbbYIA4xmtp3z+qhQh7UuVbmcQAEvWE
FJVssaTbdOALMQ88m1eg/31+OSW9PmHxewyhxYmRFQTPZdfeoR91v9W6B/SYpU+w
4YV0jMcw83IH4lKcbnGrJgnaZIsgut+tIFUuyI+vuBAX54yrI2D6htWQLEB8rs8B
6QBBnTkIvwcW2kwtfZkZUG0QjGpY41JOsWiAiHOFYLVIMsfN+7PqmVVkZyuWWKWZ
0Ct+TpGL+SVadQF3+W1KKHOimAXMu4TAMLMkkKNY9FUJFq+++IS9syjKSURAS8bu
DxSyWgTTV818PBrM0xhWoUqxXTkl+NsRo2eMLuhb46N7CZc6C16GdBjjLkWEQllJ
zeRZJnVSkRNObI4r2M2I4HtFRiE1uJk7kzHrfcReEH3pXpygtSqEbenfy4RivGeI
fm3mnIjViks8x4hn/WnJLn0uF6xC+Maoa0dATGaKT7lpv/P8Oz+bnPWcdW0OwFKm
4gTmDTGXOEKersaNQJxppDwNXr9X3fux6b/JFFyafVHqvHZ9jDK/ILea6EdQ2YA1
gRixZpQXEEGunTcrCGCo3exoQzG2YsIzLSy7ptQ1LKYpOWFNknqvUIyUZE2aZrkD
cGpViS3KNM+g+/n20lsW7nYkrCLrmNA0iKMEO4aLzbQ9dmYbZ77TinMDGfcOFTnO
lNVJOSdCYHxBgueFVevvr08ClXPHtb4qKaanxyYi8UeHg1uTO//0iEwGbfDxGqIA
Uw69xhHpjpMh/m7jWCOkFUF+UPpgp5uvrb7OleR7inAvryYA3NtTl/1xeuODxYbq
LliI34Zw1hkwNuhMCsxLHm08VqxPKaLZi2gh5ek5uty2FdcXCGGARNVs8CHtrzXJ
BD+16FwCA1MO9NfsuZlvM8qaMGVBeKAeZvBLApgRe0YA1vkkcGsNmlvrtZyl8kW4
ijU0X4wLZ6NYxPv3HyDbLGsV9ORWBiyW+qCGlhPGFZTK6/6GpapQCh8ftqi9Qr8s
uWsK/sKlkniQ6RJ9yFpefd5hVJOZec0nqXvAc1rGbpr5wo8M/CcHwhU1Jsub5zf9
Gjz+BNJLTi4aiVvpOxwNUExaljXqpU65FSLz3okzftBefzn1b7C6/CeGqxWyerlA
aoYDFUwXaTbjlELWyOKHo4Fqclyu4SpuSNKLjz+nEatzuaVjdtHhleoR65opT2mt
aeApwbvl6dikono4Fc/bXPC9a+K3QtHLe31M9S8Whtj7D720u4Hzdk90SNpk4vhE
Ljl5nbOZWf10jipcM40s6Ksx7l2d3hwtCY4dNKaXc3piLoUP5GH0WD/k5sJRsOzO
I/3alQSAmXj0Y5LdfHnGyqgBh1FMfJ08kbOm1wWxbB0J/8NdXiG1qXdK5EIY9p0x
kW9cMGfJSS4BzQ00AZrCFoieZXRJdoeQvuNfPeyFW549a42ZD/R5mElhqJCMz0pO
oM5oqDqa84EVwfGBOxjZ8nxvRzVsBt9IS3MsnXuK7fQXT1ZZGDFYFkvQ5vsMlSBM
N8/mfDGxVMM45bVe95aAG/vgK+Ss+S1P9nhKtIq3Ys3HDTXNUJnzbJbq85NFPQjs
ncwj7gNoqFJzihMV+8McJGd+76JHq0i66yJ/StpsiyGhKaqpOBXZ2NkrPiFRRuid
pPBIL8IbgPvaVdKpX5PViYF2AnUUBk/6DADmK0znRWuhGMkQzXS1FWL6LqIBJZ3G
zSLzSVKJvCxRF/uPVsFdMvT/K1xBcfaAr2O9irhrNV2+bIYaGy8fX6Czpfh7Vilp
CqOcp1e/kdktkpHobvQQzZCe904nXqDdBQavKtp/cQq6WEymx2iA2YQponQ6rtlq
idZ6GZuy7oGBW43J/Y4erijPelQHBomxcXS/xn2c2yimWJxcFSFNFT7iN9CYn9oW
+v5d08QfRkfxZqDJgs8H6NpS1Yp3kQJHK6w67YDldcHGDf1EzRZiFGxPzYQFZc3T
eTaA+BZ0G7yFe6yTJeeoFN6uQTK0V1jMd0froxtUkbIPMfcYoWTE+4ZkZeyIZdx/
OyMOxdWdtjTLklc4em9AkW5quzAN3LNMANQVC05bMthxuwBM9IIVo5DhlD++Sczv
U5g2IHs3ljhE04Shzv0hZIV/Un8SN1VZNz2cM42X5Y6QRDd1e+PEDxbJz9aCfIfe
2ixJthMcFVwNARzxjpHhXwlk4MEdOPQ81RIGaQPVqajtTMQNgQ7mnOx7G7m4wR4i
IZpVn6oRRBk7uKdFskEY7h0Fj90Vv6U3Q0PY0X16h0fMCn/HbIn8xbshBfL92n+A
EcIA7lNQ5ChAhfG8M6ypnIFnbM7mNUwDnNk8slX+pIlpNpab3Tgro0wgMAg+/EXi
JbLReenpFz3cF88qF8uFuoABhRCvH3qgoO8cXlTI9ijfXANfG3vM5pbsFW76f2LN
TUJ706aj3rit19LY7TnT5sfqgYWMGMN9lVgRclq1U4QLmKCCsEhPcwmYU4PbI4nw
69EogzmbJO4SNkM89IyRvnoD8g6Id4W1etrOOl8aeKXbCAXP7+ckxT38ZSyHXulC
XJrxFlbUJbsjjJ81p9CEc+tQ7X5yRbT/9Vrt0edICta/mUt4XoZGnY4u8/5H3ZaF
Dk1+qMCXk+/rIIE45K6rxmgLjBAKSV7NUOkIGPgwAw+C/x5Y6DPHmLZem/YMxmO6
QmkM7i+4LfjO30e6ymYVgLgATZAd+WpZq5ZLFolaL2NNuux0zSboJbXUs716YOfS
XieSSjKKNDObyhvZTU67PuxNZhS5scyD/6q930mxLHVQyqeEpFcymAAH5DqBoQTC
QKT5xEWBTa6A8CHOw04ud5kdsX4PCDbZEJWY/o5e1O7UM6VO5RRWWrob3u6Fud+R
Ycsja2urXptO3/lR7PNwRr8R95gcdqhEWvMU/8qSBmCGnkWQ0rpZVS9NJHfui4m7
oYn5mxVeb32E6S9wi0W/Vmo0/Ae2LUyt+vXjOL26sOcyxYqOEaY7rpvGz6iaLDtQ
Hxz7nyZfh2u48FMYID221OalZ4OIzUzzo0LfHakPDDVMj/yV+Aprp892+2fkz1MC
vEo6qZHuYrkpw8dGGsNHd5vg2S+HavfyKXp9kWQwmWsA1nfFSsNa1hgkT8sBN6AZ
ar0LQ/DY3FYS37ScR+B5+UopbcKxgB5ssJN5MRGAaOIyllPSCottSaHGofOehhX/
8qTJh4EtA8+OmV4WcZyuRrtwSbO1M7YVdSg5PCYHfCmtsDssLV09i+PncNLMKtlW
0nBr9pI7atPCjdofyrJxd/9cynOE6Cz65LZb5rVYlXMqRRJN8J/ENGxZUrDiOEzC
CE6lPK6iFAaty2q/Wq55XQvsJUp8yUfMoS9DTLeRuocjiO8B1qZhRfH3YYHDFAeQ
MLUYGgctJFnxXXZ4B6IEojK+YteFm3p7v6d2TRlji5JGCWSbZfiu8bwHdYULRUao
j855PfJprvBCzteUYNwF0NFZI0FnwcJoIKnlR75hx9fJlgg6uErzuz4mo6U36/fA
nomEd1AmRqUTc02SjITOZiNTM2qeJ+cyATjXe4S3M6TSaU8J7N5AMRUQ6ZMGWarT
okWR3SpQL/8V9CXc6FjiYK9LRISXiJxaC1ei9IPXsUmySQ5+AZjcihUYsQ4ocA/a
yESf96sJKy+EYVThY7e3bbbvsmFpaS508F892d8XNmvJ/H/6ghHxYTzFM5OzMDR7
eNDi1aAPFdrec1CVeZSijMw3EiH+XKFG41R2fQES0gabbI6OB5RGeuNHhyFUdR3K
NLQE+Zqy76UKO6ktFVdMi2Xhd0hUPHXsrTZoRCMcB6DYMiN0L6yRb01TMhT0oaE/
DcvnNKXOWHaYk+C4/T2xuFZ5pYePw1JXns24BALsWPseH/YmxZmmoBIc8vHFm/W8
48Ks2aUfMpvBdMVG1XAGCq1VUR2Cz+D5omBwGsNDmPiZM90kCtLzz8Wb89leCJ6/
lmlw63O/SAlrFRlLlsWbEIxh9lAZEtYAvC73cw730MqbpluKxeGFuDCUy+F7auGt
LZFMk93WqkWggHeusuCkAOn5+bjdpOCwUeQm+3jdIKYoEokLd3CFRSiu9HBXz2/K
X9uSvuc6HHPy2n7GDNRIbpib8ujUV0bVO5lNnFqZCkoVqLvsZjKOyHMkMSV1V9Rq
rG7XUuDm9iQ+5XESgHV9GdQbzS6YT68XqYn8zWz2Eq+uSubnkYjEhR15AN+BOITB
EazCzMDpsxi0NsAC4Zwii5IOdJyT1i+nFMsfkwzdB4VP7D5kuiBBJXqxy2TnWogX
5xuCcSh2FV2nrOCXXqCjAElk0Vf0iLUaJ+yiyntdGUUWLSuU0WEbKYrLB4j/dx+x
Y6ecD6uCvrtNlMa3LgAh8+HuXDli4bpxDs80OpBV1vA52x8oxsv0dcxBhRt2qTpr
YojEcN2oRnYzwXd8ISvhlkxcVa8fZ7DU80wwY8n0SsnncynKuwTio4XjQDY9aH91
5/JZIj0hCCwhl/p1FkQseh4XGTeL7dwQKjiy5hL4z9CWFDiJyllxZL/Cxu9GK7du
wLasbdEd/LyBs8PVbJayK71akbmFLfYKhy4ptlco58495pDmW2mDYuUPok0BX0P5
CB4Pap7aYkdvp3XMwSc7HQdcyPi9bdkEO0eDtRK/0cHkTpDa0tWc0xKBpf3CQLfp
yPS68Hn2u/MLu7VSqnsmS9f7FqPyEq4/eDIMeaN7/ffLnja3wUp8tf7Ap63+Nh/i
vMKqEbYbduygIPmLuzaQheJU03sRDZCiQvRow16LzmQlB9dHYAjTDXlFZ79SM7Nk
Z6MSx+2KBVM+MPKD9/mRbJg8a7Y/kHyIRQTr8wGvPQ3gtqVw0rQxS8qd+ZsNFncn
8zGIVPEbAN8h5pVFQfD2H8+R6x6WqN4QYJjYzdLtkR1TNp8nqltC5EV7xk+6Id/M
wa2fujHRBeR8hZh/Cco3wqZ0/G9MqPWulO4jhFdoiF38h9EgCm2qrFJsomj8eNAG
P/wlXy1/b+czc542JKriTbe+TY0NvBd/PRPd23geDFTwdfHDp7aYHJHze9tukkGi
M5smn4KWDRLzqT2JRlJ5bskmtPhu53ToK/v6Ufgs6BGaKIGDJ9bNxPifMlbXaM9u
DyE5x5/QtxJndikDDFUjl9/kskla2OepVPdKpxocmjNK+IWOYGZv/HpACZSc5G9C
8P1lWpXjSDEtHRdCTGqxt5KtOZ/iL6nEE4hb7+CV8G8e/K9QYZTa9dwRfikwMfa+
ZDg6TdMThb+HmjPDehHxKp5sCdoDYqrrVJqEYsGN55IxSZ1grC3mxtG2MZX7R+ko
a2F+yjl4OnSYnZnb/BvPtOv11wjx7YxRaHvHHn+nvytRq+Ip4uEfo3dGw47bMmlh
/3Y7C8AKkkfGW3NWtdGXPkglYsPusmN5m7C6sn/f0w2azVVbQPfqOUoeqh7HRwZA
YbEW5KRgce7lVcFjT4uQvokI5M52P3lGAF4UIdx50mbw2gHH7ai2/v4rwuoDh+dg
ttWqKeEzXaBVo+dLA4xQht+7VISo+xrZCHqtcwFWJrVIYcDdZUJ2KTM9q1F6fXZv
7qtz4+feY3Wl74Pi5Lw2uvrTK7pG9PmW2vVYeHgtDS+Y5uyrA5RvRqVXFBZIjIji
4qVEZu5tfqZH/bq5SjC9YAe/kiTTxwK50qWd2ufjdDTt+MX8TP88pb9oh3A1g7Jr
cCkZSXQrOOOGwNUbaytCPeU8hv0X6Uc9iddqx1gCpZq3o6xX9VYbxZt9U2d6rneP
qAb2QpPk7m9b6swrKf8CSrpfBONQhZX4Ex9obyrPU9OVVDW/AbtPYRk43kFmG5gT
zMJnTteR7Yz2BAPY9t38K8fwaezxkGWuF+kuac4BSDwWM4sd8KoZOks4qfTYHO5G
E+E6KxxZ3PJvHZYDq0YoC4wOTKyFfRYdTadqSaBBrW2xaLSLv3MWxFW3tgcLBsij
XKbJeEwcTWGSLBVD2xLymFdltGmxQR4MOZXBUNB+3EaFLFS5bVKLwu5cuRTQJSo3
8K/HgLUw2+KnuboGDMOLoCgQwlidqGA50SvADcbBg9aXH3cjuePkgyKYpw0Ld6IF
jCSHseAPfIAHGisurOj9QXdAn2ac3EvNVRncniu6v1xy0iBLhj1+cA8GOb7tOK+a
+h23MO3H/j66EPqjO9hQlLt/U8X6ggF8PZES6kIyA83v/oviL60Hm7t9GGevbVMh
GgZ4hD+iPIngoXTGBfrSyr8JvlXKStP8wa9zCSyhAC/dVPE0q/Edd5JzxW3f5bY1
6EWTkqVZmzvYQaOrzFANgt49poKjhqCixoWGyCZaVQ5DoHbnSndKNGG4vEPgkZyx
AFArzSEcEHAmeKdor7fJjzvVY+jShJOhb2zbxmAzSyKQPsoiwFMszxobiP5d0nUA
xAxOzK4B9h28odmsaHzBMK1rz+KwqRzoO5Q+a5JY/wnghRD7Ce9tbqF5K98EZVhp
N/jM7GccRhr/xg6VOj+rDTbw2dbh7Q3YSDMs8ek0x7z7j1rHIA4r4sA18Xg/5GPk
R0Qj9dupVUOTAvoH8/azB8aUaov67dYAklUccP4lWgD/ZSGRYG4pn+Y65eDcq7Ma
V0Mxa1C6VnxSiyupnVYDmZHSXOcSY3A65px7XpGL9NZY/+v4mOgxcQkbONRKNv03
1tEWlIbNgPBiY22kRZ1icYAvOE7WJKAMPrx80iPy5wcvk3g3dxiDAXmW3c7qO2QC
JdyOn18ASwF9mDOKBs1It1iNtuoY0LBuOpVpGmwIrORpNdA+22umUIgae1kIwJiS
hYSkVU7BdUcpCYi1w8WfmTXf3jfszRHcI381Y9T6ocKEntwAQANWo8jMKzPWOWEn
WsofSypf4uuhi6/8gMqb2v4ojTOKFdihUtXzelLBIsih849fcHXJ16THtuxMZ45I
u5+xOdX4WPuiJOJH2vfh33wt5dqQRE/MrgRdBZapbCsNFKsNhBeviRihqzF+vsqr
owortLcMFvd1XPLsTWBpyrXC8nUc5kKAVUcduspuH6KJJOdMx8U3T6fT+FSn0nEV
hldFtk+qHyHR4W9kczsRzDrEn3VCP96NaUed5bNieGWrbJ2NoZR/sHGRmYUQojt/
7K8j3rgoXW7t1R2k2PBmIouj+ZllZh3RuQrChOIpT57umyvOGqHmy1KSaawlWDk8
+jcxvjAF5d1ZLzK/j3DOn+Jos0GVWwX6lHt3kTEKhlwTWjuuIHdOfwORXsO2lEz0
BLg2fLd/owwZskoWlYEAKKMNOu58YsFtr/YmUoxRyJTiNGK51sNBNb4ErEkUyHOt
/22utVmVnncBhUA9SXk3aFzfYG5H2LLXflYvunU8suxGWbIuto9W1/9Yw1Vyq1PE
BNH3GJX85wf/7oH5gyT9K3NObYX30gRReItbOXd2yhGCKKAJdVdYVSHwzycJxYS2
S2CN3x6aJ7ByEy+Pp8GEAQiKZC8tzJrH7imPZ64/UT/1kIPojWPksjFQNr2aRDS5
eBvZ4Co/tRaGE7lZlHbrk6K55J4c7PRY5P85+vHiedfGVG/oVjcj0OjsPylLYX4M
VBB9S2h4u1F2HWfP05dXpeP5k8C49XBlF9sRwRa/r8PofDVV1S0eil4r5yHE4usc
OUhxwNDo2dc3KYzbY/tK8JBYFtBn2KZBRTQ24JcS3Q9x4+7exzNblB0ng3QbvFck
YhzNCymG6L8Q2Pkb2Aug0kI4Oh+Wj2/s9G75c25Zp3wu3QDtsHA5z1TIVDsCm5jL
3MNWxbTUSmNhnB6S0JgUt1ZUbzoHov/f2nsLDDtZfxJnP14686yY3zQsGO8gcJbX
CME83lWFrSmqelMzh8+LpwmxRRvAhpRWVf8LE9GwX27EXMfNeGg7zoqRE8P89bg5
yLQwW2rtuZqWHvdH9qGtMYOa41tm5DZXP2nFThHmKfxs7kPz+5qbYGbS2DkAnrDG
7t/B/HZSjAY0VyfX5ng8aHTOjHJjlFMExJtPRrJkdGBVruGeK8pvRCHsSpmaBbQS
QVxu+bipRdcHBFfoytUZ0qOQf73pU2FSAcg8LzW5b7Yd0e/5ljd6ayO7oq1UpRNe
i0gYiLGtNL60K7Hv3lQqansodjCuwwm8bM3awvnAmoLogRS+9e2eUkNALADPgD1q
rTInhqpCfW6DFVLPnjgeCmnzliblzCICAlRe4s7QqC5XIqvfpMpSI52dogvAm/B+
70QVOKLS4k0I+w26pLkJroy/Tr7VVelM/Sfxptm5wO4XjtY9K+YzPdOab6sJzcbL
dP8z3yKU+Lo0fupaR6NpONwBLVt3V0m5JRmrB82CnjHbr3SxC8AG3EmG9fTxluy5
I040t5AdGWs/9nmd6811jyW1wFC+TTNJ3/81bSz3GKkhdLiB2gMYQo/RFavbQfxg
7DLz9gyYFRLlQUQzPXgpyE1McpxOfu3GOhaFYdqn0ggsqZxl2nlCR3xlVq16C2UM
6boR8faX/HVzPyxRTJF7wh+CNxVU2KgTSZhwmE2jZv55dv5D89/Se5mg1dMsvwWk
e0IjAMzYeqVowvKMKzI7g0eVaGR7FGUU6XeBXCRdIdAHzL4s6z0roS8mkV8H8jiQ
pgEtGEQEnM/HHVIqVcrnGeJ8kluo5bDrPhMH4SjplmUBl1tjti1pnJeqGCCBeytT
YndiRSXh+of9JZkldsSIFBWRdeiF16H8AD4ogs0VEAzxqKhSBog010/iDXDmav9w
qVGjAOo3y3qUocTVul7eLOGz1gZ/7yydI0ubm+BA9miZgvd+XyojJPSIESTqWFXi
T5ds8c0EAZPsmyd3Tc7X7oCalM9Zg9/bB1tjm0sfj+a5E/TdS0kwqWbWCNi0hGJF
RPsA63dnf0iuff2w/v+UmVV8V+RsOMxzJZDs4muT97FpfoB10QOPdy854pYO9Hvf
9SCnO7hg541oxjQk7p8OXu6bZ9dPWcECRfyOtiuntqy1z6xsoLqzVpSpxz8zaWFu
oiYAwV+hLBsG/A5sjtNNv3kxWime5e236Wsej6VXRCY45O5MOY1K4nTKGw2RriU5
rX75irjwsjEYx9ILA1g/AiJdKOcIfyUZ77n0rj1CIlzrhynsJjO0ehKwAvnZLYkz
5XbYqnzeWKmonk+hR17GraNnC6vgEVvi1Fh3Lm95TamSOfxiNtbXFrhYqVVodbKb
awloc3b/RslHZKCTXdM/Z5G/Ge2aRg8u2g+GOpx4UL7ogdtKXqpGnD5FS1T29eI2
qijo6eCtdaRTALnnTYOStkipzaEhiftiW1QSxUfcyY+/7uvdCAw6XmII04kO5Gjq
KDIbUrDFtWR17DehYA1/2SzjhXuF8XiuEeLtWvnOuBahJhw6g/6CvYoF+NFLzKj/
QTuRGoizEixb13CjJlxbToELAnIxZdFdJ1gISuOTUiHXqt/kVdQgXPwA7XJShxxy
exzqfer1sGPcZasQX1UP/oVYefNlCgEg/mPen+ByfMq+zZ4fLXc4ZpHA/UzTT0Fb
rTx4jOHI0jICXsZCpiQHZS5K3gGTPchHBSIfSBa+s3rp6/xXITKph1ooLN4GnhYA
nT28XVfTeh6tkjTkSgbT86CYM2GPKiTXdnh1eraRTqC0dv3ZAvTXDWGTj/AhLhVp
gUHZjomblCEfnms8DyV/10irzfELRKG33OryPz4c4evVrxVmm8O8k70c1UmB14Y3
Z8g4D7gttvmImw66R6/17w7TSRHNyLNUIhn2B3Zh/1Wt661kzQd5O+/IfD4lKBhw
8ZflLXGV8TUbT9DLpp3eJW+sYyRZJCiFZiVyhvPeURxhpHspSbCnHK6yuAJGf80b
fOQZaANobAvvA/7aa+D/QLLDRC/JXx2RPyjcwa712R+P35HbRxmqBc5i1Ir0yswL
EHLBykoIgfqju7RyTLk91zs2lXD80dXFyeyr40t32OOhiy/s0PmNTifSUX3Clgbd
SDbpbHssGLXpNamfScz95X9d/CJp5DdjrQq1zDPW5aLuJueeO85+G4xMTUHtDjt0
dWVQEdncaqxaWQ/BoX5CvQt0GsnLPREAtpbCayYEmuW7nhR2LHMKgyq/HdyrH4aB
J/0LwfPiMVx5t+kjX1ue6l5qVxaJNXiWrXBKIn/rfPb63js2j1dqF1P13tpXskmO
JUTtyoSFemOZX1KyqMYZpob4git2pSVfcOpxVSI061pteQCG07Ny+p937YADic2T
O12lTxKyg3Njux9fZPc+DOVoJj41TEK4OzhZyn092fJncLrULHINaqChTEnLeNqp
8GatMo2MkHe+rFj/+C0GK/U51H0Bg+L8JzvzeYRQoWF1qUAf4zDwh4eIQFtGktAv
c5LmRz9dJdZsq86gdJNm81+udJcLS9MAWmAxqRDpiTcso/Iw0lBm/s8piDOUTsIg
L03yvTzQFkZNZkaWwP1Tc/dtzPKZmEhyao64ZpZIpj9sMrhUW3NRZsvDiMNmFVLo
SXG8INrd69Xd3OdLWefB7HxpAIT+m0v4+I7sIpyl2mDxSKwiF1X2WjlP7+rzSaq2
ISTM/9J0nCitaOJJXLahps1l5Zc1nC7DwtaTfaooF/RERPNOJHl20ebQrVxHTuxY
5Y1dUvSwaL65u7Spm4xyzD52wQq9OI2o8pwroMTlNdP8XgUFqNuE7YXleaSb3bMN
xRSEECDsMf0xITiwF7IpU4tqBlAOHkKkIV9tocraO3KOPbYS4zOxvxthAKz/kdt+
QEOEo/t4Brzgknwk54ZZOjU3Cjosr9+j0GkRBmn3Qa649BqaLIwh1VFc9Zh3sqlQ
1DFp6JoW/uQqEIjbNgXMvF5weVzcIJPG02TabGklpUDawkAibPaZxhnO1G18qRGh
v1FZRgx9kuGsDB8dfwZ/+jcmMn0ZUy1XB90whdKLE2IcA42T7gXOm/MHoBQEjNul
iRP/TNHClhWULBwR8EAcSbssvRGjKsL6qWyJH/Ic/b38Jj12T/5F6IKEk2ghwjpz
3HzFks3zjrhkNq+vaTrInJED0io6URMRPHSgcNBSgSGUxSRNTK0i8WACHVwrI9uL
lwq4wqjUBzsFwIGzReaWI/bKCglVtU0zMP/oh3rraG7b+MbWJdQNpUK9bbTG3O8B
jlyxq+rLX8C02zUiYpAs2mTFQr+M1kHPOpOzpAsPpBKtnpPqFRTKpvjcSxZgYVNW
ETDy4qeJMSdf9U3ue19khvrlS4sxjzb38CJAI/XnRV3bLKV4iXlC/ImGascV9LVW
RpNG0ekRA6UXCjWCohVeXBu6gc7+zVFzhRD/whjVtZ3KGquua4bm1OW+w6FN/4mM
Tbx5C6dS1kwXWmOiIttQxIWhx2gSQIN5Kkaw/vr+2aIe7VEi74iXp8m3y5yoqeOy
OfaVxgcCi8jD28v2/VQnQF5lAr0Qdrt74GVEPj1Cgi9Rix9u3hvFaQXRmzB/t9dX
xJ5xo0AOWZPUYq2IPojGnK9k0ZdD5oQnxskPA4xf6D70fm9ohgoxAPVxR+ArXx5Y
/OJXKjC0MFj8rcXyXxbMSeGz1OMF9BhrLV7/hpLd3DPry5PD2CRBNcJKaY1cncsF
O7PSPOxOn0a3jIfbGKX3kMhnxkAqMMC39P7uuTLkwxw6vgq37AmTtu/U50gZpNtk
BqV+6KggNwFulfXTTgYBlmq8Cz1IOo8sKRtWFOTJccg015ASZLlo+9yzC9XEOZNw
NlrDxgHSnDGa1CZsgaM4zwV4A3gJ5mqgwENNAjsq/1TRDA/nPG49ipyMrsfVgWE8
wnDXIWnaQincrYiT+F1MFhRbkBhmuKkgpj6twbQlZgFGs9GcXxQuAOiz29ybpNpR
GhXWtYUdhm1mUgxXgHspKFOXVApXzpY94IonR9vx/QJOd89RaeX5OyCC2qGaLJiA
Ly8aKGRTCjqhVknuj9cS0NJLT/r3dwpj79VPVgxJDfocNMTmVcMQqEfMDvr3j+2S
GSRXwjbYRh5ZDN1Z09Slx6vOdYZ3F/+KorAN+KCxhAPsHVmPk4rXF6eEZ0AV1RCx
d1l0HgCO3YW+htrvK4fQ2ltCs7wnPtSBvVki3P6v9yCBtR1+URj++zAms3CspnNQ
4y42ON0f+6DIEmrqeklvEna+cMViCqxGbSywh9MXpdsx6DgJvHtRECCoj7DNpbKR
xWROOhwxdmWlaTJfnsDEi9VFHLyWGR2LIcR+kqU8Gl+VJQr7xOGVEjQsKRUHNiRB
NdA/iqQp+8J09voKjgPbB/5R2h/8bTuhcAWaVID784do8j7cniCCeIqpuxBAvfG6
mTZuX2eLEZv8MxxQ3C7MsUbogCu/tSrwOTvVXOILiPUI+oBJegMypiOL7JLMwh3I
sfrNv04xVfP4YEZbwxnHNhfAhOx9slvLE8T375noRae01umKu+KMH2LxwROT/b7D
23NkK8s8MiLXcmgeY/YQv7tfM2BE0vN2Iip8lZTmUr9CcJMtoCVNSNgHn7iH8xqW
Z4yCWc5PLAkGpRZ/SZpxr8S7Je9eE22DTKCNCCX5ysUMi5tI8E5ONqhbHOGIGATx
rglUHXV7uzUoxg4jL7V3gPrzKHNp3cD813ePQhzWWQMIw7zOP+4YlI/wSlqC4XVM
HVYBYURfkg0Pzga8XkZvk0pfHPTcRCsub62OWWzzm9IcZMzcrNQaoTn0L1DaKZwn
pmjmCTJvlU8BjgaVEGK4y0DrDUZe9qLSGq4gt5+o1yx3lm4Ys1JZ0Hgqt4nheruR
FH5Q+md15b/YafsvFgC7cjL1GUvz/SR1c4rXblOXVOqUK1FZb4SJBZhIypBiewe3
irDi9Xin+fTWAHQ/nMxislGejKk2ql9UnEjFBjRzYKrgPE38xrUKo1S7HtsLYXfH
CP3C1pesDTHIYelekYq59iqEtmjNCTa7oH+GbrQ68HJzcy3QJQksdO/rb70ziQmE
6NeQ8AFZ8+WHcp7UxVAmOHw2WfWjV+qHtba12Hhyqo6Y1wdphfTinzM6p45Kkbcs
NrdNfNLIdSLdxZqwAmI4r3XZJg/V+EYJjz1upjgwGoueQiH3ODqRGNCWpJYba65Y
eZMav/Iz9EMOn9mdCmI6JGh6Az1P3ezICqFpdMzfMY5aIntsEwVuQCTMQ6uo4l/Y
FqSPI5oWxZShzZh1AL3tn6npBZqOplxeCf6isVe5TBZHyPx7izsb7ERoKsEmiZ8F
ERmli8A+5Gav5s2W/+jDd4V1SFK5NfyTYdoMHi74yU0aEKaZdGcJNTKa0Bc1BkhG
O30FfM1X/+tkd0vQSLj/gXdLiaJSXGWco9dpdh8+i9RgyGyR6WgH7fptoehZ8vyy
W15L8J7eYKbJ5qbVqGirIMsvlZ4OK5IVoBlzhVVmM1pgLqo+7A6IUES8ySWbiI1Q
asnMhoFnzWXyAuFrAOIcQazLK0+NLDL3cnjWEAAw+g0/7K5NBXZC4LfA8E6ikRP0
I5UD42/ZU5YfiSdQspKsAP7xVp6b1WenqBji4ERDdj4bCqwGbNSYYO1cLL1x+2bR
fFDj9r++PM6TYHGdGdid5iGI4MYcqqnF01AQiXb2fMunKVXiyOc5/D15tbD8M6PE
6ltv3eFFhUnMerB0z1zWwGXdxgBSpbeydpmZ8XbsWyotiKw805FYOEXa2AU0RssW
IEopE+g/eARbj1PHocELMvphr7KmsITiqR2L9bB6R3CAWh509knEn3WPmnnbmDuB
cs/f2kPz3NjS+b/I1OCvlzeVqvgv5uZKA+U2AK4XlY3nokC7Pqav2asCF90Ub4l0
0MEu4ZMemRtsIMRvoZm18nLW3saCw7zS/0y1xUvTXuqbdZ9w/zF9xuYOxcJziqrN
wUa70mLbMbIhJGT4hWd3ECB+hU4I7g9DwAlooMrhXXihh40tW9zzNSWCaBxfZTVQ
F6ubblaSykvCSRR8GdqnN8fm3WUTwPL9Vr4aKd/v3RJpz2NK3N0owYuI73blQ2w+
wNHyHG/FSF/1iurSbm6Wm37hP5qt78m4L1VMSyBDJRi+s/B95wfM/qFBS1/6tnGg
Sc01V5pBS0uj6vuEYbOvM1fMVjoVuriSLACukXKLtw2zfSUTX37PvLkJlvB3AWBK
qcTwMTv5TrYWMTxqSndcF8KjUYM807RrEemdw/XDhwy0yL/44N8SOjREKlFeunp7
ddX97vHP+626fDvopkDy0sjbG2mhvCLzHv8Wx+vMhqo+QeJAXU69qqrW0egCfLhP
ybp6+fqkB5ILmJdNKUwgG2TdXemaI/CT8K2hBnw3mL9IAeAufu3996WtHlOz0Iwe
FP1j/fDLO+djOkYeSgXwwgxQV0ERPSzZNJwiSp+kK51XrbBiHbY9y58BdyYx3gSY
8cHVisRp94lnP/Cu4q/oh73PqnuE+UE8NRY+LM94xaqe6RRwVRbuKBvbTvoIbA+S
vtpYuEX61uZcurlf+fTJjJc1NEI4+2GJC8msFaMEP4/1fez1E/IvCl3kHrItbIs0
4OatRFkwg9cig3MCFIeUmfnJKgr7TeR2F47pRoEnibt4O5QF/I0cSTPOCr3mu84Y
zqJQVuAsyXJgWZN+g8xc1pkK+CUhsBgj3Hx88nZAummB+JHml4/cHWuQV5IkJPHX
hHKsDZMmoA9MxhawxPjLf2S7iefIJ7qf5KkFpSKU+4yMapf9JfEcREefGONn4mWd
2UdVtbXkvx2w5AzwH9roDc5cAkZp/fgxC+fbyFpe+uCgXmha0lI46tMNYe8A9qOC
l0giCopYayHc9E+tzs+i9XzLCmEe/hqRNZvrz8qDOrM9Bfm2+U/fm4ykGWLzsgIn
Ydid1wf6rB9hW3JOcstBrce2zuxoeH+rQjAUUbrSdLQiMlUfwdkS3zAbWLH1g9f9
4hMPCc1CyWp5hXO1aJIRdwhfoLGivObtUOlZIaWNX1p5FzuLJjqCXIigi8cViseZ
zaG+yHr7JYpUi3JUZUIJbx7QM4PqqBhkUELQXpySXJEr3tvzsxbnhQdHwdDO9wxd
Qkw7RM2cOn704inZJjFgNnltppvU3jybt6OtfFaqUziF2wgje3nXE3MwvjtGOhpe
jXnuIxL2a8kjzsa1UQvD22NI15yRGjW8+lzRB4pZ3FElJ5gGCwzvvu+k9zOad6rv
UtB7M2t7i8EqKvxab2Hy7g0CyFKty3vh8rEMLYYHLhI/kVTAN5VgzjV2ryeXTPtj
SCHm/ce2Ds5/iRSP/S08XIuKEj1fQZ8ozSFhQUpuj4YgSF4kbkCdpMRHWNgDHA09
D6swvWAD74IQ+hYUxlRkAfE++/JTOf5YjNH4E9m3jcl73hA5bW8fTWdyvAwQOJd6
81uhwc5A077KQytc7knL1+Hsmk5p/kyc/55iHjxV5CkjFEspHo3ddwh2kwtoRXZB
LjCmWvCgeuXwTqrxVtstA0XOO1PRspLUeG3if/OAJ3WZX4tfCbxILFOn48Qx4DJc
tTbBJ9hdP/pHQE0/6/pUhoWy+rQOaRCByZwMY2aRjBz6ey90s4kUVa+wfdFK6Gd8
k8q5t0pqGKo5nY1q0gOTpIJVIuI8BlRSXvaSntQs7hFUdwqAzb8lbDuUVgWO6Bid
7vorAmlTKcnNf13aQHNPjJnlgl6bkD/XIIOF3WY9QnsZgZG/9bSMCWnQEcZVFhMk
/Nh6cY2OhmPzoTB8VRQvmzOqgLjXxO/qJrI21bPIAasLCNuMHbnzTWf4m7cF2yaB
lKocPR3ELpO3DqTcq+GdYex7aWihLTczdT1OI80026o7kW+jdWBdQqVndpdf4F2F
Qz4rFyF1xGEOHX9QcVKfym//MKmak10e2bfqFpMDGuYs3RPGd6gOZckAi439ZAXL
/9E79iCpdiOUxKg7zyHHleH4DCRz4wjR9Y4IMaIw/WOJvsUxChSXGjAwyKTYIqG1
n0TsC42jRvz3UsD6ESoZ/vKaRD1GYB4pAh0MA7T/+3TB3sRPZUWr2r8a6cpu+QSD
DQEm1+2/lIAVH/+Ri2TL8irn6Idb+n/CADvmr8xlEfFuoRERZ9dDmc7gRiG1puGr
GIPFgM+v40QlC2Ag/k4vWoVbdoSm3+y2EMxZj4xQ3NgjJgmly+Ji2QlQhX7DkIAo
fA6a6+mtX7zGyV5iKiS7jcMsIidD594FDPIAapeWXwTSqEeh9b4Kex6XKKCLg1j8
vgFqBj1OHZfKlJoW3aLIVmS+ie/s6tFY1NQagOLsH/njvkItTP5IBHNkrNR0uCTh
P+gPFcJi637K+ZhrBfvah5IW+rFkz2ASXfqJJoG8d5+i5D7ajrrpgb83upEVhHtu
5OyrJ2Hqp4fV/5Z/DQkJprb5B7c72dTQS6eYSP2lLYxsEsBKEIPd4r1NrZud3TYb
WfS5j4E+9LMFuyKZb3W4zTwEeE31oHtQeyNs3WrtSA570Bagmy1aoFEoIWaBEGOl
TVtwvya13EIRgMvHySyxf7bovAYSd+XIJUiD78+lBDcXI26+DOfbbMjnBfZSiTDS
0/I1VKJXujb7vYFPMphKkbwSYGjAn75X+KEu4sxugEYu5jrxH5q5uWYEVMQG0kM3
l4w7J19pKNOm0R94ObCUPLxUZveYK6C/JMIDaJwTQHxYC1Ljk2pp778z+oZ31bHX
I9bd2Ylz6gdU+gHkBfqubreZapv4nzhXfXkud+sSz/vy1tKizn+57vh6LgKX90MV
dgW5SmwEZdd2X5DuTYRdhAA+hSeZkfYIW/1nPvHiTlWCd4ex+mszUb8qHFjp4mIP
KTs7hngZYCjYQsvpzBqjt8K7gHJ37JJz4RkojPmUdaAIcid7uyGUN/a5dmIKs6pY
5xtB0Yor6Q/r0JEDNDsGpz0YjNVxpWara+HVClgTi8C/831zyux8vzFpgUkazxk+
dWR6HnhLmNsY+2LN03L1VccKWYQ48bihzDGBkpuVixzbyfYBaFPwYjuDqCXaq4X1
vEJOpnFlvBGn59MlP/nEVA/N3tMHLlNU9F7T1DcHmOOMe0GRHBL7sOEISDAdJkEj
OH3zH/8vd3e9j3xujWmhIl9iM57MChXZhnrNNrJk/7/By8Tg+lWosJYRjSRSjNXL
0KL0f658nOCe2LdPR4f38lociwKijL0zbiPymR8vIQrdd/F1K+n6JYEjray9kCdm
LIorLYFmC/L0rnMWXtBj8D54PCiUYe/pFsP3kzS97hbNbfCEgIwEnGKlwfNQur/o
fvgUTkXyNDeuT/lMN7bLYszOkPeQal/CGizWQxBpAQJ63vzS+RyVaNooGKmBuLT/
9YErJ2Ded1FT2ZKaQF/EigzTvqgmPIo/sVpQWPWMwCRbe4vDhOgy4FkKMrBZ1AsA
4JWH3Uq+d+z1BBpIkKACcQax5ZpxDFp9ItLNoJ3KnjesVQ37d57K0yDkHqhF7m2J
Dr7/wPrK/4Z121G2vStI8Alp4/5ikDFKyXDXs038qqekkopgtWzUQ4ZRKBv5I6lQ
pSUzL3lprHNy20IESiKNv7yiUCb5kZK9hi5zHrj8orchlSQ2e8YG+0+CAvyqs12J
gay09baNaeEF/s0Xi5SuZtEZaeHf4Da7WLh/A3PgH8FDbFPE2HDT4toObgf5/hv7
pi9lf1aebUgZpb/Zvq9tZcoLuTH61nTDMBxOYL2bcBrMdOjkfjIhNAa75iFmXCCw
S0SXbj2koPvtCaP2bYR3VC1+GlafFEhJnkDRTG+NOIgn0BdRSzKDvioKVxeujStl
UJhhg8pK6YKlSGOufeXB73bfFiGBX1slRvn1NXPqpQ3XpIfzc38ie5cMFZ9wqKnN
OWVmf7eT8qjdADPk2hL0d0kYkrhoRpU94TGX81M5i+DI4LUKMgtwNUO0G5cNuDNx
WeYaWm047mYlj4JQtLUkRRnnt06rOFRKRJz7+D+lFtZvYD6go5bOfLtxnLAZPsHE
0t2rVx/OpfgwSKPBh+zJlpCulcn+0JGua0jJwXs/o9bR1SfJUpr7wwJrSs07Mv/n
2sNVk17KwgvsrUig7duim7V445YIZgRe75q6ZGNNHwL0SjlH3MDhr/DW19h141GV
kunp150RPEeXgqzH+k97zQF0B8W+ighHcactfxoa+3no+PKg7C1JwpV5OZ4DX3BC
4Xg9eoyFE02kTP0cK49kuOhupx/vofG14Z6gQWr2ySojoc9kQTU20diXnCi+jOlk
KzjCVsKoKui85Bxc5HIGJLtwsVliCjYVnyqs5DAYAHIobhFYCwAyNeLKnSs24PNE
4e/ZSeFg3tiKOVgl9MUuDX8uzHjfR1kVT4FrTedOC36aYEJbFoIHTOKJA8OcyT4f
C0rGwlDqns9GwruhYwvospJDSDF7RuSZDo1d99gzra9umfJrSfNAoKv6xVd1NbXI
DAJUVTHCf22SEzqQJu5foxKqLoO2rWf2AoXez2o4sZfIWXcmZY8Ir5aM4GmZMxvT
zvm9U8M+TU9HuoCJ7Ae32m7k5G7gpUfDi6sN0Z9XKhPOHKc11j2c1LdLLEIvUpCv
LsUCPfCPLLILrvyXLxvXBCEoRXojHpCKNapTtB5OXPKvT93aOto2eyWZ0sayM53h
Zi5n9fMH5gh32Yp6fQ/jHI3YXv2edxr/U0Krm9lolwl/ajxIVpDBxBndSK65uxi3
ajHp8o/wtK4WChPrwAJ6y7MBpIsjtwgVqMUPS5jrUjZ+iuRvGuKv1ETeqwMhJK1F
9yvie8clZt8cpb8nE5ibAuVjgRLQAM/3Nibvg8eHnOf8JkG4J1TtZSVItl44z3yu
Jn4U447qOe7imZfbKq1kAvosgM1V4Vzbqbmb8kU9Cebo+oJVGSJG+XO1lHs4AxTr
AFKUe4M/CtdBbin0hjCzvr1a3V1B76mBVdNsEcR9edEvuNKeJsKN+ymAOAj5+z0e
CsJ0pguqyzhrZyyK56XeJRFJGVGmAO63lHxzh5hb3cEAvUYiW5DWRms/FLkXBs9U
Db4LXT3T1oUI84XCMdCTivvtq2PC2DOIqLAGnBWiqeUI+7d0KURIR0hTVh8GTM8+
GAIWMrIC9Cyu7ngL3GNYuwQNvAV2Klscg8dTZ87krsayr6FFCaAByzkg9K+3Cx3u
iUsp5H7a44Ca5xAIGeQrfS+fQjfz7+97RKj7uThnqQ+lI6gIEbL/H0of4F859t65
w7g52UW/l2X4FKwfw0Mz2Bh4RQl+B1Biq7R2pOvwhVYSY1eDv831+nARcL+aEVrW
Gq85/zhsUQZaUWShC1oC9r0e1kh/eJDf5hWRVSEtnFirHHNENhxMd/qTEaYV5zDU
F5DelCPwfTVxf19frK+TpzDKYOouT5uKfhhXkCq2QtdMaNJYDXRbtjTsvUmafNRc
7Hsm/E9gzk1Vb+oNtoseLFlXyKewWgilLaHm8I/DlhWkZRn3Z9mZ4iDvY1cDtKd1
71h4WtUxia4SIySbTgzZfr1CvID2usVcMgLTTbeijIdu19g0hCXYy4CumP2c/LI/
zqs6tP2WsFDiRLWLVu7mEF38f2e6kT96bUmQJV+FSS3MSC9doCIeBIwLA6PWc16V
ROZ2JdbAWuL06r9THl2JR6HWbW//dI/fkIoApC8NAUSNRnwu/lBEel+I96RNpivz
yzDf6dy0l6brOzDsvHX8kzOiMPHVDAXr/HtbJBDK0P7R16/wyiquPaC+726qJYWQ
8vVLaxINjEkcdt6+0yIgrWrpM9ig32LbkfRNfDIe2o1mulEAQWAKwnKNT8q/qLmw
XL7rPDonZLoH37rlKZigiCBzAFL49eS2eN8VwlIJD69VBUkJB+lJ7UcOUgOk75+e
CVVL1iTbqidKbA6OvmDMBrYMiz8DRe5PMrHB3GW+VwgCsz1Cp4LQ0jvx76gDvlZ2
IHwfJglXtKeoG3YaVFPEYA0/nJlTp+sE3AAcOqOESTVXHoi5YAbJgPNKLYFHxJGb
UWqJ7xMrez88aHC6orCGR+nuUQCX6L7KaUAnBFskFav0/pt7wCja5BQc0LdqI7yo
o3Q58VO2msHmMMNXUfv/4/digEqXm14gOdWrwU5x0FZRisql837fnjMFBi7qVnpw
jDGtcAJIWRwyvkmJdM3LOqjlE1d3RBcxrkGZzxaYYb8T8ayPLl0lmoblyRl0DRIv
j5RqGcFNCfzzfK0ogPPlOYTimYmWwf16a5+bFVWdfQQsuz3fkcZReeF37UnL/SdG
KoIg8V2lHrCq6PaOkuOOWFQGWiOK/cJ+x+CsSc6MR6iNFpy8elOUfKiYkwl+nJCA
01EBM0hmZV1wpC5tE22ann8FjVfEm9bwDKRuFq/A2IYTAGd41yKxzwI0KQ3DwvON
upmD5GEkBfYmXSEy3pHp+GatA/Zlg//cGtWRLDaXV44HgEnMGSRrh7ugO/6Nimfi
i227Xy+kSyoo2myjyBTYh1ULYqAF480UNMI3a9atJunL5k+NUicDxdLI/frRQ4BZ
jaTRpeoq3nYUJhxvvP/oyzuUtBXrjrIzApjg+MdrXsjbBo5lrPZeVPooE5edI89x
AZuk8cYKjHPjEQxVdl65EtFuVAA9UF5Lg1Yv8uAr2W9ZkH/VZnl6kNbAdr5CRPWO
KEze/zqld01rCJwx84tZFzBLyhE/gCzoC6vGLdmrXnPBpjGGDdm+cHs1TFp9+wYI
18+sDH9sCrz+dyyNvfGfhynEFQw5SGm3cHITVDi6e6q4Gafxv8Kkaa5uSDOHEzzH
bhSTPDbN0vfPmNH/H4r618NGiwsEEaepejKOSxefO/2oTSgwXH1WZrXtZ6RG3PcY
od/fswnoK9JpBndrbeqTMIuGkP9gb/nHoXoirwY9b8Rs2+VtZXlqhB6k05rd54n1
LrSpu2OLQ5KsaHvaI/jxB/uJyoSFjucQCQXGHnUkf0xxBux6VSRC4gC92ZLdJbak
QP47pFSoJn0b2kouhZOM7zoZjGeLnIcP0YB76GFLrNS6vYRro8qzdnvhQg8tPPXh
2l/h4RFML2miMRaVTQ+g48udU9JVqDsXRk5zsFUYE4RUnblLfo4e5tgbAS1V1KDG
bUIapnz2GQQy5YGW4pBe2AW2ydA06g0iXlAKKnNjHaoD+rZz6TCdoTyyMk1jP+4v
uvejRnFCKx9lnd8I8yK3VAVQfQlDmc1GHhCTdemAhrz7JtBx20TsDdod1mBxas7D
kVhmWwuHCEm5OSkHF0UpwNdvLuCFANwsanViZ8jgIgchTroFilnjuODw1w8qWGUc
yd1OvXUqEh45p8Mhr3r4oa2qe9n2mILDn6G0jHnz715m1FraCFsl5xozi84wsPjr
DrRxpdSjaVSzyQBS7LZvriD4tsiqd7x4QAsyPu9myf70++FYrrByaGMy2BBYzvDg
nF7gyPxIq/VcifwvdLdI7bW7vHPX0gqsapTS9EiYHU9UC75l5SnMEw6gEF8Q7olo
+0mb5uHRud2dQ1Gf9rGwJiYTXgqm8lQkF5a9iLUGiKVh1JEWWKc6+i1AvfblxpYc
aL/5U/bkhx99dHqbAKAsbDBuFxn3xxg6cryppA6F7AM+dpVhIzKh0NO/Y8yRB7zT
ja/aSbOajFgARDFDgCqiNWLB1C+SvnKVablzH0ZgG3R4VHe1IwsPwyAEWK7ChhI0
6UbDxWptI/XfMQRRTUkqh+9ZHcnDW797jDFUVnjc/ejQFbrmiH/z1DHlYAaF4iES
utoFhu7fruu5pIEZou+iv46aMqpCmThuVTxpClSdox/6klCgl4BbmlcwA3YUAGKR
urklxJCUmLQ2yL4yPkSVRlXnXlWHBUtFaS0KEojDMr15OQh4VtHjjvyHveqb3t4k
GV8TgUIfUsbRDoLwJwSBqANSiDz0nvIx5bkstao9dPu0nRhCjWIz8SkEMsy5y9P/
Dqy3I2Ok4IAweEgcuUrIVsbxiwQRoXkvhjPdszQzFT3nfvP+8i/A59ebBS6B1Jrj
KGRXGEQ6HwZe10yYF+EMJkFUkZ+Fld7Jfw/z8wheoi/5BX5vXnE7/Ag3k7iA8olq
CV7B9cpXNcYyoPpebjpKP2+6qTRru4uCzoliMUU/uBVZqPW0pQD+JFMuG8RH1YiS
ABnbvAV+p+4XnySlVFKTwBYTH99JJ51sD69qc6XadUpeWdD2BCZZ+gJc+DFWJ42k
icDrGIuWxB/uX/ziFfx8suEALu1gzLLZs40S+0eRSdE0mWI+6F56bpy1TqjYdFqB
vhdGzlnqq+WpUxEEdxGXcLOBtCvFJDxIMoADob3x3Qc0rjeB116DPZ20qyOSPNNv
IYo1NlwJJmUKeko6ZMfXusH2kmj1HMqSuhXP/ICA2vPLTTjLV5S6mSQLRkYCpc78
g08sx5YUNNtLL4b/ndGF97Pjo1oglqyC+zSWQwGkTvDJQgUbUZCWro55ANHb98oF
or2UCl8P4dExRGuRcveErNdWr8thBLkD4SigF/RI4xzZHvTKdT3/qh6EoT/d9NDd
mFZLUlJOMkC7kP82dDW5x3WSWBhW+anX2z4ma64cgZcvzNszddzUpWRKz5MW2MBa
S8AWDLQPDd2v/XeTS56mi2ENDaYxdgTf8BAw5GN9FSneRXGgr8hzS/FPxZfDYdIK
GZRH5PKdCucuC3GXQvCf9Lpd9b0NBjBw8q7TnHSDTevC8HuQVUaFm+pPidRp0sFA
q8vCXh3jcI0OCox7K8+XyeU8v0RrgELGFUKH1IR/ULwTAQaq9+AqWv3eMQ95YE1O
H1gA/6Es4pnNFwoJ5mdGrVqC9mVTbeV+/SJ+2thtl+6YB8itgsQ4RvhX7qMldWWt
BRXgAQnqihNJiv+YKlL8FU5dG5UIQlAY/BCHGII/WojtqHIFRMRBbrRyFUoUtbHB
8XFjZEOtfu3oswy4WlDPtktghBy20kiWB7PTicLqwCZFMCWwbMrzd9xo2ifIMowh
JJhVwAgE15ijWnUEMJ8eYLuKAZN89pFWoWOqyXC6QqeoayJO4yU44JRjznMc27/p
56O5WeDyKN+2tlg56+ceIeiqR8llcLm7GD0/uVGxZE7I9iX02Mm9mFckIYqvBMNL
vO0ORKbGayg3ZVQWECQJpw8GtoKSdKenfAU0yvM29YFLsssTlXrb/V6MyGfThtbU
cxAwoT64S2dEV7NabF8VXQYG4lKYbfhaqbOyJnDIr/p7BXffneYJp6AiqpNJgQ8v
i5qDWS22rYJNhoa9v813sueqPwQZ9e1pF0TiMxF3cn+wWGC1IdVfKk/eFkO75Ip0
KnsKROKCa6TCvNVEGPXrX33qprfAWKfrGXoywS1k9S6TLPpT7k38DqHDgxDsWRjI
Maz3DzuvjczDgwnKpe9ZsrarcM51lx5N5wBHMR5ZOi4luHaJ6kwbA7SxCadmrbCR
mbe6HOxJL4wtzoOcFXkMz/NRv4EMy9pu+jdk46qY5HGu8Mn1hRQnrW+2NJ4U5AcN
IcPt227lnfRpkWbHq8hwbPE0SNOSvm4609W5bpLpSD97zrCXqydVIwspBzj59FHY
cphNmVta5zdqnGR8uNvn9iqFTYHIweySK1PMoS/vLndzo29N6Eju98Oc5IPQsXsw
v1tDgVyfOoYJDtVppwV090rO5hJ4+i5DgEbBuiGkIo7Q9ZV4TbXTtf8YiTD7y8gE
DQGt9BdLOtX5yga96WoeBiVdniz0ibzgWJlw9dgiWfJdGpTm9qKvIYPaGCTz1dgv
8cjnr0jPSw7zF+3T7SkPW3x+UID10azZHu7lBPwP58VImUX5zwSrNzg9G/DBNMIL
lABC25FG7rlfxC4vf1x29mrcrd3ZpGMrzSXYb8o9gCP4Q9uJC+HZGQkDpRajBQHc
flCo/s0JdNrgJXF1FdtKfYTi21D8jzAkldmq6V2gndr/bX5tGlzv+vj+3OcacRZO
ty092w5Qb6wKTzNi5ytZiF8rvneUdKvzlSZ5m9J2oqQAVgMLIOEAXma5BEVwAFde
IZsDXHZt7Fq2PWvJ6Mqu5an8tirKOhqMDWDYntMu45abDgHX3fpK7aGlLnXC2AGy
nPtitTodLe+7KfeHBOKPciaA8FpF02s++9/UjxVJ0snzVgrr4dTR7cjwanYts14u
waX8cge2ZfO86I2UVUt0Sp7JbiH9ZF2IiuGpzf/SzAQVfmqe0Po8YcSjp3bqaYnV
kycwGpAt6xCIuEZEDNZZlC5wPCGe88HJliQDQFsQTtCDuZq/UPTq7vERqlMNJlsi
5kDi5dScdufGEfXl+199FUya5zALp4qpctFRJFDBnDKS1wGTP06li+0truJtPWiO
bz2jmPFdHqajtaFMjcbQhiJ0erpDpfMU2lj2dHnswmEq5Rpb1V231yRc6NaAVBjy
g8MysxEbGiRPZa4gvr+8gLpJOPtYRTSB2L+4/jcJxE5LYXupMdKRJaffokem7iYt
3zM/hIKZr6/2NLtEF4VMvRCzKKVDG6Xl7GLRbSE5KZSXXvI5bgrVDPafx8CcJSMA
dNrua80wYm5sbZmBgilHcInl3PbFOQJI96lVWH7qEQzEJEVoQbi3Jf3SjTFMF99D
W6EaHOE/rktz1Z1LHFGwfnToZiTaJpfxBuGgteKK1uQ1NeBy9G6BijlTImUqAMUn
F2Bdwc6XWlMcRLhAIhqAVcqZEJc2/QhiCu0qzB9QjtJ+qBm/fvA+C3Vdwpr7wPEz
fT6YtH9gvs5I029MDVF43rPrgdZkZdP3uR5SYQL3dLKEWQD7c7i4VuryUmBGF2lA
wk21krkv2X3GapdZXdj/CFQO5g4625N/TquOr35MDjp3Mum4FUftBYINOjeQu0yz
kMlrjlt8ICGgx3g6yfUWnwxQyk4QW9OHTIuH7s64CNebv7ybDk0k4Zs99UDg8EqZ
2HQ6xuQ74ZlnRM341aY4gNTAqIRrcBWYk08CXoqfubg1GqMhufarTw7yXaZbeSUh
Lbdl05ZBdS9tuZvB2QpDlOnpUHF/Fhi7JgLvl4q4fdzlSdaOfEUs46a0IrQmo+yu
A5RCljYDbK6KetuUPIAJ1QyllMLE8rSFzBZk2Suis8raU7rHunxGKaYrnWpEpJzx
DoAtPD4kZcbbkmGYGGUKmUj0eCeyC+Meo2J2FBJMBBQeSk6o4BmFrDMXIlWuhfDn
vonP2Q1C9DZHd+GwbT2HiHdE9apNOc0PGux3cir4mP1z0gmPzYLi1GK6+DHL5NZl
ArZUDXBv6UWT5rqyP68ayyRsZw1mlTj+VSlIuX+3UzCCNVw0l8EID/Pcr8Qg1qDF
WqmyqIaBCwY7BdsrPo/qDNA1TdvBuU3ZFuTv3JH7LED1QnTSogyNiA83rv6x0cFu
frWdgC/4Jmr7a7QwBudXzGdIbdKCRMB0fig9Yhb+cYrdQnRzUj4L2DHbuFqqExv+
EGBlVjjY7DNpMOcxaOIYfoc6zFgoKAa1ud71/ZkdkbBpY7udUskCKYFiMJnVyvuL
gtiJKp7dg3wAhF7+3RLP/fEXN8yKU36r9oYJSVlB8jUtI3e/XNheGEzJzG99eXI4
XVsu1YVBZkY/Bv4Yhi1wd9gdcG2Gqst+zjd1sZMjWU+/jrTCSINb8vpYEaG5VGIW
hUqGbyljM4J2EzB48Bbu0aMLTA/veKmquix5S1HelTa92XEwovrSNUnWPFNLS8MN
D4fs8jIB+1jt4V1NHMAAZxX3nKxiwMQphZ3lknPybxinW7TuPHkwQy53ihGl9PZQ
qamGSfcnFIJNKAFN+GZLDPsrLTlSsVEHe98gTE8YZmyNh/Hw48FsWRnXJD2epFuW
wtDkvC+2jbcpdmMGp7MPk7S9wZeoy6goG9OQc8WEBFG9jEf2+/GCS9oEXy0EcreQ
8H0aKB+uesGJXP2hNlz+HrhjJVRTxarbHSlUHGrm2MO3oUaVH9JUoU/udbsWlEqf
MkBwNTKVuIrhO+XdMIIx1kQB0qHNjkWFWqXdQy0S9fCf8jRjX3kA2+KgizJD7q1Z
nxXXmyRgv3NITJ40ryr8BCvOVah6fiFU8+YBmhC7y4tXxye7FeAbJmgxrZHsdvSt
bSF3Ev0ZporaOQAaRBXRY4blTHjBj4ehsx6aqXk1Dw/pCQicOHl/pg90UFNHWjN1
Y4yN6DSjsY2FoJIgb5rVYHn7aJ/ABcati72xTUjvucIu5U2y663HJTcOXZy2K0Gq
GQ4m9T7eJBAZZ1+RqGvzkKGOlJRlELj+J63eBaRDGVKLAlboIS0lAwDIEfoVAYi0
s7gXLy8zDzoDhv9Vt8fcv7R7sYPaDJuwJRhTGk70hHVu8ytirw/paHsD2T/rz6/H
wYwzYf9HS7uwMpHTtuf2zrr2bdEmkoxCQDCILDrfLJiXgAm5UjMmbfdgrI8/zcyc
2d0lVjIU3wmlXtXu3sngjJKME0jGtrPEnXRUYhrqvjSShva47QilzI2eRjyI6UUM
AULZLEL6l6D4SMO9zfvfIgPShdllpTyqPydRclEBjOEkOqWCqwvBugLpRnVFNtG2
X4PqaJbhW1KmJQkQ6VgbiYIevPuZ42eCXOWqzGJ7EHV9dh0S4vV4nW+gV+L7BFsQ
ViBYx3/TJemTVbbSyGnhfRiHTz6rSTZcHEYWu4y8XtorVrItpa8smx2kDINPZgJS
jugcyAw9A+g8pcmmQ6mlFG8kI4EVqeHHDmXvWmdun8Xz5lPE4pGM90fUY6qFSp7r
e5+HI9kXerA63pTBQk7tFuF1tZdFXE893G/lFxy9P3vpztE70H/IEEnt+m5wyy6y
P34h1NuYYNkcREgwL60T7cpPQQD2LJopS4PisooeMq8CjQvLmQal0jtZCdNhUq4Q
HLU2VYbywb5cTueYfy9CF8GtTd7Yju33MCtk4FeVWQ79m2MpeoNVxL1z689w9tY6
bggBI5F7bOw/7OXRNtZ+diU1zU1Rw5zXTnLPQ0TYgzVtOOqgvKboy7ABwMtijIYx
esGhN/kO2LoKaBeD5BpDYJslGncfDDjwPkeCFbXJ2HURrqYE5nSTDPG9oplbh0R6
+w5ucgbqkXxKZJ+wM/So6HWKkousXeqbFew8WxYnNHLXPkpxNYAWTnmgFTTDbXvG
5LN109DWWqE1TMWvFwcBR+U5ePEjnlW5UktvFnKiHvZS4EHZtpRg7qYlfTvD5DHS
Sr2NjknOlhOiXYvVq4FoNI2lA3HPom4lBaUVDlMtok4Vk0nWETPQ6MhONbol/FCI
em9dipx8dJD45o5J/Z3uFjjIPJErspfERbfozikTXKnQaaBI6sKcvLfQktm/S+CU
vt2QBEOXcSiwZgJSub9kQ1p1qHoOFjxdckzctEa5RwaqrLVzpZ4pzClnlaZ938TT
cD57yMnATBFYi+YJJ2/uXhbwEZA6pv5DpbwHqBMjzhyEInAHIdwQIywSNoYDWwqV
+lbaDJyJZFvmE4P7WHEjmM25z/msatLN7clSnRdYGCjyKsiOSgxALjujRXsy1GtG
d3uAv6R3BgTeJPi/G7Cc8CvVG9HBNusvXA1TXWQdzt6REcbzNuiGVcDYVlqdAal1
VtPc5erI8ysS9ekGixvrbzl/a6fI2qIXYkPp1IiTQpLP3j002I6v+NilYMBFqc2I
3iJE9hxgHNNjI3LX2OjNPmkHH7C60Z0s814NstIUpvd1c4LiRXOQx+22TcE5nsHd
9klDQZSTnT4GsFIiXFVN1Ea5m6BQ6Y8EhXx7T1V518QIMjyKwukQcp6iQwtJPJp/
RjUMz/QKFwlBQ5EPSTw4iepE74+gfW8ov0nMQyidWB4VuhrelJzVrCaIDasIQYa7
Wc317c2ewhdFpTwInbBBByQsRv1+cJSMfQsH7O4exVXBzLRx47te6FOCHflvoHBA
7ZVp4ufZCazLK3W8A1kBIrnLicgxj0J0CFmIkDPelpqUEAUCA3K0eixGD0GtDZ8J
plQ5b8TzlPTqMf1v2LlAPu7eWstSXnC9PfgMcuE7KJEUi9+yP7eTN+M3qekIdF8t
FT7dNTQLGLAbkGNOX/FNKZyqTkgcAW1qC37LvKqQCXOrEbHV9WY6SHVeF7qPTz3X
cwoIO0St1O7+2cJWaj/nlWHwv4tkjwF9LvA8VB9TI+0QlfVR8cuO2fEv07yL3X2e
9y8kjp0Y3xbyXICcgzHVDOnwspOIsz8w1jVP0yvXQ8/P5hB9Xct33WraUC9lePov
2UGB100xGYfpdKj6t5A0PwPnSBONbMRAKBgGGo9vRaxI/NIxm61zsFcfWjn+98Vt
h1W7tLMSk+NyeiqZk+lTuGSTsU7b6qdeU2MKQqDoeQEIWBc/v3+zRJ+OJixq9nQm
XAxezI2naTQtfdgBbThIgn1zyh7RV5ASfhrTh52Qq6Vyehsa+Pese0FNvT+6+5KC
+6cy/H5FoaFydNWNCJYaq+l6ofrfbvxN+6RQZbGGrjfXZFKa450PPoSCiDn9s3/7
WSftczt4H/NUFNC0GviByDCdaR9y/lfDV7UexnCUsV8c2QqZIURgopdpgLf3k9tK
iE/lXTWAcrDWt18y9yil2BPPvXT61Aey2UzMyCBHRjnq0DKYDvIxf/1kgMll0hRZ
+nPpuUweO8W+Xa0C9SHxTBsCYMcN3Bg4ZxIKtF92amVTZxk6YOTVWcKefzSbufZF
INLp5kH+3+HOEhEktQ5fWsX2DmHkDvFAcaw+Aemh9251oZHhuau4fEnzClqhDFPV
q25I2532ZQEu4xq+aPKW5SONYAhzJeWhAhE+Cagod86fExBw0b60fvypEl6H4rlS
tXyb9/erClD81vFNx5b8Kov6fv0/DmrBfoTgB2S5TRcXcsEUdwPEilEV7qNckAhb
PgLKQ7b9KwXLXgk5KU1CDrYBUMDEGjEAck30XMzEcIku0FphJMwf2prHkD9qSAKS
G7kn8C1LyTVyefly2ywwftbOiDAq7FPAfUn4PiSeQm1qPIkbRlCkIBHFMXmlmYBf
MgiG99qxlGrVPiz8O7LfS8Q9r2MTsF01k0VTStbq5OoD2L1gnE4OjPN8e79DOIqM
r28uhScruBXP3iMqVduN2zkCOqW9LVCaN6F0hJGkQnZsHrCwp3kA/q/PCT6bg100
PWZQvL3F7IPlF6Qs96JldtzVVK9B27eIrSdbU+dqY6SeJmEShDwDdaNkSgXgqig/
PXlkE9Jh4LWa06FHvBaLcO92wfMj4arycOVn1D32Dra/p1ZHETAkPvqstf/mrQHZ
9BarwDIPIh0aLNhI6qSPRE+qrQYg699yZXFMtHVlLE34LrIN9f05bG+qz0tOG33m
a5HKMmm6dZ0fpOON1m9yxVZ8YS9NjOby4oBaLuNcBC7UjyUXGI1hoAZMWI3czEII
w2F0ZG9Vu7XULeXGBfHaFTTTmQdenycy+uTsNh1XUBIzB7EpItRgZtQ+Lunu8CUb
Nv86yMZnW8+VsUIQE5hCm4s4c6XYyApFseHvMMWkg1jh5EBzhg6p7yuAZnmsCIcg
1pM08dqSeS6yxqUjDlZX6oue+qi5Le66kmfy+sZEPGdS8W2hNRg274/8KKJMvqfI
v8Pgt4WvrrgClFkGc3QU9Ngh5vLDnrfV1om+GPaAWbuKK8xFaxMyQtuxy7bMz92y
fIorOEra/aSaK4Uc+KLY8so0JRwTOx+wC0oLyMrPomKfhIrpSXtHxJCNiYFlF8Zd
Upid9UnlrZThTAycUpMpl2l0idKgKezqmK6QXqOAbOBhlzwOOtKf4ETBJxlWOkK6
yTnse2QZMs04fgNdx6KcacDN71MGRecNySO4FDtX58svp/uAcEofv8zyg8xynT+X
NU9Hy/dXqJXW8yW0semM1ErTvZqILVeHCRWFJl993v0wpZuj9Yj3ewCYMSGAbxiX
/lbqBpefdpSKw0hy6KwAkMil0eKgwR3Wyp7BtVZIbOJU+bGBz1WLo1EYodmycPG7
ZolJ38WW7vwJJtT+iRjYQ/umQOC4x99d70TnVNUvnhHtxiZ5tBccDYHgIPW41ATh
muhzcwzaPA+6e5ZPSaNgMZlfgW41oePMnpG2uPgLKO0lrD2lxy59vyrecn1Tzcti
SmsVWo03LMzT1xhVxYsQYGlTayKEzyiSjKfYKhXTzasZkwlzDPimFzoo+t4T9F6g
Bffil5BDUJFhHsjTDrqbtWD6npVuOWxar/CMYhsYk5T8uq3awL/ZEJYvjzIPEu7f
YPLDvywaZBcRLrLIyiyIBRvHTOJGr5vJpdrGD145yRqVz1eBaSH/94J9ab368qwv
K+FHNEB+Em03KKrAKU/tZJDSazIJ+578tevpaSX4e+LIytB1YZQiIJNXTe+BzgcN
uIiA1oRK3cBMYG6ObQPwdURwkS+HzXagJ1R4is+iMLl7XJKxEv78rNp5Xo4taWi9
bbrSFc6CRN0LcoviAZhPorXQqGYOlfg6Ycqn3WB1tW2u54+eJSlUM+Qaug3jikSK
tB1POGX2mQnkJ5iwUcWT/D3yGWoToD9nnFoGhkIOxCF21M9uDsyAVyUuuEe/XhJ/
W8Uqn1n6iM7unbVbQhzmXgAY/F54e3vDsvk8Al0WF76jXvRFswJkks1xgHrFMEN7
QmzNmBIF9JCCKxZzT/SzHT7RYdSihOqwE7FyCD/PTFbMamnm/9qz5PHkQ7UyYJHs
MUP3jo+unAOb9HOa2mioeUfcV9AK7m+1HGqUpbZNfx3+9IdpCR56bLuZtM8Kw7Mk
4OCwr2tLsVmR+GPnnFr820ajIhpuGubT8rkkhqCPk+xIYoTXCfwi1KMuUBUiMAd2
zaz2ZPKr6yQk1GvxSFNeb+tnnBDndt+GqB0pCBezor/TLbaOV82FyBQZY2V4Vtgu
KrBGIP9ARfBEJ6zEdXPN8PX7GWuCi2Fh6LfwX9mHwEsRl/uajC2Y8L68yy6fsPzk
+Go9UinGEKgFkbU5Fttz8+wDRpDlx8OR2KTtHZ2GolT2AEKh1tEbCEIvuO7v5Umy
74Z374z8ZylY/mzAiqBoGO3uYHuraf1wEfOULDzCxHuyvMNU3q+DQ/SkCzQixaDy
nWXsLFaPWNOGzkEMQHnPpqYoNQNSFcydzdGlo2QRN+kCq62fPYQPDyLboKVY6h2c
AI3g4S5Kebxc6YuQ10d9UMTkNHvJCEcIjD0rx7Fnlc0mpwmPrm7+W16T86NGlJc5
dhyAUJEydX8c7bDF+nhOoWWG1CLfFnXj+3J4z78PYVEwMm8CbeXu2yQ5RZJlKyZe
XAH33SO0ZRPMT+z045hM6N2kxbWqb2CoTgbO52Y/yQTYPIpy5fQDBl7mPK8YnbwH
XXRQ4ZskXSLR13buGxmYRB+lDrz8qb1lnEA1bUFF1iijzeflFtTKJc1bdgxo5NpM
cJWDHd5wXT7CWMTpBo1No2MygCCbun7Y3vfihL3Z9x8Mj+oneTRXB9ty9CbNekMN
FF5NANsbKqFzWREL8NvbqHdZEorAkqWBKYbqLYjtSamLvlmIz5YcY8qE3GMAwG8s
UT23wMiUiCe23qxgIJdjMZ4lZa2OfQj3NPBBeelJSbfL+8LOjfq1dY5mYtireRlW
hGwy7dkkzOBphmJvStUmqJJkXxvt6cG7b/uUBl3jwHn9zdAezlSmXLSlgGMuhG3P
UKfho39+5ejqJneEp6I8XPqUh+bm4bc+1Aktei/RZNafN8q+v2wQeXxY7K05H3P0
Br3CWo06t5I9B+wIW5du18tkjsHF8RLLPkjXW5s0YqvQCAPbQW72aO3eVCqhRQr6
zprcVh+SxXmtuvbX21U4+SPuoKZMr1c7iB0S2rcRX3srntGfdF66YV6l5xINv4zZ
KOu/0uIdZPe+cOwE2zy7MJYKB2jeLJ3ZMVQugZ9TnX+mQIEYSpC3cGT9qlJXZqot
WxMJ4wA5MwWbAiaPchXFe2XCD9HCr5xmEf7UIs3EDRvMp97Ocg8e3FrQEM/xtGFc
WR4IP4aJgaxM2S9WeyIiJc1JRC42Lc6HWIFz0Y6DA56mE1L26yWtUqeQkpRPCCE3
dcg3DZLWj3q1nb0gboqTj3Y+QRB/kcaljdpQzie1UXZ74DeRGUUVlZ4LHJlsxwKn
EpWyW8GexRrfQbyCwUdodUgRv6uZWSh8HGEMm31xhC1RpJ86NRAdxK3+ooS1Vawh
UAikhtAJcCEX1TnVcNfq5WC4P3k4aKWcr6KPJUFKfxGXhLl70+p4+j1t/lqwdU9g
bqiwfwGrT2lsLRbInzvqDUtkisg88p+ev4rFLaeuhPoOzJ8jzRH/5JamHwgZvzVi
EVFEiQBYMh29xIQaHk4Df0P3dDuHJZv6G0DpKIEbbBm/8ed8U6I/+fiDfelqclnm
2kP5wpwke0CjX59fSWqSGiIHaqiJ68As29SfEXFA5Vd0J1VNG+e8OBdCrnSS81Pi
F1HcblMzj4nV3Qiuik9uHjjDeHPKC1z6H+lx2Tarxi1JgImnowc5GHa/OahNPgNz
JKZ1I//vCY6ppPsesPHMxWGITQz7VMPPsa0avr/PPwe+4+2LcV6jn3N1lEZMgs00
c+GH3rjvC02v+WHzTCVmhB4fnc6wmF1kYpMM1hnzAuKgh5sqDZ2hoi2xkuz0clH+
zU6kiK1EgbRVmi4oyza6/J92Vn9yI7l2vbq8toLlFboaViuyBCFr28P48D+W3whQ
nq2i49R3g5mhStOFNCHT2g6xRPp0EzdjeNSLsl6+ZIyGP71Y25yaVWlNNoT9D9YW
ZEAFzoPAJc8+qx+Uzth/zwgiQvz/qYmyNXYd11PWgBCXrS7Xt3f03Vg+H57UvLFg
rV0FXa9Z9aKgyN3rHdvtL3Spaz9aXaUJwks1JW8EMAVZmOD1Vl9TzNOHo9+CSKQm
LGqV+tHl8G2mCwXtYbGBpz+JKWYHu3IahPBQHtgL9Z1Y0wEyhDQjISDk94askumB
12k9l3i5K9E7xWTfZCt7cWeqJBTuEj4L9yFIyfVUTBrIo964Knos4IqV8UyomPxn
M9a/nPKusIQBXle3+5LyIUt6mAYswX8aaPN+np7TQUFw2TB3kzhMU6XRijdWu+Sz
414wtka2aHoBZ0fsMB600JQakIlOapO1SDDrdGg5SzNmZtAtX0aa7wQshABOnavR
lWb1gyIGvyT7Rj30u0a5rOdXlLeLkLx8Qo+Vmdurq16lxJS3cYsZR59KmqRbNHeq
j+6dR6snlRZKvnME1arqh0nTCMjOu/dNsv+AOX0V2+mW3qzNBE79UPRVQdX3IA4m
Md+/VSry4e5lb0PF6BmXafuAOgrNqIlImisasF93Lah7HFCwvkH/BhEuqYdtRcMk
4DRjFqS8PGk21WW3vFE+a17bUn2LUFa8AwKxahaFDEZTAbRfNsadofjThK6S7ElJ
DwFr5vfahtL93zIoBXIPxX+qxB0ab1gtHaz+gUcKWAwuC6eeWW0BEDEBOYJhiQZo
dmXSe3TZjnWvMmnGdGPuLMunulU2N0nIkQtxyat3MtMJHGyu0XoW7RuyuSqjTNLQ
8hF0pGdFaelbi+HO1lUVz46ncQaD9V1yQ1Fmus634QJ/wjd1YgrrtJuX3jc3Csct
7HOB9WI2l5yVUvEp3W2vGxkeZWYg+4psgZKOdty7KPzlPMcDfatPAnRoilbrLxuR
YC9uMhPNqkB5f8A6oqblZQSa8qGCbQmFTZvkvSgsGTdHcdeTXBSka9eA6MKjkqCh
6olQtdrQV+uhYyz6Aauk0ZpJWy0pq0wuLLfGNb/B7Ke/l0qbqkMqXDO5R3VKcktw
aWXty7mXRDqzsqqvuIJU6+oohijH0r0zPmvRcxBKqJxCXWXXRfJ786rzzVnGjZ00
MTnd7/fNADx1xaZM/rV+eKELx8l0wHDQke+utXNBi1MvQR0MLzqQxk0l8d5f5b0g
7SpNZABY6sVYUNHfdUjRCRkmW7sD4BwxkqYlQwwVhUfoJwGP0X1Y9vAMWCEFNTlv
6YOxpQeLGywqTtZ31UKAT+HnF8L3YpsLO0kld6KoNXQo/u+/V3/0xpOglKhtFe3K
EGpO/wDnu7chaEyPeDcE6LyZuqgG1uGgskjUpkOygvIrHWIIH+4lqFwEcBwBBfOg
ja43GoR99mipx0d4Ewqm1PXCodPwtaAGsKTPApaEvDqDz5e8Kj7DnoFVNiXvgs28
bpkH7i/fKxAr9lxj5O5J2m3BU/Wc5YV8HIe4Z1fFSjvr+etMuzroqdhYI4ZoGBQH
dKBWIUETDBOxsFnD7Da23Bi8UiKUXOA0WndZc2VBUMQA3e4lfsrEP4Y+cyUAzr5o
FWjme80ceI26LzsFsZi4EedvmGDvgo2Eo/Ai1PVzQd5UPetxGXKjLtG6LK2LSbNX
v9YcPozNPKspv+qrxt7xEH+Hw3GCFDsTViAAfSc3aRz6UVcmdEkSxZ/pw25HOvdp
nmAbHreb+rioyGRwiHv0fHP26Mk8H/8L5dfmbvziKEw0T2PBEdwVXu5RD9syz3MW
KXWpqKp2sl0SUyGmk13Cvtx1nDAhCcrfL7NLWd3jVb0ibuzxsEuTjIggDP50nM6M
LNXJWlnGVctbieaGksvrX6w4Sli6oWXZR/5nZUhRlBmxd+LxWGaaciXbvZZ3F1xJ
aNue+CNBBQTkq69GyW/3lYB20Nx+04Qdy9+36031ILM4unvgLfMNdjBOi0odnWWB
7bGSjnHtrObkdeN0acIRPrArV30zSInWfd7++BxayAT7GwcvOfCx88mxw2cGfGqA
6ZZDP7Ig/T9DF8pvi1PwXG7Cc6AG6ATd8Zcik5MOybTO+P6SL8YfxkjR8MlDjg4r
wAyYAizhXjPn/kbYSnZnZ4u/TEVPzMjsptsjOT99Pyg+/CWSIUm6Ox55eYAZc51h
2yW8j+6PpqhMsvP7q+Si6xTPy8z2dPeIE7iE8NhJ7ZxlBiceHjedfRCsp0W954Zu
wxbXkWzWBBlK7uYpggNo7HPQok8q6BnH9bbi7TUeFH8J5AP4/9v3Fysa3GhbqNXP
skfVuZeNDCiufV+H3F+n/Yb2v+eTccJFwOdFi7Yh9GY9xcN2kfzTpF/Otr+FNgWk
Is0TLMH8BtIvIs5h/ahFnUiay0ZjoF1AfoXdtpbqASlpLmPqVRAKKIMSCbw5clJ7
Kh56qnu1o34b7JyHtvd7y4ZRuVjXraw7QgUpDHGnr9ny2UJN4/sFBzTPY7F9G3r/
JZmFzHjnqCdWkPH2Tn4LUHW7phvWM2T4+Z532mYeqhdhEluoXTlEeS+yrK20P29e
iT5ca1s8lOUXnfijD/gGcyIbJDgRfCdh6OI1AxRdiOCsg5wOUDmWg6I2GajlzrEr
37poX3ENtlfc/YS8wTzrCerRSxRFEgo+bl9tEsX69ziKQJuapmcgdbby4bjofCGQ
bld4xHIZ+yuEPHihtMm8JIP/KxVVwVyDxKn19t+DefXeUcmz/9OhX6x6J7sotduk
VM7Pq06r4c4pb4dAPMketczJ8m9CwMuZZDxBXkUUAB8MDMWOYyNk14wZr7uY+g/w
ettkrNintjmutmhEMb65OXu6imU4XjAlc/JBQ6cN+zLbtyLdfiTXEysvrOigFNGD
fUnduH3iDwgeoaGDDU21gzv1FgxUFOihIQqgoVInTRQzy3UtSJO2k4/SEbJ/qXR+
5OTgf1mmy6tumxLquE3p6Yf321EyEJTizEdFtZHYUaVy4ZYD/HdpY6UnMt20BXcE
X3DC1pkuTH5azpo/11l1oYDf7gHRTo48mR+Td48kiCbPlEfC2brxUcCEFLpuk5Ea
GdPw/gGwcMyt049tPZ9BDhbb1yGKZA5OpigbpVSpxw4THKejpyJlv5lNeXi+qRvg
UtZSBdm/e2P5P0lvD2+DObO4uM4dwj8JSI7y00fVTK9+LTTj/5nFG205M3QmQAuY
iD+W2koH+6Du07RkNFuZwNVev9BucS5weE7BQlHlbsFUaN03UdNEZN03a0IztCGe
SGaUkwiOExBD/uMQrGIY1XaewLVj4bpj6PrhF1qVUzwF9OoJy9Y8nXePvp/lZYlo
LAx3U5FjffFo776/xTvi0J4djkKDG1u9qdBHWD4MzsOwvgwkpfl+rZ1U73QXRl4j
YGVGicep4oZQfSfIKHWSveu9X58oz6bcmThn3rNIqQb5qBQYqWOWRmR5bGC1lxts
WhVmb+PznSuI+gJNBKSSxBkaCWyMuh/V5HxW2BjzUVcLNwDcqWfMWlQ1BasUjYj9
1+iMRq9yHcJ16ZOe8q9PN67X9IvXg39S4vAgG+3wgBfiv+2sWhGn6C4AHwC0eNaY
q1dKr/HYI/rc3eEMCrtzt+Qj8GCKSuFvAr3SrNdAzq6H+Vb6siZugO6pIukD6wZD
uj4KzYGKYsh9QEZRrGi4dGCUPRHdZkqR/lkrd9o2Ue/7bwipVeqP7Q7KdJoSNfQ4
goKxMItWKuAR7Pk7ICV/uFqZghfBd9MZDChgSdBz8Qs+Xe3dsaSrqCfHouDsmTrc
Olk1ie9SxV4tmUZNgB4TBscRRaKqosKygQP+SK/khLOCFhOmsbrrXKQ5QiTxMM2d
sCzra3AqBzjXa+93vQAt81Xa4Mtsbi6yd8P06d4Pq7XKwRVL/mq0t3pSio/T+adK
XIEafyAE33LWdsW3vClFRCF0LgQ/q6WiPcL6+jzkfqCPGPGBsELpWVGhuosWmVTU
D4RSvDu3FM5XkGZ9KD/UPFtAGnPRwq/vlju72FQ5mbndBuQyy//HQVWdDGBw5yN9
ev8lypllBOzxpcdPYnSDd1v4RCTUd1RXxMqt/c2EThQbggd+6gnvpNBMUu+RUlkF
zMXz+npyMOvHPNWpS+3WNIyHxAU8NgFG0/GPPCc7iHECFZuR4NSq6f0rlsvDQf3v
Yk/lssJ71ydIPvLztmF3pcZx4aJZfzOlL4KgQT4bfG5PoM/TFZHM1SIUknLFW5hm
CX4wIj/m00Fslk98huHBapG+OXre83AWceE140hSCyl/tveDGM7cqRypoqyfy1yL
JRRHig7KEOhi1QcL5FrT9F5EFWCzzVFYt4lLRLWIw3K6xtjtuYIdJjLvry1OK5TW
N8SnJtvO+qh8Pf4SBCbXOpdWp1uQgIZXqS9CwHOV3+v4PZQYhRBVzNfXS7UBXpLZ
EPyYli2DGi351iYUzv9lYQ3WX2erTAixoFf6wH8BY84G3AqYZZIIZ0LUeLZsdtTY
im5Ww9QsFCZlZf/+x2W/K2WMJpQQpvWqc7jk6Tny1mvod8kBHsAYNZexpC//Q4jY
Ap6lFg+k3HYe58Tx9mL3xtWDmmcZVn4sN/AaLK2gvMuQz7dq3i8sB2pMrROEJFtO
2R1pRodw0J4a1sygHB15fDc+CxpNZVaMsATfcaHbZ4Py4voewRW/w712MZkr+ejD
az/BrBLEawFLwhSzfRhinQfGuCYWMtvBzJYgEVecaZFzI5HTtTSeIBUd6fJ5t7SX
VrgL1nnX3/+kfLYzICKic8OLzHOjgvgE7zngSFQLh5NF/8LaotcBIIJSec79RYJw
SVJcKMQYE6uZFjKNNEoMg+DglKRBJSUN3cYmGStTU+xsn920NnJWls98zQjJJKvY
doXMdlu03bGBW/VR7uq3PIVjCzF6nRb8LsKcWcuEb3SU9gZpEBn1zRjKvY/2DIPW
RL6nsoq90mkahlenvg8j4imzQ7Llja/T+lhPIvZMOdbRvfGDyQLj+iPcqKsitEfs
cbXkgU4T0vEfhgPjLz+CDNt4zkLv8toVKet22j1aawKEl+M3JjZtsA06DCd2k5QI
VghSN5wT+qDefggZWwGNiGi8avSRESqYu8I8DhbAo76QDt3f2GddNIEErIBS2IKK
xJLwcZF310Yu2+P+vVr75zfzbXfASw7byctM2pvjiFrDGolEQ6UCrJJHqUUzXi8+
dqSK3r5NzE2eUvSOaxrsIooVSy2UQl664N4Cqsyv714FocJKmm84qbv9uSjGgwXn
MX36hMo3bm19gjRogetGIcFActLXNF9OSg8mpZkdgrLemtOvKjmIdAnGh8qsUVrl
W7JbR1hVelqxBkhlZTbL3af0/+fmob1O34Q1eyw/Y7/NrKnwwEtA/Pa0O5/OR/yx
qKmnCeu61K1xsFwH577CLEy34uehRGBeINyof6pSzwp8iG//WMcbn3ZgN6Kd/A7I
zc6mc9MYkGTE9TrSI1jMmtIefwlmXgvRys3U6HwI0MKMnY5vjvEZInCNHK66qwAU
9s+UExMxyWSHSnGUNAyS23ZQE8O4J/3y8WPm2r0BJSiD3B8Y0FlHlt8AaOtimuuj
rq48Yyhw+ZsDLiipUwmZJIyy2cI6y8h4V/DVN2kL8mflMja8rOb56BspaEZ4i0vx
r1ZDQrSB1utyYsSV7LU9K6xV2cjMgUAr00YDvUCP9z1h/DmXrSGcS/iKXVVn5jo6
Vj2o43f7RCW6wKulbhT7cyfAIrbsKbBQbVEoPCM7m7fvZJNtAFWR3c9jrcpiMP65
wOUkpzpcAeJmrvD80l6/hit0uNNTMrXpovXkrXQPN2MG3PM07f5uhG53Jm2f2k7d
cOy9Zjh7kuvPhNWP7CqLV8tQbBlP5d/vvzNvcJZ13V8/pzNTgyTsV8Jk/0ABZKPN
X9Tt6qIcryRxOfTA1lQ2xU1c4Qi5/3PeQxc/EzCCyqdBYKxBBPcHKQC+0AzWVSqG
kduTH4yAj2VMoomZepuV+7LgefMt9HO+cd83rliffgd2NozFnwGuru85b9sSdDe0
RTRWyWLFgK1/4WXhD0bfMxeGBKbAR4Q1MuXA1iLVZ1crH0UhuksgT5d7J06/kHzX
QlNCLBEvyhC7D7vUAlf3Tw4ut8hk12VuqZa9FUoOA/nPIGj6qcgsx6fCTEuzOWRy
y7bknG12LGAyRRHvvmF9zgCI2aORcYJqe11VAHNxyRm4q8uUwn/+H/hHxnpj6yMn
Xg3B4kjAGkH3+QnEIXsVn3stTmmr1tOZL9WUrHL/axtzWj44carfk1dLlOPf8TZ4
OO/DgjnUBcBf6Jt1yylSIPq2XNxcF8+pV/dE/eeICoSqmQ0OfIjoO5kP/wc/z8VM
kLGiUtgl5Mvm0bsN8Ug+w9RR74i0hcGnV47YOoWmKvx23vSPs0OgNEECygKfC9v6
7ZXN3BoZVTaXGfIyw5sFkthfNiu+pNQNlSIGjrW2HlwXPwDaV6Y2cUK1Fc2fLk+r
x85bSy0fxoKAhWGsIhxOfcMzPXLfLq6a+ORX7Hxcz8fjPwwei3Fl2B3l9EFKfiER
iPg0AXzgeSQtRd09R0PlU0v4eOL553Wtb0dvin98xg9C+3kzKJC2Hvig+6+uVpd2
eTY3NBA3z2ZuSuq3V4lcJ+J1wBIUvnfOtLnnNYYKFjjRAznu9QVP2HrCVVhERaN+
K6PKn7mdkbDF4UJ2oa/hLmJ0v63ecPlxa0bshwQajrjAyTf6faeSw0du8O5ZeiY2
OT2tN5CkUEacmqFTedoKz5OZpqlwJEyCVg368aLvZAB/xtaPa9AsgE+qEffuav/3
vcyddz+YRvv8LpQXkmvuUWs8pqzumB1wXWZldp/GlddK5UcHsJzg2V2hlmggAx8h
hC8L0Wapig4xCGnmkh7E5Whkgz0IRir/GovP0KrvCAV8LgMJ7zEJqHMgYCNYLfr+
IDQjUw374GOK0JqS38LweFp6Om97QsvqIDtS/+8Coau8Q0ZmxvyqBj3kao0h3//U
vt4IzsWIxnNVdCNKlXP1TFkoTuRRYlHDlc/zUXxQMvcbwvim9773UbpWaep1BOgN
nR1vFVQwXYQK+N25YLWM7ZM9e37ydp+pKIi+VpOjypg4en+SBsoDhZBLbyOQ+9B2
mQ1KmX2AzJHAX37gDra7vmvLwhQs8YcGfAoDLePKwdXPVRkV6K9EtbQ7/a1Ww5/F
RrE6nv4k5sHB9oLkGRTCfEqWZErhRLLMxa4ErWbYaQvJRdbJ7K6mGlyE4h6Z+KR7
qPsI9Y9hYTVqfF6RIk44xfD04cQm/EoWYWxsLxySgR39CQOMUH3v3Ggncg5pUGda
Xap4x39uWHHnKkalvGD8EU58tLZZyisJjSYBDKC8ySux07IdqtDtLA/9kG1LAtck
4f7zT5t2TzLQAQjh69/tPx3JsBX8qiaj5KI0X6GYHHNmnEtD+iYmK0x+uBM6XSaO
OfwjqZz90RNtXL/meffKD1GW1/tzbhNKsI1YRMPIc2rw5DOsRxtlDNpePY+kLsFj
w6ur2PtPz394RBC8wDeOzleoqNE5oWXbms4NCyxXwsFemvmCtnc8F2sLmwZKmJ1G
6/7fnJ3R77R6B1CN8pLtZzyARyfH2n62GOcGBpcP6V5/cUFsh0c8JMfMnsA+DDEf
soMSiVH8BoEONoxbsfPD7vNnlwNCQRhpE1a0pQDJBtUYZToG+8nHEAgMKirFWp4F
oDURn8SACieC0iK8Bq6MtZq7nyXErDRoY7Ec3f9u9gl92jDre5k0yPpMH2ny7aPb
OivUnyba9TdcBapdqtrCIhJSqDw1jzIra6svGRCqV6XRdb+qTSj1dl5QdFn/DcQs
RORquIIiSmxGZztVjzYEClvMEZF/VmvbvpZd8OJOHnpdcWBf0t2lTM6Cr96YHgnj
Y/87IwNFoAHrMzBLJJ+aNrLYnm50NC+q5LGQ6j3hlO7yVFJDagr1PdGlGH410L69
SL8D6TNRB7txYkqAeNgI9S8k0+PuLl4BvKtuAiefIROErYyB1CSLfPHefCljHumm
aFUODZeCY49htlT1ekjgY4XouoKdWyD8zh72TneOWurDBztl258Zzb8JXNo8lUmy
iyHqjy3gDBNTvFujDUeTqCFrJ9kCk3zAambvsIkDD/sk8PbrEVpbksXMJaduTGDF
05+YI++Loq2dx80llfwfs0gy4BQ0WZvcLG/naJEgj/IAgBOTTQAXtdln4i6AWPyS
I3/ZZwVVydkpTVmCAP0WP9GxYB01lOd+s3gnzr9x83lc3Lrp5NX5cqJM/uYNWnoq
PXVRV/KACvWo6cxq76pmEcTrMSczYzwQw5+IM6DFQ2NtMoD355OuKNEqMuHHFT6u
0RZigMGqP8zNx+l80umzBRZQkDIHOVMJ3cm41gGpPCTpB5YMv1OAiNFQd0EWsPy+
5lUd3RWuNNWU5JXG6SXRp9z9jxB44vuEWh5bAdkq3Sy2hkmc48vU4ambHGR0d781
VMsuCCki3/tY7I9laIJnhujWdF9oCXUoPWSUeEhR3ngpCB/u85xqXLfwcE3xsvz6
TklRmvSEggIWCuiJMckm8tohrGSXbs9JPBxTfrxtCc2dOt0BteH2MHX6jHSGwKyx
aqipRSVO/p4QHw9BwjDXOWArv47dFBMf6nxuWTMIsOHVJgYBnNU1v5P3hkW7xjff
JV7hcdDJCn/Qzmu/zysA4lJ+HqwNfmcT919s2Egb+3vDTCT/0haljLKGYqERNIw9
TmYybiDrTbVVWx3f0PAeJPGH/kGRxyrjiScz6h2Tt8gcV4HyjPtkUTt1fZhPEFzX
gCQoKT0RFZftPP5VcKXw0GnZFrpf1gNC9kHmAT4rmmO46Wu6D0DRGdYF74Quy4vP
Nny+cSI3L6NIRvAkm9DcCXtW30dSv/MtzTKAGa2OSuGIwe0Gy4jVQ1vAJ3nE/iaG
UCpgoQBlZwQaQn8rM2yruYWsw5UnnArPUeOMY8fVcgSiTwsv7B5doWFeenFqLcV1
exmYlB6apUo7v/g1OYn3G1BsWrSyrXdrp2PNwB4b1qUsKYWLEt2yBEdV5ywosqEr
YmnFcL+GTgCHAmRdnklHsskDFJEW2S+0ynnpdRVZg53hdCE/cdCaCN3yHjJhxGIR
04M735Opz/fcKxTYC0KEwdKG877F7ZBWU7rvuMyEpOvwmR8+sBCYBu/rBhHmIb9T
XoPTzJYncyxX0/h9c2UI2QF9EL0KW9pfQWAUnynaa2PfhjRTfEmKkaofs46B6OgR
jrefLBmgEJsvuuKmcI3+uvRVgYVpP9g3aAL5rggaJw+XaBDwAVfwK/qopV/1BG0y
bpUiU2Q19zFjrWn2cXwAE2tdsD6ozDD/K6W5CvJxv0D2nsRBowDTBTTOISqtaHzk
o4GPR2rbOAxPSfB9ZEsQxypUGNFkOK87LirD2AgcK/YwaC8O/myo/CLk0PGmxXvn
xYjyJONYIzMg1MNASGlPBI5UHkapIqnrhVQtF5mRTVwYDxPuPQ1Ru2e3AcbesCYS
va8YpQjSe7PQfjfv6vy2T3kCo5ylSGiib/d1djIXxFKcxN561bjK+lqvmHSk6uT8
SG/8NIVPv4Vt2sNyPpPEnD92EhoNHMvXyC1SINTfcMo1S9Y67zyF3FoGp5vRRu21
Xp4CdE9IHvjV0FfVZqJtLBZKaAWBNPixJQ4WxRRGKW/kKbuJkeSGKDohITwgYO8d
AQ4C4kTpsvAgkFHVqMO2EZc+YHZkIMbKJqIrLEIOKcP5Pv+hL9MQIDuMoC4K/pN9
wOfUbAx7NQNlQbjjaMKpIVFg81GCg6uLqsWRMXewRKmG/WSJ2QfsImKpKyFSShBx
3Dp6OXizFqZex9Dx6/od2Eoxc/6WzGYJE2ppg1YeW4Ub7eUG6vCGK3vXB04X9mr/
2GTqB/3OuXalmFzAz4XbIZW2/wpfDG48AqkBzwtED2UaF6k/K4DgWHQinYGjgbZx
RBAPd0mbJduFMJuVn/e7khxO61wmkKc82PJ8iSf5BxW4mkYJdI5cJcecH4ObwZAI
mweWBgljrYHo59f99ZRMBwRSXj4Z8y/iEX2CYdsF4PD/aX5kZFje8s4gubPEm+Qc
WfsxCjlyx1K1aEF419m1r7VU3JQbcy2fsF6gKozeELb7dOXrV79+PROEhIO6GSUf
pV4MOQyDxRLllGzpBFKyPpAScaVQ6HZbz94R4Pdmb58yW66712wrr0seWZS3I6Z0
ny52KRDPfSqcIDWO2QvDl6YvQyvKhjmLuHI7XWMk6rzVCvnH/jaKIJp2pMVthB9f
CPKDK8WtZ19fFU7G8BJmXP+QV5x1yMqSgCk7FhiHwsjkMVq4x8nWSj3RpDH4Nfmr
vpHUoYqLk8nVFfN7JgWWSO/ShjVl8hV6SUKPy2sk7okJqeckOek9Coa/+B0i9c2f
vwYzzkomsJJJKaKS3HsB7gYPzNcqvfsKfuGNmPIa0/9rUgbqcRDkpk1ebWDkHUC+
nHpVmQHQOLAMDjOBKLZuwUR0+xP5Xca1BMgwij9vzOpH76W6pDhhUgAIjPOdZ67h
dA57wMxVJaVr4li8yQsVklv62ExpvXVdvwAerMhhvtTx5apHUJVdxpamCr6jdH/7
5Pcb415bFStT2Rjywlf/xftGiSPP6imWzSmDvcshT/x2ni8krgAvBwxe4wOUo8ul
/7k9cVZ8dEFPKkak3BGa90ZjOyUqCwjjyENbl2KmGjpv3TwtpgkoXj5Y1U1OuBwi
d1qKo5l+IXXshnfc/WX9T3fOiS2OZLJQWu8O2m3OHQKRchMKaoVPM92fjbBpHjKi
DnV+gydxnTyhgXd7sYmC6GtuTfviRR8TJcXjYqNQhlQjMkXr8OJ8yBCsTlz8dAPX
HtqrcNYHbrYoqUwhsTVEkdSe42R3LY5hfhCUcU8Bm7fUxJGEJ2g8siFW7PFOG+fx
7Z8BYx84w0KQRDliuq+2Bji8mg0qsraVHeB7mN88Ywb4nbG/whadWqk9d7szzCi0
DMMDyRPyGFzkublppiKhINpxNcJwOxET8D5b5iVfjtG6yk1Faag+rTpH2VJ3jjkx
q3axE3IjkCHzjI1RnMHOemqJImKM4eud1QiffmVG/OFXCpydFfM4Poset7XXrqKL
CLF9/iAJF9bNEdz6p2gJSTtRjoxUI7Dzbc0IQqymu2/BSO2blUFUXseH45VwvHhG
LFbZsshGPL/crZGGemqYVeZaWKCcgvzmLq0aqgIGRG0+XU/MzJDrHBF6zIPlI1Z8
g7xqv+7K3PmkSCdgOe01FD4Ao/6BrRmW6XroTW+hkN04dXn49aBqp63NKuWnlnl/
f+eHEAGJZipkmM7p/S0R1i6X4I8/QoEVlnThJE7PeoAKIq3J5ZzFMExqS95JJgwq
ouPamBl4RShMB0NV7BjmkLdjRxmZPim3+cgVWNSl4Ciu1iyMaYWOUClg9TB04B7x
PyRlvrEBaDLejORtTHnaPREBriAB/IimTntuV/cJWPaHJSd1NQHaQybvdJOFlFU0
C+nPkBzefv5WuEq/2/EezoQGYEn+CaJnxfhgqQwoK9HFQzFzw5D9TL6fgtONUwy0
TDxHDxbSGxJtpEdOtrPlLJmKbtkvydfAfcvlu3uxGZO8/Vlr3TkPGBMvn9FTm8kw
hfUgK3aHZ0RFTysRyzU1gMg8lLq1gCmbyI7Wk/JLXHX5iY9lzr4Hc/Fw21tuj7af
UGWaYbC1604kURqv9YgN8kwsitqbiLbH8j8vEsZCEX7DfGtfZpNPQsN7hqFeP0Nf
d95NBA9D9yDUkfiMc8U2sTjWkzZl2N9oa7GesgqMvFsgIx2TdI/5qzyU6krI6IE1
WWy2ZMpWfadfl3q/BORkMGV4Pi1uFn412ZpDUM2wIKd0CqxE5JOey+BivrcYzFmu
D+Ra31jIVOUAVeY5ByG/HARzBf9cxlH6Nn6E+xamOehp8A41q7KhLj3Ub2jD413r
W0ESsMxitBng5ZN+WeGijDDbOhAKWLp9hX7iYGIEvX0D++Wwl2CvSTxddiyfKb0Y
MJJUtQtarm4ky6PqcCQGQoqRxIlkbPWeRosEB0Y9zCQ8ffLpw3gZDKr58oxeF6P4
CRcTQ73cD0jte3rAdw9pTqBskzAL03RwnmPts5BNI5H7SR97N796JO+PPUIPIfNb
HyK3We2pdhEXHd7BZxkeAWwu3SF0AtL+f2HTMmHRHLsajqGhUE0BDxR+iCflMDfW
s68J4Atha4DuyLzup0n1eJYrOf7PipuYMpjsfuYPNeAc+raSgNOdZJ/VUr8a59Vk
ego/vaxBd2gTuhM41Mu2Z6uVhvc2c1X/I19kRQ2dkJfk1/HpKJ2/TpqUg24ijsJj
1xXGMSLlaYVlvBbe401BjIP8pWEUVESsEctAfDX3YaL0yrFdTUA6fbz9zhWtiPaq
8N0Qx/A4385VZy9VzhHi1UZ8IvXpM1J1etjWnaem+bC795HAAez0DTyFi8GhtIT9
JBu+6OrdugqLpQOqqawWQScuCOyRsvl7FMrTjwqzRPrWO8T8PmGCpQZkc6aKmas9
USuTv/xZSrb1UCvmT2HeGzJ7x9EJfPbH4m8RKAqeirJv5T1z5jeWKPPOCfwrPBT1
g92W+DM9TKc+61VzOjxz70yI+Ids6Ylh0MoE2V+/bKBGUTtxGMi546Kua/ZTeaxG
03nJhCjsuiQU5AI9iFerOxaZ1kzCRad3/vT3wDhedX/bQ2mdGZDCgVmimTvuV1hB
wjisKcE5SiLtf2ph744whE+JkLPZr3WoU4iwxxCwJ6tt2x2vpJZl1axu7xhlDOJC
XayNpl8rh5AjpGHEFYp/GU5ISrHTXhaLtpQi7CkCp6KbuFu+bHxSNXyopla6s2xK
bCgBc40Nz2ARaatK45j/KaZ4/06trln8cgH432g3IrD8NLYbOZTzBbGBZC4s/bT4
ApxPSplBFq4g5KZZwRs3crULRSO/R/ZICF9NwGll2DWDXTf2/B2i5SDuofN1dye3
Rz0zj7TESLzZbIKY4pK/eKYcYzKP6jzWNpBXtOHn3+ATp+buMsax4KFOQCamxZmM
6uvkDlQAuwjGZcywj5IaL2SKE5DtReOUixuYaxRd+r72ci57HJo7gGTpi/J7A2Gm
cxI7GmREtpkthMyEBarzXLhLd6RPixeeLGIt+iidDoUsTx7F3H2aUo/ejCBFG+L/
Nq55+eRrVduek9bBNbus0N6mVjA/Eu/nPPa8HJRH9dbJyHEeE8VqIuJ0P58bLhPh
PTG/cDH0/LbptfY5gojROflFfp3UDKznYx7ZpMTeWX5Jdr1VfLO3fbrmvTGpbi/7
XzBZVAOn0uycKMIX5aqSzx7K1Qy4D/18cTws4rA95P2oCNSx+BKFnwyQqyv/AAhb
Ro9FylWEFIZEo0XDGP2Nhb2nyVp4elgGKxvAhiGCsutLMxYhK7/lQzdRm+J+tyse
HOnVwByR0DmyHVnO6csX+Cdr3skeJEe63fEyeiwOQ0B7famAkQ8xwqtsgsdehxbF
Y9B4oeDyEBlscDox9YvZ5fqEyvgaOwaTVRk60UIZdM8rM25lC63J4EaHk47gg/6Q
FXiMHSXaFQvAyIf7IwXmF8aIFZLlCiqRRiXv20Gy+r40GiPDWQjsdszSzX+r4ZMe
KTGzwk+4nlcxBXv4bgiKIyaI9I1iyvR6jUSgu81WrsJjBPTJa4MYYctAGlii0Sn6
vwKla9VXr5zqLkJTdkgYZDAtht64E2SIOVihqS6zCGGFNr8UR30mtje+JtHi4CEI
xnUw+Du/QAzMMRVufP0ZpK2zssNo+9yBWmYOEDTpcmSsAg9pBidN9vQEuXWc0Rea
d3pLoSSU1IBfPXRur23uMOoYaMwa37AYUoVmuxBYH948A7vFVEQ0L+o81WYRUSrp
PmLkveqfrWiFTUsz6kcXg5HaJ7turMC8f1ujOpN45rXWdUbO/xbKzDn6TwDZ15NS
6ry6GuB2VfvZyDoa0Mn4mTyPFob4HX9oCeGNPDwHIZJDCvc38otJQZFfDutUVc2F
2v/K8IN0S9+PDUTRRKL/YCkcVsfS1xvxE348JHfaF990rPERedYwBLXqvVjrBzXv
gvga7GNiluNmdHFcVf6fESucGHYRDBXe25ntq9rtjrDC4Yqe1TSgulTqLonoJXPd
uybWLfKbjYhzxNsy+ooxyOLzVXjDg3JUDX0wDQA4WqHVy18TW95esuigcoWzUuAo
CsHxvB34M0eQN4Qt+gsxkUv6sAsFrZCxrnGblRbNTUUQA7iMdaTbBNQoAr0wxzxC
yL8KIUaL1RYitbCEN5gYBFT7xXgryX5PLaqKCQX9DnOCsc9eDt68svifOC5vpirc
VQrxnbEct0srywBNqBxHsksa4wmNv98HoPUCWj9KXiN4hVNugXoRhl8ArXrgbdgy
H3A3mQiqi/tv9taUq9XZZN2eWhXPprHA4PyNIvkBFxDCM3+g47Vb25fQ5N7ss5R8
InOMZzxBfZWvlumkKUfAK14fQ9YxgjBBLKcxB0mUDcJoZxFezwHNh06gYuINBGjQ
2tU10VZ0YAvp/bqRasgdnj1nk+w2A5k+9BklpAwyf9ZsTZhGJwkfnWEDlxjlLy7o
jwj6VslXa4OBFH7+CeycRKRo20G36TGKcld6T88y6D0qfg6Qg3IAEq7K3S/r6aZd
lHxEqE3Y1kgyycbeUuvXtVL3WVNqnEOxrYxqSjPr4X9efym7yem7B9BknyVg+5Il
J+NHuVqm72gdAeDU3Luuu00lfNYNLHPrycJp6xkX319/x9gzrltNVF5Xx5s96PgH
C+Lma3tt18IukCrzYpLuW6bI07MGhVTcIz/sNtumG7t924Ls4+03UHb/PrjpuFbS
LCLRYJSxkrAfdHuivaSzw/0XnOWHILNXS5mfqEC3UfNEDe94xbPrAKOLbi1bouNw
tceEo2C4OPHMOgCFVwH0tdSDDuWg8ZZ0q7fvZRFci/htlVBMWpaQkyDUZTW17aCE
7HU5bSsGT7gNMhWRhcby3c6OrIzqAwFqTTgOyTjxub7DDQRkk9zyoWgvhZUxErWu
RwH0eXOxeG2katdLNdYrJ8VX5g+omA2xgXIkDViTgMVh9s3cysQDBvJhqFjZLP3b
fRZaiSwjrc9Hxi8KRntSua4IZDR3ruXfDR1j++KPMZ7Tl6B0fB4cC18nGFxx9bbr
HJfM+aLFJ2UL3zrV2tQYSbFEOOPBwljz1PhJRDNIESteoqaVmECKqW5iLOFNvi9L
TD7GlIn5ybIyUw55tap7B0pcXxBWMbQ09gHvUwFMowJJmnx+yfY1axyLMO8vFq+H
AzfrgENm7sWnr1z5APEyBjo94g8D4fxxOyAkTD11P+t+hjYFcluKDSYU+sVnEEs6
s4DzxpBq3XbDm4riX/7pBebQvwC82BA6ePvAEy9BHIJFdkOrST9bwngqEJ9s/Aaa
+l70XwnVnYfsP5+TVtFY5TobZqlw1QtzVrqUzAjN1H74j5nYIo9U00nxseTojXmb
IdH2/RQEhf3nkOFDRHxlg/U4SMJSBU42KFNtO8d4vdrUxEFppqTk8balkrGAbald
yseWtnDnfR8i8F5jNAlpEc2BuT6KA2+iVNoVSsQQ95TOq2b/PD4GHR/EfWbbdoFO
Z+uTzO6ST+2H5wc732No5xrUOgl3bmNafZjLJELGqcbVuLYXWYD7fF+qOmcpazSK
4iCrj/Kg5K4NuHhqIRTFsI9gkKtc0AfWyOGyjxYfstl+SK7DW+qtb6VkzvdXAOFY
PloijVboe7etcZl64sLL9iRjWbFBZRzC0FoQ9n1+BuXzkwebEKAaGllDTXtdUFGC
nl+vASbdkA/bdQBYyJxLDRKF5+LtdvXTSghnj5eREk/nqzwxihsXAnfD4y58/W2o
F87b6nw+WEpFibWsPTxOjlCcgtFsIVH4yGpD6dTFwSG07BWYlgYUvHbuZgRZ5pnn
ETQOdsTEH891x/TCGIUwNr3QPyeAO7EMiUPa5TSa8k+uOrqlkazWRvLGoMMQumNi
7/04kDUWqThl8TfqvGzmBKEReTLBnG532S0R3JfcOfTLsalKM0fouksEH0DBOn09
dtNBshp5mvI8yPvSeLAFz5yz8Le9uyB7h0TH2zyJRNKTei+ILI1MorCS08vxE/Js
wOrMCQ2U2tfmF/QnyRqpHESqXKprwDpqVF/XQR3bTqQigDa3X4+67wZbEE1oQcX8
u8/jzrzAAMqGe2HqY85QM+hb90m8QutLfcBkCBjzrlk/YPa2ktAz9XUbrH+jH1fH
PVb9yw4W6b2xK964YmS1OUTDxLQvFlSQ6iwxRVONhO2wiqFlqqp7IV5OG+CgkzhJ
pg8oIT6Ibvef1fWIrLywOX1TM75d0kZq5SNwX73vyB1uuuEnFesXxSTQgwHhMvl5
7/JztLI1ahGssb6KjKk0dQL6eJILuwn4y75fhddTMvxofTlHKYYbsqKFaA72VxNm
pwx2ToH0jQQdiwIAFLDw9FPOJs8KKtBDAL0NBWwIvDAtWUSNUxOdPvEr08DXEHZw
FNF0RRhpaQyYuSu6fs2FAFQhYKYCMJLJ7x0Mvj4XmI5aORDrAguOA4zj5DimuHKj
jM0GkT4KfMEMLQ6PXEzA/MHcxrJM1qELFvrvkJ/JlyZ8UIAOKqppv11PmPt7CHrc
e0X4yWPj41OTChAAOZbowjyEesix7XD3SjarqMRYlGvYJc4SakmURAgNunJROJgr
B3clT4qGnDYr+ZVq3yYZjy25jKcv35rgvAqUKXvrdzPSt0Mo8M1o/qw4PNA6U7tE
4noxYk+4/kz+PnQPG3M2c3lVvQSJ9CFrzkNhejjiNMCbh0eXyKlLWQDX9jYJ/sw3
0lUdTo9ftqwWcwK3ZIi8ehz1Spj4mqwOza12GJvK377vO74KgYr9V33Rn21XYDFX
oTxODPIqOzmOQawAKQp8QzNFgZYi6ppTY3xs9e5CerY0b0ma6bpi0b1XHDB+vFcv
JknYQgbISQ8tNAR5U/YeUqLL5EQLLu5UcCyMgf9okSPQZV+52c8gDfbPGOjpHaHT
ciyAO5su3OcHEoA15I+Qipa1N4GbaAW3QBHMv30e0N8zWyqboNLP6wEilaZ0w50A
cMFZ4xO76KgI5AunbkSkPyUF6GYC6MQVoO9kFFtlo7+VccluipWD4LyuAUMLxQe6
SInPP7nLOrigEjWlkuCZaUDh7sWAHETyjbtbb0cZ5bV2OCzIvqQ6Z/+4Bpa8h8ye
DTrDriAskNJ3YPtQ722iRnz07gGs1K7FiL2+BLHi8Er9fs5yFOh6V/L9XA71UXem
KU7bU61qGPdJuxnlwZ/3SNwTKMDjJTuyOui6Ok8AVvOw5dSDmPin6OSBujy+MMye
udSrhBZO2t8Wz5nfHAU5X2LwcGjFezmENkTQxMF0TLK/pNJacSTJ6ifknszvk+sX
MtAdE2EnYzToPCxDnv2Fp4XDhtxcXFXSNwRyUOkD9oVuRS2/j8hPsHGmTWG1kFs/
AdXrfwqisl/sA4KuOGmxqaD5oshekeQrHUEyl9QxhBP01E3Ut53Kyu2GS205+3b4
uPLI239P6bvESB23zal/hdc36OmGy6JHWp2/E9gv9SNqnt8LktGQ0hC+wjXEeTSm
VgsBtYS6lI6IhKFuN77CQs9cKARAekeNrGSp8k6pQAC1anpv2I5pvgDPUWP35ggV
ogir56GBxuxefgPOtitPA1SihNkiSVL0ogQJO6mL2+rNgVKE3wnn5GQ2njbPOEZo
aIHvps6XMKghQK3CVmPSJq/JGVSalvJw+BoV4aTN/7Yqfd0nwuZXPoOgxAtbYyJg
h0+P9D7Q/GhNVRaIVEzVdZwuTdLGmVXIgm/cqn2HPpfNGRvVv8n/Rnspbqoo26pr
q863bkXDEGdvXoMCuiBXdNUP2EL19oOyzREECbzOyPpehztHGBgTZB8939cZFqqL
SAJ1D3TsUtPqpXSuEX3WbR7IS0s4f3ms3lQSBOyZYwYq3y7t3Gh5aNx1dSnwc7i1
B1OrKhhATlmXlf7unV81VF1ScQ2sjKrXin58+RZmhjNxKbZ2xZ9Ock9+yML4a6Ni
BqfnQ7hdnMtWi54eQ0cjjmsYFmQFTi5cQR1lUQE/RP4m/7JJDHYQdvY0S1OaLY5i
8/Gexmn+ik+lFY1UNce6I5LTDpSwW6ALEpGIb4o0tc6R7KtcBAsfMFoclJeRYQ0l
8ma8WczKz6CoVBm3vNZCOoNsIjQ93xMSbVdEPruIydIkkRf7ltDZj9UZWfoYJSk0
vZm51zOBSjpFJvXYkPcBW9JuYri5isMskM32Ny/wxvYmrc1O57G8R0ZHhR2ySUFe
E6RmOSYncv5tOhZ6LO30iNacirmTteH7JfuSyP3G4DLmntLsuUmfmSS6aDIhe74H
1pJ6Rf13oJLj1NI7Z1WhaEgTnJP9QrdUGLOc/dtUwMqCGalEdF67aqTugSiPaDwR
iVYqfcV11nSPofvh/pHpdOtEuP+7ALNxgZPUlnx/tvPaWgpqxw89zwX+UCWjuyaF
aHuO/MIUMApL8EGgPyASdFPtoBpA5u/k+f0UKHT5wf9Gak9l0LHqgP12cIJ+Oqbj
BVwF3g+3a4U67aY6lEzA+9Dh/NQPAgyo4Du/kXxmsWgDPuNBH3Xaa+Zs+20f21eE
wuIXLD9dDOvcXEi7QUryd6tPRP5Luhh53OMillKSB0LdK8fokJkSeTmNMIkJ/Hf1
oV4Nzo1CciRAOK2UAMlkFynbNIXDRDuLV4P8NRFMB90qI+58ojPPdRJ+8lLmeKgc
ZlVGgPTCOjYSX6uENuTHi9R/Z74MQ7eBmz+hpD4W6YBLJGEPJViDYpEdWZJRdQw7
HQxbocOAzy0fAoJKfV2EyfEvict21DLweam53PtEMb+knhVgAVPTL/5H8LLtVeJ3
C2mlo70nbE6wQzJDOqCRQlBilDTBZZf8xPv3gSRCeskJ4p7s05nTY8ovLvukD+LZ
fGMOH8+vxAIGe1rv+a9/aYGhhqWe8iZA+tkKj6DK6Kn7hFu6EUKIuYHbbm5mHJj+
17RxRjmJ540jmt6oFfF+h9USdZ00P+nJYh0/4IW+ougG4hPWxG/wAhFwhhXsLT1k
krErUYkMMYBeurp0U3NNfJ/3TJMeHY+3DHHsfoUXz2BHeyORS/3TRg+ivvhdDJrH
5577CsCfYxV5dVSI5yKNgKhGlmka8g2pXeln57dyDdjiicQFcj7XZUpOx28+8mAj
GD8GHjW/pBt8LMtCHOoJ+0zbGe6S/vJoKLTc3o7Jh9X8jrfkmn5zX+vVs95xU00+
v0cx2xWlcFkxsx4XYVpvk831UuS8A8V8r6gt3M8vrp/2K7d048T6zctq4ghSIXEy
qTJFWRPIyd1oUXrUJrux2KcBIFFcKGBqVpJRtQvrhhXv/O6XNS+OQwbbCrEzHVWz
0WXQIvfNrWUWCBXGJoqvGJ2o1jyI1IOwBKwDHxSRGSGgwQpmaKYgDDedHfQ7tFcd
+39sb5kDe4cDqNHrYHpTMrD6y/BsQO/0jTjehhtxfpb4SkFyS2xXXMrXGidMgZn5
J9fjRSssKum4Hv17Hgeww3G9iKKRE4GEFC7bvUTS+NL8wRPNv03RnMtI0y5f8Gch
amUFKNYM0hf4ncTM8LXUt4x6uKYNZnmMdb1WOh3eoXoY/wYKn7LAdtuVOI0xDuTy
UyL1iIbYjoxqUxe/llog6vxvxGPwDO+awEacQkYQNWnxseUVVpZclyCyzcdP5UVI
7zqueU28/U2yWWqdPeB9gVZ3aiCoj21C2xyQrG6tQ1QuBikivdlWx+KlteVybv/1
qQgNct71CXJwJVtHRa6Trs6ti7Nk45NMcN1rW8bvfKe9eDoqcBqIDqLUcCkvOH6A
wMpUUrlJAj1u0LNcHOYLVzsZ2qMw8YJTaV+njqm3kDyf+XW40X0I+5Lo+NaW+GMh
F40wDMYIayr8pO8uoZDBMduFZf8Iji7HL/KanKY8DY52C11+gRmGjSfzEbsNZdZ+
vwAP4Wfx/oWKzg3JMPdhN1W0GKeFwuH1RKnv+o9Q7IH8NR/0oEaFg9wSi4NCVazd
x9zrshqtW37Fwb4j1n+wYrrFa1rQ8Fy5jea0YyrwW252t6LvbsvpT0RiNWpvNjmg
qtptTQzvuDVY8RGg04zG/NGs3jhVjWHgRpBoP6RJj8zgbOzi+6dHwh8x6qOJZ6Ri
KO+K0QFDLuuDaiIDUKypHyMJwwU8eJAcHf5SYCkWnr1UsgOpXaLbDuw+XNX0RkYd
r/bT10P/B81yYywqeP8mLESdUXd8Pyq7+AEAxSIpL1ZSDaj5xb+jjYYSH/khrBo7
74+5cd1LDgweQ6nbGQ1FJIe8O+ss17QGh1EeKADz4S3lGmINk9hNYEyxWYh1bK7K
hK3XSXyPrxCpjTqPr34ujao7Tn2F1N101zHYtVRiKAPBdVHzVTWyNKAaDBofnMe8
6UmO2bYMAL8g8kJgD4rzLk+77AseFemStJIO9BB9IgSR0kIS3EG4W7qw5PJ5pb3d
W23LK+HsmMzDOXUaOSTaULX7pTCxT7MCrrf0iQec1iknKUz3McGXZOy4xwLdizX5
vurNlt6GRsOZAVOHBKjvQEZnoBsy2HgZr6F9jtPTPfyVHJv2Krs/L63N8sq3Lyzd
KsEj8qOseZCldsvNVhXy2anRcCwneUKQDeSJ+pIqbjbGdMH95Tf6okdQRMJZBb6R
BcN0R+qwiIkuYMrWfey2lc1crEhvhxWhXKu9Y4OAT2WU/E0f8uXoZDgW7co2YSYz
VPwuHRwP1K7JOnf1WPP1PqUiFBGohGIFxpn+zOs6Izq4N4zmPVTeeVCSwE5hQJAi
kOPSIhgFKO6nFI3gRTW729CrmbxLTHSNepyYxo+Tu+Xh5/llbYUgVDSdL+QmHxIa
9TN91zQLg6fWS99W8hdGB9MmmocbnYZu5vTG2AdSwZJb3XbWL14RzNJph3Cs3WlU
WLGeeIC2+9wweDcaX/B8/mCUeQZDRc3wEpMpCP0j94loajl/7PNrhSpwQbckZW/M
RMUOjc65i493ke6IAjdvDF2j4cJV7KT2oc1i5KnZJLWTQQ2DgPZoLJ7X4hD2qhFt
vMRY7gJWoJtcopdRSw5TpT2TzIVKAUW64VcZBAvy2r6CpuW0a8y8erF2/gJnEYjI
+UqE7nTWgstyZ7GRYZn53sdBFrd8wmyFLYwcKGVdhN6PWFQSLPcPFqHFLWZBdVjQ
TJ3CiYhbhycORFnnHcFCyUkrHLgn7NIdFQ3jQDqWaXGgoG0DV/kFWXBH6Jf+RjQg
8M4+6DXfJS25UU/5yFKIcduyVQNC/P0kEElD1fF/nLnfZ2tX//rlcDfDsVKIUzug
GR9rCmfSAMQLTFjTxUBhzm6HjRJWVqkNDM+cABby7F+Yv5lrag/6C1WNUpx/G32c
2sib+UN5e4/sBOTV+ju/aheduSavXYizNj6HYaKGY515vWbUiriuE3j8Um8jx+81
7Q1RvwkmRGGAUXCEZ/W6uiyDJckLVC+5xSDwJms7KPrWJYAwfDcOo0IK9Vm5etW5
ZpSWdBwYs9QhROatN7ia15UrsU1KcslT49ltjU9jbfOn5Y8+C3s+jqYl0REXiL0S
3+4r2aWbjZQPFBCU0ozLPAzWtzne38XIyrh1tU7VgIaR6kRld0+NNSeizQRaIIrx
9r99TiUyKCI+u7nyp7XHTcAD0ZNUKsq4ICHDhaby6tYB7Wi3oWjdL63XDLKDrxSx
lDY/t41lynmHJCspnYr/qPm2VkAzVa2PSeMZuRcZw3avagYOY6QsoR0zwzXrheiR
WI9PuVU4a+jDyIRAvgM1OhTdr0Adnkcc6Mk9W59NCG7Lradem0Hwk5ssF4vdfpr4
9W+2ebsZTEEHreyFjOF9YRLePHCCVPpUYKpp3S6xR0/eV2FTLm/bG2UJHPyN9mwN
i4vtPwTR32EQfZ/Sky9KChaslGxviqQF8A2snpTFWmT03gQex2qJH2sRBqmRdeZW
eKvce8aR5NvsEOGDvjN/MnEgHT/gtZp1O8u+nGU8qLDYppph5jNuvD/vMxVMucxE
SIlJFZfATrSzm/WMoamioOdGD2toF81o6KPnnJ0AWRevmi+qPln6DehSo/JHdSYZ
n7lyfzSDofcEvs+zPtuXbsWEENtuUUDDz5UU7jQCqabXA0pWIAOS+oYqIBG6Tbf8
ZEL0jTJnxaS4jfpQA7MrJgD7SLVLwWLjkxNJdw4gA96OkJkGWu9BfVJYv3F40diA
khnjXgqHHh7G3TPAnXly0873uhYn5on7LrdMEqB8qfRKLM4NF5WqFugwbpF0Yken
6iyk+iqHl5XsKmE+U6WQ1eXQFnDN93h56r32SQbferXTuOGxsnJmNBp0a4UtTgYM
iGdnMRF6O+ROMz8dfIaoI5dejAqRLElRLKbyJ17OGFss04k/s1aS74yMuI542ScH
cRMkEGOZRDqMcWWydr3E2sT6enuZoRer7Ikzo5NCLfz6iXdh8h7sxTQuao8CfjED
7vVwkxx+2qJSR/yeKOBcx09BlM+lmrwtPl5qrXIXEdG2AhkWQ/T3x87NEkXzMwjr
jLANO4zO4iwNiRrupVQdx2bqqwZsV4LGrVHkN3DxLX+rxRsvimqRRWEN8m9qsc4w
+PEMDuU4PFMPL40QVzwJivlW69YdBrmhL9g1m7DQutvwngUl5RRguUCAOXaSZHHX
BxbHAlIIsHq8KTPWNp0VFpLjxJmhAok1c2hSyBqciI+9qb6EZquwOABCtaD7M6mL
YzG5OCPmxWjjCiWGidTBxST7NcJos293fYUyfUFdDCrizzprFnzg1R1Jr/2gdYo7
00qP7QjxGmJ2Il2+3nzn0ssd7hL+qRH/EXgE2tMrTuRAgmHd+2yT3eA2yO1bJSg6
Uozbz9FQ2mXcDOsOBzSfu1+IoNFjDHYYnCo91ioRQlBST8J3d6gaQ+3q+9BTpqm4
OQ2SD1RA7QJE9FV0OusCBCrHBFI5hpp0+/IEHfql48/BieD3tif2RE1cZNhCHHsD
xQtgyot1KFnq45UmNUHQKBr8/OCcCZOGu43qbJnLsxupAzjFzIT1kcFM7aHNbCNP
5IEpVm9cTxoM2DSsxt4cbzdyCJ3ZkVz+KKUUhgwtBmNsB8hgTn2Lknkkq+neE5dK
cl29/S2f7h3bEkrNmutMc5LNmZj5AqHQNYNWwDOE3d11NWX/CU77W/oulZu3z/jo
LWR/tGjyv1bhG7T+L/O0wEJudrVZc4CYyzO3b6ztf9shsZRzc2kg6eJNW/DjSkqT
BNqXRpkajhkfabFMprBss9NRMcKYHWeFJIWrcvX0J80gHP8TYMowA/l6FFIygYzy
I3tWbUIzFVYEH0h1tabBmC7DWMIPCCd3+SJpSUqA5SaQdxhcd5v4BHy5o3F+iFVO
wBxT0PB/v2pYGpVZPpBx7N0YaC2MKPNDKi15QDQI280kp74OuOPLZUKqJoluMTtp
GFzt+j1rHhCMgQT3LRH/B6oIwsVNOUhDUgiU/x0XISMfUEHOYkA8+u5tosI4NI8M
iuGnqY4PAqtXA9Cfke/eCEB0gMC5AN8P8r+rqOf/+2qMbW4dJyihmM0sVMMEfWau
ebrEZZCjoPonD2/D8NRD5DdEGRwZDHtdDS7jKScfEB1b2SlbRCbBhDhDPW8IUhoL
sImsU7vmEMaA9ZpGMWFNMNa4i00tVttqHAUj9GAC54OztHMjbhqnk+m7NgNI1rG/
XWzCteScq/qHUkQts5azSp4kWIyWGX2IHZd749bfcRLbo/J7dVH7hYkBx+1uwZ0V
sWo2skt5plLx036Bmc3sPOuvsdGhBcfKLHmhsfMnFdOjXb9bqEhsT7IO1RKH3dMP
ecezA1g9W2/ELbJ/FjuzYsg5KYA83PXYVjNW/eeDuiP7sUt2ozK+atp0zCZPJ5PT
/MN63Pyj72gazGVErTC53+FsHuL+easi9fe+IpBn5LaH41zXBoUMrgNDEY2zuwiU
CZdtXMIMNVYOEt+6NzR5h4y+0jRic3hCT8m1ufUnIf6R0BG4IUZnpwlE99T0y15U
3i4gFlsERWDy2Bk5y9uetFsnZiDG4l3ILkS0/zXKiBSsxaPu2VxpcBTBQEDXksx9
6sWv7S9TKwUbFhib8Yi/yXlgpBovo8m5zTwI688h6L+HEieufG8IaUD6Lh+dwmUg
B75l4oryd4j/mF5wmZ8yQxsDIW8rs3/FKfrgX+/69t322Nu7s28fIg7f5XxYNANT
yNgrV26AG3mgbo2BjF5S8b6IUp8gMT9CBB7osup07dlFt4YCwCMna0742U75ltVP
3V53gS+SK6w+wTaDIX9cBkVzQOInNn/Lh4ATYpJSuKoXMd6VNoqBZDvY9DotZyxp
GkvuC0XiUbs0OJah4JbS8eiK3m5ZTnfevMHU7yka36YVyTu8JXv/6NxyIEI+evDw
q6Xe5JOvWckoTDBdISdMoLPXIRUF2wV9JRld58WPha9JhQ6NqZSpgjd4meqNCoYS
LxW5bxwNRaMOKal3C+azG90kqSaKt8JYMt7BjqIZwUkZ4AJniYPd6otttwC3EF6r
wSQt9mcqsP9dT4A0k4MGMop4odAWce2geISNg4HyaoavhWYVDS/vtd8nyPGyWqWj
mOFWchcacIcdRbp8mvDvZVzXywcvaR46Wycf5LXNp1esduHAu8OrDHseODq8h82H
3TLFrR/4k8vK/06L050FkI2da2aTaUv/YNsaGSKzpxGWJHJ+MPD1DZhT2lsk4ywG
z3mIShrscgHDBO5gxMcrzrS5e4XH56Dftwmxuzr/HDCaQl8gn9A3lNDvBgSdEsLb
ZdYWsnjxsoufGH/rFr/2KYhiyJEjJT5sn93/Fh/0kKoDowTfF4Rdz37quTQOqGmu
zEe1oThFbJ3qHud3OIbVnz77EU3RVy6JBUqJV6CvBWRGUtUHDjeNAdGH5Qc1GPnW
ojVTWQgjsaXarX25oZ+vDo9MSqiU82bDYkVz1/Z6viS0NRH8A1MmqF7Lbg+ERbAO
kbCd9LBNts4+IvsIjX2RYCIvHFctFNqnxrKAzha8P5MBeqHJs3/vYpG536WRyFi/
+c+Ia25X25KLbRmGo/X6JaZ9kTPALNS13VU7PXOwtALkg3zgEkCnTF4hJGJ6Kfry
FXJyT9a+hE0z8vVZrN0Unfc6XGs5koGZSMe+yIfVC0TpKdgvToyqFgeX7Sj/7HS2
KmjkT3o36P26AXCCoXQu0xSAl9ugNpzNluqS+3y9lJq3qPRjm+jnzWHB9PQxOKuW
LhetNKcM9L4cxd6nP1UzG4+1jm4m0KOTzZZUmeMMUXlIK39iplfwbpF72YKl1Lym
BM5GS6kNGVfK95DhOalKgtdalQLlo+//0ibibmX/VjEvCeHFMPKsjWNcdO5BT9tP
x2OPSJ/HBjkDaN+nkM1iePSqAL/Anb7OfH6FFTr2VDkDE/AlFyzWNqskd8tf5nNb
Cz8+kWhOaiA/3LUfnJqc1uEaDyX22OZpeQss+kxql6PD4Vhv+UFdElnNMmg/CwG8
5nbf+JgviZUnS5C/bLQDbz5Y4MYeoLG4Uy870fkRRKQCaQ00jqkJ8mNIERxhQY4C
TBp+KNhbBkkSJDbxJeNnFzNQKNfCtjXWLc5/1Pr2Rm8MY5SYzoP8el4ftU0yo05h
p6B9iOdtw7OtPWWmqRYuKTBafwtz+hohIItTIc/QilVkAyQAScjby3IVoNFDRKv7
+LlioHR/SX9zv2iIp8iDp4RQz5IlQ7qbxdUJNKXR5G0vbycFKDoPxIoj1KOSWbNO
wm+WoU7l3lCws51bMtXDJgSNj47tRmxva56pdoOpEJLVppiLeGWX+dZj43ueYv2Y
q0y6MjqRiO51BsilnZw4g4LsHxTHL2/H5mSF9LAYW/IgvaYXpeP1TvxzPcRViyDE
+Urh6y8456LiuWNM135xRtbP9twInOea2xMIJBuXhxjkTIEy6iUppyswesutB00h
lu0sW5VWODDnJ3HPzcZX9//F9jZT+gmW8cMoMxDxIFJ3vMKgOcCTMmTUHFvLn+VJ
6W7BW9HvA1vUzFli+OK77gcwCmitS9cmGUf8MAW+dk07tHBQLY/XHC+MCb/0cYbq
rg2DG6m2UYI58lUF3/VkYBJP8x9ctN0M9J+Tm38Lrox6FlGT25UrAHWFYI1yS7Bq
AuJJO+YB81vu1rSTd6kJxrrHLqYqYF09pN2uHwaxwVpOBFfvo4mUymw5aaMJC9me
6Ws0wXRY6zlXH9N0zdBuOAVNyCb+/XJ3po8mhS3rs+Bw8hL5vFlYgM3SfXgciAav
cBtXABNNZsjxWXbPd5DkkOymuSMoOaZankaBlMGu/z0wj2yb0YPsw45cOopIc8UP
y+ufqtElcVwqJq6XFCnMBa9pwH454sUHdFHZjvQJbphLkOpzTGMR4DhIryYxPDlq
hcQHrvHY6pIYk/J8uUrICvkx9huWSP11rNFC1Db5Xxmd0Rah1q5JlHxr2CQRAQLU
KMbCDeFwVeZV/BI+eE2fEsIcpOx5klaEpIMCjUikVRphsUWHCT9C1k9lhvAyqSyH
cntaBENDDOMIS90a6nK3hcPG3QgSq0aYmjZUFC0w7a1xwIRLi47POpiJQcceNrcT
beLTOw8YZu4E7VFu0TPFK7FDgxosRJZ+I2SZ1jGWUevHJfoWO1oOezNaMtoIbdRr
wP4Oe6OocAbk9pNAsodtynyDtXDjLmVK4zaaf+IxaZvPJiXmtRCTTYOuxEbfF4Ew
+DEKyy+WwnZLLDyB8M5MmxNPeBG22m+HmyLmoiGTdeH/hsnq4R6VibgEQC++sWeA
RJuzWTEg6kcEkC0xxx9sw0t9umFTTGJoKTlpwh19opXhFsce3bQAsdKJkp+T8+C4
AJ6uBvMUZTDZTTWYvp5mbNXsHuyOQk2Ks+L+F91r3vs/aw8aQjG8LA4DYfiEFDj5
rzWhwzXXgBfgR3ZB31YWIsv7tmvxVTlEOI8T06Po3BLB5T5jzHqZmo74denLHOrG
xAOMqrH8b9XoYx/LoHjCt6sEZTNAQrFUkm5I0/oEJjdDj63RdteoEO/m8ZGJhUa3
2TGRhbXz6A07QO2To9JTTNEFlwZ8QBaDs8Hffyri2DwmAtkO8+Z50RA2Tmbnbe6/
nnrBLsdAfcwyGcRXHNAlQF8MQQXxpGPquDffD6CwwAImKxP6rfQjtIj1U2TRdDIs
DWk10KL22ZzQIeewCYZe6qkFIaPgQ1PCLe7VgEy29qEinpwVwfDc0vSoAUccOOBF
0w1mIOfURSCn91V9pPo+lYLX6m3ZPeO5yoc0Yw0jNgRw4HTtUR8NWSYqq2UGpGDH
mrcKz8tB3m/JQCXlVQp9vHeuMPlzkZpYG7ZFm45ZAB8ziFe93/OEkPcHmU7GKIu/
pIi9T7X6HdTzTR01N4bH4KdD4GTlWY0+yVClw/1Dsrut2RqukKLkD+WSe5k54qcq
Ft1rvjDtXEREhnt9pHhNXb5318woxSel54TypIs1bXB7Ij/LuCw//70GsSdoG4iI
XkcenmCSer2+aCfsbcpNewSlXxZgTIRzCLojnjZJq3ZiqeM0hHSrziNp2Zlicfyt
4A+3zlrS50rbJsXQUHivzg==
`pragma protect end_protected
