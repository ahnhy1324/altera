// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
A8AeOFX68e/7teXPgW6BIltU+1ZEX6J3v3KhBeyIqvc2oVWHqO7G9o3Ow3bvEqVW9L/qFDNBh1R+
rJSss7W9Y52O1XT4frlsseN9pf2/TzL87cWMg+Yo/UkAwo5AUSIvDYb9Xtm5KRgvqLoM3Jvu8S61
4fDNIM4Ms/+lksnWjRK/sXUzqS35lUt+M4vW76OpxgWe0Nhyi09ddbiwRzwtH/N1KnFCQnVWdzQ6
QT/SXc/OupjZbFHKmzAlhAMx6Rj/TVXgNpNTtdwC7W1mKRhdTmYTAXpGEFtdlLxNp8js8m6jcuRa
8tGAiDJjLBN/Zdx8r3l6WuZyIMC1baK/nRuRAA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
mYvmSQITmJqZbUgkkdjbPa41iVhk7jPPMxc038aDlESTfMMbmtlu+ZzqHZ53FaYqdjZKWZwNl6Qn
tSYnzEG+8ylZeJw13cc/azNnngSq9VIuDTGtbQ9zOXhnPLQR3hMJgSRSQ4PL/SPuEhNuf3a7GBXl
ZVVS/EjPjsLRkdnR/Xul7kJ8T/2y7BkYMVLS4efqlLgAfnBzU5968C8wKKatV5HH5wESFv2Oh5lQ
cyyUrsxXpb6nbr+gBx9rPViIowbIttj3zfltzCkgg8VwFeSvwDGIvQ6QvGJLtKsQomfsOk5Unkkj
R9VxN94XIiShVFvfgIo4/zYMUdJ9w/Xwb5Q88DZB4h506mNT+HmceF+itzn1LbvhW7DPYovyd6Nh
LNzKnDamUjnks3eb3eQ7XoyzOPY3XvWh9EGs9j3Y8lQyx/o45e7AqqqMkWlXapAoRGhnhz9WLUZV
0HtYNW0bFf9pDnxSUwugyJ4h8puStWU7HtcTTLGub7LLo8u4LsveugCfYR7Zk5EwmXk6RVC7YCM/
1zyPZxVOSOITie3gvm8f/4RjljUd4tUKvPG8izGBH4IsajE/7iFsV2qk/79AfNsuXJY9EB70pbKz
fagcrrBSee5MgWo756HHGz5GZyCMMYemZQs6iNjGOW7kBql+cAbL3dS/PxRy2bBMBB0T56O4Nwzc
Fq+I4xG4B6bTNBqVaQ086faOFL16Ijjs72pEBRDwMgW3Di07Y2iUpKVSekBr9sDKnX6ZypszjlEB
+IiYlgSESePiH38MZ+Bwibip1RsCINJE1LpwVxQuMb4z/ZMvgK1ov6scf+y+Yuu+3uXKZlA5xbH1
uyrB8hHA2FwKwvVfwtsIn/AIpCxkRqfXMu9nS6OGCjp4MDqLKbj/apMfCHrNTdNY6UR3b8LTh7jo
9bCqQOBjsduUfd8qRqO7eqA/KSkziIGI7JRoW8PX2ZoHGTEoGmKhbHinVOFYgXb1B38g2hRoADGj
MC1tOjHQo5YM1BPLnBtAQggR5/XMSuhX8xqr/PYmIHacmWYR0hM8V4i0tbw7CJMrZ7D7VuQkNhLL
Z1kaxqG+CZSjHgRhv7zcYkuT9Sv3lSZgU6VshVwsyosBIyWCdrxZ/YETXX6XAw9Wol6J06bxaGZp
f+5LHEoJ864byn8jIqEvaZcILL9qsHBeGfPvSLJbeI2Fzh1WOTP1Y2V9dwCLl7hp+I8IcTy/yFrM
ycrVmct2l1lxjNcPA/yVPwbRYf+Kn47O+qeDlbFaIYtEx5IiEqcud2hld9UbdS1rJpHOoYf4ygl3
RLEurTz7HGM0JSnkWP/TbovU4njWXoVUAu9FXlLS2S+rKzSLQK5Mt/yzvK8fZBpyNDln8whG8Iky
uVWHTqNqF4xWc1lo8QgVS4p4IkEtp6Hc+1NXoGBCM/xgHUaH8loVVtNFcKr63CMIZ3R2nM4BYcMt
c+x2BoZ+lw9+BeEEiQ1j2FH4rwEK765umFIAkPnCwQEV9phf3uVBLuQmXNth1SbQAn3vGhQ/YqWl
zvxlnjIIQbPbB2OArb6eQOcpMdwTLtCOBsLyAWUlN5UzZj8lv3TymwtF14A1becFnfLUI551lUMr
LrQFL8Y9wPlTl/0SsoSpzBk+x3Lkn44R5R1oIZQzVsq4N2z52q7DD87wtYZnaKAZ8m6Xjah4lAMc
LMpEO73CIGKQeC+tKAT02jD1h+sz0gG2ySq1Q4u4KxWU9fPa6wSZehqCFmypMCguKsQUxQrH/XDD
7dA9C6bT+K19uIn21ENoafOjoOq9MzwLowjT3+F3HkYlVKbjv6qFYECCCWMcQe5mlxozIvLj/8o8
vMfejIPx4B+XnvAOZBcCcQ511ZMLJ51rMhMw3s4TkYSodgFVyx3aJ++Ezi7It4GciePP+px9surK
YJnsRBo/5rQuVh8DlXFreBGgkO7gQCYqpSs6X/5WBg8Dmby3IowkH9bwiyknl0CVCKA0lRKIdCj2
SR03V5EnhDvGoydhDQghRRqd3R+j6eXX6E5/Z6YrfnxrItT2upALAa563p98/ZVb3Yyzy/51SuMm
9DIJvtOfWgTwWQMNKyZnCvxefghgzNqQrrIZyoqafjBAmy/iaqmmU9Ef+5LFGAz7kseouTMKD6MQ
RZa7Mezy3X5ZFb+I8fVxSJi8UUufVOY8MshvESptzJ+9ZgRR9wgDOr8pQqFrxcNvnI+EDY9P1ZVC
0GgNRgx124YecunnwC/bF+s14q1YRwljJwFLsl9i6thnsepaftfbF+1fx1LiUHkqAj37ZcZRsSmu
qdUeHlCkQm4OxrBzgBh35UR0Me0oHyDB2IgC4VWZDStkZeLT5CLMBDh9jFeiQZqJ75dCCYZrUcVX
BNTOdyXIe67USGVEpwXKBYzlB3y444GaOMtGye6WVTEvUPrjhxDB6vy89Yjc3joXA4Yrm7RvR27n
ijzQuGZOscpN7CVebkjA4hajmUzeHDCIk9MUerpRW2XJgg4c4l9N+Ppt5yBH5aD7gPa5yhICxrry
2KWatvkMU7AQ3bmNQplEGPTCJIsRR9muWMTg+5dp3rBpZ0RYJzMFIi7LjR7PTgAzmqZsbJ/WKyMI
/zbeYCT1o7TCOcoh1Xq1VQaXZBT8SnYab3xA6dXGfDJt/sF5uuaB8uPjGR5etuZ7mDX0mKs3tGZK
AxNGzmk2QetHahCO8gcbyOFDRph3Fd3YXfMHDrwOxttQqyOeff2v+S1H/zGdUNROBvBDOrNVS6DU
edkS01fQSlsYDX0Y8+W2lWSVcBecfb+smJvxC8bKhz/0YMes2XkJSFUI3bD/0Vff0MnI/agWWNAh
NMmqDkUH77Ub5bZ0kuFxrQeYKcOlf9UEezW0Qdldz0NhoLyIQbDXMFmy21I8v274JFocWL7ujhtQ
AfLq4C49PPQCMftfW31pWwXDYHdc9d3j9nuVsm39kbwydhmZip6o/QWbxLHeLS9AJ4/3EQXRS6ln
gI1rSgPPyCLFnJmxKNorrdEp4ziQ2hGXT55BbVpCYGWO8UV+1c/XFzgG2rC2mB8RK/Msd36JGC7J
nJAO93uEMk9nioW0T0XHvuFe5U87fVXp4sgim+HmYtXc3lP4BoCT5FQyZGPvtduWCLP+pfAJQ+Tr
NGL/8ETB67NN4RX2bhJ6PpbaEwMSjHMyfzVwi80s1UXDO1BymVeql/qttSt08a9XiX1Cap+O+iAQ
swRFV833pieBVj4Y1+jlWaoA3/PQokVHX38747/21xdBmBHj7Y5rpeBbRCwja3U2CZdb8ypJkyYd
kVeIokqZ2Qz7k6yAXBxlcZ8UfkGaNZA7utrMDAriSnBMTbMRLs7PotQVtzaklngNDRggdEmPxGTj
QrkmcrrySc3XCdx7JgYV/Ec0GPMvJOsUXEWwX6xxhRwteg9xXBIfRpxpsP/2sNEpmqM1Wq2n4dI6
hWt52fbnSEexeame8hjLDMJp5SYoPC3TNmjkf2yWyxHRAvhky7JKPKRX6oMgybKbO4uoUtB2O8do
/Hw/e2/KFJUENXadzmSU6Br4g1CZLvdYMZnZi7ChmO/gtKFtbmS2rKjlnIAzLlUzO8naXkeeo2WB
BU7ln9yaK+DohwArFfNlVBR0neGE/ITgNJ1mCNEZafnCNwiXih4ceo4DKaEDiFrryuxlak2Xy8hK
XWEpd9L4GyaJvGguTXcm8rvnFrYsAJZ8+zxZVn/dKFJO6CUGf5GMY/Dcd/AFRRiR157k4zPIEeX2
8JguTgNiSfV2SZNrDuJaC5roZujYquIL/vND/A1Z/xYJt0gFcc4FjugEqrbSf28UZcPBxQZDCCAx
vnlwoIMCfjQfdWl7/miB+7EJCG3NqQg4jmOrjz2MBwy5lu34ncYCBe5ZsFF+5cQbcYibcVlQrV5C
T55J/eFQFDcMlAievSyx5G+0nKH8a8O77etjRtV53E2uq1zrkrNm2AN5lQ/LO7DJOCROjiDFUPpw
ZQcjGnhETgIJIGT6SavEia06I3Or/GBL/RDwShX6roG5NpfaeJdzcGx62FbqDOzQZwpmzwCFlngS
ZPD3djCyPgkPci8lQdlPcJrt16FzviSvFoE5PO+sCIYlSfuZku3qx8eKACq3biSpymoFe73e6I1f
fNC9vmv82iZrZin61iqaQqY9aeqOqEjG7YzyJyZjIRPZGXrGT3R58yWmIthW5GJdoqpjcTWm3LeK
vIBL0f3MIvqkfc6kbdjHm8K1SbQl3inUULfOcfv5QPMyuh4D4dCj9c/lCV7XCDrqKb/5iQNJxOgs
Q+l/CJioKmGdlUL/U9Qsm2yGA3F0MHXHVjuLCv26jE6Op948vxBndbA4+oRnbzrJFb6G9vUFD3tZ
D1Hyye23gVckgU/jBGoF9Lju5JiSdvlWdrz+BCcu7bebgojeVMVnA+Xe0sEJUx+DBq+Ol1Z+JYRr
prN/HfAIDCuMBZwo5kEeLd32FBLNsaRECiSrS733Ck0hZCuI+NRbqVbaG5zmTwe9BYxqCKWR3pt8
AnM06hmtrYfZjYqv/7VS/J1wjTlR1srtCK8aTi5OTn/451o0vNutSvRgH6Rh+s1/EMX+NXuBjj82
5Zs4pVOh1T+9V+v/+AAP5tcvkQuTbxMJbEpy9YbDfLHGYC7Zvvvq1nUwt30ZO05W69TERRvIMWzg
sN8DuIZWhxpK0lMJ+b5GSfVp1MzNpAVJgg3USV0JGedou9dI8fRYHNe+z3TvvHl8zPyHCCyBG/el
DbOJNqnHCbgzE2MSEQ1DyT53QXIsCPwJZqMMt/kn3/wX90NCold5y3OgAFs2kSdj0mLnKePZLKlB
/4PEJ8QnWWGxnYB/PGZkSn4hiPOgPEOftdufOSIksHTp6U81kB/f8Ngcvc1Z9v3ZdYJpKAwDy3UI
q5J1RX1rsgpxNzXnxV4RtPtHgTrppvglJEy+kYQE91WuqqyL+5XjzDq7NLmMxCsPbNAjZiL+49cc
MTRGx/MT+0/zY+a9/ZAE960Mk718UeSvP6TfHqLzeBq40WQOZkSJrp2iafn9AY2PIuMsg0e/X9E2
MB7Lr9abEucodWqu/OoVNrfnzzQB1Dde3uPdeZ3YAavgdAr5NdtRiATUFlhaoDKaozS14Wb6o+QS
GWx7cfvxkrreXquSZSyuvBemxYtwZ2VRYDxnWPSZKVSwOs5ZzYs1C+a+3nUkBrBmgjdRAAWwItuB
FAmuidqZ44/zGofakHFaFeA6pCopYfzTyGa7011ePIu4HaxFYaX3KJP5zrA7FSSInOtfT0FpaWVi
1edP3PT25xieX5au2U/tDBH4iixpLQTrtK8NqWFATqQALGya5B7yYPe3LcKypv8Udn+shPhXxcPm
ZKbbOkSjurEspznnvAnh6caUlfylFkvFefs/NiwA11iUedRrCRxUyDSpqjVp9V9TJEa7KTJK4Etf
cQAZZN3BM1WWLntFVbF5JnCeKFGEYoUFL+AUyH6Rsw4ZDO5qXK+MwTb3IlY646saigohmtSIAy87
dKkoCwIO+P7q4a6Zo/MWsenhvZOnVpuKM3LQnKHhvk2+THeDmRG7P5P0KMFwoOOiL8dzcqd/GI6x
pvKr8bMBKGktfPFipSDjQOGyB59gRZVGHZqUMMiilrhXtqj/+EOLyvsCB9iUpMdoidZaf0gkmeI0
IgwS5Ex0n07FwKq1SHAKkzRnVzDbLEmU8txqUA1dUWOtYwSyPDjh8P9j41QnkIdY5d9m9lTlfHxe
RsyZ57Hzh0oiLEUVhcrIIs+Wxm6WCoJeZ0Qw2+QgeuubZ7HcprucDnQ02HfLIi8/gG8RvvQYxJ9I
uOCDDAkrYxeXQR/OYpXhch/XGjPdxEkYFFhN/KsQIJ5XxNFneUoarNKDWFGxjb+3/L3Hs4bT0dc6
hiLJMQ4Y8hGTs/YfEWVdocZ04R4+W7rvwt10aC69Pts2Tzbz/v2Y8Ro6OdlAjka5nAnXj8VJAojI
uixBQNpWE1s/FbuekQ53uMAzTMN7ExsuA3ujhl5RFTkXx6/F69spGfXsYr7nx4by4RV1/5ZcgNWY
PEYZZp8nUZW1wUu4SMF+iHhASS1QneDIOUfu/t99eq/pIvcF5eWSex2K+hbxcc1WV8fGZqm8Werh
IoMa78oTN9QKJT9CENKuK7r0AX5ITF8qhiv86P7/UhBDqKIM8fzEVtZSufdJDTQycJGcjQTROAFY
otcpzSOmjWH/5hYfew+q+xzQqQZ+wILOZg3S2n1A2XU6eihQXTv7Bl3Kdti0yii0aijaduHkgzOw
f4j0aEdXESBkiHAp+lgri08fBzV3FhWViXYOY3gm+bDMnrGup16b/eSH5EdCwyJMBOFtzBqe0N6z
o7YHqtZyZs0f1pzdUolhMgd7WqQa9+38QIFV2023fEmKtFQ3cWpnm5OCW7zVzmmIoo6h6vaOJtDb
1qbh3fA6cKZbt8FmJnTLM73Hpm64OBJaBSQmjkVYisTiCurBbffQbUl601OMUfavj7Kh/YHWCc0P
Yd4KxOf7tj76byAqijoTAFlVYlDlQtH6hqk+gzVLozs4hGYfsAkDJxq6CR/7h1G71xW3MAxRw+NI
Dasx8pAkaLSGqDs5uQOy5/UbHdKNf0mF9sE/iNLumhMajw1aGQqfSUacgSxmmN5vyOBYbWzkSMzh
frmdjo/QfOkbDDwt4BCmtQVaQlr4kfoEtO6MmxegI8bpPCMLC0n7bNG9FgLU094nd2EPbiY/bFTi
GkvY4DkmL/ozcFjRBP93h1JHvToU5b9vWbEzLLbHCZMrt1q7EVCp6s91dX1Gp5II0hILeZHmARqG
xcuStOAwN90Pc7csdnqbmnPEAJxoo4ryJ4Pzlq2hvnm0IlCvkas9ghF0kAIElJ1NqAB9KA/ziNN0
cyOrZ5lnBGjXaCvH1D6Zs6YUWgTN5tEN/VZJfCInGud08ZLM9b2KycuNuemGI4RagpAOpX91XBaN
nrp7NqEr7bodKdkGcLiU49GBrn5lapmYH/YPrlwJiMEuKu9X+s6C0eadd57Dx143ek8A1aQ8mikH
tJFcYH0CYqYt53n5+uOFnx2C1XDRlfp39cZggauglj2d52rtfptmubB80BB6Gu4XICfZ/fAhCbdh
dmcO4hUmApAn6ujprmoNctDw8t0Cj53jyF52mns6HvkYrkusF1i4mB6qCviXzDF8g3ymSvHyLEMd
7keUYF9VGcOm2QWxpYLpE2LCms0G/NHf5lgWJec43gfplv59sjaSvDmIOE6qfR2S+g4HwJFxscd9
xmRbTmRoTAQZlcna+13LY5miieiDtmvB/itdIp9zEfGSQjFaPUvwBn89cyKSECrVyZGXORSSr8Of
mxj3k3Td3fKSrt1e4vSC/w8VRo5fp0ZZ1yHZdaLuOYJOoCnpMFKXVETz7lrhP7XOgBF3XDeVENWw
4EaYpRJmHlW8LiGjrkOV9hcD5HBOc+nc6/LS54cB7cAjOAIvGpGgNG8tq/ZJh+eDc+L3L5dagOo9
HusFC3ylZGGqBN/RfYILyt4+BI/DG0oMIGn84MOFN7gJiWjE378taTfd94suvGs/rQ5LTWSu+jWZ
v+NmWzvmEfNrJYKYxw3tu3jDyDbS1HpndtqKV2Uik3PhMX6W9/ScZvPBjAwcMJPxpGvDzQn896lF
nroUyHvkEOZv47VgiaXJ10yolFn3gJcTgDRJJRQLcXg/Q8we3JSTKHfteowiVW0j4I5psfsuaI5V
9DWDnRcZjean3oH/SrpvOugVgDc7lTt9ljDPlMWuVKejI+mzJq6dogQ0zH/K9ZIGjvR5xd1dcpbu
rgzRpqxf+dqjhEP2dHAzYNMK8TMRSNXlopM8Z5UajpFrN80DQ7QKL+WbkuhE0YH99xZ8cM5QmjtK
vnUT3UZb3c7vqMkzwSyW44LTn+6AsU6YRHkEy/JIXjHxBIUij+X8n+UboJb3OsGEWLTuCaZBkufV
0CME/emK3KC1CcZ9I/sZjwlwd2Sav//rySjyfFDTKritgHv1GPtZbODgI7yMl0KDBNbMzUHlaESq
Uy8tWwrTcTWounYiT1Cn2JLbLymvzzU3Kdp2iZUhz+ZG1Hugu/zkNu2WMcUUuSB/+LPxZyEsYNce
mK51u+CMcMRBWukGW9/CICBcBAmTWZsIH/RBAqxKtMIm7LvUg2bqJnz1T+5gm8scSIQssfStB3e+
Pu1hn443zc5DnfNIMdTWAWRM8QmehduYcbpnQh7kA0q48jaCp/X4PhTgigH2aZzuqmF+ATVd9uJt
k87EpzYAPug4RFTgsYjN44nU0UKNYc7ZM4w5xrSy4uQ9eQQaIGpx5pX9ljyTkqqapR16RC5HwSNg
3Bs2Qaa4/nG9BvtIm41Y2+whXIYgFX4yrVX6Ofg0gTm/GCU5S7VJcYuGNMLQuOKFOaC8CcluqpO7
UcZh4petH0pqdEtjR31AMhNiV/eeAIsiOGpCEEr3fXBCQzyL2nfEbjQqyc5Insx3RxfwiRhgGYPV
N8pHhDfOotQ9RSUUTEl6WTe3leD/q/RaPNPY9j8dUsPj07kblWMAgsEj0Z2tJwcnOipPQt3loz/h
kpjHzOSt/zH/ag6MB24+6kSnfrDAc6Lx/uosHc6lqQDY9m8Yrhm5ICDtLpLtx5YJDLT2Z1qLni1g
fW9kuBVdLmacs5y+1IHvD4cahMAIoanmQISm2bc+KBfUD/+KKCL/09pRveI9UGmTBdsJuilOYQMk
FMomR9U6OAVkjnO76MO9edmapjoA6gHUMBh0mrz0EXz9622TtwB65krAGBZHrc/y4WKvIbgZ4r3U
5hhRdB7Ecwkbqtn9fmjrGsFGL1wKBt6BP2uR63AQApVyFxMiqu8njYpfnqtKhuBBvTGUHJt/Mk38
q1XrufBo6UoWgh1meaaJ8s3TCW7g4UIHpmexbUiVwRJz2e+HAH8e0fzYhJVvxX/dlMGX9YvuxCtP
rwz/piLA+zPl85X7KbF98PJeOJDyVsWxLlLkMiJNNxj0YCbwpCq/mBccfNZoBoseePoTJH1n6KNv
pvLcUUy+MGkgtZNDHFFoxlBb/PprlUStx+s9EWte50FVyQG0+r7ZHI4ncxjWdmrMWT+WDt+JXTXr
tqNwc0W9fBFYcEe4/2ZgfJlsy18VYFyLaQ+qFhO7eGJib6+4c0sfGP9SbevBTqA+so9Z27ywmJYe
ws/tAq8ecAh0KVW9S/xIkL0pIy7H6nPtigMuc6xq9x7D+sVYS8ZWZevSw8EpmoiV5BA1V/OLXa4X
3//mjcQ4aefWxLx+H/9fXsSsKkhm8JdU87mpdTcAdmkC9I1bMkJQxcmiyQzcJFTTnph2OK3+opxL
8sgXPAo+zJY0D4p6THEkHU481q/VIFqtmEpOUFuykGLlStD38Q4T6AOU25hVYC0N0EJBN3ZzwRX7
Y+/imFtqNxMHClQCJPfkgDCA4f8bydX+iXWzvOtxR98ALe0L7C2ZfTubg8CFLQzZegJouCV/IG5O
XiRncbMSACPJDonHMjXg4vDtL7gvUSYl/qlfiM3PX5sUzCNKcE+uI6aiYZqDd31R06qp5jMyg8vo
E0aZriDc27BN4OI+nWB2lbGDnE5OVjLFgfb1kBkT8OlWdxq9qBiM+zkhp7DQb28uhiEsHFV1vgpi
tyYBEKHez4PBfI7qn9ZySaGnk9pf0NMY+MHgQ53IJgycWStyoSop09+QMlYUmrKhzKY97av2cDsW
XVS+OkSkmph/R/ZbBuF3zcgkjQbPta3Tkk0EmyVMQhUvM8Yc7xXa4FVRRuis9R/3BMUlDCR1RhKN
j3eLvmSEcEnoWCwRn9cMlGbm3nYyfJCMzxUXKmvBcrZWdk6waba7i5LFTZMZ9s3Ouz3zgmpbNls+
/NmS5TgviwKdxdC6Auz9/3DoG+BVSue/9pNK+b5SkKcEJnKt82QDWsqPUzkwuSAi3lc/cwTCVWdc
1WZTkcYEozQ6WaQ/UyJFkOhrlhaMy4J0I7u9Fkr+rozB/Gap5C1zcN66bS/bSlpE00DcMVprSFwb
Gjb7qYgR6OoqRJZz3xXC4pUk/EgsZF+1yycD7N/LvIJ8qqzuoOWWwRYiL2Hkbrc7lOY+sGUsJyns
veG3et/XFk7LAjjWR76hpFf6XXW61fQb3DDUqD92nrOx9jSFK8knAbb6gfKciHqgCsY6kuJbDVGx
IWbiHr7DgWXiWKo1hkvWDoLMiXvC2GKnnDAEXLiGHO9vjI9EiYknvCxULI11PXXelZ5WHIIQ+PiW
iu1xVFOdHLhU7wYHxYlxFgihesqO6mceVpnRb506GNcZ3HsmUWU3pm0+Rq5D/LcdOYier8JVL7+E
vGfGd6FXOC7EVEYbYodIlyF0/k7fuEb5NotpbtHEdimM4Qv5suCcRtA6rPWt8qR2KKqnQn634Ktp
kKbby579rxsef5VMrfXt60xy9Wjrs+DwZqJ6AjF2hsUwIDY0gXu7+f1Bw3tXlul4jhnHOYOHK118
WPzW36uyPJMgNZdo0S2o1ZZ3f+uZWeQpr8QNYt4rKxE7gcmspjsKrUcRis9FnYsRsbcsInVvGf/Q
ocSHP7P/NAZoSHJXontx4gvIvn5wE9QAfPU1TV5aMUKeqzaEnGKrDOZrVeARnkSnpidBFkaX9vWD
6MfZyHEtRsaKjlawX+H2j9M52gGC7rPQHxDwz8/xGC+fyA/BOH1O48SplXxEhHNKZOwCrPl8/N4I
OVtN3Gk5tjHBcjT+T84/Goz8jlXCGSl4dy1/e697zgp3cctg5Z98wQZo5K1bWE7vr0i9ULTnbDDZ
bSKe9CEE1KfeLyXzVbHfmDD/PxEewMSADyxh21D+Ae+2MIMDZXAws7mUYjyFQjp6xAto2uwBalQp
g5eRSvV0JQeYFebI9oMqNj1apeshK3YGJpNXHLSJIQy/GpIbzVAEjKbNQB1kcDdt7/CH3x6AB15c
oN/Vzxds+yOQ5ztmlbqWhZ2b4mzDyf94s3JW6fCVEOdwpZVHpYowfZ+YY3WTpR2XYCK2RWtbhaVq
OBq344XEDyqDJW0dEDdU8QNx9bel/nB6q4wOyIPo315M3D77Dvw6lqPs8Ajiv0XdrAMMSs3DaAWN
XIfkYI4EYu3k2TUe5A0WlxjunaHgCC6V3zckfvpWxaT8IDhJANOGFj/iY4dhx8DHig9nUbjc0JeE
PczSU9TuJWIwDrpMALW8K3w0uGw7GcVw9LjFlbt1YIBT3WMR1/6kUuG6w7xRdyjzdwdsgqTxqPVL
vYJMjROoVN0Md1e5YFS2F/IUYyMQQpqvQocOAccBJjR8qtZFQUBdTZkwfVz3rvzEwJlTLOiXEflU
cENZ4rvcPqIgPkXjSQKVD40pkHedSpVdcfQMsmULHpvwQBNAT26MLzPTBy7qHeEDwbpJNN4U7C6A
34iSKiIzc8t4lViLf/EpyyMZavXMox214c17HDApRwFVKJ8q1/oKggWsM+ATi3L1CMFpsWJREeMK
RSiv5aUMPpkVsF80lD8k/HdX0QimJuZZ3ZyAgDIn/HHhGH4psljpC2AxrdXsbI2IyragtIoz2sUp
nyMYsJXe7rFYELIXARV6YiA+JYPUHNiGHh+1dP6uvj50Jm8FuSKBscZCZD9F8bqyvya/WkFZIJFv
l+gsoXyonpPzpHexrnQ8kQcbx57vZZuUOBWfqa0yFD66Tka/0Qbj2kCwGmw+gXxxgNTLhfPjizZu
1zJASvFgKHhJLl0TgA9wH+HLSWlMpaZ66OIvJj5XimZvWInUsu4NWBzoz6ICY12V6PiTG+rt+Ckx
/OdnA7Pmcgnlavt0VfjMC6ND5g1FBaqsUDi28qH+luo40/rsmFSgSFImj6jlLPJNulywyeVvg0ZA
IDwP2r4VMTjSYbO5BXuWkNJ0T8bU7Dj198f1wEwJBOsafjUY7CctiZpODog39Z1Wc6z+QzoVuG96
doGRCnCL2wH/u0/lvjw/k+ia7A0vxAOS9U3q9Hxa5Wgy/5mkyxPWXSDUMnOp5+gP6H32tvpNE0HN
spLaCFrcSCe42G0OfDX0TH4uEJbtACQi2T0WHh6F/oVjP2HtWiHykurLL7DJOx7474jELPEWZEYB
Vxvz3wd3gatlz8c+sJUpn4AzU18bLEclHeslAtZu3EPL1rWymkxaSyDU12NFWcMcXnSw1dXJPPpf
tkNSiPIi+Tq86mrAG9RaU5iB6XqC/jAcGUbTk4DR5b2IUtlSgdZZkAS4Xsh++TEcte53vskgINQR
ICoPnvAh6B+KNRYxJe5uxmQpWQ1RNOWgp6+3xlR56CZEOz/ZFv3/d1lYM/1TImqvgf2wJzMzuvK2
avPTEpiAeRvUvcdWBFcxIezhdXDnMf9LfRUy8NQKnsmCMV1KXaxswWSZoyCk5swDv0A6DRwyMQeK
WOOBwn9E9OUQX5pCyzHP3Eq9MQuyq/xhQzmtmAXVBfKtcZydJklyPN277/WkypzuRmtuRYH+/k8n
C6+xZ3Cp+xzJCVFPMuIl20fjTSq5AXbM3hLiAySfYVVrpRwetLlwl8Tjt+fSk7Ep8w3sFD8=
`pragma protect end_protected
