// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Fxi376jKmMX0NEByEIvtFn2lZ2BfBnPMfLTPc6fU+xfEhi8iVKwPDbI+nRDdfYYI
IGTRa7DJLYPwkX1J0y1OzYMQusOCzPr0mtvfTDGcCtMMcTD8WJG2ACuK7rgWcsH+
QZEA4ix5fghpVti7OcihB9ZxuN2klTJMDNgXK6SKvew=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 62144)
We+gbos4V7IlkaWh/xvn+qUXeX+iy+/VASFxUya9YgahlvgMnfuDxgD9Phi1+AZ2
pxAcx//lr8MrNAnz1ObyoCBSvK5GCJc8y7i5JV2tiNWv57eAJpQF7uHZ7mHSFxzS
J5nSqMo+vP4kmJFpOUIUROGe8YsPNuNHGGdYZeU8WE+HXcx3rWMZTmEZc21PzUKJ
KEJhFbwbrN0973VaB8nKiJEIUm1KDmJF/XlVRIZD5+qzUiyncxAgBiOYpG8CyRpl
MJi1WY96JxtIm7Vv5ybpicCpPN6cgarCXI61b5V8LjhP2i6FR2FcbRsn/ODE4xU8
9CqK5Q/aSgdwpiraxxqoQmROEX9mBJYfdxRNolSNIOwh7KoUC2wLxR/TAfxKHNg8
f+L0YTzMpana53C0dgcGbRbfjaU90E/PrKiiRO33vx2GWMrQFnKWC1ln0T+eQrA5
OpiJ99cpq8Q9W9ffvHrBgE+O2cJ9j0VP2n6YFtBvhqjVKaNtGhSIsNIdamvwNZZw
ueUboTbWNP1M7RIS4Vp1+iFOlMhfv4I7HOhTYecA9BgnyUJ+1Z5Div4B3ltEhsPK
txg+MkIjKZFC1QNE3Sqh0LKCGwAfsXn91B6nLdN8gfsvhm+9iMebNdWXE+XHtd2a
CZrJwSZ99xX8B/iBR2Z4rkTuauVY/7aiKnsP160phCXzuAKtfG9Pzqf5qBQS0Aiy
ThCjW4zNkQ9x176JbikHMXzSaOaYqQYub/eNnBp8nusjZc6Nv7Z7sYljYLRa1yeG
nB71p39N1x5RwjbA3j223xhRSJ+8CsF8RjkKOkRMEkspLDbNHzOzMQwJBHwmnjX0
vgA6rUMcaRYqQjUgItzDdL7kZg9LuHfpD0R4ah0zZwrI25VbBak62SoeMq3HWLM7
BsM0je0GcogYsp9MoVI1ZNQNdXbI1XWPzzGhP01Gz3ckF9q20u60kxzX/BFK3LbS
ZeCezMl0a+rUciPVkdtJAd5SDXwLiq0bjas6aO1mIbAZKW0GGy6IWnHv6fmtIQi/
TPUIgeyeaCe3u6lXI02GJe7Z8flOowH/hxadAlOXEBOhYnzxh8htmnPnW+wac2oq
SawCWoGYfpINWGMbv/yQnSidHbIcBUuPxS6lGvFcWj3qMk9A1Q5V1UfijWJRHBu7
PjYuBLqBEFjxqu3WX/JHjIuTC2AWvckdOSjqjyy+8uUYC9AyFxUj3lAlxKHpKVp+
XQ8009k+490NpMDebaiXkfInyw+UgNbYEV0NABo+cps8Rk7msAYLALQ4EY5p0cLQ
LorZXF3kiTcejqCmEzD7PbQHs7L4ClHrwqXrOlXKdXPT+n9yDFqvr54WKA2mRpOS
GSDOrwkMTX7rjyg4UrldPZByZ+5G2j1B7+jnjW38tHkzzzwztVwQA+BBxPJwW8FY
+KOfdo96P+4UugKkhqr7LMYFu+n1W90gzwhDMYMbXXzgBwmIw0iJNm2cuRZi0w/2
MSOYRfUQnWmXeG0ANT/hlrgFZDeNBbpZ00fBTGit9qwAGvuWlmLDAYK/ymZHF/ad
piYG3L8W7pbgsYiNbrVDw8xhE6WNjBJWELaFhbM2EmmzCVbJYFjcQj3VRzgJw/5u
8biaH5s2CykrgrkfEuizFeJNjWdkl88cnBzkZDHFtRB+bfG3Dh7JLxusbFTohc6C
2WoJhIU4GXhzqdcyVEWPS0ZsZOOWxwK+JnM9RsmS7tM43/iAFpMyt3MdWVhoTYF4
YtIqt1FKHaVitc4gnWrl+G+my8PGCi9jegHvIHa0cALETFmSMbggeeu3UD3lYQ+x
lFJlGho6OUUUUJILwewxro7FJzlEnOxfL0N9hgdP4JcdPOCOw9IRBWG3/dqe35fI
jw/tbu47tHMrI4/0KZz6QBok4j2BccAk8v1BQzg1PVbxHzGWoEaH3nYnxZh+MEi+
7yJmbTecV8U/72XQscCLGrBCOKNUQwNBZ7C9FIN6qnNO/EEUjb/wxGfNwsLMSfty
n0oLuXQXibnO7Ydrr8fCsqlFdsqy4veLOFYAfq1AO9N5N4MplNrcd4HraKGVYw5Z
NVaRhQmj6y4H2rXNPF+kxGgFbdj8A9wywv0xOAB8fc2kMgyRiuqwCHBQTlfBbUEE
YhwubtHGuwMKj9LgK8RZBzWFHOBnluEY99viSf9EHmgd3F8oBmfgjCtX3r320Ium
vRNMERWDw/aPVEIsDv5TU8I/tZp2kg5JS6wTIVHo6P9YVT+w+ZjcYI1EfO7g+soP
8tm7rZfTvQRcezqS0bUz8OIoXav7iOVRt9yfod8/LOiHk+A2p7IXaNgApsS7WPzj
fz/Oo0tJbCMQ1szE9dTqKzLSH1teJCqmg8sGxtQZIu8Gnx/FSIw5xt73oXaKCTop
ZhhcqbvhUQEP2tLiDlxsNEVwKteZGE0mSmiNGlxuid18ehB4jwjRZ2mjJOmTywFa
BW6xBQkMKfOMoD+ewZWWfhAIlLXtDgVBPy+PTTnM+zX4uwgmS82C2Wf4krO52xiv
GMjZl36hZGRBPOLU5/NyeWP5BkRiu4cG0BLQJXHO2S56kRtOkcjamSebJyZiioTQ
3fMU5q6sc9sADCNozNiPRV2n0LiMg0qVETTMNg47TMLep7nQu7cuL0nv1hqIp5T7
IkSMKi5nljDYJv20dE/69rozLGgoFoNzVs9+LfPAWT9mzsigjl0ypsatmiOcQ2l9
rlROad4atDiS2JuJ3DxCT5Es/r3vcd8MsFf1HqWmPDyPAHZDru4wh8F2TvSiT3xg
rpiS/zma+pd+UPk7gc/ja4CIJler7e2tyGAyYW74mYoWQJPB8yhEOJoBw40ZQur7
R+61OH2uWnPWtj2+R4VQdRAKj+IOhSDRRUtDpCGoDfsMfEO8GlaN1xUUtyaJzThC
mPzkmWHSMxHFlRRndeqy4VkPinDv+l5upXtec27s9z27hYkdpQ2yoWWX0c66jZGk
gNE/ZCuujp5iVmcYOSKpQ+0uRujwAcTs6oB69C90crxmJNyV83Yu5hgxrTHFtg0K
C8Xka7zkkwivkCvhv/XnHRlHh0bl0kX/Kkfg0KhIL1qrfQGW/Q0HSzBJfc2Dyy6a
OZdJYGnM+AI0UDIIjQwOjNfUkXHUBRikERcnGcKnHBUS46sIsqFJ9Tpzdih/QSqf
4lGVRCX5sOM/gYzLY5cW2SUPDFEe588IQl2BbZkai3gK6g8aG3Wlr7vRdwpCJ1S7
RaLf9o2s4x6BtB92AMx7KOSoqV1ZMn8cmQV7hl4RbGXis7HzVLlO3YZK6LXUozFy
DVEcD90BDn5x3IuK17ai7BtOF6R7Yj0H0GioTEUXXhgSo1cDh7DRyny7msjSUr3j
yqnw9WMFIU23sl+vk2mWL6WMBSENl9MrIMbP4QF+A80c8CPQjFY+C45eec//Ve/m
73kYXEjYTZBEOF8GjPTm1iEsfnwTsZtWgskchwsiztZAOP2PMTRWmfOpUsLcTIgE
Vf6zgX24rjOjsQvy3w26+8GYPWCRuw2JiehQJvMKm4/2E72dxHCjH/32xx0qCKJi
8gY9++6D8OOx0H+JG3Ww/adicvfLlzx/V4AE/fYJ2pXG626PCHqYn9yjavarFrkA
l7qbQNVieJvOSse6cBZ6ae3R4GsRKS8BcKff6iaXHDmEveBPPt3g9bfJeptKho3w
rFdwG0oJItYv8j8fDM3jTz+9J/a6EjALLgIDewLsYgdRsTHst9ixDhNY4isCJQqi
pDOwY6dSjRjR8GzYYSXb4UF1+ijyeEtXlNfRQowdhBmL1z4nRH+vDmkrBCoOI/j1
8iemShxxZrGOoWhxn6xudRuz7PvuoK1UNXdANXU382XEwLLMMBJpceFu3aBFdj7r
z2D8AOaMlJN5iHBHs9WDF7O0K3sBSkIQ9Jbd4NMN7UleRf2MowjKsOk7wmd0nC9J
U1xMyD3LCWnkDT1aWW3sgMHB1WhS1aG5TMXy0ECZG+Zm6lO3q08wqW3fVPxD9Aii
rNt1hywqDZbkl1oi5EDokzrmt8dAj76UnAqy5jMCD17QJSI7qGRaZ3tr2og4TKS2
k8m3Wd/WLyQfY32mNR3JghCIqDdAzBzRj0P8/JNAut4bRLC0RJtS3sLQAETKwyZV
6jDRB6t4d3ubaINBL0FU2+f4Btj/g66O0yaETcI8Wp1qcN4tiZ/j1RJ0faWs4y0/
RFGIqZIP6IzjgJOVAuPKDAH5IblfeSv/3YT37QoSHMwkYDE8xdvGSWFEscyVZRkh
jhkwUfUSPymcgLFARmrsMeW+0nsEPp3siuTDMg9Ky+3PkZpVHa4fPtsJSCJpn24T
QPGOFzxyNCZtk6XqDxITsB63cl4XgOb7zJPoOKCb71Q86j2+of4qBiEFST8du4lr
xAKE9Pxc0mQOlj4IqoDOpMIvptv3vrKbyvvLnLrBxa6FvT20nMDv1o1pAdiL0gh9
/2hTQmTpqpPnrXzlpAKL1raU2TT32ARJDjM4UV+alL3Z96dNJEK6c9liouuxcqKe
eba1HAZ9YbDMyhRi1mC1VN132fUbIxXKTzlCDrkm1xUUJmT7VpiZcV8ZTNmN5Cgt
ErQzGuz4A1Ilm/FiVwWvwIRMd34pvzRuyUiNYJPT5f0rFCVN4hwtkS5HEXn30yFI
+D5MBTVT3I1w55gH47FXS4dMsuUuP4h5LmPWeZ50g879PJ5ExgyYuWnRXZgMpwgM
Tnapk6qpa+MO1fhc4VvxJfhZnlcf6lVwUX9rote5s89rLXVEpI0SSgfHJm/XmrMo
oixfG5/YV/wQVAKNqv1BylwNfpNPnQ4aaGQN1CqJAz3iUx4cAvD45w5HqX985H2+
u+Fzv/IbqtY3zizcx1weF9l28Dqpr+pvaD1Q6KSPjqDQ9e22sVAXUQmIRTHeuTNz
peRCQoUwmOXNCHWBon3pAWDKHCcDe9BQv/dLer2dyiDeEPIR5ZLETPvYO1c/tn7R
jTFmn+U833VSOuzu58ELxjTth8UNqnySMQnDIaCHqFeiAEVvl4TQHqTioVOPoTot
1fRtGPUJHbQt8etle9Ufne3uq2HNZ3yFtB3FixlhSoppPPcM1fZ8EI8p6IB0p3Im
6hFxMpxOX+dnQm8yXhnUkdLCYbTDrYvcoNNv1jF5td95buupLGMTntyEcQCMBLys
CrMGVn/Sfi/hw2xmvrePDIcL4MI/Mjck5fb/AIeRK5uhuO+QKecT/yMv3Z9jp44P
rBOLImuWjgZX903H60K5UYeuMug4Fzrs2zEauocpb0GfHScR3ZiZxOJupITRaVeQ
mY5kAbA+J8h1pAfcDsU1t5cJ6nKGOwF2trXMQPYk3FH3xMC2u20/SVAbzKRs58lj
wMxMRWUeMS2yLY1Hmj6mLcM8amQV+aTuYG2NNRAH+qM+TyN9yKC5nVI3nxMdMWq8
2ReEBf8u0uaG7llOn+Toberl0bsXYvIIBJZdThK5uSgZuspf8JxuGG8bKLXb/qhO
3JW3Zk8uI3RahNDEX5Q6mCxv1NqJDmEZQyww/p4ylQ1b3B7Y5+bA/AgTIERcbuQ6
dLznPnnY7L8T5KvyZYbK+8Lu9/aYcUI2aTGo6nK3viIR6n9QqA5tx+gnqaa9O3Y5
9WdUSO51C2Uv5eiSLnt+sQ3WdUiPSIWzRkLmWpRGxUIdIyZ9cVqTlyXj4fcN6MWl
vDi+/VPgonh0Sr/RSh9HWNQdXTOuxfy0uu3QP3K5MTXy6MHxhBr8fXEzROYguoFB
yzNssCot56/qfEbXWu4r9kLG8mi7kFCZ54WpfYnnJlyZLae1KRWVzSb6OnCen2GI
rJh+VL2408rE1h85xjYRzbj3ZERQzedNyMgLLJlztAIEC6Bt7D6sJZRR33RsPkNJ
K1hdmh5y2y9xGInolbXj0StPXTLAc6Z1ydXxJ9sdyR85EZs1Y2T+1D6NvvtEVPPQ
QGOL9IqcXZbqwlnIe1K3ub3/iss32hd1R2cJvnzPMTXFnnB2ZwBFdYUW+QpIsyeo
zrPdUCYc9vYgue3FuOWCRTciZRD4avqVZAZKooZMazA6b8bsiBpkOCUDYlnOCGUl
NTN8k5pONHqqCsvsLofA10LFPyRxwhhBa30NOwFD0s6XjNMxoPFHSURc7Ww+Y5um
UHY789Epv2ZdI1yWFSb1sasJ8QFQ8MunnaG7D9u/d84GMo3+EkPA58Sdh4MPfOLO
zogEeGMUIeGVpx8vsmsJ0IfriJdOBWxOaLbgp72n1LW3DPQ+UaLKGx6e430+nnnF
AFQNwSdPScP9LdblaJ/wNqT8XxU7+EAj03nutPBxpO6Sbhq+2rIG6dr4kbALHDEB
KlMmy2hK69GshOgmkBzhFm5u+S6aYM9nGQoTuRKQSVJRt5bxL/y/48fcG4a/iWrp
tDQKcHkr4xdnvQlPXPaIO2lnvWmaXwml+/n72ou3E2E7DfC9P+6WXyB3R/FxjivE
IqDwu9cB0Ku6rUSym2oIpcwU//T2orJEW5KkBaHXhAGwdkLd3qNhNxEhms5hHcP7
LEwfkR56bgK1mSVALIwchTrGZz/CJR/cCuwSXOzy97ikwezk1GtOvwAbe5DN47/E
j3GBdPFcHGj1h4reOkf+3wR3Lm+rOnYWf3MtACvkjeeOIeJO4IFDf+qvVhff8WJ9
6+8kvnZx0bnIQzlcTJHyARKMTe0L9InhEf3gfY+uOwPJmIbVjFlwvGPelR0n7HS7
5Rr0ZYJd0vDmWAi8pGAiSIGcdXgWkozpVVLZrXojhOoxTgpugt8UrqaoR8D0qZ8E
9tVBY8ksIaQHYyWNxYyLvy20orqwGa3S7Mn9dPI3FoZUh39W0fyOuFLiaOjjaTou
RYTkwa539CPNi+2pHOUb9C8H4tX5HBLIYRhEG0mwrzFtiIJOi7Epeir7wlGfbGId
VMrD2ylF26nss04Kmx0GwCzL6S81RFdzrdjs6zXAfWir9pPuYDeuYs+SYYMmtNhU
TIYUQgY0Lw5uiYguztilrZ10H5jYfx7GkNnLCD2eCpQbQ5vI1AjkG0G2L+npEqQU
pXYNkvZ+2nGFzgiU4isuKHyD6F39A42+pIuARt6rz1qlmgN5rc9muHI+IInE8xdV
Kv4XGm7CnGN3H/MSekjmpDYttIpRgEvbGZ0doIXVduWBLDEwf+ws1H3floXmvaE4
VdP/Xnn7NPicmSBjL7Si1hbTgoHgN5rcW2FS7l+uCxbXNKACdquOzB37G4VP64ua
IyCMxMPQ4zUYjI4fTzwCcdCGa5xTu+aXEQfC/rZPh3hpwreD6EV23KP9qqWxPukv
6F3KMGXnRO2xlkilXlrnuiPDj3jQiAOF26e7I29IVfFWPy0502wu0If2vZKK0mHV
WwU2IvhTA4lWjWeWHnq+J+bP2uxPEY+LBsCxrOkzuI31mifz8XOoQHHasXxIQgNk
Vj8XXdSMG4B7mY7CYHNSfopQzhQViIQBatykCn31RQ1ofALxq1diyfYGRSGQ7Sq/
xpxhJk0/cXz5AAxG0zRWBl0IN/qmFqiveqCmaSzFSf7/nRL70n/IWAYjN1kTzOr8
14OAPWKRg/6xFxXyKcoO6rRPJc0KrGGvs19foNJ54qgTBALjeVAgD6G8nmoEZ3th
Mn/oG6KCI/iynNPBs3yPwycpjMhAborAvN9LloDug3ZKqyq8JRRf5kNB9CKZfB2S
zS2HM4xur+36rnM4HSF83C0UBj0m0soA0mtiSTK2lytYqiLLHalpr/LBRLwZpRm3
K5+NDU6s7qWCdufM7aISg4bgyzkLZSD7KnBpUUHadPtafVi6BioqRDsiung4M0oW
0us6mvPAh0aY92R9V27GK5XUHUVZWNCbYnMViVHAX6oxmHYSQ23hAbOxzpzvItR8
eQs3cs4OI4iPS22cVrGck/hOp/NZEfh9yqfxsgRk0H+stmsnXr2GNq7eJ6PXnHah
pzjs/yihD4dh+0Twdi55LxqQPqmET5nW3S7G+EB+ezvapXpFfK6wUBc+2fhD+DB0
RdPiFNqYT4ktFJsygzpucNU5NJqMaEvbmQsqOwV2h0DI9A0YEGdMkH5d2Y8uyTHz
XwTo1yOmIZGkn16au1hfHjYEyJxkPh+ahZVFeeDtm2iewqsk2XUblFB2EduA7qaV
o6MUrUTwmbF7fsMX14GTp2rJRiYeTE3/6p5DM+Ekgrm3m2g++fDEjmeu8iNn4pP1
F4+kXm3No/Ztpw1bGBQnJEsEuLHQPvTNWfu22EOQkjNTkfw6+lMuaChrOY/716R8
DkvTfv3p5QKajtTtB/aC+50uPDjgSeZ3aCbtvjnWAvj0S3+RlB3re9uYt0PqwBLv
b6bHJiOim5UYdx5ZYSypF4Pgf+BfkS2z9ncEK7Kyk9+GdkIgdnmY26ueP0+QAfYh
s5sMPyEueeStNz0tQ9rOeN+dKA3VU5mUAOmLG9cZXFbmmThoR92qX+yagaM2xCWd
ib/rwVCNbDozGewgTmstgw3ubflEOekNmV8OXd/z7ZRUSVjQ411+su8B1JdqQrA7
2G+CADdhjwKMVDb5m02D8lxEP9ReFW2Ys2R+vXLYgw6ucnEVP+jfF3w6a9cmOjI2
sVbwy3PzTpDN61t+4cVn6ToLoRI4cXe3P6LGV8cDIj40mOWET1qnaBP1Y/yQUOuW
gj4JWFX8P/EXPWgMBDLCexMibGK+H1A182jYeZR+zXGqGhDX3UQ7L5aUfl3WRlGv
v3MbPpH55E1CzM5AK4fMDqC4jwVFKnjD29aXJRZRA6a9bu8ubG/wHmFkjc/e1ZL8
8d0L5ZUOKfexO/V00KiRqh3ysuAU7WqNo8hyeQJKTxpnT+N3n1RFFl/SkNKX13PQ
D311psJGiOGm2PbEKo+ePuYItZrfQdgetI4pSmLUUwN2NEDKAWarKiLS01Cvf4G1
ugWtB0up85R1jQWjLPZGs67eteg1h2sGZG3KKvHul0dOP0+wi2jYrr0nPzifWvTE
H7946hzS/CL6Cj4yW7nVKmLoL46bIc72cdnl5gdLiaGhkM38MDICgJGn2Qiwg29v
eXCdVoM6twxd1tkofx2Qv0PZtTBIqf8nvi/mUWyaav6dISnuyrk0pwRq5tMGS4ob
c5LZTnF/DHWkimPb/96/wWUAIqA63QOP4gkrSrCEV1EzyJC0fNsh8XSocjlq5jf9
ItcFVEDnOyn/3CZ1FVMMv8vydBSRJnnp3e/5Uh+BmE2NRDlRur4bo5iJ6cLABQDB
IR4fJA3fE64/C6bhjun0Qu++H4CVjvL8BLsyw4s6GbxAwfhwjzFZvwvoteTrjZrr
EUo4F2g/DBqc0Q2D+IIR4XAnARlg79M2pXbZPe3HnI0ykUyH/7mKjErMwSlYvuDg
YzEVzThR3x7adTzCZ3SJgW7rVogJsAaRyH/pWonZGxDg3TahvL6oyZsgB9vzwT43
33fcuEQ9oITssbnSYvbA76tLlmuiJGRC3WGJF8erZdIj8zhjxujEj+u0AAH8vwC4
bcjpHp8J/Ie92mwheWJ5I361fmPLl7oub92j37eJNWKlpfvlZWYAmeOPbYA92Ryd
dvUgF1eP4Yr35MxT6xQJme2kaJq13l21Eu9EFwoWJpx5t5dN/QUqRunPX88SvmzE
kFYszqfsuj6WSrqJjzv0k0bPOP2E1PxpHXRVJVxlNrpsQy1RGSC305Q1Kd4mCjxJ
u81mK1StbYl2GM70NfL9kFLH+ZMKq5Jl1FHsTxOteBsGKfidGWqcQHPecb2TzPU6
UjIsWQgQ60rWl/hBKYw8R1PZJaFOpIVrBb/a324xm4mMtAAWQHBwQ1W6E4J3pOFP
tYIkL7lSlrcbjRB7UY5icyIm/+FXVCPfPjcOKCJknf1RrVsrc4xnLTxgKFuKn8vK
P2TcYF0jB+lqCYDwHV5nDLt6CIpi0hqF/dCWTxZr/txB9y1eHbUp3yCw5YqBAnN9
k/M9F9Ss4FrQ7xrpJlP43d90d4opfnEOfu3+L63LllpOxxcEfkEBTeUE8B5XRXZC
ri505AVN/kJTIaI1APdZH6Vq72JLrPZX857r1tHvjCCuCBDAnqwcB9QivDl0GDUR
mA2pe/MMATOe8w43KM/syjvD7e6FxvQg2pGHZE7IugYv1UBtkeR+zZlpMwXWjY1s
XNU6XyAoAtRaXo3/GSqvdfkGtNDR2Dhljp2Zrf04ItwAmKtUM6X26PuXFUPwwLvi
EpgcPKA33GSvXGphE/Bp5PA9IDYMKwTMUNlkDD5nzft6d6MrpExpGYuu/97IxLYS
dyt09MxUoZGuh2soA0XKvrNZR2qDRXxcN2ZUrNfrwNYzNKRUeYXtwsFvPCB1GrXa
yveD9OXtRLrPv7xL+sQ1vi8xhYe+YIeXDN9PjkSTp8Lzw7qqDmz8Q3aazlGvwh+y
53fTzPTvlt2Q9fWAL7ynIxTCe9ZmEYc5PSeGVeBSc83Oyio3MDr+EpEhRt9gk7hK
Q7XHFA90rhcWY/yN/xEI1sNM92jQKM0RsYg0uCVVTbU7lDzE4ATwqJHmrC5a77P0
pbFJK9tQy1BbshjLOubOk9lgbLTBB3rYy/WFNY+3AYMSoihKK9qECoh6OlamXaOY
8nGbCCPnuCpe5LYkdfaP5+p/PioCDDb7ADbXSJHP6SsXwsbkn+Vp090fPYDuwhQh
qj5qNSbDW5CjZcYMLs7xEsaUqqMQjJ6xdi2ftT6eoy/OlGT2mBKjSC3iWrr5fhbN
DeyEUspB+2U1Y4K8RVQEqshwlmBSQ8hE0Ki56aPMvhsavmd4PxFrinFvKSdlWz0W
wCutbw5udteqnWOUyNoPCsFtKALmolBhS3NYVl/0hM2Y1riz+BFAjYs43Xr2GVHh
rgwwdIYuDSU6gHmH5zmeQq/R7ZfZLE8kX84uDPLYex02bMESqkueKngdNappJzNM
CUS2FWPE7NsIAKSdMifCllNosIrpLQrRsXsQIhKdMCQB+d7ApATGmHoFYb5KX2bi
VxZTumGY+eX5YMQPuMFV5w6AkP79tcaNMErJ612NkVIFLz9I6qCT3sdx53xT9bFo
ESRs5wHh//WItIvqW04XDYfju6yIpKmY+rGtDSg04MPBzbr6kIrW4EF7y1bK+gXK
WAaUdF9n27CDHj7vHqM47cl4wDxXEkr+Fjqnu2HF87zLf+6gaB8CEWtQAyWKYCSg
FuOz6+UnDeSwbd2NUAL89zfs+fe6Av/EbTNI5x4+g4fvnh4mMyx49UlAY/K/5iYy
O/bpxjlmyIWeoN+TxnhMYWU4DRSLQl/1nkFJ2+OlGUgD8NZ1Zs4HSFWXKqBhYBUx
/0RenPgPSwKRQgVbggEAui1+Upu3zjHIHDHZJdhKI04HHIBMPT0OTZDJiUiMeR8A
fHqFmdoevXTbYAX27mYjz6nmCBm/UsYVG0tVk52EhqKW4j4NJYNDeLctmCyRm2Ah
uLDaX8zOcePIkML7iKBbdUiRkJQnhBLxsdvs+CqA2ecMxwhVXsi4sCQpooxd9vrr
YNd3N6pup0RckvyYaBd1Yz6T/OlgcCbUwmkunnzJZTq35jt/6yafIIOZt9g4YyPR
UeW18zkP75poumRWHsskjJSY62ptZZ5W15Se9/QH2seUBBNjVuiRdXJLH1wq/c4j
rDUwVsVTE+JV1Ukg7lNw7GJfLyFDCJ2qIzQL3uGy8dynEMRE6mRDEPZv7gH4NjBa
WEOTqagROaFcWxjZDw12Ho81pcZCL8HgxD5eqyYtRgiDo/xwcC+WSYKl2wwK9Nt7
7JCOe7TK0PJ1NRyRzGq0TtLhIlWP6xbTQhtNC0t779M8CsqsleyhJP1UJcEm79LZ
kGl+snZzR6yQ0fNUuenkHWA5ObryvISWACrCmi45G3UE1Bfjnv0knyOLno4fh22I
HaoduFcOYM4DrlX3FqR4wa2WqmOZ5lIh4giRnuoEwZ8p14AbzB+tlVCAWeH3aZLj
H/NgM7KM3KdMaKDrV5JCjG/N4LhzulxnPT1/wzR9obkPxEikDQHd7tj572Xa5SSd
+skSlUaaquQ2mDc404Rr1ifhtNCHIe5D714fpDerboh6gg29RdKIqYlCU+1UGJ2R
7GQApQvU9VmG3vctN1GKZJXXquumEWt0+xKCyp18oQqe1yXn8LYppFMdgYLUmeG3
1A538kmg/X/LFtllYexht3dI1d+VkUPPeRlzhi9QuK4oO6ZYgf3JHWj+kGcYSMRh
kaItNpIrKDrUZAPQc5PrSj36JVzr88EPsaQhPcB80v/EsRXBY+WQ+jKQYiB/IWDT
wBZ6c/nhdkf8m9r+Abri3+cn6b6l7eqMYyL+5Yt70ZmR+uRCJ/2PPnVtoJW6P2KB
Qk3o5S52hpkjhaZfWqDSbJRejr4eLRYG/3fkjhIZjUYezJtGWl2J1gJvkxACS28i
euz71WNSW5OlhKJk4TuWJvTf9oqe1kZ/puPwcds1mpGuLKK+HGnnSjkvLX2YO0hL
zOr5dBmdZ78Y/BqK54gHHrv25pFcmRtmneN5K537/S4AIyvcltXvZDO04/xzOzSD
ySUwnHOnUJ8InQYjJ/yJ2Qd/vTtlz4Tv3jIySQ8ANyZK3a3lyjZOJXQrSW4wzwMV
7MyLzR8QCVLl4v6mKU1QG0knU1ew27eCeT7IB5hmTH/z156OfKDSZwn4ZjJjvU8V
orU4qNMYqdMNqaEg0fwvgDDgwr/TSWaLczUMLMYQ7D9nBDfBN0SfSWYX36M370EW
sEZ9u2KqaY8bq4NR/Un85HWGblQd/T9NNgJ6Nv+HqV5jwyvCIgKj8BlI/60LjB0d
3Mtocht8kSKT76lhQa7ZNtDcaIA9CfqFAJld7dWN2oaIU7VfyNtIAG1zIMwQmnfc
qi4uVpTNWn+Imhi7O1NTslPIPYOT2qY/7h0xlHJka6FrRZFCoRQA8ViwK1t/XCwb
3A4BAsGqrK/FV58b/y4XpVdWgXc1uh2x3iHDJy5ddSXkrrhL88O72EFQ05ZiC10X
MLYXa/azOzDzsiWt5TBqM2uHxf/JVO5kV9RalUzAN9HnHHE3ih/aT3Uy5pylBiNN
KX4p6Un7Pp94wNoajkHxUfSaQUdPXw2pgnTQj+MhW2ydlQsI8hZHsIr3TOK5OtJl
Ca29C4zl+VGRj5sGStcIuTCs4Jqfqonp0vqBSWCr0N3oxCrD4zDgbKfwDyjpewOG
dGpS2IDEhk5CJI+KyBZs8f/CqPeP61BbIY0JsCKnDOkI7de8pS15ZenUi6nKuZkh
klSPnjPYbt7W8bcE0cY66VjvMXh5jfjLRLof7w9xZMdiCHyAlv4p2kohUEO+cgCq
+uDBGVUOODdsjP+AjPfnAvleSEbc/8hcDlSwqaEqREPjKHANLK7JVvs0khw+sL7X
qtRZK/Iu3RCZI6Pkws7eXiWLUoTAAjorO5vzYEUkg3gdzhII/2gsiczzBPO6tZTR
my7U+XXxbfq/xejAuzt54G9DCoUdEWxrwJRjYDVx592QI87Fb6UKhv75FKusfiJF
IRYP0ueOJRSLey4rpq3Z1ztWrw+cb/XJvlz6k090HEXBgE8S5gDe5wM7fvpdz3dZ
VpS2dXS29QhFGsezXbvNi17D7LHK4c63MjMAhe/kCF3Hhn5qZkg03kMywQg3F3vd
RO46GlZzUde8u9o7MHVG4A/YIZlgwR5+QukeIRauKwKA/WE1ZiBhPR5tSPtbLEwR
xsfNFM4zKsLxLWOwV6ZttuYcrnv6tdaRfVxD0lcuIrKmwl2RbdBLX+qEIbVeMGpU
Uc3i5OYSU6zFBoPQf0HXgX+NOMPTXnKA5AFgODI22MKFZRGEXKapRy/Aik2mh9LD
cZ80obnQUHFD2HrQ7IG2A6kXE+q3aTuPgV1kmmJURkW14IIClhgmcL++MEJtdyxY
EhAEXJ3NieV/cbZ4QApUVEZoNIFnfC8qnNvHISOUpo0F0oJI9tSwUViRLx9hxX2C
U2G40+yUA9eDLXYY775yP4lrQF5550vvSV0inHJCIwvoT5eyqgn0Wcsxo6hlvGFN
/4bALdsT+VgWUwjsIK59lGw4swsltgtGwOlyx6P/Hk2eJow4zWBcCgXBF0fuuZHW
0rkjVIsTRDXdgl7fycHupDcxZxPo4GIZvGa5pPnuKMMZBvqEb0EN8k9radMggyQs
YNWr8lAudCxsLVSkrjm0w0F3xIj3plg8gxKosNDMMujVRoO5wrhCqkJwJEtYxOJG
1m8LEUoaZVMEHAt8qc22Bahvk7H69kOI4nyVkgC8YYc392HP40Rfd4Kf9vdK0lmg
tzuSpyXOCaXeUEtU1CHRvMRlbThbH9xK9tohnLitb7zAaRtRnqzYO7g56SjGRRL2
o5wsaGRLwTc1OnynUguvhvzHT70Sc0xF3bb74HReBRhvzpLxTJZCb/yO0V3ktOb4
C7wtOUfNGrxKcH5P0K9MUe9FgwGM8MWGPnyycMEk2eDP0LOgRNTnG1PqGSQqIlTv
pqPEjztkRs6sDGOH58eC3Go+hHoM8zHpnPRiGQ9deFsG9r6Pwvk+khpM4+sIdL5c
0J+D1ZtcNxo8ka5oVyB6wjTwTLsbnu3mzprQQYz24bw0sz5moBnRuwxVFHJYl3to
WUDRL//w1AM/n26dcDzfjbo3X5g7j4LKwdd9QyWetOykv5vZskATXA5J3st2klDz
tpsc3rHXr6PJqZYOjHW7YHmyiRl7REQf5BXvimHviMi7QrsjUCp6c+vPJR/fFZ13
wA9lDYUYRdEJ+ATmoETHQVOaDEdL9vsmPyQDVh+HzI/S6QzvIs7T5tq1I5hr/Xmq
NKyUCkHk5ALI5OhFdZCcsh0HYQUUCVw/Y1gQH2f/pZuYUqNojB0q+ExhDHgvOyy2
p3Peoe/21QM3fNnZioUZXyF7Sa314iNiWWGaaZcE2o5Z8u0lHfVDz+gFdzMNemkO
LtJIVHFXBimgv3USyXVP0WuUGPQDhoWdyiCWChqbIgibMStxVsLzg7dLglZyKcqx
ELAVzf5OZmpfnE+sPbNhSMaUQ/KUb3zC07DEOLaSSAw+vYGGtlkAxvj96tpy6S2u
qHzh9e6nrTjLV9jfXROeGp87chU0IXLcXP6q2dJxXrTpHYi2asOutzyuvEDw6gIN
D8zt2+UV+ugjYbE4ttDl1NATDnEU0znz5fDjcGGmlkGdmry90VzRTKKv2JTBqYPD
uCI20W1XId1YE7efIgfm8TgcEEkNHp5CtQaaBeJwYG1WmCgqltTsQspRPIdMU385
NqyTq9f/4whanyuUl5PIR4KPQXxdhK/O+zAH3+nAb66agUqdnqNQz2883zddy/SH
Q63k4jT0mPIoZ28vb3Hjd/G3LgiZX7cQgLafZErN5pFXWfjpxMTgc3mloZ9F/30q
E6vfRCuU4aq2I7VegQiWT/dl2UXYd4BKoiqs0N8KwUOS5n7YIYNi8E0t2RsYdqf8
vD3VWUJiPbsFaJ43MdeHrlSF9UbLh+iwubzGEYsp0mWFo3slpz9UtOr11My21vRx
+RmmBza7TKPYDPdC684hGmuxPpuLE457hQCY6KqNIVXV6PncuwR36S+j0FhqI5Kb
iBrIcO5CoWgTbvS61ZFc30EIZDK+JW8HvbLO0MBsMwhyN7+yBMZY9qMG+EWvaVML
Oc/LDhppl2SGzETjkJNt1I9BSgVNdq98qwEsAGR0STCxF4ezCUavKcYG7wdR/zQ+
frU+9y2QLSlM6gjFbf7ZrMJA09lkQajmtokjhKTAoh4VSDqPaC6qWTbYoRfw0dLW
4HgPiFfORvjbbTg41X7LHGUsDtRgzfKLCpcCfvlDn0GpD4ZT/56JZYCrV4h2Fj6i
kJZAHpDXyBJ/xkDTFf154iU9DXoNNzXl9Yo/F3ZvAla8rFOfjAr+Zn/CFkK+DFMX
aHWwJee+gk6BrexTjD+UoT9YThijKNZV8GRQoKunnRzAVXqJZUDY53rLJvyisF/W
CpH9nLVE2+ekNArEA2dZQeX6+Xr8Rwy/BO0XemzGuwChqhOEz+FhIAUOzML5bJEI
6UEbGXcnoZ1pwjaiRZS4Y0yMvMgR1hDKDKyTt4B4I46UrcUsUBguNYvcI5mlQsay
isazx8F8ANplEQDfSv3gWMhCvHdNbtvO3Lq8mhq08PSROX26rhBqZQDUppYM7c5o
fKAO+oxWx+dnTJIKjpUaTCuGoz16FnHzUSuPpeCuESKgoHQzPd8uKx0OMGgdANB4
udbKoyY+1r+kw8CVeHzRMcieOeVKOW8crCnnAooswQsTU9MXKtLuupykB6XZPBDq
32NQu6NZq6MDzUoVeIdS/JkJLBp0DwswpGebdK/BSWRQImreQZHegdtDu7aPBF8m
JDHpIHhe31wNjgfeU9ld/QacWlq2wStHSTJgNg/Qhq90Bq8VrpjVTeTnLurDXOMn
v+T9A0oKSWYqwQ6z30gFt4YU0OSz5G9nGAWFLGsup7VWbB1CO3pGD5eLX13UjiTW
dBMSpZsa5HbY44MkigYKunLnCiWIvpY9S+zOMluXksecpX54XtR8eDf02QeME9rx
7iJI5v8VrIaWj/Saohr7MlbeL959AR86oRG53XJMVCGUMKZ8XHxMM24zZlFer/KM
BgSzeXiWJcTegw/NSRaE+02Eyn2Cf9KAxrtIm5jcMO+Xckae7iqNLyuJf9OnB1rz
oSXvwJrfoycyDK65afsvYlACaZNQbln/UmIYnrYd1AoBURh7dlbDt8Q9KlXEMsjD
ESvamd0Y54l6KQRUJscUxIH7Gb181mG8ctK3FKYQUHxNnes9HdRhd2Jo4i0me72E
odeX0SUHvfeJm7tdz4uRvVXI0EtGs5vlBeh2Kj/F9rJ2RtrvXp4d1b87sAYzw160
pCzoqWEamB7swsPJ7QHBngk5bJB8KgH4X2DT3GR/hKMuUx0FQHmWvILHXBEClpfI
SLRfQlc6fpcVmberetT4cf77RYDqAdoCSx9rJ7T27B9X3As5LHDshNxPYv9D8BvX
Ub3PngRcYizHy7PHrFQ2d8PRiweGYUIYMmu0Mkuj06Gb9DvMOIvywk6mbJycAAj9
aUKR9Vf0XC/qJNyPVxj/Al6UpBD9XoE/D5fgBm5rTS9BrnRfWhYCxpjrZd1uRzsh
HwCTV0gDSGlC0FJbZ8UKYnUqGGJDhOl261J4uRc0Q8aBRqIeJMqBKWQdBQnhbzLj
LuFtJiBD6Ta//VbAFXdCO3VIbv6GAKBKU7wK5FuryonMKTfz2p0g5GrDbH8r2GvS
OumlROI5IuveAXjKAsTzAMa0zjunKj1jKPKu0RB5jmGPo9ljIzVYLmcdFflMevMd
QP9B7//+lF9v6VqFPqBX0ACIyQef89hfj5qKQYsLxOngClxOzuSp7HKxfbP6OgST
OFHxzpgQzaq0rWjrSDWeryv0AeLnwr9j2Jgqr0jjnULPE4v6PxC8PaQkLxck9Yg4
R+G1UUZC+iKTY5Qi7F0srNGxncaZwxWQ889IDiDEtz1vqt7w0QXjqvsFc7Ppwm2M
rMSW9eqGGvMBTGNT2IvfZMgMZqSH/o12GbkCfQfZ0+rBbdd6pWPMLz+AryW6AsCp
Ubf2IKNIrJwonRT6w8xWRHbB839Y5mLFtX24JrB+KVUKnP7fZe948XbiAX2lMezc
5htBkcYsHZG9pLCvV9xZRKpNJc77lTXSfy4o9ROMxoS1ZHNEggY/ClKVQd3jjX6r
gspesPNVJgMKmxdo+uWXzFJ3dZXC94kidKkknr2hC1HQT/hrHY76s3u7UkzqokE8
ojO/uELCwO2+0nXwI2Gvx9KGbxrmkuaNud3gAOOV7PF6E0Goncc1T8ydNzvGo0qD
GDkOyYuCXwAGee0Tvy2kmpoMsJtKlHvSnfyxMEvTRRvaqUtpiSwGGfe8PprKbjxA
QpEpBd2kUzI2LaNj0OqI8gAug+a96aOSdT6Dp5savLOUN8oVjrmoBm7W00t98+4P
qs2fMToVjiP8rw+MyvDGtBAnZroZoSmI6Nhs2a5VBI4OrinAVRkzdrCg/bMw1iS1
67ol9q4eZgncYdDTiJXcFNGtKGo34RmX4hVMqxu7R+G4QUM7G9L9WIRJkjpDJ9Fe
lxqoQCNB+qKNb3X7tNfzopEqZ31GoDHntkOOLvXkw/PucxuVM5LoVBZA0n4mN9p4
FO/eZUS0mUHeLb6CRFOjZw902DKWxhOW3TB4sPCxKBJeqLSt0F/7G+qR2HXV/KYk
UxC0cME5sNOQwOPflj+cK3mK6NX3FFVas0pOhpMoiRo2eqJOcvnFzLntpmuWLnum
wxJ+mxemdUOLAqMzLF17OSqF7im3Lk+xLoS+VlNNna/qR4k6qAw0IuOxsYpy8+Zb
szDyXcxTLSWopMFMyGGb4EnnyPQtpwpVBVMHmMXEqIMpGhDqEXgD/vB15TYaYC90
KbBOpR5hoGUnJUQelPEsmepKlJTQzOrULaibGaqXRyjyJS9Ld/AceDJvWLLZQksg
BqM1hlB7Uxms7TicDeB1hmwnFNcKUCIpYiEBgamB6gilhSduCEq+3sgAeGdcVb6E
WRX9D8c3UGRGK1O1tS+1ADOT8j1tMAePvyBsTi84/9yKt22Ox4xWCDdDhjQLYZKZ
Yz24T4bF2Zl3mwi6GLYBt1eHxxHLhnoMnJ9IAR4XJOK/KyeVYIgk10y4AV55h3Cs
v85eS48LUa9qNtWwNCu7sYTHrzcZuQZtZJf1pmepx2BP/IXxEzIAO+6+eFoCACGD
tcY3JGAI8T14XPL/5GiPQpsUn/NjYzhA+zfaRwuC2KWqaSKwjPgtb6JdDSR0iwQk
upqhoudvFRN27vFAOlWxXFWAF0YdHbPAIWuUOjVp3GdSCTQ+UkhnqZjEiwwraRPU
/JfyBRallsHdjCRJ8Fb+lFZ7gqWNhdi4sfAgLMkvdCpGbiFZW0VXusieoe2uPuXg
ZSuJQcRtl6OxQG2htHiSdYGjuEX2sAbokGQ3t3xoTLGQygoe98CyuRYsU6pAAEyv
2IKxA4oqrsWzI1QSwzd8sMWhcP4w73Tln2N8ozX1xt8PQL4ebA5A3gg+WEk6xy2U
5MgQ68ZX8kZ9mqmipCt8Yjv5JxkkNIzJ9Iqpmzm9506HVzR/QtPgp6uPkyyRA7XP
j2onUAhbBE/a2LiRgOYvQRhntJZYmTo8viMbsJPEwdRNRCL8zGW8iAkZsaSeJBiw
+oiAbjQ6phTj8x7BQPK5Id3pvdDbBe5AXRoYH0w3NanmR+lv/WLoxTUZ3kArRdGJ
9pLdB/uGbWYiZbhEq1tI3ATBM8p9u7of67dNvSAynxopja1sXlBOLeKmOuA1ad+p
RgXbZ5yHBIgSDOSL5nAN3bmXMDJIxsIGiXqteJZDpX9K0VC78UCu33vxvkMewpdy
gqptwfzwAe3F78/fXGQ+SDCA5M23IVrWGUo6VkugS1zqnnfHcbHTdbGBY+gh8sc1
7MgFDR09PsWa36rQ3yBnA2kWj0KgLdwJj/TYKLwlF5hx0h/eAkPUx5bM9MAf9dUd
vYvtkjMG7Q4qib4n2Uu49PECcXr4IrXi+O40rtW7NkESeqhX//ql8S3Q0+BHfbi7
x+IQOKwqmzqYbibhy7aBHjT/dDgmEjYym1DprrhNF2VhrteMzAYRA3nSRK7PwR3R
0FScbEHnCdJWEpJHRmQEfCAKonOwVGgHy+9xBFNm4DLaEGybavDI4AuIDN+SO5OV
18xSD0xQeb10g15jHd+4T5H6bvVOLWD71rN5WvsGaDx5HXyb8d/KXSyvqgQTkmvv
l7ZjMz8A/GiS3akPmmELY1siK2du3gwuSPEKf+a5aonpgwTke6uwyTfOFps6AeNy
zGSWxtPGVxdrP41xrhxYryBtNOPOB5mg/6O4gSW32y4lQqWPs7JOKf/qYh3Pkh+A
JXosTJN6QPSpW1BnhLALM49GJnP8hAhcjKu+R4H50HvgEoGOuq3aW7yMWAwz4dXz
t+Fc6Ftw4/i0xICkPkPoan38QQNUlFEhUAg6T0GrMWy6w2HXiRR0GcpxwUav+U9V
EDZRAFDCdTXI6VVyoHqJLOa2w0q+VdJyZSZTlROuiqN1dM0W3EIn+lceWSZXYaiF
7dKK2lRh9WgtOdmDcgaRF5Su+E0Kk2K+3ViFNltWgXVps6AUuyQ0pfYVlLcvg/KA
ks7Ew4cyj5xjC57vvify8Item7kqA509dLu+Ay9kEC3WMTMMGXS+uPrX6zuBJP1S
aecs8QzNPfZu57pZZmhJj3T+W2zAfLAdkbi9yw16GLaOlyLbk9tPOs/tHexhL7cW
MXjMFPS2SQ5LbTR9o78ouGmPmJdo8wUIAOpuvp+J0weQHtSFzbLhu7dwOpHocw+Q
MMRkX91MNJ+ax31Xb5qqI3Rg5TXOJ2NgP0hVVKcKEJSKeE2mvYNJQn/HgMpZct7i
q0WYaDxE2VjEqByRi+OkzJwB35yZvDyDVF940tiATZT9qCqSjuin/SRSgTmiqnub
QwMJj5SYX6Uhiezk9wiDvYfPkfSp4sf/aQqmnbsDoL5YO+oc57AMbO2wu3u+ZiBR
yUEmx9QNLRw9oMiT0HDCKRqG7hAlyAhJoDo88BzEBxDH7AcUs8n0ZZwxj3LmKpEH
mvUO0XWBU1LqjydGBYgK7nJ18sdaJa+jRSOLiCsxM4qAStXbfLbQYGPBCZLuvtyM
7hErmIQb6Y614Iyt2XeOkVqkrg95B5Pp6ec1PNFMm/hBSZatZpZk4/Z+HkXAQl6Y
EnJvQuCwn9aKp3lAqx8sNvMibtKFiONDwaKU62uvoCaD05qfR2QNejn4KidL3MFN
gKe/0x/rDvCVO+SnNRilb1L3mY2vjeEGQRNOKj/CVQgeZ7WmSCJDRlmeFQMU3MiA
fCCSkiUyZbsTNiAYifUFa1ANgQ5x7Bb56K+fStyR0BbP8ibLYYfXDPQ+UrhjfwSA
BbEsQpUc9eUdzrRbViz+HmylZ6HbPBuKkGt2aczzE/zzlcrhYMGr0lRjwv8z86Ni
iHVMTu5h8S1r0MMc5dgFoAGAGV2+GnD5hvihzycRr3/ah83J/7XfMS0MzreZk4HT
MXVQMoVPZVyt6gg4DukLRCN5sZCVwKZS51WWmIlcs8NkOQofKnAQApjaYT90TFU9
XJk+DJ+gpQ9EdFgezrguRUJGauD1FMBz21mkX0Rc2xdLUFzmumpwBInjKVIy1V9K
rwWAaSOSsYWP4S4q3yIoQGIFgD0Ke4bEC0e20fK7VIkF+z5mZLThSdJjx90rpeDE
T8w+BiGqsJTxcU71zNzzCFb7eyYzVhHWCYXvHgQNc98UihHa5/WeKWIWXeHpynkE
SAwt4TTZ4lO8extZH/OcyWs5db7l3YvIciyMp9eAWoOU7KV6SLwJkD4hr36TV4f5
8+WumHRHM9wJqFRGhnTfPDUuMS81eb9VqdDrW2ez+z3z1Sb6AGSNcIyscofRT1tB
ZzopLuQIdCGXx0WYK8INV8/Fq3bq7Z8REusB+/lO8ZW2tLjwFnUogBI8zPl1/KS7
x/2RLgKJ4C1MhtVelq7qce9rrkgmr31e5Hex2oTBnvpLPI2+rF1iD+DL2+jLJmSl
o9Tu59/cryZP2eIVi9Om62turyqJvwTDPFHG4ezQaBca1nTmXEy3i9oL4WnZ5I3P
1CWu57yIoi1gzpn9nCX2Qjf4WLHQwC3Bf1VI6OFYjwBO/VUiHdXMBwcNjIGYmZki
OXICRGhb1WsG19uYxkSq75Lw/GZa+9iNuBPGu0ArNAuqT8SRrhNYYO823shxhUTG
gYQB2IvrJLl1JAqk4wKRJdLupcgHKCPJEGGTFNR8R3hO7YBoEu8GZtvuAZWzEHCB
o24wmXdo94NPFxmSR25kmlPcWTjq0CP2Fvr5h4L8lF6h8IuPtqBQbDCqKycrO1pY
tmDPwVNnMIBNH5OU6YGsMYDeHx+hA6eEvGLvecdcXlGy4AjPNchEyNPGv5hL0n8A
P8Wf3NY/nPwfEP03THotq8PFiyRtClqer6WLpO4lOf0n/jeSpxdTqewPG5upyWuz
6BFbW8tYt2Wrr2ZqNF1JBek4kZMsxc3Dw6s/okU6lYIe+6RfX8PbzxcrZ9GxKMaE
QLJBffJ0qL/N4epL61uVbpv0Z+QKWN5ez1rzmvrrwlPVHS8l9BIqP0XXnBTSl7xc
uvMXJ/9px6r5YzzFuLJMVwXrtLe9x/qX1SZN+QeJlGrEPVBC1a1MojXwy5FUrfqh
wDnX3QCpZDhmyZCwECo0apZFT3uXArscnqkkER3LIutWb6r0cDyiYFuv82oOTid4
bDmN4pZ90pPCMAuntyDs0Zw8R72aLuq1FjaiDH9cflAzCTlLfpkBeBuC3//lQa0i
fAaKtT5R0FMxSmRvv/D7OqXNTCe0F03Zo4zGonrRKxOAmWSxB3fTJkhLwcOYeixy
XfwtEB4ql0H7sWlJ4kh+pdT35oQfd38ZKwzkYcLZSeZdgamErTH6FDWGXLc8i3wl
C1ugoA4rN/THs70zkILtzCQ0A/2e9mXrhrQwg0x8h41rGb+3YWxab1BwkAJEea7k
7q1Zg9zxdD8KCGA9NdDVZn9UdsMv4BkZKhuzGijrM1SG/c0teeFU8kCX9nfBdlC1
nA28ZYRfmcELEY3Qc7720uU870jDdOKRS1cfOFeSI0BiRI5yrcrGtoWJlYWxejPE
5hdmK7z3+zQyVqJC2kHoOrW1qRebPDvda8HjtM/WqfZ6tzen7NevuXMwMjDHkjlo
RTDUKRP/n7qb/9ML9CFLlzwx81gfQYEL4FiLuUIPgwVtJ6kGroCIrB+Bj5FISMgp
F3Hq0zFTwJrSLxboRV6g8sQvi/uXV0B8VU2sxJv9MB7ADTSfc1xnnsblz4wXn0rO
A0LxBhJhJ/JCn5pherHDgHmbq1eJlvqESuTUmc0/UOiyYp+5drnWOHnpG0LeHGAU
2XBkBs5mqduwyvucgm7/6Id9tlldH/8DKLztWMHIlFhBqdjqRxM3mAhaJHV1hdJq
ZuGG7pvue2Sv7H8UmfIDMZx/1QVaV153X3mFYzINYHxOaStKOKWR8qp511XPMTvm
7xYF7MuqDaE+ZVaZ7Mvo318uBQIkMki0/ikNjCzyJSM+4qO6OgaBs4m3lkvr00ev
DvgBX9sIo7GzxNgFx+6ynDT3jBLbtOq2G+qVRCUJuELXsIbXPsh8++rOn5KYPn/t
lFqVc1KUQTVhiqzpeUFCmS87cNM1lztGIT+Fz10mCXvqFH9Iu63P6unBlIQfNPJB
KqypTYDSb9QGRLvTBE6/+L+xEO6Mt5BSB6ElvCa+QqwvzSvxsjVribR5OBpim3Tl
kPEy4Nrqzfkx8Zx40Q4OqQl2hD6IWMs41jOYrkCK8NxdH5pFI2ilSYM9mummv8PQ
cCy09Ue1y7OILojVbBCG2qn4smZhSPeze5DH49ZIaQ1hwriv60m1ZhtGtGx52IK8
nAyjhDp57T+Hk32tTRrHOTBYqnx/OefyivN0NtL6/idl8nA9jPXmmU1+PxgBRdpM
O5b/wSqcKOJxVIJ/FpuM0hwkLBL9C+zeK5QLsurJFFXahIQz68OzHzAZoz2BsU65
fzmHWWiXBUbGKeI6S8UF5mUccGAkx5F3YF6Njz9gndwbqt6dzJZ0wRgK39bRf/YR
Dn6Ck2EgEhNLkIuAnqykCK7RwbvF4YsRJagPsCcZQvP7kXV2ufx/jw+6nDQ/t9md
C5eiZbgbHjyijIXOd8qBJS2C87ud5o00iXXkCIRf0BcRFl+AT1wtKTHHqbbU2twC
DCkCrlBFpBdiBAc2pyryNqf7ls9XG8ULLFQ7D+FPK4SoKR8EcKgH/yaQKnePXVLu
xmUMHJUBrnEpbBikKHSJRRfJD3s6wzubwyBuX6RORD5zKlsgYgQhIwuj7OTJ/r2a
NABHaPTTv/AnVneCxj+/3KzDSXfULgRz9pMRP/SwknQ1l+XQD/yEt2B6WOfgylMG
lr/E3wt1SGZ9PwGPjmRVMqDXQDiOPVnoabZprLlRjf1t7SWyY7jbwHoLsZppbT3y
XxY9FrDVsq2sgeHodCCRnGdIOEXlu44v81aZ+EEtkLCoa+ehzNNIwZfBTY0f8km+
xFQBcIlqi6EkI2P6c+BkoeOYh4i29CPrbQSxaYnizqvIR8f7DicAeUA1uujhdnS7
5JB2v5Ess2Gs7/ThJEvi18KjN58f3w2kMgl2gHYg/KIMw8fBAGplyJw6xy0nAN3X
PIo/pUhaTYmUJ5hElVvTBBgBVzgIxecEVa41Ivi3oMUDlifMFB/hYWgi8SMNDjqD
PbGJN5WiSKqbMgkgG4dsb74uvfKNynL4zhFRwAT+ctb5W2AWxzHOqb6dh3UPKWQ+
UBCW5e9ibpof6RXZy2J6jGgXvLxad5shAgTA0S4ScEgna9dYlnDrjU6jVbqzUyFA
rXDcISa24fOJI345vIe96c9BszzmGFBc13l6EaioA5xM8+bX+zWZnJ8CWhRzp2H/
QAdFBd8esLCDD8SeS/M0rf7d8KAK5/ZKQ4+ZZlz6gnvxjECy7B/UfJISAGEhWBkb
2UIjCIp5gNbxVkmM92xSyuzM86DBwCemCE5KWMmkYtN2okhzz96lFscF7fBLqU0F
AXZafUhuQZEqdPdZbBw3mH75DbBQVDNRHlumR1414qaQo4sVUMTDrMCRbR3eb38n
5GOTXd0efM9dTYbQRA2jQGgJjVIZUjNnDg9lYNu42yjTKz0Z92dxiqqChbJlylYr
v2OWcGN0w7hOS6tDWk8DKjBWmo37nZcECQ2noGMNw9Tav0kXJ3snJ01ClCD7K/5w
92pinz188jvDXZQfUJMVNrio/4SoH+VpWudMnf45ECs0akROLY525/kpt4pcJwN2
fQ/tiS/AIWZ4Ph1He0weVWdj+xU8n3Uyn3KRD76q/rg6fBm4mPgPAdVE7DYt9de1
siRu912SyR3JOc1X1ue7oiX3dh7yhZAUw7Qih94JBqsUgNRq9fYdaj04kSGz40/3
Op9EqZtK9UjgtvMa5+z6cmQr8XAQXg3dpTKmtWcq88SMldu8+sqJ8kWh3MUNHpvt
Di+Kg6fwj0rmd8W1B4YjJgdEBxwOIEU+VNo6kEPJuosO2m9kAVvZz4NtxrHPwgy/
hfd6XMl0BHs3TdeOOhlPsJR2nzNOWv7SSQZEO9IFkz/8+poNBN6TZHgitDRqe0+0
Z6GQhP34VxVp/sNuqFIp7uIEY+tYTi2Yla/pN1Shlj1ZKhvdtQTl/YyXfusI/f8i
HjJe/+0774dwwOVVoAy4AMau+E/DoVgbgvhYfXRFmdFAPKJCcEG0B2tr08rcmIJp
cmONZSfBs7is2IswUTIwRTKNPe5cUUUzzdsHOZu6mY/yl3TL4RCpfvmi3h582yOW
SLAwjZ0T3qyi/4DtzLjL1Y43pVsxx9X5fHGeQtRn+KvZ88hTTcr9mLd+ZOgz8e0X
HV94Gxrp8sZqVuLsroIXkH7BBFTHuT3jZRQCaPqX8WhCpJa+QcfbGH2lxqWl/lu/
cBbBW57cBuDeqfha6blKa4hJV96WEsoWI+8eoYbdeIbzMvHf4VtWvJ3ppcuPmUFU
BomuYvueD3IXc4sZtQB1iuI0VN+XC6wcDkTni9WUKlGUA2qwL2N1lvFprk5skgAm
ri0T9p0+AOjTmjXU9qVSwlIyc2t6C0bp+ZGW3M2JAoyBkxyLpPO3L/0/cUz72Aj4
oavun45qgLbPSsCvOI9Xx9i8AIr8NLUQqIB6Hy6UCzM1hu47KNJGh3Z0JG1F5JXd
Lpgxl3LyL+JiDU2i1kZJZCmvYOYhyeQUmVTqXc//Vhzzdz55+aW8kAXQXW+Vc1Co
YfTirKJ+w6ndcZ4PTLdFTzYNwimvK9qVTZlKp2Rb0JHNNL863iFE/ufcwR669ik2
ht7Wp3KXdysSqRFKvEiEwz8x4ofb7+w0iNH97aEmbPD0N/Qh7ojS2zpu18asytOP
0nRShhh/Wu7iszcSOEe+TuqLYxrvBpqOYZJ8Y65v3yhyfbRExsSQ/jyTepUB4Pud
ldh1ZXJSoRBX8rPC76Gqix/N640HQbKzAlOt5PrpnB1lMWIuMbdLPsYrQF6rgiz/
0NRqvnBMjkgUo3eGZFFTWj5Pdr6EA8ofHUmJ2DCFsVkTMEZ7aWdlsKZ5o7oYGY1T
gvhP36U9UoFyZnDcV3j5WsvIN+cRoaKxPAR8cMVsRrfBjKZ7dbUM3tgnRa2PNNQi
iknPypTBqz7U4CFD/wIzRIXasR/PEjZWXf7mXR2bPpsVTZF+9ENOmTkI46UHoUuQ
bLcgp1k90pnH1QiWjxjFItMstm0ym2U/R99f672WuoH2pM9JmHUd+c1TexrJxG+z
5innaxN3D+35pbuRpxDf33h3O8Qq5882HUQDKZGfxKHk/FR+WqBMtw+wyd9lyUIh
1KP9fN1o+wVvwNiJDccFSBQLg5M6QoifMRvy8J3HvyIM8ZuwigXQs6YdEQ2PYMo/
R4hQTy10t6k5aFF6Wmo4aLHr20lbEsfAuG+mNpGSaOERdrh9AnwCDnoymKgjREpI
ZAEmd4yM4MTBQEg+WBQUNWDDBkkP8YD52uc6q821gnC4CBKz8C3+OYUzHqOpNi+X
azCdK7JlZ8QWLBndh+OmS1Rrpsi6fABGF2e3226nFwzcJLDDvbLoK9dPAIwVlE6M
rfNhopt6Ff91zBlZd1TmiqtinwL1Qm6OCbM2GQwtlEFDqYtq/DwedwNdYEipdaSh
LDU2Qcf1ka0f3CFMef5rXPJgHI4RF0P3XiZQCXi9pwE0kqluw7j57pQpWY2ouVqr
NGTTuK/35CnLUL572W98mwkCQyeb7EQFpueSY0MIEBZnaSdw/0FmvCo/+SUjwn3s
G3TwNlW6Lt+uIx+YlPsXtljg3YR0mowQZ3VL8Ak32eOwZqjNFnTgHNDylmPh90SA
i24TQwPBrpFf7VbcGzgy/Bnu3rzVoot+g5QXJcJszcAovswaJxZNHFvqg3uo2rTf
0OOX+Ylunh5R3l+GfMwxkG2gqrP9lsRlEwn7bqU0JnWgoOwueFf2ogHlZXkV7101
umQ/j/YptCtN7FE/N0VKS73yTY3xvBL1U/BtUBF5Dte3yGA2UNKe+ksfjbuAXit/
5T05Qcn60bXle/cw/h4mn9d5I7/JdL7IEZFgQYid3sVpK6s8MYW/2Bviz08WPqjW
rCsIl/F/ROPtdX1gG+F4tRt94UFOM7Lzf/8a+ZcjNg/R0cJTKV4u347cjKbmJ/Pw
ShvI248zLXIvlFWtWtfRy/Os3IeMUnYzom+ZT2ps9ymXjc9X5ksu4kKCfn+k5LPR
MUOpF7mmiZBtSSRnpGH4UDhydrKIzdoePxmdeaTbX5QfNTOja4TvhGS8PO1Nh+Zn
cFqUGYAIjaTy1+F/dRmf1KjlCICKQxakVvbF/bei4sSLZ6zfR5Rp3s/qAQmX0u7d
3oaDcesFyDs0PpOA3wzIOiU+mZ1n06r6WvshmHRTGHCz9h4m3x3ZWUfNYZZYjGmD
cPCaFvmA0GdMBqY/n8IMEcngThIypw2iuIBhsmH63bX58q4FGO00DDxhSJzAHfgy
kn/IoUwUjO62ruqwuunhMIim+pftMNiuCYDqllRC9/BReqroWC0+C06CtKMgL8LM
BpXLh/nHOzgfTGCEY45Him9nsbYs5VY1ubvYqg1lkdq9H1VVJuWGytBsR5Cp945k
p/XzGVoFPqvaxy40Nj2v81s4LCJDFm2jPpqtxFyaXjG51U3qQYVSZV4MBqaK+JiJ
jWdh7Rx/MEbehfgHGY/2iL9SA8jZyeq5jzGmSdkDMxDwHxyi/Cxp+irXzI6NwJQb
JxRBH6bbvvLQCkuGRVIP8FCsGso/2BfHKWmAmNOWhVPp4OdSXippVRdcTIzIjm2l
SA98g1TvFr88EAl/g7NrcXo5kRGj+nmcY2jP7jbM+n2eozHFdOVT/1NQ+nTkc4lN
os7xq5V9FxQq/BpWei2dy48YEZJ2/yKSoRh4cskbVw64WA/ZIgiKaXhE+mgNKXQx
qeo765oGK19dSooYpFuAmfIkoID+fUn3TkeqYl67sneG70LWNy69edmNm0klt8Je
ybwv5KA+XMMdsqUfDPHkjRIZqF145JjOvXB8IICw7pXM0vMbbmH1iyrPoL1OHSD5
br4lLXFbjVLaJfgfYXhNJZn1X5tEstjuViy/9IA6YYl/QPe7fh2HyeHnoK1+KVCb
bekNvjVQ06wwOXgMIJnI+OhFkMAS8HVLFlIV3B2noUCqtogmJYN5nkzDg0Wk7Lyr
oDR+JvFM/YsV5e1YgWwHExY/bQwZwSpA6cYBJnjRx+5PqZofRdRuppill3BRP1Ut
bEfjaHcPJCmK+kr8fJag0kOYV5nP6T6H0iPKrcxqJ4LOyFzUlDD3QMupxlgCOmLw
JPuxX81Je98Z4pN4yX0/hfQta7RZ1VGtZSujVObZPdUBXyUDaNnG1YdLlW08OGBs
GudcqDWsf8yC4h3dnT9JZZzIBnq7gZQgLjJtO70GF+vIzo5XPkgW6ZTVLpJxQwoN
UdWWnJNo506TMyQ615SHAywr7VbVMO8TlPUn+vM2GG/pIxd5Dm3RKB7Llo+SCVe3
5NqW1dxS4+cuVfc6Nf0Nbszp5Tw6u/ybYh2O5W3c8drRLrxSMzLoE40O68SXrU3g
YsfcnjlkP8ddE2v3AYJHwP72YvFWpAa4UbMWU3XvkYcQjRp1RmaKp5wa+mFC/vTZ
udEfvuLjq6v0FMMOpqfbctlO8/B2XIE4pV5xTb7dx6RZFVq7Q+BkQUdM9uiG0QnK
C31g/IToRUMOFAusNoaw/ASxbAUS9QkD0p7FATJ/EXnNzIjk+rZWGKqGG2EDhhD3
nhl1Ha/AiNhfdtYlhrQiKblU1cjeAXKutk/O9PhTwa2HjlwpjENLGcEzsQvL+fQw
AA8r38B7NnYYgOfjvxiGdVh2yZxUbKLYHcDB162iFby+HF0lSDhkEwnEipBCRUHP
qg1kRAfvTENVLF3+bQEtJkDqNOtZS63dwwHoIRd+/QI5UP8/2i7NlgukvSEHj0/8
kyxE7EZ2EbnuWRqZLdiWSwZZyUPDKPiE8LLhMysYYcuRKS1sVY4yhrRIFyY8b7g4
bn21GiuFn4V56wTxWqNAYFIOKwa+djnnMoWlyFVulDKDTXmO/70zjyd3B8shsGvf
CAGvQS4lsrys9oABTG3EV+NCzyUNLyeY+KolCf+Jd4djA4bB3eo2c0ULOm9ttcmr
/CfKj5BIzwqoc+LzA+L+hPsoUzMHob7jYxm4oig8QrbRtL0kwBRqZl6Ltxo+xqQM
90IecGjn08JBlq1+sO7viGDsfJELqCkjkdS3E9Hddpjxc4lZ0gTXiB0DJcHc2LQG
9j1BWcIuA0LZZu670mjL2hEr8FKFXhJmPqYuMtR3N/cyxxb56w4cTjJUA/fqahQm
O6Ou89SSJYodkBj3pXM+LXkxPGUuOmWInH7aD9QId4bDNr2k4D85cf7yyNYJe+WK
xtfsqL23ORSjJEEOLoL62Gsf5SJ+gOVKzH6hNpG0fyCGR+QLwTRkWG6v3c2eSeeE
TZzLi3i48zBbHS44DTJLVwSnelITtSB8+1nirx2bVjDII+T/UCkxL6mEG3Woximb
MsifjmkLrvt7Ibqk0X97JOFoLZJCYNFGmrIbSZed+GOUwGVbUoZWvYSIhiIsNs4h
WVaeNJO/4G85Xugx1SAJF7YzU4cOqqaRHTiqDpfG/VVQP7szOZbP2BsJc4c3KxbG
or+z5EfDeUdMkNBN7ciU6aFt6IjImAS8M4igdobhW87F1aNVZv+/VbdmjfB6YU/H
3D3sqqR+bGpEIbULj0hvL2Vnh4jnMuLALD+3rZ6fGszhcrjAd2lefKa2+G4wcw6V
mARGytdZIudL5nfZzAvBqKOHNMQ5cbQLe38y72HhGy674tEiMkjJ64Rgprowxe0w
WXMbj2uOY33M7muNH0Adai6/LNV6wKUnMlNmqnhdce8rpezxG7IEshxW8z6+UmSr
vchz3Aet/4JVXYHB/0vC1nOUIt5iEdnHEpEobIwGAlRofEaC0ol/NXy+BFDyaUe4
mVeVUworJkb3lJhSrDYAFaC3MALOZMJ10PU/+MhMOTbS+fOm27+1tJl7hIZR4JVu
P8ZjpWEJ4Q540xTt6vf0zYTTLFDVnrKZVJ7w2wPoVi570qJfPYSB2dlimseOg4qq
4210SvbjQtv7KimMy0SoP+uiloIBVVqI22K0IWM1eAPJjOMhIoXIiYmdQ0R8pgTb
XjPhX1brx0mCBCaci2hQee/cy4aMz2fiM7GCLGPIFnzLyYizL/4xpL0QTdhJtsNG
qmgJl7+C+LGXyBsL6EKACdWX+JxQU5mGs4L/PbhW+nrk4rGmTQ/kc5/Fmfru5UiK
d0seLSyTCNrse8NKKkPUsucLMQ9wvDZiz4pK3tgoXn8xsugt+mtFAgXwUdd8XROv
p/QhKGFDluYTkWoKDUI7mUMqYyjz00CmHSqFJNLQBniJncBwvbJOVJKXVretYW9I
8Rk9chWSPPk4Jhyso870h60xwQBMshKGnxw9a41NIf9cQFYqRDwsjUDQCzOMRWs9
f5w9sMKxMQMiy5MB5mBXc7qOwoKDjUYxPktDN84W8ytaeq4TKyQp5uTnNuH6Ivqh
/kBlVaw/Qb12dNdjYi/LF7WzvvdzRje5mMmujz0WXd2rrjEO7pB/viwAunbZYpuv
lGG2NtjIEm5cN0dqKxBth4EVzOo3dSPu2UxwQGmmXLexLI+4SEjqPmzKeS0SGa6n
GW2BtyXrtJFNbULivbazys+8IvY9UjFR9ENU3acsLi8eaw4pTVRXezNkmzeC6wlm
gtCbh/Sqq11FIYJrRH32JnfxjwRpb+4LR++QFsLzBDgwXXxFLpNLqyOmG6+x/7R1
1ekDWUCNAnWRCuHkGTQBD7S05zpkOxW8h6dV7N82UssnYDK2QoObPDuA/KgSIw7m
xOgcDJJKZtIOCO7tKmCIb0atxipatl6NO5v8CLSmPuyAsWpgQPLt0MVUa0ftrwqp
n6mK1uUMYB+mDv/8ayCova3P7wXipwy3SyJoOzLn1XPi49knozmnMP6nZXRE3FYN
BAi82Wv2Bw5sFflYEKFQsr5rCzUYtUPENocTwUcu6t3ftWRF3bst72V02LL71vOA
N3BA8VipfjHkBou+9GA1+4RWLmhO47Dy56Kc9r4hMjsahuubi1uka8xQNVJch6/P
jiAFwORqi8WKJM/jBMtEnX9dQTpdglxUh/SUyqCXUbKQvcq6QGbEGlrhkt6pFLYz
4tkpKwZ1e+0rvWAeAcKWkTp9VdHiS4SGsuH3FgarES/xKgYhtrAJ+fY3IvDjFlay
H8HHtKykjAMhjp4NYD0ATajrQ6+6TUWNHN6MWUMKCOqrSIp2DbbASgvHfdVuTH+r
NTcHQSd1DHUOkacMhdsiVv5HvMUFiDuTuHMyGWQ97Tz7dVAmz6apGyDk7GhbKMj5
cmzpSOzUk+39XFO0pj5ovCbteEtX99wsn5QDp/sBBZnCMd9nRnF0z21ioCFry8pa
oKaFKEjCJIsSQD8umFLMsl9h+gLdFdBEeMlucQbZ+1OYrzqzsNi6MEVLtPNcQjCw
98q+X5tx4ZGcOik8Js+9wVMeuhk0Cn91nNcXEP5CXl1sDKQIU3r6X6lQtiqBTJ8h
gKwgYmF4aywOoePKaXNLnPsiDMm2c4kS7Orp7I/EGw7rOoERZwbcqU/Bhg/p0o0l
E/uTOuF3puPTAc1ODsV8lFAht6P/q4HDDJcsX/RZaMiki4sMW31JVWSroE/zmAv2
TrpKpuG7Mjn3zoXArT1HJAZxWuJL6w3EADwXum0y7Os1uXxDCo2oQhj6zMXt36CC
3JdDMx0aaq3fw1hUAsrWrYyai2SXDt8mxR1OBZj7f+rHZA6MVPtW7oDXpxQHGrBf
N7Rr5zomZz3MNcjiWm/TVhAmJsPyvn4q/wLsDpa/Z+Js4AWK5I7cof9/f6rnx/zV
45dOkR9dpPlFNUOzOi0Z67OXKwFWSKmqubK6YSlGPCRXDn+VsAKisdHgP16QMHhC
Wdf0ntWDYYb1dxnT64pxDMTSaS+K3j9X5k/crpgPphkm28aPu6+Zi5eDJmvmOkR3
F4la5XKGgdsfMBLoN8Jxp6n1P9lWHZFXAW7JX+WtSdlQYb82YkaFTXZMEH8SIjg1
q+DVmWTZy2ZE0ptiKjeovuiIyPvMCOH1NAFvfkIOJSiutEdRzIC+zmqxNuTsRDQO
vfuZwd3U2pNLxkSq68EVMHcvHqVn+Ww4PnhaJf27BYegNDCDNuIEPPb1z9ioFR9p
BBMqAVSk4pDQz15ctQpu+6jIbbsqDZweVl63ljlCHfA/6rtjB8wjYAeQzx2enZbx
uidkufUjdpvDXKfq7lyEg3kZ/7zuYVhJ/k6WwZHaPpr5q7ccrRHs/rr2zO1U4ylg
zVwlS3Wg6XYTFqHo769Nz6/fArANIQq7CZnt/0wzaaU4gEaZ4bmmIZB7zSpAjSuN
xdkF4ImiI2UMGzQJGHaazSWMFF/SYcV3BPwHuzNxQTbCIe2Zs/w9woZ/AO6AlNq4
4JLz+Zg4e0n53ptmXZvvJMGdxt1Tudkla71iGMZurEiCiO3RTOQBqTJet1LygotH
U2GFh+ezR9SJPRk6w1C6jeFvkRdldKZaw1+iYV9jPSFuqK9A9hqPA8NY5j8sKc00
ONj4EGUm8a5oWQHJPfen0diaDKTGyJ0moNngpSkz5YVUkjdrrbCEb/tI6wI/SmEZ
xMiXWLT+Mv2IKh+kVSr0hnfk6E8N+82uZNJS72rJRuTTLRc3TmiMc5T3ZTamnz4Q
lVzU8MGmgD1i0NItfTBd/KuS/+OgLrF9/deYY2KH8MJ6fA3I1FQgZnrhSAYS3Fbi
rrzmPr9jCP/0pSXdO2HhpXmM26pmlU8jbCYnMANDtzHcVo2oe7+GuUL0suR8OVN7
uM/AigNuayrQfxL6LpiJgb6etu8ImV8TqpCyWbfdGszYrRyw1KJYtS9ZXWO7j6bS
NAqd7MShHqts5ukeRbt6caipIlGgZ1dVCzqS26vRieTIsRS1b0tzJqduTGNajFce
zFzTHLjAkaUK68eq+lq8R91EJPMDQhW7Nss3X6GZ/QK/NmKjGas4DAPt9Onvc489
14BVKBzURh1KI5CnHIb1uVNH+wPLLXjIw7Gr24pOFEczUZ7G3KZrBkB8MlFBKBaH
HRnw1Zi7HlC3zyPPQSPe7LohDNNM3jCcGhinx9Eb30jldBVOx977TrTjuTf5It3b
wS2kKIJovMloHIysKxt3vHo5ma/KNjNzufiDTFNx6ODRYuq+LuhBVv6117cNgkiY
B4M7Em28HoRnEvmZJJNXIv7L+oRtHPBIA0W720gzph3ykmd1ryxJPEfeJdixPEQO
C2Iai6g1jocWFs/OyxcZYUGpsDVEd5oJF/0Od9a6Jhp3kYVSZkDO50LX6Xol72Wy
ylTMhT9wyrsSz1Fh+TtyYVpv/A7skFMzyEBnWBF8FMOXXXsy0QdkDYhf8sDsme/N
fl9yIR4066QXI3TqP3AVkc8K/cZQBVay7CaKBKx26+wTEDIRs9z/Huprbq9hkl3d
2oTGYw5PeYDqSvYwbtCwvo1Ntj1jVzNSxC8Rnd6LVnoj9zMTsTyAf2lMGSkrYjya
mLMi0506j1RwiePwaDF2VwhvfHSnwH7L5mSf7BV7p8CC/c1Idya6ea3xqk6L1Xv3
NOUx4hXYqFx7lVr2ood2ZR8z9VObDOTShbLPmKH7K5cevKdrrdlb52mEAddbQtqI
7MutFZURYllEyE2cCSIQNrg6V/M4hR2PqBu2R3z2uYhlfo3Q7ATpwo4D3JQGArgb
oddQ2aw5bjvAVoyetKznvLs7k5N/rOGFyhdD5zYAFcz45T1r627cxYRavkC+y7d1
toalB44YxdCLh47cNtyguA2fLv/bGfh8mHTJflOuwfUgRKFX1DNtzvPoFaK/MNDF
pX74TkzQxasggl+XGQZDtox0odLrbBHVF5Bnzf2q/gj13D9tYI2jKkwDQNbMl9a2
8KLTj5QedZxYNs+W6tO2ymQ7UaEV4CnaUO89DnrTJ9DaEEepGvzxikiVvIJLCoSR
wK/n35wEvNp4oGiatwOaNlUIGNvtjM1gdUvraEVp6PWGj31RVHwmmQw3ec/GCyQ6
6wbDVwXglvdUDwd31onjhXJaS1G5GABns/vlgEOsDYuvlicMLjYbBR+QO9RcAlDr
gnMlmceqVMPXD5FAwcua5p6WLpTwLD0E4HRMcXZzbUd/m0kaVDLsw0ICftW6rEVk
k4waBJtRJvvOqvoss3LBeFxzq7b57jCVpivwiVvPxrUHxnm3ggC62VZ7k41fHhuG
JZ1rBLf6ck9q42bQ1lw2KKy9ETBTPtQMNDjLa0u4a5ga5ozajgh7VcuHPiVT6A9D
xkoLyUXklSd5OKkae/wvFKgBXnE9/Qn0A++WgqGBq4JEBrtE7i1O0DPwtTLwrgy6
h8ROE1TnPWND2U+qPhor2QJINN/0esGruzQfKS8YhUmELbS7dZ8U1bOj+6e67weH
zmsmE9A9GcejT54uiJdC20f/ycVCMCZ+flRyfXyVYaDU7h5d9vPhV4p4FYoLG+Jg
E64raFxGB9YxNHtBGv8f/yn6+x0F02/RAww1XGgK2IaVuLjz/jEjMzVxIRTDW409
gzrghI4Eqqs0AD+5bJ54sCQqev/8PoPU+g3udAR0Nfa73ALjjbGjs8w6sXT1LKnu
nWSzJzqxoySRq8bgWOW56751TBYuMy1/JG6gjsg8nJhoL8v1c2ob8N8TwrijdfJI
5AAAw1lKsZpFrxIb7+8PZVKzsSVqoGU51FZ9ideN0+ovSBstI8SPjMsPYQcQa1gv
s1qgQ4osc1ILB3HAnSm2Z7hkv8JgHf/yMgUYt6wdHhxQtLVujdEuTErovIZbhuis
4xZTUWMAc+3malxbpzaiXcYGQJpdvdRPR4EMRXPVe0YhUo2ijCaK9UOJJr0lfJXb
6biY9OXXDLXQxQ+GGOjr/BcdflXXynmQBPPbXA3HG2FL6HZ+LLjKrNfB+9tl5/FE
uk02fPewj7dNcYRLhIWgpJn5ersvm5BAnOZX3/ebUIHq8uDyYiz65OArj5jrLg9L
6C+Pa8ERzuVGZeZDOjaK5UZqS84mjaviv4BVqvUQZDkN9aGY/3so5RhDAiaqk0kS
nHRfTqrlJ51YpuwSaocU9EmQTkQNy7KQXVBsU3ojOZDo+32XC4vnoCunlJ/r1VaW
H7VBP6IdGwozmh12ZmBhTgXIJcbkrY9g2m0pySyhlTKT1fdDEzoYDCyrlcW5rzLD
+aisjVDLkDOmt2A8//FN1IfXnoTVeWT7UeFR4uLKEf8rPEpkvOQxYgDHsNTggpF4
pb41+e1DAUKKQnOXMM6YaHF8qCVTbbmbJPZqfKF6PzEx8fcBZlrlrK/FB1oi721D
sG49Kt1QcKe5QXNoh2n42HzJ96sBYbB4HULVcqQZ0oOUpHTDwbdgjVy/eQTQvfAK
6Wn2Rt0gxrZT2V3jSpOJz+oVaOgB55ynF8G7fuvhMCzwe73cIWQ3wkK32cFk3F3B
Nn6jQ4wLzz6Csswr+gvPg2C21biru5RLl5nUDzl5gItl7X26G7shfjdyqddKYWB/
hzl6ZRSgayPi3RIuWRIySQtnPY6IWPhiwljk+GiehjUT8YavAP/2u7Xyocc6vDuh
VurEX/bdBl84HVFaNrYjiS8OVS/YP/PA8LHipeqdxmLvothDURp5NT/hxeqWzLvS
kpiI8E8gZW2LSb5cMNc0u9gxzHoDLnza6GgzTRpiMP/l0Wb0EuvTUNlVXl6m0CpD
PnxsiDVOSqaPmMLNa/yxMl9jEMdoUcXep6g6tT2u8F9TpwmmhEK5OoPTCM8hrvit
1uhUamwCVl3JuDESGWaGd9ieURpUS7hvtX3ZGmidIk4nCCpqw8C9QyQ111k4vSBi
5QCCumxTfUlOz05Uu18OfTwMyPh2Jo73Ka0jNQOfyVJ6UbA/nJQip3TMpmdFThT/
3Bw067bI1k6IzgCAeLyAfoENkpQtR/c9A+rr0CbNezgfF6smIN/vrpKXMHwFRQwn
jgdBlgH3WWJZiT5YX8BJQDEougoCxi3AqDWGhD89OON9zOfG7gfTl9xCY3rboQwC
g6WAA9Trz3S0X0oiORKmjCJ/6bZeJiqQUaKG47B1n2vXGJh8AR92fiMHjmFU1/qy
1R9VvZdmGZw11sZ1TCxplHh4t/paYiDMWlVAIcVKeYfzsLx5FLtrJxkYrubTkeD+
chv95e70IrhlEGoXCsVn8xxrgoZno/W1/UR94gg5T0ca93mydxIEukBgbdb83D5H
cnkM7AMddnuyUfx5MALTzlqpRS5dJ70KvH/R9In58C9s8Z4hls4ftwZzJ8vnsa9g
bbOp767l78lGNSsx3GbfZQ3icl6bAt7J7ISFW/oJaUIv6nHcdE5ewdljq8jgu2yl
LXmq/ZkxGmu154eJuML/g7OTMUOZa1tMnUGF9uh/XQgZV8KPVNs11y8AHSO69s0y
3woG83mGNcxW4gxJRQqku75lHUqLqEEpJviOnY/qjqBuRglcn/YLhRTJSZ+wagr8
PVrmGedvT0mWS8vrDulrLAzlw5Df0o7dr5o3Erc8TlUEUz3CvIgSz8j9cVKXWk48
xUpiyUqDtTp8dGnJT2OKixwW67JS/8rqA/0cqXR20FosjymrX3hJxjS0pFciIxrv
53DhR1O7mOx3tc/q8tpaHAdY30CxrqvCwqZikcAvPTE4gX1jzHLm5/PjzC7Vx8Od
rKZCSi7/sH/9vxY/Ng47EMduJsl3oXcg3CFmJKHYwnWJuPQde43YD0uRSRNdTeHo
6JBXTkp59puYnJpxEgGAkhp5Mx8XgL3qPGrsGs+DEkz0+LbkOtlpK8IfsyY4aPkn
nVemKtMidy0LklkHjPXlWo+onn6SNb1oUDvaV9TLcjKFz6G+8DUaHeqFjoV4QUEd
CQ+WfK7aqsmRckD/BKw2kSwLZaTwkKSAzMOVkb8RgZoaCvEfideFrJe9v99mV6ym
Kmj3Anw6KLCYrU/Jvoi3jBpb7iS0vKP9yZJFj7FU9TDSswVHazCKLDdg7XwNVFTd
KCFpHkUwTn3V8KfWMo7/03qPPstIL0c8DCtSKmc/WESHOiPHfFcbOYfTeWG7jRvl
A4lI8GP4ReTf82e6vK79fBJMlYHxacv04MalEG3SGB5BIw6eCkDgkYxdv+Jb9LGf
pcpDti0Jb80oZ5yZrVw5GmGScK+qr6io1oNmXOTQr8Hq4T48N3HAT0dhuqOnY2d2
zWT4wCR4kCFgoYuw630H7yDm1VeMalPrPGYmAAb7/5o/rJraaAClgZ+vvz79EGg0
zLz6NVdTwmnEED763x/z664TRuaShQdx7nAlDBB+uSPC/blPuEfTtS4RkZyqAnLy
SIjq5yBw7cattNoS0cK1OetrQqrTWBiu8P/JqcUOaQzUb6f53+Go0u+fK4zUXJNH
tzzitbq9l1FxmCdPHjbD9RgeYpbViEOJU7JIpLSsuA2IAFNtAj18rn4/TbqIN85l
yjpUfH06iwghXqmTEVUVq1cntg2M2TaYKLSsQN4LKGGTGRc0M1erHE2VFgW0taQe
mLTcbMBiKQ0dALOmbAbaO+L2WbdJkDWeQbJgNC0OxIQVIzLqMR6+J/r+kn9614r3
PrsMCJIY9BnU6DCatqDKLUPV5Mz5+0f2q45cbf5I71VLDz6fNOFPolmOIoA4FY5G
XV+am5ZY2ePFq11U6G2tObL3c3JgMTF+6l5sf8lIrjV2qIFoLT5cyYuMFwYWPB3E
HUggMO1ErovehYPJ1u3mSBSjBtpaj7uwpHjsxXkE2jxdV2dJLE9PvE1R5WW3ddA3
e03LSzXK1kIzMU80esOA+nlwIs4Gf15FLkJtRSJY3JAkfXzthVEZyEsokRr6HjMj
XydyXrQMW5kMtLtZbDgabIjoxdKPtIupp64Nz6h83XeSenaQyukHjkpoqt4xM33b
UykWg86qKWiA1FhtN10srzuw2LFXztzPL1Pgw9vrShv+shy8Nktyf0BAzOek1kc6
038z2JLNQpm2NTQWiWeGRPRoZuYjo6SBGclGdajt43g65T76nKZGLeUj/8pW1Jr9
TK0cDbKJatqK6VunmeX9X2XcensDHeThJ+hz6eSnU6VGlIe4SDn0tjQs4Xy89D4y
f08Ih+MYOF0O3niEmAKcVRdEAK56gpA++ndwbxalHEFlzPyFTsVxjNrEcic1wmY6
IypkKSObFX211jcG/QJK4P5oU08cCmUjHYzal4EfiB6gLeZaNO3OrjCBDS7SzKxs
xGwQLl+d4+Fnd7J0Im5kkPF6BZxmIfPLPJols99gbAlID7470JjXHvqw07y/nVki
yaGxuPLz0iYnDui7p1TO7+WtnYF2P5KqE1Mjlw0f+gzDikGDg1wgPU5jMb4Srx6R
u04/Go1TjxMnX8bBAhnPMaBPraMW7GFcgbRRdq4K8l0oa4SQo4lvduCabSyvLUbZ
PjmxePm7K7r4lhy2TBNw049etiwTD9bl52/0jqJbRks8jru1T0IRPJUNOmWo98Rt
qL5BZ1WgA6D+Bctzh2qHD5ltg9mHdXiZ7/sUk3TR2/t2fI7h1YPnHwCP6CowFzks
7qfv+wJrsPX3nmWYNYSnshzMOSR+Wg0i3WOq8oPie1ne+ZugNGh8FjZjdWlb75Q7
Npg4+EVlogusQhVSyILmqpuB1jcyOyJyklG9g5cQ2ssRsb4Y/5XnJxod25gA+6Gy
6VBOO+qaH15bUvsrT05joMO7H6IblxlwNBbY04uk7bYtP8k47PvbBrqFPAv64QWH
+YXo2rsq/QednhlIA6XBD7dNgEBKztkMHkWYRkQg9oG0eUFf8MvTJdNSS+V5kehZ
2Sz8gQ4geBYvzj9xjs6GXIETtQi0aiybKbsthUdFY500Au+PGZsBu4WXYovYt/mB
cDzmpZdg5p2+FMqhyrdBT+f0m2T7aNRSg0D1kYz2W0TAB78+RbknsHC8UwTlNUpl
W3UHhqzpT6iBGXOnw+dBKAwxIl07oNdV2JhWPtvnWIo7Lp9u55PZ8xNVlMDbELs3
CyTN1wxkzITrBIbi6xSnJq3M2znswU/fOTLZyGrMOiaEt8UySEJeQuNjX3BXKiOy
iBMB1HNx4ODZogIR5WPoMq4b5JUJ+YH4JV4QQ3Wed2IPhRSsdihNnos7pBnvj38D
90Y5nBwRPi39vOlubdQ+PUUA51cJ9fbnmrXY02vUqmqHk/sSCAM5ICwz5KxzyDx5
LjcCX2yAHgZ5R9nfEDS5CbdeolLyiLbdPCytE/kr99dWSrEg2Gxr9uJXhSpGti/a
/EK1SJXJsuWbOBX/SUDd3fKvdRFd7H4l7CregJIVkPzun2nsq2kXesfg9GEzJzjV
aC9PF3mPaMbBQkiLwHmv8SQLol0Ptg0GCisk5i0tdW/A6alAHeMmkUBvTK9U/+/7
YojSlmPlPPEVsdLsRgs2Nr7Vl1YnmNruA/U31z/yyb45Y7Wxmgq95wkYTRO4irGi
wnsadQHmTnp034UaOFrUHI4ZPDzlLP1uwPWrB6c/G3yoe7A6QUMAT+VBUtMT5yn8
9pjD3fadt7xXcRWuKr9Yi8yOoOEzCwGV2agp4p6QqeT9AGo8sSSAOQXynz+IrLBV
jS/LbWxox1t/wE9dLszyjN6oY1hNfF/KII/iJoApNfUC5Rg8pSG1sOcnZw4ZJPq4
dLhEe8eeFLSl2FqgjFet16Fg4jB1axCossYjm/bagszzw+X86S/3bQJbWXJUcvTd
BMzer7bCBrFqj7PhLbUdjccwPDbFkZsaLvuP2edXROwdxyRczvMn/76PyT9M+e3W
01psdk6Uv4LqQJKw+0w26dvhsM5M1NddT64y2MM9fYmgSLHYHKzQ727609kvE5mo
MgJ34FEwerX0HUms+A3rVg7wXDGM9F2RZDo7k3ON2juQojlR9dHDvJrGCZXTs22g
XVsSQ887SlcC0ElXxiDS/z7mp2/RS89iLCk0EfoUIQgQ7v1KswmT+0uDJwwPyCNm
yNJgEM4PgvBEEVTGKxJpsfQWQx9CTqexeCNB9Ht4YtghkL+mL8/FPlRpxTixlEdH
Fcg9jEvBfVLIXc7g2rDbNIdtldfeMtzAKBfPZaXsVYWRJqod9JMG+nVF/vN/P7Q7
ksktyPLMU0iUUFcHQ8SsoPA1/TgW3lfaIRttXcx5cmwUkXyEFAf6tzflDm/Q3T1O
gBrt08EvzhibPYUR5t913HZlK5AE/HdhuftWNE9z3qIC3ahG2ce0oYfX6jSehMVV
AgwhPgHFM3YTSYnHyZxL6uSfpV0pLv3IE2r8arZo3zjnOAgLcacuc68DoWF7RulE
MWa+PmsshfKFBhAopPKso7JuLYn0Ul5EHV9ZFBmSN+Kj2oC+CoK2Nk66sKN6MDGc
sc0SG3CBmfQ5Wg4j8xmJtyML6Urdnm9CZI+ARCLDqqNjNiqgOazWG+uYwx1g/Mgu
fBvjqSpwWx4ZGmC1WPiK6V2muDzZRDX2l0ioU0KA2ZF3vW+8QaKXhzpBFyfMkRej
fVf74/CkI/06Oy/shKx0Cku5dxnl96OiqdY1GOvI67sKx5EwKacCncJMn+o+3eiu
FHHgjnln6FUTkIioKAdPKpWHrp7cBdhmPkMO2NHKU1MtH8azmielxE67FRIARSp1
J20OC1ovrs+GS1IcM6SlgsbbP2JkGwdxTsQIwME0BxtWzayZ2I3KzyFaNsVum7N+
G5FSst3TDZ6C5N8XZ/Lo2ECfaSPNUAbdnoca4geWPqaH/nRdteUKFq/l88f4eY8X
A15IOw57DgyAHfpjj8FauJcKcj/3keYiuWHzL2J/f9CJfp2UDE3mGXatDrT1bSxe
vqmHfQiLGEQ64NPtYivlEYth73vsa1lRtAdzvn4H2gR9SIk5OepS02QeJwyEMPCW
edXIqh4awdaac9L4rB1Ff0RP1hSzKWIls6IyZGIKNdcdYUJSZVgZB0O28TU1JPVo
d+tNQMzY//es85MGuAVFaz4qbcMV1NmadpxAZssL8FyMmWRWCOvxDxp57FL6Lc/W
hVScV1muvIQ9r2Sj23mIXbFVixVP2AhKCRPyxgFe134S6MkJ0EWZeDM65+G76s9Z
jMTQ4qUe9iAGTs7DnRnJcFaXLKfs85S2OSpfXvE2qZgtq4NoVvsUenXAIl3A8Num
vrPzkH5xLzn36Du0YJPN0UewoIKm8sB1j6FDQohrQVR59+i3sr9GtegBwKwcA3Y/
BOi6RfM5fT/b2OCsGZND/OfwALOKluK1lC+okNBZiFfCoxLvbkgQPNskZ9/GzZVA
l1Vrh9vw5ejT0pKfqSm3bMNmMzZKoGLijfN7AFVTYshB0hqRjW9DX/FyQ8QXA/27
dSW9bCGqUbKrS2mwTx29hEbniEMcxi6Ehci7bMyhg6SHXi6wK8vjGVzINi2nDdGr
UystdbBZ767eDz03R4qP2KePEdwypWz4XAUHfJmdNf/uX/p6PwpY/2a35HWDnEir
FkiezVU7QrmSWqBRAKUQYjQqVy7FnBSwOm1uuKwxtLfdq0OJJuTuYUxVbowV1Z2R
CrvZghBRHOlN8jgy/wDcrZP+9IBI6QnNzampItcJ/tPOlWj8P865FzFyjwgdzF21
PrjDdZFmaCGjF7CgllV4zFn2+TveVoPp8RGEjV/57JTQwlFUjqxAZsfcE5jAV9xd
ODNYP2oesev+wT2oJZhtbdwMNkwb+tWkV40Xbk1uIaQPM4FXxkg/Ajfp6zRu7ywB
2oJe8iyJHZVP4OLQHzrvGjfRPY9r7ZPZgeViAxq4JYcNIy3KRsvGLFLh6X7dPNwM
OSANLB5SwKxp6F02O28zE7uvwHY61sri0DNqT+QhgPdh7NWb29/YDXy9oyL/XS1D
nzXE2+JhFgYhLc0oUt47NCROWAoTW0WXmKFrukxeiFOgRlEK94tYUC/1C8L1H2bb
G9W2vCzSMqEBrfvXPsH7HVH6LknGJiPWJeFhtIXnil7hbpB5Ttz6reARwHh9pZ1B
NKs+qib+EwiCJYsX9axp3uy1I3LdBJ3sW6LBtfFL4aKxslCkDCPmnKt9taT64Gtj
VlyVxqoRCgezV9ERCc4rohSobFs8fYCX0Bf1qOpoR7I53m0Lpf3RyKL6WPyvU6LT
4c5o1Fq6RjKr2OvqZEuRKP+JKjPTZwHRhWrJ2XrUtMaZWWmf1+y3oXh14G5Mjk1K
i0Nd+xJTXbnLhyDuJwzDPs2Eq8wIbg2jctCZNgaQHP6JamolRnCE+7cQe11vUsqA
/bnnXJatYz6BqA1+Q+AFEf5sRMBnddV1IQrffbJiQMNkUm7Kyil3ddNzA0jzKwAQ
n0AYUqllRP+3y/2Zl1Cf5Nt/3LUPD06HhLEdBakgypRnr4/WO48eb//b+nQ+NMC9
OTzfHDKBYs/6z1mRjWuo9k4f0lPyJBNj5JWVLHz6wq6K2QayxpKmvH+E3GsDnkAR
RQiwKvqXEqSDf5GA3aG2H2bU/AvWqQ/9rXV9yTv2JkVDqzNcRDlOZ93kldQqmBRv
OyO3C5i/VyQ1m1Kp8tJepq3vOWGXVu9NB0tKty/g80FAJqKCYIMd0Xu0n/KsvqAb
Kfhk7vmewB2smI7LIvajyqjda1Ef+olDDz26BOHOkE9MbXPgE17xckqCzhSsyuaX
fIXOs+6pgB//feFpnSOqWhh8lkvXDSZrAnrXUN56pdfJW6GACQlpm5lKjT2dgU5z
L5OU07reV/bRsg39bWQqSIVZPDJ8Ey4Ybspq2DjSRHoWpXBUJE9kD9oT/TadaCok
SeDObjmNna6q+ZzJtJ0W9/y3shqHFciqLAn/s37sgzgFYFsvCsB4qlfdP+BfjlPQ
x8whjtQkEgrfhPEuxtIpW88zSM8dJnFVbF/GY4N3HwQMyapU8s3YSiVyEcs8Mlz/
E03ztpJLh508ZzmgwcZr0MtW8N+edUg5eaAar1Iyzd9YOSA2jHUTcizjuNk7lIgU
vpbHtcuKulbk2Fv49Qhx9EJe6IYMKPDZeR8yxMQg8Wa9hBZJyaGHrXil/wtdFy+X
A5U8E1AhlMw6IzpCpCTnsT9skYUhrWhb5FsxtEtrzM6X8PwhDS3zVo2ie2Zt3u5Y
rz42Jy2yH204HcUoOytavBAKKaMGnK4P8Qm5Lor7St3dEZdL0hrm4Gcj5fc821QA
Qu66h7X/zPD/5PgtIysTy8ymH0dUjZn1Y2B4V8gMnlgiY1nadRTvZVZbMozTyBGp
p6b2qRzvqir0ODZ/9Sv320agUpzj1ASvNIwk2tBvjwIDXEjGOh/xQ/sBIYbX25Fc
7sJm9vqOm236vbac032OWOcwKpOKwlGH2ygNZKnchp7H135z7RuVS/lOfDuVuaHs
Q11L4y/4h11is5Zu0dDh5q+mHsVsDuDQsI5iJlAgS0Mf+m4PHiunP7DodbPOjEI9
QypV9EoZq3gHOK5c4VLlOIEUj3lr89bzaP0UQDmR9+q7pfnN+mjDU6HEQhC+sNDj
VNWkWABsmX/kKI1OAYkrmWTJjfQM/UmarzHuYRYe8+OL8tQMcrXyE/HkvAxJoR5E
qJB3GGSfujDCfxnqhVofzUrme0QxkUrApCvnzStLg6GMNXhOc5Qo24thKC6eZC20
fcWHK2Tyg8jyTTTWQQfygKJOJTYZ3euey8I8/ALFU+ZUIHzp/aBmSUjjKCK5OkCu
RXXxu+bY1ivQo4zVKN6fZ8FEJIakKf/uk7hKmK2M+JfPmkGxU1NK+dlB6+Bhicli
BIZ4xZQpp2+pOrSEUfgy0OaIWo9SVmOpvul980HFk6apFMguOV7ZXe7TAtxdqDMd
qHM1b3eazyVXPjCD8h4Yl5+wx8dbz+VhWo+OAgMOgif1dLb/wYoZ0HpG1sKH6vZU
QKcip5XNZQPXv6WbmbvAkhlNcZErMoVhgz7RbaOUSTG2YzEWPv4orRA+sZD9o37y
vL5wvHr4slts/5LVFKMwm+QT1Ekvqje2a2jwlnxBzQBCe+VWkP+u+esxdyQIdELG
Fpt2t1RBGkM/xhbSDsZlS8ThRH8HkjEG8vGuvvuktvgnKKcHQYdxGzBM8C2N3APP
9JDdGzSTNNZ9MlnM82mpPkF88K/b3ge8CrfYJzlMcNSP5S7kmYoTCJVhzV34izPi
wx++j/JpBTjIpFGxmo0rZhhvsZwDTKOCYw+25THB0ch8aqtl1LDdiMj+k8fAaGlF
Gn0jFxe5JSXmZ5sgNUByFmXy73vnrhvvtfXoBpYWuCMey1Pg13PPi8FjeuYzyu9v
zS8brrATIGMjZMqCJnKH6DO65nO6F4VLOC50KNQO9kUoPe9xUOD1ExFu/5LwChTU
I9XXl0S8afceUk3xD/Tqc8Vv2hy7uw4uuHn2KwZsx9pcjoOWa+a9W7zG3WV+4hrF
RqUvTVYAnTy7QncKN6t9DJlsTzyDgphBID5QTAdphPgLuwg3q7ij4DnXstN34ptP
dPOn5FMxKa43kh35VUr8nm/O2ukTdKC1vEOEEgVoSStsk9KfL/F8uqVa/6VOL4Yl
lVcZwDwMOzgQ5pY01gHqBhDc0VSByb+o8pjn5dhY1Tjk9iPmPgw3C9IgDkl+gr3Z
oaSe0tguG1bm9ZnZe6QgkIA/8ztbZbaPIUIThf7dIwVwqosoMswgrsKgxPcdh/hH
TiuHtK2zraSiDHxXiFA2I6UOOFv2G5VWL/HjAP3AxU+OeGQni4qWyrie/1bm2e/A
ILt9FH4QLrUPfhPHxJ7YCCtEij+lF1Rt/lNEqWpwnav81K/hciwP3BaTZNdkfZdb
SL+rGaOaSm4/F5AEQ7b3xwNf8yoqQdajFgJ38882ds2iX5MYuIu8YgJUALzNSDKv
SHQKqqfUua0z0ybOG6bg2Zr4NFHxclJe/pyFjqZtumvdsFDFhvMN0ePpBth9B9pA
rMUaDkGt3uwKDoAcTmJjdrOj8rhbDe3MyX3fqqCgnL93l0L4INa3582426AadD+S
fCvJH2kFrrxTL9EHSB3pYY3jBasw6cFqj4IlN/nTmyueyt3nXmTUvhQ1s2ECxAwm
JwW26j4Uz2KvPi7h6RafjJF+JODxGGOxeQBB+gvk/WsgPAztyKdLAPlohHzxmw5X
hhGADi7Qa5mpUBoMKUutJkvQTkfKF9G5LiA2L9R2IPYeLkjjDz8LuA8BhHmZ+bfG
jeP+XzTS6xHI+qePSCikkjZK/zwP/FsyjGkEEGnmRfSclw472HOmMjZGerEFAqMz
bEYyDDyRC6gCv4ebG8VohZuPNhGPFssqTkH2wEOUkNR+6ETiUfry24aVOS71VkpG
retsAwOajoEk4t9apkrvBgORqV0190sXwRYcDVwkYM0a7Xv3XOEQVo+PTFk/0Xrp
e6lhpc6IjdqC3oAxMN9kPTH0MRYNs0tOQ1/Ab8l1ySysA15gmdokwo7i30UN6Z9N
afOyz1FKpy0RzpGLeHq/fZjOhGxSZlm+SQO0vcIgJf8JYk0fe9x91CwX51wg7TTf
l02QQI99LEu4RlKKwtLDjzKfsz1mpJxs7Dwl2DJVDGw60JHhVghIKqnR/LozgSoo
4/pYgafNPiJqlJ3cDgihHefNkgGLfHkB4IfMedh/ZBDc+TC8YmjnVjYYes++SHtq
fYSpCsGeG5ViD2esXmxKLs/QowtMNRSpkNKFYDJaAmFxRTj1N4RMAEoRVqEu+vJv
rpTtAZ7LVTKb2OH7korJfR4xSFDekJD7U3gsJ9C5wYnTkgcGJ7YVagaJjmGV8ai3
jH46gQU+tLUOStLd9WxgDuU+YqoTS6qzjk6pc/MTzWIndzvEbW8G8wclL/hkPwUC
uo4n8lz2RGBUclvMNvWNFrHWYjFyeI2NqAj+ho9rHnrwKuwtJsm05LOplAaH274Z
ZUXV//lcJZIdgReHHtPjVT6QmwI5wh7QIwTEGiuxgaUxKnPW+xyMvR9ZkyGHIOAV
qPYjzO4liTvG5IJoEXRhaTotqv85Yo9Ctu+I8RdTuPeRad7T8dIvZCPLLXiPHsuy
hBj5rMUoBNey33qkgx9QAQGD8vXGlytqHkIglYpxNXbpptZt1GORVDbxUgoc+h1f
L9t7UU5zEy2EAj26nLS9eEn3JfvlB591F27xYbXAgtBMVqVLoh4q9IDMZT0u9WBl
PChK15Di+5gZzLOOzf3o24gXpoATDGspmUBvdWEXnrk/wuGlbcJCexmdNt17p/pq
eYZPZVxkqzLY79Q9gyU/LmIoCuwq+A3JqhFmVeGNHaPgg6PgwDhVrElbbH4GB3Mk
A04o0neOQ1xTKdH35NWj4BW8QO90mRxm1837jCsjQxuKL7KtEVvVyc/n1W5aRRaN
P1RGHrM5yfurcmS7QtyViqRCR7J9xYjsDNw9VxIBz4jdJd9jgwz0Q+f7rWx2yUW+
jEA995qJl5O3CuWNP/zm+RYWZK3oRLGrkw62Sw4odyHdh5UGKj4b9ViZpgwZB2Wb
pDiWrD4gRG7JTLP/mS9bTRyrFNcxT4BGGB8ASlBkfkM1BXgLO/e2Nbql2Rr5nvZT
jaS+sHVbc2xdvU4hjzGZGie23jPI3nMYjJsyKP5/SFAQ5DyLjexIQANQ/e6FgiyX
UBWq3a9YxHw8xj3YDRc1Ovsf2392AYybKANQb0zS7htohqp2KlLma2ueCFe+cohv
V7ZuAB8RdApZOzsgrv5a/kkdxEJMIsHRglf1AmxkAp/1savTTgadGQInTTsArBsS
j7myj0GNd+6ruhvtd2vrhVBGyPC6O1uK378WkGqKecIm1zMGSOpCAJZuvTi38DhM
8wta1TlzOk4x43VFZaYKJwtmUkywW4edA7jk65xN0GNd2yU/rqmR0Yaz1X3IJ3zF
gyLhg3uUa4EDR7Z7XDV0kI9gHP5JeeerOjHmLly5KtbNpb6vd+TDqFVCbLLQdPWD
vm4SggDEneWtmuB82r8k9laP2iM1GIS7ZdIZ0lXcKLvWmY3FOZYs3X6g2hAwZXCs
/ChTcOHTY8ze/6EyZyLt0Ss4nHWL4pMNKR1dDiqVzc0tXfLAHZ5+37/3p5tuHuNH
no2nsRQthli0gq7DVAwlsC+iuQDa+z5OYaphEtsbrdPwQ6+yKyuEeLcBi7mJH1z5
oGdG0ivsMtQzj7YK+t9mnhrltS58prrAPYhjAJVj+QDkSjZGgSNvxJmjfueeiuHa
OWfAhBlo9qEgkbo/uLEVW9ZvoXNnJUSRt3Bpg8GzuwlHqOyc7VUERRj8IpAkL1SH
DlJrF8DivaUT3X2s5FIr6zZxQugbU8AAFJg6VVMEFxlPqodUEqXkeb65FjwI+wM1
x1vDyh9XoHEcxnnd+Z+igNlVQqLrPt/MfA2gGZ5DkM5DT0BLRV14jb9/m5RWSEF7
LmtGM5QKnTcRKpa/30wJjbAEC2B0l5vlip4BnbYxLYjUDDd7jFFdR3WPFhCYTXYE
0g4yt+Q/rThxs5cTupq3dxfxaZiW5wL9IHy9dm1zbFZLA91gninEGf9U1aGy+zE4
9rqqT4LlgUZ4UnmQ8F2U+Kmmc3SKFGGpZLBupo6A0YvFAMYeCF6N8kmOxpckGTC2
ivYvqMFfpgr24Ze1BPASx3pb89vRRnvVQhrpoQIZESVdbWsk2vaK5He3/VF8nhvM
UIUWNX/xjdd4g/cCfq9umySXkwna0EQYDmYCOSOLjNdi0SG2POIJeDckq57jBIdu
k3jN8Tyb/UUuBF/wjznwHHVFXVp55nXpLtcrcUAZqFSb2ZYwJKbp5BtJ3ikuiP68
TTNG6jqT5Syv0fa7aDIMBew+/fg9K5/rM04coJ+n7d3nl8CBw7Z/7cUqnOxgDbif
lpdhF5yjpXbga321XqtolTZV16jl26vd6JC1+6F+Z7+/gRVtvXhit9lWwZtV3F/o
qGkANLc272VB61NTa7NkhyfMbxBXYqr6DW6dkAVdGeP87aB4P+KYKG/pCDmW67W9
GLmoKp0b0ed5QFo1Q8mcwTDM6k4bltLom5Si3XaUHrr099xtCPuwv1ipjL0nQPSz
Kp2/fPH5BELuUnCHNXfhMh3e/g+S60F8IBWFkAarI4g879h0iSH01IGe/UWOoKRT
PO1Vh6a7qw+bIlDwJLlPuqbyweezSOk8naJoNkwGVyi7qH93bFMYs4WuwoMTCas1
BmOH/FbfDV1M1sR98AwwNibbPczKP6ClvjiQCrHT8JkMgATDyhnwDYXdAsddiARe
PqB9T3qbLYZlBExMIflVjGM4jaN1cFzZ82PXFMiuGSTSPjzyScdZvAtReNRKoxsC
MxjQPmQSAlCRCAQEX/FtKs5+BfYMwFdzv8hgAyhm07KDqTZPal3aftvegrVPUFOv
4ycI0+7f8RZ2ZbsRPaYmee3g10mpPxqmivZhL+91u5fEQvHeysvjtYup4hs5dsry
vIig9IVr04cfTh1QY1OhBfEJtzJIukF3/aB/NPyxDs2tU2Zp+EZYGXSZIpJ5acKE
u1yVg9MF8nzN4mcf80FqBSyPfDz4irpnQXIKVtw9NTjERaIh1EqJKR1ExXe3sSv4
aCsHXPY4yiWSRckizjBqWYY0j8cmDoFM47IqOAIm+g0/6ARY/hCl+g3F1ZjH2JuP
WzJnv6uSLoR7KqWFuO+G6xhu8x/RfOCT8/DQo7JLaGzk5OcZpD356Lsh69trCBC6
rhynfOvq8FQjOBhGRVwGkthOTG8cSm35KVFJCyXp2qb++D+NLDoPvBES92Flb4VP
ivYi9s4At8wWO0Zw30EzHwObRBdTYYessU781GZXvXbJstZGJnJUEYVaiO3pXMkc
7QaX/OFYaadTeB8OCDTopGJK1MCX1Vdo0sBAV7L7jc5KobPVIveKJp1VyVAo+qnu
tlqBnWfKn/DSS8V0t4vXuQCnkxh7ICElAdptv+iJvNzi+l1bpXxTqhcijGay+qkW
tXTiAhXSR7J+ZIMHbGAfzU5Qmp2GBn+aKjQtjUHcsyPxMP3tNUWm+MyYnrkiC8o9
cYaAob9oT3A5dQHzJgxdlkrvCInBf77Ee5hy1+ZtCNFB3R08l7M6LnAR8Dfj2RSA
XTbJdm9jZeMQjVft2csUeaxLNXF96OlpnhG/Gm+rT45KfD1L11xGOe+TSylC3jgH
Hecb9yImkt9R8GhdRhpLhSPrmaYQpKqzCSEckuVBoPBmr64FANBJh+ip0h3U0e5s
oGyrEV1UGbzpcvc5Jzh45DFJTO0uwmm2b9Mhj0xxZMmeGIsoMNjWNXst+ltN6VLS
czOYaPqw9t59B78vowmps5a2N0/eZGwMrBVQtgJvXjMrr9E+4BtaxBpKq88PtxJE
vd00ugFFyTkGXLZSzR8bY2TFRMJrobxL3mDs6gqVMZcITPTOAw8p5E39L8MsSamh
dwK9/dtZDIwnj1BLZkZP0McPBZlh1ZgyaTs18gvzF/GnWU06zGDytIykGvdKM//6
f7c3eNbnvLO/xN7pWBoMRqJmxoOYuuEX2x0yICq+ooSDuhbROyKQp6g1OtWwaTjC
8wla4jXJwujst6Q9CGFIgTNW4qtxwChitnjpuT3ot4/snkzze1s3TE12zgJfgDdz
F+y18MmmX8PpFBEmQGQPmYXaQefoqKQgDfD+hYRQw50wLjp/mniJo1ApKOg6tMVh
c3vNnK7do/536sH7CyogBjbi1neDptBGkTsioWDOpdd1pYI/2kRlmsjT2nvghirR
WmKocaKf+DRv4ww/OdDoIAQgpGbqTObfmAXd1DnqSODc+B4AbwE87f2F4aP0dTBJ
srYtTbu2DMWl1SOhxtFbGzNR+fVSttE+rSHxjMPXxnIBSjm7K1xjznui5v7NawYB
yBqeeiZ2O7dvd1IVgkBQlQvv4ffSKcIY89ufBAQ2G1L20BpuMxlUlMtYpyd27wbg
Gpxta2CB3YuAyS/j7Ne47bH1Bg2R9U6pNlvzY256pvv25f829v5OZeTXFX3my2Ua
v1OP/0ge9nbmVpmiKfnR5G4Z/uYkO89ffgEvVGpMH/OImF3JsNoFmkqtwUGfH9Me
OEznwbdCx6kGiKPV64Z2YGnE5XFxUtzqBG6Tx1H7xkM2tjhLOzdc93wVMfjkR6kD
utldYQra87VFhYjJKVnV3iyp56+RqiNmW7ubaThq+y2fif8RrGk31YuZElkX1aZ4
6+C47xJlZKwxHGZ5MiuSrzFYJvcfORSkDcEtQXsGCv07kXoCP1I1AEUstF76Vd+6
48TzGlYKX3Isp8/N5w2jw423GchJgD91FRewkf5tAz2KV3MtwqsOht7cSLN8Aw/H
VN9cZ1HUssigKe5fClnJzLSPAdixm08kMN4nSgVVCiI21mY7AHecpSzyIyfFtx0Y
5Ic9yo53kq68snsVQef+ERRotljOmeiBM2GJDvp2KFahYL7d+79cFSJI2iaJ3CIZ
R+dDSOBgBOuAWYpzkLxrG9YkD8wjkLe9adSoozn6S7ZwQrJ7aLfcgr9kyVNeaVPQ
/NaiFEYRMyoX+fOI41pPLNSLPHTvetao5+6ICku1MYFQi3evSuMYmXDD29n52zQ+
PHVeT1GWA83Y7UCan2/3HfaWQPn1kfJqZig86CfQzGoBE69ydZ4iOkDylgJfhoNO
bSIJnK0smzd/ZqC8KlZdPkGTwOUvSuBeAsxjRACtFm7JlGF89Oy0VWIecM2IwwqA
VYYj/6p0u6eDxi6rcXWB39GjQvuq3ov0b3XAObDE+Ll1IqdNKNWUlmVh/hR4kdaR
qzknSEt8Fcm5WOOCn5mSJzErEzmaKoX7yjst+YXogFC8KkPBi7upHcqvXO5p2UDc
IH6wLJ89H6wt017jiE8sC3oqAnAXvDuHtNt1QjuwaDkBhQajBIMV/TJx14S/5dPY
eWDes+dxa2mk+kDiJhUs1oVrzSMb2proK5NV2xbUraKAVN++mV0ZT6C640ul407v
tk9S0IDzllojK3JV4aqjAhLY2ySsUf7NhdLUkwyBH1kLCuoK9eRe+6FRnUJb2wCf
vTFUmyNEsTv/aJvZIckE+aHjifRsxr8kn0OxKNrwQKdmhEwoo+j2/k7+8hMmUFWD
+P+7BimNJ3y0XrKaVGqYp1vlNZYBWD6Cmvw7gvItvnFPaO6JXRUABQHOpAzuci6L
Gtl8ABUbZwyhEsM9f1u2hLtbr5CT1tJVWby2NRvL6Ip7tag681HGS6XL+7aKlm61
889Ighvg2hzMMPNR6Kvf7zOUCvhTYWzQtUhZ+hJtii6Q3b+4W1xHyqVB9Ektuph1
ZMzXVxL4wQca//w802GBtMtuTawraFw20+24xsB4c5SYKHH0oCH4PkvRw/GGlmVi
WUBGA4+eWzRo5wEWgxj0MFQFHB3iJB7dl9+LjSF5ESEZLvZG3VlWaqKL/Sun1ixZ
YraXuNKxs/h550wtR5FahWG0OSm85zgQxY3QpoXLW30HrNbCz3JIQ2weWx+SbWgC
fkivgXeFZTk5KHNojHDa6KVgviVSGLGgmhL1WnPCOWEw5Yunt9i0LfRAPXiLoP1s
Cs/iMc/zlUT/KV17nK17rLDN77t5oc13GnOg67W1LGGM+ttq6GrnBlOQ+FUQAjs/
oWkrjRLBAztAA5D13Eqhny0ARK+dJTM75vZXTcMe5RZxEQjp0191Zq0WaRdMeS6t
g6leWjF5Kav2mMt/6fec2mzkaqKXZDfMc6us4y2gxz4Hs8ZTzq4BvJglxiPx8ROt
cOn1o6MrenmNtBeb6PVFPC2CiMpJN2qQ9744Ks7eCxDaKrGFZoqtjTUfpy5qL/4i
uAiBdCGUOr7TyiV4mBQcY0E/1iBNoyrbeuhi2ZBr28lHqNcqLsPds83EoBGPxgqv
pZXLNM2SyhFaN4NkgbVVwVg0Mme+mBdwJVh6SzY4ysVeqzFN66SToasa1IeqZaBq
hqg8KvjfI+7SblN7rma7ncV+5x0IqM7aS3ne4JktCUMxmYRpxCHBrOG8OgvVHYng
pVVX/IxhtBDqErZhtnJ1g3tf6fg2UxK3FkvxZqiIOmHjKol4lMu7S2V7Rebz4StA
sx9YywrUORvkulrtQv4wQDK+8a+f6dSNVOuaKiCLc8A/o9fbu8x+aW66CorocQd1
84RZcompvoRBqn6Q04bnIwo9ScQwguCUK3pjIGsCxUZ79ZLjdeyNFRENNo/NiNnk
c20OFhSKdMTFhuTDN7d+z/bJ7N0hiYVTUgO/EcQD936lQOAFkH8+PcDUFdRQe5uc
A8llPC4LyO5LEobuqejQvCOvw3APJj0yh2ej+klmGdztxpu+UQS8dWHuS/l1Ckzs
5gWd3eLEKCuBfJt3DBT792bBDbbQIAdoNaFrHQRXEckxq8OnJ64/ieg9zL1qI8Km
VpraRfACDzkSe/kmWWfQXH2vFnPIOYNT0uv6PXAlzbxnxJr56+S+16oW6+jp+rW7
MBFXKLMuRxDikcjz2453aDD/Zb3yBV/9I1er76Mnw9cIHbJB7IG3Q/1F6XpLBr8D
wPNbYnGIEJkJsElqSxvA0Qv5dhfEd8WYjAvIE9uGbDIiOA3WuHagCCUIJ9tO+hfg
4G0jpY5P8ZgWFDmpAD89+03EgAtwb1QgRARDjWRVO1q/NeqE+dlQN5w9OlvGeaBw
yuC15y0iNVUU3Uoql0A9hATA4/AnFD2oKL0I8ysa/NVz3WOcYbAtPQvn0XARNzS7
DTOCyFw7V7xo7DsdwmKSxSaft5wNEoK685xQv8t1vnhJOIpUOBVcmMKcoYJRb2ER
l9Gj0fVw4RUWpwuO8GQGMHMfJfFSmUCIbBEnFoGpxFBV4v54zT5YOFMsRxPYbA+e
zjynkNmPvL9xJns2i8rtTtOWjebjB8hFBxJTL6xWWccyeFDR73EGIw5PANia3UEQ
46RKEDdzDkNZ7ToImTo1xGvUrYnI+EOAs2au4G0zp6PP6muLMcOpIhgimmHwz3Vw
LRvV+hxt/fQuNKHh9s5L/5xzBBdlWV9XjI00RBz1jfuO01R9EAazgmcdVwqOvJXR
u4pASPGsvJfxBAmxbhA8YTVtPsP99kuUZR3QyktlzRAIPBXRSKszwm3WfW95gAdA
/JZrLjw8Ku10GbxaRGYVRYUD6nzrFr35hkqNKw0YALP+w1+EGEs5sLgTFPxBKhQh
1TKaNQO3oOSAQrJXiYI1CGrFE1U+G6JMwNiaqQAnpPBwUXxNKQptQEYFNDEgwV2o
HLpp6BUxniYKslXN5M6bBpqqahWXn1d2UuVA5P7diwFYHBauL0b7+pI3/4lr7ite
N11qSzUrk3HD++9ta4RGAms9/ZCJD9oPnsJnVPc+Pjl1czH1SMwBrRVR2wyMYNSN
g7tRDYZZOnBwOkpR57/EKkpTminteo8Tg6DEfQUjRR2c4fi6u9BvF/ZuquNje+Jr
4gvvT32pycn4mIsDzOqTbZP6yuq2mtF0gc9pfWsPkDzMlBT+ETlJYX9oZ2+Q4yow
MdE9i5XI5VpM3TUZvBrEG3cU/FNg4wd6Hfug22TZq9moZmQvZDHCaA3/r/K98KBd
sAvZ00no1SB9j8VkYoTrfQiDJJbsfNvfhj6p+YQz9LG7CxJm2q/3cQgGCtLwD4ok
2AHDt1lHTa8BQTiZCbMZlAPT/BRs+Rg9o1slDNLK5gdYy0ykB4wD9Tld5IhMzfTj
yU9O7sA+rHtKJWBW+kLeWMgeAvIQYbaM4+rRT1MCuUNOKzHoFUA9NzvJYp0pC9p7
kb8IYDj4BfrcbgXY1F+DwE3nbxOl5l6QTkXDWvuHTMmQps98lsKJzy9eJAfh0D1o
hXfuJUjyl6NaC1kMBh+dUERUiQ4Ga4i25wuM+hSQl9G6il8UpEu5s6jlcSZqlHxZ
18YESUufTteuycPjeZ6UqO2YFMoFkWmjjPJLqam+b5J4sKYPzZX/kpcY/2VUjNEf
U/vvhcRl4+sBES9WZ9uJf2qK0xDDdY9JDalMJViPFjXXWltjUgA5bQV/MbGQaIQH
rpwF0zqOtyvxCE1Gk/Jxk7utUcM1ZWC+iRuxxWguk1gzWx2vD9XcPm3pn39D99zk
h8cnzIpTLxZsZ0YF7QsW/dDQeXUSTTXV1KoXCe8AWOkmlEx0MbBSwCOlQWRYRjmR
3O7BXM/NQp6n6+pZtGFDlU2q34Fg95lGNURBU0FoxVQC4NHcg/RQ2VbYMIuE6Hbu
fOHpmszLtsrXIJatic2aibRVPZWaW8GXwi1HFlW++sg0lILOPOF17pd4No89R074
u3PU4+ICHXx7JPKQUGxRzHo9rdcAHb8DdvJsqifbvRhyCDhwRm7AlWLnU66UxxHi
ERLSN5RkBuOyU4iVWTI30FTBe3zkW5seXi8kZTuS0yXKPing6JzidNQjV2yThBRb
PX87uMkNffmxjCv5ZaDSjJlhuVtcuNaYsBYqUtuWSii5IeCv7ODr5OuZLbMl3LkD
IGNF/dati+hkYNPXVC/M4+icqIKHKxm7Ntog5kVbPs+o3PUW1dnympS8dMhWUFRE
XX13y6zVy1xUI6NqaWN7q2+Doisun2XIDoPu/iruLj46YJ/mvEYY1nZ+VHd/TPBL
vLqjZBL9mPy3QglKwwvPXy6kRW1UDVuzVe02cahIPJCfaubg7tEi+nLhPkSs7U4v
BcsHV4fZl0C4/0mJI5wtWoyVrBjQwHadYtM3OoyHzyVOXTKl3fiMtcY5H2huQ3Zi
cQew+/XNU1T6BBQNc+UjlzzX9rfSo9pW4k4b8ey0vErzMl345YbVmPiiTKqQp+hT
KERz3e1E6I8qmXSSLby1zUK+umy2hmJcD0l6VTC9ndMJMT+4aAMsu+eHSbOaDfZJ
PqabUOIiwXqz5uai9jZdVi5hXt48EEBPL75KVyJHd7o9sRyaAPXYw54xa4Ws9r02
pSo8fUBbTYKyNU6C83dmTe8+gtm9xMGIFQX9A8paog9aXpZwZRbpqCK6ekYQVCiL
i5+tukBHSzhz51k6gMUugU483ugshkTt8HvaS0m35IxreUm/N0wGm6al2VCfYwrP
nakVjqRFt4vy1BUodkyrTPuEhNNTX3jmiGSrSpXx961bYo/0/9htEbBdsuhzqfT6
lHF4oGpykewgGu8pjNBk9JbRPjo1h7qWv9ZF598croknBhy22NG1NqNnKTYMWPdK
dYXHD3mLhX6JRfQ/76TUFl+juJ9zS36Pw3zFGxt+md2Grty2HsBAesJtOjzouiMv
Or4PLAkRdxD5L0eWEQR4mdmDuKQigJX0opY7LBpkEtdC20sLM9e3vV/EEBtuRWTr
Ef9EQiTQLFbSqjri+ac/T+GALuC0OxKPdQ+KHWvoSndrax8pbgXTtPj3QHXPtD/G
bUIk+9XL0rOPEAyUh++1DFzYTBeE2aAvtSFDhnXQAoQDLu1cL4gfvHZu4SyhY5FE
ND2oXcwzCUFwrnG6rsc2kQ7FcRJAuCtMEXOj9f/T7g5O0feceS4iROKecr/mj/Ru
1JHy42ycgY+SCcahtVEOO315jpv/6VASl9C1J5dNho9mP+SMMSxdIAKA7H5DcAeb
DEO1E6YDWykwQ9lZZi2dphyDmzJSwCqdXIa6m2PmtyZ5ldrOd6MMjT5MEkI54LIp
G/n2OyotJPTVmsGwppm0cXWzFE8mtRaT7YRr9iuw2xOVHGN+eLVanQsPoDC9EN/o
siYHOv5HXLkQjO8Zm3lKZJlbZ2TG9mnwXEMzGieYgAKKkodV0AnmATMfJyZ++psv
rgrCfTzehlwesicCkgCZHEmxHWDKSCF0f0HIqI3lpDJwRffF7+oJpdLktinaVfZW
ghae15VzW7kIdWLgOq2hlZ4mQtQU9FgymA8mPVbo3pohrtQiLCXl4jrAJ69a6mcR
qbyGP3Le7LVf22flj6lQ9+OSOCj5bwHN3ZYFP7pm3f9dRzhEf1AALplRv7srbiCN
z3ewncYbwYFBdbuuYceAago7Ebb5sFkHIw/5guiWhkE0SWz58biT/74wOs7WG5TA
URC3rdibmb1upFFin20hZO9CO3U4NN1WhyCxecxFjd6UHEstO2TK7gjqboKULu6R
t/57fZXK117oEpossdx56ZqxOlMyWYZsJTiZO9dJc8fpkfJbpD17MPAVjJdbGBGz
LIvxFvukzkr5VJ8egHwto/nMg55pSatahK0xAC2VAtHaDDt9ZrUPp3/9ZdvNZr3j
Kg1gBst50WZ2FClRjTXju/kAdx9OOBb1UIQ4S4JD5effnT/SLNdKaq0/13LN1yR3
rSldhuO3wCz1E+X60grqXBo/m3CSE0iidixvOMLTe3LeHZ1Duh76Dxx9e0yHKpOZ
crkl8MN66qY1FbcWFkODZSDR1k29zXuBEdmUvBEyR9OFE85T/TymGfM3/Ku3EGpx
FVLzL0Lya+IV0Akc45LJZjjYYmlSpn0v+5yyy9oJ/Qgyv3BUpwndgnbuDPuMwcDt
EFrRIUXWqP15f/v1vm+dq6VdEAazls3SIEPVFY7DZaQD5fALXQRZisPdBqPCYEMz
lrhiyuwgetraqvI+APIq2TcrQdD4tDbKyvlKOk4eI846r67ny1kPna1eWKHtQtVR
IQ0uO8v84p3yREXxU5LQ3TJosgXy55cw44VUKlMXj5JVrJsLYNyUDGYJtnKWwi+D
4cfag778ACRUOu2syP+5RbsP5lUXKWmzOtnvoJz2lcA5n/iedZ8RaAilZMP/bhMk
gOwYCYDHwtDiZ6pQ469KJA6qwJeJ9Dh/U3WM39G3SqKupAMasmBxVTXyUUSf6BRM
BRh3DT9phqiCSbyRlySfAKSiazWmgvjAiWExoxRJ+JNLYDjmnfCId7a6uNvH+zHm
4lZZNaNpzaAFmcGQDHjJOKAzXL/XllU2AEPXM10PsZhjrJaKYDoJQSTtXLEYUgG4
EKvmZHbdyNUTbAVzXJIwwKPk5lrUFJ4uL4Y/S4OQUweevaRAWlD6Gr8SbNnggjI0
gevDC5tI0j0YC/Fb0pkWc8XIs350tLN1sQIeP4mp+GhzwRNOTKlRwRshbXREMe1Y
THLtKeYL/eWd+HVs59SzNZZzU4Iw02aJmuaCRiB/doaD0MsmlAFumefo1bU+3ziK
iYCqA62jbbasnYCoUlZFFMRFcOw+AmZelJ2NGeXuNd6u3GqsyzRL28ArAO8WATCp
Irax8fHFvNeOhb+NgHLmQqQARzcktVI0PB/5NCTJ3dhn4sLQH8jW3vRDXfGOynRJ
tP0wRbIs4bq/rVu5McZV8eYeCfELgT0iOxLHMLe3jaf0E6uhEt1FlNr4T1VAdBv3
FeM90Wxt3u8pIScGzGwjXAU8TIDUPQiruDwBknownplMNDM8gdedLZUQatNFUWCD
0bm+RPT0ix3UaE2QV59gBiYDQ8ECbK8dmU5P4qqTkhI+xpWVJ9DbTkI5ZbvmZM0S
UK1/j7Q1x7wqGbwAHJhZ8q2PfRqyAaJwpxdja2lJgPizLdDNmcEjcGpdg27CfFSU
P5iCKWwp4vufogpDyGdtOeqTWbpaCc3zEsepc7dyxNYvMCdtrH5cUybMIvZykR34
XVhme/g0JJ7l+v1nA17CouujYB+psfozCqcvDnz1Thf7xW7+1NF3mZ05n2vmxlV+
jnzBS+4TBulPysBcJJW6I4yBAOQvvs5jJbErY/uaZdKe6M9bUJpjlEVGGaNji9G2
4mLXzpwd8qurWTMKq4d8q/e0j6SgiVVnxf/1/6K096q/yRlUGaXNXp78puBNfeqT
Gu86F9jXUQ/YjaKkzqifiMiWlafdD2TvOVZ1T9Gu/+D8oS83CpRjuoY7mvx0shIQ
Ww03tcN54ZQXQNUoskB67BJOpIh+OHAwa9iAnurKVDZOPaaq9F4VcZ2e1tsVPxrP
shylnU6VOiuM2a8dXeZEvhKYxLJYrh386i8KlbTZPICiiBKNVp/IH/DPHRfiscXR
c1XOSFCyV9VvOGrx9XmT2C4cz4hZfJtQKL7YDPIEcnwWAALgMYsQ5vOb/SfVCA3X
V5dTZOCaWqP/H6MT4JXQRXy0qlHqT5pGnl1SRMvExyB7D3hgI7B2McQzy5q81cAl
0Ts6xigKTJwPQfe5jNoc6NrLJHH+vuMasRA2TOjQlaB87SZsdJ3HAEQFff4n+weO
L2HUY7qs6jA83n+T1Py35vURUkf18bwXQaA4TA/fdwahx4Bn3m6+3o/BhT6ErZJs
Y7Znp6hbQJU/Oab7EJsK6CzGKi/rFi5MC1ZP9Foe8jgIT09dzf6OstyD+wmZ8AuV
IgVZATO6B4vVweEpkE1+GeJI9ZEQ3mWkDARrCbyvgO3tdhHKECJSf6kmdGTqnYKL
gVj1gGtCKgLBpVRhhVlrdCE8fsyjj3i/CVpb6a3LeBeKd/2brX0zdABg4S3FTw1Z
sIiajqHRnh0yShyR0Muo+KhmjZn4y04AeKKgT0Id2YBBtDC+ICbUJ4zjtVMaMUaE
BL2WTFXVWUARP+/6Lm7QeKQOMHT4O6bGQUpn/tSRiZyx+kjh6BsbqofV6X5sQr1F
tpqgVDPc5sRALs2zbBUlKDYQtt3u/VOMQPoecVCJmzjM1dt1LOxfqXXuIhwWyGrr
hEyFTObU7WXBydTpeBvJCiLm6d6dY6oqs36l4zQL0d5CALB4GOVIQS2mzIpG/pX+
rk5ryyFrwBEAMuA0n+gsdVVkMCeuc5aimTdNDYAA9fUWpdBF1YRoXGzafv6qAc2P
KkCtkzhCe7zstbzH39vVmnlqkAeEnn89jvoxrGzMq4gYrzqQNSITBfxbEytT599P
yfJuUZRsp5wc5tYxir3L3dzh29BP7n6XolB1wpwCsX1yXfymwY6/a+CFORViOJzj
7vEXiTd9P/lBvf33YdbYnN/2UKUG4LLRB8GPmlSU1ff029cdET4ZGahUOT/Ni9jp
ghcAJWClSakbch3oLaDEp1QCnz/SldAAbYA6OFJK5KXVDEoeL0YlEGfzdhZH14ck
KrQqB6FPI5LCHI+kTqwkfWuvv+oIPCuywik4ew2CNlPIuSdyphEhaZm6O8UkEShl
7306h2b8zK8kFO9aoLQ38mPMlb0HY7SlGduacVbGZbOAUGiq5/MpX2tTsR9ISoho
fqtOdwjF4Vd/JFb1eIZSi5vNgkmAZPcvK8pU3Gdni2YPHVdVA2eaks9DC8TikP10
Ig2x8BX3w0jEK8ZGXcinqiz21h6K8TP5wq9JaJeClxqq1Sb3nr/IAru096219s7O
M6WOu7bN+tW1M99mcWkiKNGNtuJfZ3GVYfLOE4hJqzA6H0rCxivmofnlCaUD8Uly
MWMTaAW9BAcKicxdPn1ExtMWeV2RgpRu4xhl+yPfZJH7zfCBT5csgIXnsoc9YJ78
+HZIb0VUdNhHaLPwba+ctGhJFGWFv7x5FKibH/Lv7o9D/oAuUtUMtuCIoOlA7JFy
+FSdaxcta9XZv1kKxl+C4B/Q8LsukM/brbaGRUGWjE39GXGiSQ8hlvEUtn14zy9j
Emxc41mOfK4Yzwy+WZyYf5QstHtVVktyCNYacg+ybIa6lN62DakkFrBFnY8a00OP
jNYRDT2Q7Pf+AVvpzsFvKQal0kgkEQSNHX2jaMISPxZO+v+uSvo16Wk3/2+qlKBO
Twy5nrvClDOQgpPryGRBDVatyVN5P2es18S2tt7PmqkwCuXnn/TzmNBHZ4gFUZPu
SAkTLkj9AFPzc5PpznZ+0dg13FdAdal7BxJj6lwXGnYCjw7LU5apMBNOSrafYt+D
ywHw7aEMajCpPsa3F2ogD9SyiaUXIE9XLeddAChojjdLLa8Veug84a485NX0WnuZ
8tbxtUcXyXmLbQuFSgkWgWWzIes3H1i/y9cxmXoKrbqpnrdCdBpzPIRdojStC9rz
pzqDaVi/E1AgwSuhFJJFC4pNGja0ZGuw5dG5NzQqUZAAEetS/TC0FcpuSKMGo4PX
RfpyHqxxnYy3ePYLQ9n4n9LDLjSASjyLJc7I0eCBuSL+MRFub+FreAwv44ibvlO6
6CrdcRDB54NN2I76oKgaaoQzWDcAKv5U2M9+RI7TdDdhpT7QISnZLvbYQnt7qBiZ
v7imrJa4Nn/kDh3mlRkRK1OGWFohO0/ABQuLY+ckxWZCDiN4HTtXT62n64iEi+9J
Pe4dOY1fEbVdKubZFydn1pc5yD+azVtsT0tF8bsf/nxtw0VYK+5btL8WpMK/Yoqj
8KT1djPSo/8YNR8ySVKchmM63TtGjgBPXmFTC6auZZvfHILCjfjVJ3MB9kI/uS3P
V79zSN6ROm4JVnK8NMvxIuinjAxf8EJq92PUO9CWgSXLmY3CRrZ+wCB9a/uk4A3c
xjYTWbFA8y/LFHufHQJ7wGSazFQKLb8khwBJlyOWOxF6Fjdm/ZH/StC/mmfFQwPL
5wiyAk8K6wXohRKHW1jaURM4+SBydr2dw2bJFkXBhR8u3yjJVvxl1A3uukfdQTBx
bNSn4t/gYItDUXkWDlGEjB6G8vBYzesfHsQZxRw6YqHauRnDNPNiiHSi6lSzVVT4
p8gsoCSgfTT319eIl+jgwKXInPRo9HpoopLguelRcvKHVyebW8Svp3bDhyzD8yIB
tmL16uD3yH1xN6DjcPOaN0ddCFkacBjdns9U1i3cOpbVLYbwQWusqVKD8VSemwZU
S0+M0fgiopbAw3JmoBo25ZJYXm6lyvjdcmPqYha/Xlk/fGwtI5EXbPkFYynn0WWV
RSrVspS2EHvtjXhuj6QfWr905q1kIhmJk8yhQRflf2UpUWN150Ak3XXy2CQD29LW
PyazMMTbcas0K04PsO3JNxyXnOysgFULhVNcumXxek9Ol8iS2s/zsNlU3qCc/DeA
6akpnVtAgxZe6U78iHcYY2oEq/mq2J7nZCt7QG7u8VR8EUS+T0xnlBHnecPlyqXC
LPqIRkufO/sG1oerYD1ZxS1o6Yxd6Y+6BFyectYgwmeSpAd11+u+KkIExtXJv8EK
mVppLky8+jlThu/yxTkgMIudCXEBHW7Da6sEAhfO5gKswGD3KK4wEstYUynNejZX
l1YC6pkiMvG3dTcOGeGjqnV31jl30IUppC1MB/Xfa8XweKggkCv12gu6mm2SFNmV
Qtrb0w3Fv2WURgw2UK2yN07PqNGAOE+Wu1iDHjcOa9VrH7WIvR9RJZXE/0kV1N7Q
wYED9nJkR1/S9wTMFzYBuZWkjCN2cJM04FAHHhIdKHm22lrYUc+eT2AVZ5q/8RIy
T4UvxNKbQOEO+7+aPhzJKUlFJmafHFE8R2bbYJL8VNQzkK0ldnv2DwuhdsUmiAyU
ILEgTmARsguQVF5cOCwb5j0nLBOriernkxJeXV09D11KyeOnU3vZzga78E7RV2oc
yQFdOOGR5OtOnfshPENXpvdEaRc8CPuiyIVL9EOP1RyXQDjmiiu0tpfJpN2aY83M
Qmktc49MDRcYitOo5VCfZJulLLohURMLZhCh6IKCeDlSZqAULo3gVKQ9zatKYfPX
B0RgNrls2e8DfELJWlaO6tQAAjzciitSn9EARU8ppeQnnDIhyY3JMH9N5691/g76
1dN5cKChw2/gvAtzPhdETNXfafRoIAnh47tfmJ5hoggYGs8JVUlLuIs9SpznSdg8
8oVxFJTxdZPe/226g49Tj4zWrfb7BRBkDkDU5YFhjiReqjyq4kK0XZ+WgNKEr1YB
jXpbYdsxFFAyHJAlPkIDhOKdebL+u68Y2iHDaBqaKqWFownyXAZ9JeJ0HiM3X22M
Wak+xrF82xyI2eW9iyXsOyrd6wd+yT78sQK5Un7KoHNmldmoiw6JzRlUhdHkXq+F
fkv5AG/SyXK8DAXWUblmvjdoaPierSJlq1EbCItjF7u0AmL44WRTDIgMCyAacgp9
eW8wy31M71ky7YRSqg71IE16onuFWXd/B7ORein17rDQcd2wIS3sCw6NjAIUJq6I
CnjX1DGFEY+k8jkhHn96Li5yZJ2eLldPkPWjMG6oMx6OH0FXR0H1SPB5TGY3/+H7
ho7vxqezlQy1L66yE0rrctjcqoMPNVHs3Yevlrrg1Hy3qoDs3hCf5y0jj54/EuvD
E4FLRk1vw4dyCzZ0/1KlJxDmCRSe6gzJe3SxjgNVp+j5OOwzradtYW0KVBFWtEQL
3Zy8uYMow9Ndi3EyXxF4gMwNsD1DXfLOG9TjmvTnB/UCIVy3ZiTXH2Jwu5Q2/IBy
hn7Vy6TV5x0q+3JKqo4ci71j6pNwa+s0IExACGeIgDBUEy/eAiwEKrO3CyXcGVf6
LZGyMRVKynIpWJJ7TkgnPreM3lvLoqfplHQ9uSpoNld5XsaNa5rLYkVtz0nRaUHu
w0YB72lwXksRYUq168qJPAs/V9b0wamt4u9PAKYKjdEkce2LHMQ/2z/9o0tV7aAU
em+zACMqJJXFuKHszm1W3kZi3VsFMSf9+LJ2rz1duPHhKugtyvBpElBERaAtjfy1
du1B6hkPWB9dcgyjTGu9NkRJQK5kgppV00b7aRuYLawTJrDh9VeNK5jddDHnrjSh
ivnxDPJsLkt2LHWA9Iun9N/UdtoaD0mCdLhaddCb74bqW2BC1MskbU56wynD9CFi
L8fpEHpCjvZmfAyhTEHenjMOPld4m6M9SeFYsPzbkrpaC8nTWEKDYZchxXPkUuXL
0cko7apVS4op2crDTt1KaOptAUGKNBD+nQfgn8JC9gNN9dbbEFVET930UaN4hFd2
rVbN0K/bXiZhIQSKV1Z7AVpWWu4OEYuVo17rngfW4/lMaT7hUiNpVsIqcJRxKn88
yuw1MQkIXmbFRphW3CiWYL3NnZmqI4kQyfH36wT+0f6KIlBA5PVcl6fAo70TSoMV
T+NyxNALZi+4yPVF3jPXV32M1a+b8W/3S4ud2IogmLFuzS76Qz4UUKCWA9iPjNt9
DnsmbyjZccatd1KJ9gXA0GMzV72QZWEEitPvndy8djPizyMY3mi3uU77+ioEiVmS
bT+jp+DSIED+ZthYSTS7l45tG3DaqLb1VfNTImBs5ViNyT1MO58KLwTYeIvfuJDj
aNaeq/MGmKG51gh6HmzL2lRjYVvyAWZ5Dyflq7NkLhakKRxTm3Ut2Y25Jrc0zK2I
L7mZwCpL4ZK5C9G1yPy6XFpUMajAaPi/p4x0u4pk7tmO2M5AuRsn/hJqxyUuvOGz
D31MsO5oBKC0dC9QN/IcXmQ19Yw+/raYOYtXFgBezSdx9M4tZ4ZWi59fhYBHd3m0
sc8TiYpqYoFDmZxbaE9tuExuzZwmHg5yd0rM4/ilZ0iQnKhEpOf8DIGn6oX2mhpH
3YF5yrX/3/FYI2ZGCiMDDXxRu2hIDACkHYRE50T1k6YQZXWkUAHreHYepwhOb+Ts
20R6l6YsSInKsib+TVBL5Sgkyg14bxssKm0Tla27eIvc+LywOGjDjTgJCpQEueh7
g7AOYhFuEMeZh8IFHQVVXZQAobnMsXC0GT2VO5x9HhYccLlfF9q0rgxpfhl1A7Mw
3q53huko6G5aFIzljZXHCd+++81Wx92ZiFj+qrITb1gewTZMDzBJvyDbKQLdJqw6
VSwdxTnYIHb3FceUaXf+3e6bNWx9/ihoFo2oQMjUY5AKWw2d37DRJ0t75ymDMQ5d
O0e70SIj4ITqF+zRTW2vHN9ajqAS4Qi2SD08m+JsSBJkQ1NQe5W7VPVFqUahJQpN
qTbM8c3iJi4Vh5GNv9IslsD88RQOqGfYdMZn+FFqfhsUpeGWJ4IotMRG2bg+3ZNF
dTSZ3zb6SKyK7kdxyOvaWrwxRljihfUfgyS8500ZpnyCZlfFSac3QGzKkm0JT3cf
ggw6Io6QKAUpd80o+CzlmDf0kP05LdbuH0KQ+hkVXqh6gCz71SKSLT8abbRHYJfk
zIJlTYUD+60AV8mDZmwoirOMdpJdXwkY33XxWttjY2wNmlm19Z83zqidC8vgeT5t
0U7Xu3G4zpyw5+J1VGrGE5ihO3aLLgzhcwICcCAAhkj3uX5R/UfVF1oq2j9mo9/G
u+LHD6l4as9PCEG7rK/oUQjziwDWWmO20pbN3m3b2kDWm3V6JXK4TzuaxNPyIzBE
H0leXlIz6wZWm85n6HC5KpJA/ntujpFxFD10QvVk3YSjDA/ZOdiO7kQznqjH/mX1
WvONCY7rXxr3yERvIf6a+LvsDqy1lOMxLsYMF7+i7TznNBAin42wr2JJ4V4v8wOM
Gow8HjIZ0OAU+P48O8muMKZ9yhmuToJ7IgzNh5RynXVL1GWSDIimXudebS6Am48/
7PNy2R4H8ZM7OAvW2lJ8DPnnCb3sDkgdfQZ3bo4vIefhabqQq4bmu6ks9bwk/KRI
99vOQ7/y+AARx51ZgSCviKfkors3vv69NKpTm8xN4Zi7uR9REam02DZsyitZ4ocv
zo7vHUuim3nWZtAT4gVCTXJgPeGnt01Q1o1zN7vRbiQZqqLyvNeyoIrvlROXh8mb
FbG3LfPlInWwcoSVJOlxpi/5e0P4x+yRiXAKF2a1DaS9xYlkWwzvyl61hsfspb74
XtL/z8+U0+Vp6ivy1+xLF43DGZAnUcmgnr7WiZ5Jlj+x4hGK993X//jlbcA6LmPw
5rslDvEDSifN5udrM2XgDKwHuKT/MX3HdL3KQg7wDtU3aWCkiGUe97Q9qHfcqBXB
4082XYtyDNSpangAbNu+ah3LhFCjExUbDea+GOUe9z5K9/vGFpf3VgNohPaIAz+3
yo0GTYe/YRh1/ajUQ+iHDufxn7gwWfSWsRQbTXinfI1jQGsBe/I0rjjC5KNumK+p
I9xujIY8qgDdnzLp6vpXQuM5BqLGe6dyg7aGFbs9HdL+PWnqTjS9ZrOt3VVQ9etv
YirUIdNwOSOV7fQHV/Kr/FvSNPg+vEOf/0rU+DyzdRwvVl2+C3mWKQWSqSru6D7l
E+emKRUK/r/Z3lfrtYA/JM45tPrMmjEF/6r6ikajKphp7dNKqUGgmMpi2kPS2cMx
uSg9K6/vanjEubjUJjZAKP1ss9zAjTlGUcmR5DoBQHqdZQ2iIFJcuEpFLSwzt8U0
/tjOYHwS/0KZwdnD/gg5M4sZBgPXD9APa1k8EsrTdTcnirU8uG0CPn1h1820oCPB
MWh+u9UOULifxqT5Cuwh2f2Xn3UBCAlHO592dYn0lVoOjJUz6HlSfFyTmbYGyurP
/T3/GAuURRvDTIA86bbN4uaid7Fj40JuynPahdZCciAmppRoOn2qv2U4gPpkI/5U
p94+DH95KbYnEy2NA4SOHDdAApNHIvzb0ZeKf3EcgsACpjRMtkKdI0QK0N64QU16
gEsx81PRGuTrAGJJ4kupuyS7mvODDocgLGjbF8cLfKJRchjV5XNJC0TuDD4x1Zsn
NIYq+lU976a9W6iCwX81BjsmP6JPz2yEyNB6b3A3rrGN7CPRIVVR2+SVhytq79Ox
yos2+iAqIJBmer058xrG4aOTVHxJHg+GcJO9oVv9vRr8t2qr/9/AOZ5f6ZKATUAX
2mkkyYUMZysAS3kSdlkny/7qpXLKYB1BDUJyivGX/paf0QXA7JXAiQAAyf9CesAU
/Xkmpc9UUrXe6ethww47wgjp8DNvIu6G+77h0zGL1dyeSHwst4FzGo/X56zsv6lp
b43Z99vpGwC+SdEuRXUCnl9PpTZHmhBvHyZ4DIjQwpsV7QO7cpB4bbkxA2qiwjoR
V5J1nviBamreRj6IcMHPW/oIl5LDc8wuJwIqTLrrSFKMHHm45fciU/IRhLS/asO3
I+qufR0dueneeQzqZOxv+cP7FXyVhNY00IeZlmMi0b9mSIgIgk+WnAMXinEjbptM
qieSXsEHNu9NI6drY+uKXzsPp23Ilmf/g7S0tlQ8/q80vCUGIfUI6r/ygQ9b9fM8
I+CX7Gfm41+cIJrxf2w8gxPcKQCNT9v/wrH4w+dVnYl9JyhmAZ3aVuO2Mbwfh4Od
GMMjbAqBrlfKdX0xOELYlvJ5KhpfRbaRTIbhWOVf+TNacIWz6gE/yT2CoquO4Qpw
MvSHIwKD6oH9lx4/bJjwTjXagIKRiRvxbZHWd/4ZDM/4NEMTLlpxTxKDczgW0F67
QTDNYlvPUgO+YzQfYeAgls5Onk0dZJPPahJPJlLU8M52zaUIS/jQHHRqdmVl53N/
QaxYL1Qs9Mkp54I6l8NctlPgWndDGkm/TQ9i/lZZqJIqDjtEmmpy+1BLPPt1q1ff
oBm32bj/kBL4XRhA0SIfb8gnC+rzXbrpgxvf3sr4hypSPkLuai0Y6AkWotayOwje
VNhnEC/LpBTn+R2YTXz4NFJoS6wTiBM7WM5D9RY7Et5ZrSQ/q6wzltSnPBx8qpVU
9NDttxngx1jZynB+wkINxr2Pfod2Ypib/SCSHeIl5/VyYPyyoidrpyUGsilITWzh
sXyffj2d9xNMS0Z4PQCAhj2WcJr36WZanJJvUC1kgKBcxSMpjWAFDLknMKBsPj2Y
OYsnVBquIArCZdkg1KCnal0aBJclOtdarYyP1pyKwgGXVqzzpsrBiMGW59isFa+J
pUh+Z4ae6NoblTmQHiIvBajUz5zqTqpMzIFiuai6qZa34G3B5lYMnnzKZdhgslit
D1nPjLiyyfDXoD36naT+W7JaqH/IRmRff12SvoMq6UGaJg0yaegStDFvRvb8AFwa
76S+rsJSkPxOc7xRdjdrQGM2sStyi0+pp921rSZ1a0cCMxuHXoho4AHxkLtvzKOd
fPco58BWKqdoWBBePQSsRaPw48yriT7Pu6fJFxveDHpxJdCrpxI4jgcPMA0tBG95
BpNvso9AXZGYsvcnDTpIk4uS8d/u35fWR5zdVwMnElO2N4aONdpOzhWlU0kNNIU+
hi1clpZfTpmoQD8XxNLNSi2suoANNq6TLryiHJ/nAwGUk+nCKugrZd8DlPiANY+X
QvtjkTA3b9yI0pW3OG2C8622+3qfUv8V2C8LqcLNDcPrmextjTaYgOqoblmf97i4
oJ8NbQcflzJL47ZpQ1+PHO21Sq11u9Q02+NLkDlXFsh5NjDDevFHk87j5Cho9rj7
3Zi/IQK1rsbBmudTSmwf6tCUHCXKb9WTLiznYNGBa3jRaalTqhVLFkz30ImzO6IF
U9x1GXFz4NSVZaTN2icaTi3rhn5Y+GapIvZ4xD+4BYHFUf0Lgf5Wl1y3VQY9vLsC
kjxEOkr/Bt4l4ysotvJqZq4jtpQOKY5vpQ7aaaPc0ZoSVcamXcQ2XU7pqo2FkBQR
KYGPrf/c69LDg7SxtS9oO4W1cFL4TChCHyotLdnKBTDcw8SBCQk+ne8YTgbAPJLn
BNyVc7x2DGcj8XBJwY9tWYNGuyif8xqvG4k4TMSf/+4zrjLlhKdw7p/lOPyNCuG5
NbmhWdAI92bg9iIo5+J0RIUfVD570CBUNUHIUqxoKCPnjEZvnuH6L4cH7LcPXLcv
B9feehQ+QQ/Sg3kAlVk0oVO9uahLW2+2MED6Tr0Znt/1O6MDHdFevX8DsWT3SgQF
6uFcPOcdMeumI5eNnW4Zw4pZzOsExTwqOWm8s8UUu/Q5S2ohqXe7E7FG3aTQS6zG
L3Tn7eL4wR5DdXnpcXLLLos/9X+TEG0+3qJLrntvrT7POe8mbyPXNVOcxEAzrMyM
Dlg/IfGEpgn/N26Q+W18NfuqlY/Gr0BBMWhGhcT9jOj/wkrDuCVh55KukpqdbEA/
Iu5NimHNyPc0PWk2B2DLhgDpcUSJqhzCyPDyigcTJdKnsQ45R3/7HsbOLQ1172dg
GDp8vl0+lO46ZLQpZQoYJJ7zIHSAmwLdElk9QvGqdRrwKj1rWu0vafq4HCsoaQ4+
iOWBNJcVIT8Kiox8gbIS8jhpBOIEQ9MjulmZDFV/f8pShUQRN2p9JWH5/7Wrznnp
W2qidriMSj8+H/0Rz+WVrG7cYd1E+084A6s37m1l3nfrtt/SsiY8I5RVp1MWwMmZ
fJqxA7gCXPHPhP/j9X8vb7l0NazDmeXlo+Z4QtOzBlNhsuF2SpSd3hCaf9kVG8I/
HZsDeWQ+Yxe8B/oOLvkzAUNbj43hMVHi5zAkFPK5eCRmoIzbf1yDEmzEFUnA3n4p
MEA6O/xWuiSaOzKDgQkk06ob+nRQgXtcfgSO7ismBEdO/T0uuTNrbmtLDgUC1fpe
CrITt4Gxd9iDAiVPAE/lOFcffI27ywUiyOIIJRGN6MLgeV13jtWokLfXsg2/6pAm
7+lgIm5BcvKNzTn+qb6igojkGnwsq+D1DaqwrkZh8LilQa5mByLauu0rpC/6PjBn
ioDFusbBKqlbga4yVnWwdahsvbDbPVFQHOVsx0oB7HjfeYjev/Y0SQiJdYoSq3C3
EksXR/QtZESOd6p0XhC96gBpPdOyT5rKQXLXG6j5UxAyuoFEwFC9Hcgp8lYDJa8c
3e2dsP1/J+0ovAyeG/hTU6idiZBVCCLdayXz6CRQBEISqQxMJaZ/WiU5AutzttNY
baFumsce6+MGAim1NVURadTiU/XegOw80EXMNM8yPKwFuwkqSOrXfHjjLIsNPEhk
TSwcrhtmbKx1+Smn2HGSz9tkT7TJ3WIHnFQyafIenf9tQS3ayFvs3gTnHzkKeShy
TM1Kd0FpY/WjquwMKLeC+7CjXv1tUo0NQcv5mHCA5+iVgIGcnQJ7L0hSm0x2lYUA
BbNvA5YVLnKN7fC/p86KISXu9xBhKtenqphN92LUBAPodciTESaErFQKt5N/UgVK
xNpEqULnJaLTcDewrTPI0XHTnWZLndZxDgCrQfBLUyB1UIQNzyJChIcfZA+oDdkw
QkJEwOgQMoIwI1xEChavQzmAxQGRrYBInbeliZpMUA7GmEpDzp5bYhkPY4thWAJU
m7Pf21OWnAAUMkmUjfTqQ8M7q189WfX8zXjhyRWXg73tdCtsYD4gwvTKaUA/eutC
8NWK1rZggBZftAyEYIopbgCXDD/wugCo84TDNWihSkkmnFzMnot6siQrUNvwsSKM
WEuTibg5uyYCA/fpV7Il5LsMH32QQ8BKvjcB0ZBoKL3ELYshEwY7rZ431XsxKSZE
R7Hi90amifYZlS/vD4+O/U8Or44jL0rfTq6ugJspGzhwejjzSBl0ys2ZuVrR8P7I
e2/ydSmtvv/+JWaxY/7h+31FC/nxb/0//MMKuKijOzKAwYEfrWxT958VngAVQP6t
Obx+X8fiMSw3GHSqouW/xl65zkv2Z7qz1pdGQ8JrGUaPUl3fOF6A8nEr4BncD3Ff
lA4VzyVbgdN2ZF+eDzkqWKi4dyHlQmiL7xU++ICoad6XhQ3tZDYpD08UDlVM3df9
nlluQ/gCeKxOsfNEnj1dQwMVPHDcTODd4GipvGsDFb848pGDLw3dJpxx635IdUBR
Bbi/DdpoAyrfJL8D4P7sSJcttWYKZOl4JBZ8iZPK/AJRmB+0/JLY4k6308V6F5AU
LEf85bPxS/TMwLoE+bDEDMilBoWE770Hh26S3mh4D55y2QGLVELoLCfLnOIKTryp
rgc3kOW19U9nMOp1gPkfjAUMYPw9UWZFO4ljEY9W74ZJRsoQt3I4nJKG1ZzGA6QF
9fsBCZ6VC/HocPrYfkkt6tW5pbMM7pxH8uUD71U2M5b2qZLRWtLDaD31XHL3EJJF
GUS5iOLfdcPp9NS74nHfeO4AUjfvDAtcB5pIh5jEdy1SikgjlYrWyjP+5DoGHOYe
PQaAHBtIH1MsFZ9OpqubBgaOLur2BvDUfc7nFFBAIQA21VWBjsCRPNWpu/EGFoGt
6aGyYHQz/vI4OfjD60IxYKk6yWqJROGPkMd5gRptRVn/1Eb37sxeLctW87CCmsBz
YjsX8h7cAu+6LF3aGRXYYZS79nGv+mpiENyRwi3trxikCPjiJ9UktWop83RtmAsO
+tUkFgLnEwx7GOXFZJfwAhelSwmDk+kHxbv/95KRin7impiwdO3/5nkz0TH8oYjh
pO63mufPtz6MB9dz8mTT/HD/xc7DLFKvl5zW9YaB5XoxkvOrMobv1bxVHBuZEHYk
hz87TWUUy460K1S2DJmT5rEszIXEqQH1T3ueS6JXScw/3JdMJPDr9PYeG42JkSRv
ueg0NS4sSTiLX7b6Phb5wMvAj2sWeqKm35Ki7JmqYQGywTMT5apNAS57DHtToAI3
Gm//YAzLtEPtpB1mO8gelXwnZzQhdbLG38dkxvIYRjdk8FhNWSI5rDfvs18cuuTm
6M1o1BVlk4zf7qvUjV1d5/yetXrPWXxTAGRwlixwz+653ANet8xs4PtiYeQf77+6
bjyV8VfgSBgdKsBtYvhuK+7iK3w6kM245rTsAFKxmbunCMubha6BtIyGdUZaypoe
UHtr/AVljuTNBx2ObMJAps/QxrznTTrZUO9QKtm+tziVOrHuExUntu69Cydz87Qt
7dJt8mMzLaK2y4I0NrZcbT0/wMzHDMQYmeFoB+qk137irO68Hqg2x4S9d5O4AyZ1
lqWDdqWMgyKQiEbp+9aCl9VVNP5tQ0B1QoFmOU3J+oVNUpW3MEDjCq5In825t7re
3vWYFaz8JSyNUtuy+ve1kta35t+LhPLaogAD4dYkWe3vjMOHN3FBOIcPZa0SmSBN
i7KLSXPPzFrd2lfoNrAhGCgMH1irs3CoTdVB8gCh6gB1qAe8BL2tMfvTAKOSp3vF
XcP+g1LjUrEdOO1UAhod0bAdyhNfjSFNwzn+R7uwvl+DkfnjkKX1K4J59scFWuzZ
31vqQte8SHse1pIXIKY4XYjgDlrbOz8wB3AwmVrL9MatWcmRGyl5PQa5lRaKu5iZ
iBOlWxKR6F6YA380s9rSM2daDYYl2pqcAmwozDfQDAq3+gSzBbYVp0NDMpiUirdL
kCV5UhVuVFF/5WBAVKJB1lINAcjDfIohSB0ErOnjbf3wfOuvOX7QkZl1UFbzg4Xn
x5MlBxMtIgdVgXcPMKNCK6S0eJKT6k7ShPj1pFh+c1hRkkmGlbR3YJYS7MoMHMe0
7T7B7+KrNK4QQBhKjGNUvy5Y7rfnUSOANzgFP3hm2TaIO44ib6XPN2ok+n/5+gBM
QlPW/TDwqOuuoEP20FCA8V+LmP+DOGp9mloOr1GPTO6vIF/0kFY8zlFfooXjpOwE
7MuNT0Jpnsxda0qWGBcMCR4lxOyKLNwjzIni2FydhJxAFBQsgsoyqMqdDjH5MPOF
dGoMsuv6dOnLZc0D7VHmTBOHtGifWLd1wCgw8LTlwGi+UCW3Wgpfgd7axjqMMhpA
i+xCmi/v8Nb0/Gh1zG+ul67lpjZ93MRDTEP4NFDl9jccPcVB60VI17dmS83TLTIu
onZYOWZY0swTJz4aR3cOHNXLsrtOrNk98fUra6qrV8NZUDlcaC9Nj+MJ8iZ008qj
twN2Jnb5umxyRJy3govlUgFysyU5D7QqQEqauvmbk3XACQQhw7+Z4F4xsQofgRId
Qv6FsGfmOUvP3b9rBMS2VpighgWkY9BCLpcUGeTVYvfXsMp+FSBsMHbWScCo9+or
85Giqbfatn4QLrV0n0zwpo9D2xb8r2M+JfFnd6sYiYmbEDZYj5h4LnR5MO0TCU83
UF2NJ66rFLa1r93+fJWGDmDTmmOcLJ1FVHb0Y+BFbUpR938jxD2MfDgGOSc3y+DF
OQ9XPqXmRDj+b1YyyJ3xrTfyrPP505SBpdCwoVq6SgVu2iEA8xJCq4ujjPTRynW9
gpgcINDUDqqLZ582OFcD90Pw6U93Xo7He+nOL+gGKJGrSDjHw2bSKQ5+iA1Y31Gf
ERiu/gW5qZqzzbWIfLr6OBPPC6Gln47w0hiT/YpagASzCDahzlBUgUAiCZRuuOQ6
/3d7fyXmM9L3IYY2zOwyyZwpfl18uShDk3K3zdxHZktHRaw12etmR99el2h1vo2F
+25RBUG4N+geq391VJgcAlAnBkt/7dCwv8oe7hK96Y7UYJ/02y2HpKoOfdkUOU2X
s/4QFVm/Mbpaq4tIp9vD8lPyMqcatxYbPLhWaTfmIX+FwwoLQtovcbcWsBdXrmX2
70YKABHIOeOTSBfa+pZQLSxdWTl29DeFhOv0hGquQNWjZhdNtQfv5JwBZU+NCngR
XD1ZxgfWl5xWaFFX6xEP7LJHtTJb7g88hIwYDhKH2FGkV4KSq8wDuS5liOnf7Cx7
8fBW+yTE/C4x+Lu8v0SYi8DX4POYcIN9r4p3DH/s7NjatKQSaWs2Lyk6oWYxXlOk
3KK7aBYuYmp+7WXwwopa8tWmNWCKBFVpKYPhibPpTc+Lg8AQYVDJETsWw0Jb7ZOO
IPtd1n3g4XTI7kXZBWbnw7V9ap+7fE1HGs5GOfdGUn1eAkSGqA8LzsWy9lQMhE1g
o0MEpgk4/OErT9fGXVYUB+hGKnYLfLgL5nxwnb9hDjAkReVyqlg8ELTo4L8qKXAL
k5N0sh5l7m2l8yH35qFFmDPFjdKJm1GF5UeBdSw+Cpa2AVuJQevXSTFpygNfcNUd
TKlp+c7lL4SWJ5Q1MCcWps8mycEVDbxfsTMGGJkzErB7n2kqHIonAMsd5D9oe07r
pp3iRDuFYClR4/OQXzOSUHCvLghx6cWl21rOrY68xioRglR2rEdDSRmwsm/QRUqg
Cok4VLGydHby/IMuW+iKz4ZeURz+R/84gjR9+ndqrrYbYpR8ZA7exWhae331Annf
mDBb8vjQyUAyjfO5RQ2zBr0xvYbf7xuSu+PDPXHW3d5IN6ApXcv8qaKRA63MYMtl
UVcMzojqgkxAcNWGbPDAA8u2RpJxVzqf2MyvlaI6scykjP90djLwINGYaozftihe
3CQmq2qdaWJESDEXXk7UMU9HelUYEcxU+pFZl8VNy+Xt8bQNYJdWQ1LdC6gprqTx
zX5rOj+TKKTnw9zVEcGqkX2TT0zmdC+P4oQBXXcCMPQVWJlR7t+rKRoZnXgqP28N
32WWU/tGyEpqFfEf+Z7ZJX6/CZXH/gdmSVwiTqnZKIQ7y1DtPilFJF10iF5i/vyh
UOj6OhVBiNqyYv8TcXeDuO9rKT8lla6zSt+uBka8z2ITOBfH4dSYcTRxUtkAzOZB
dzlA+5E+xwj/VAbS6iM2ZTmPzEVeHJrDdCouw5il0aLqK+QJtFYDEblOQtlo54Ht
JwjCU7j4E+1IdZzP6Pc3aXzje3M+yLj5haYLbqIGNrlkVTJfsQqGL8zzBaRpNMJV
EMYCdThdLQbudzvpFS9quzeTu6hFs8jGE8JqffxpR4RFb+swZJ1eJ0Sfp3m+jtQC
MRlL34Nqkr6oAmDZsKPQQYtanSbRHKG1OqSobvgaWQK3MzDOLiYaABSCsQPg4WuI
MwgHk88IaSgkAt7KRJP+u7pjSb8B10kl6T/3UYeIfZdLtvG2RvU0nz5w3A4w9ouf
pDy9EqYZ2rCsTYW1vu+lrCvhhu7761ZsH+kWoc60AIR0ahpMIDGIgoZz7HgzBTw1
LeVs3ONaLBeOWxDCVjOlbk1RsRbr1MJTGHV+2JIV55aFv8rjolhyExds1YJJX8YM
Ju6x8Gk9lE3tSDXblO9lPSbTKg68megtv/ZQe9/2cVKoDfViOiEUkJ5t9kW9pnhE
HLFFbLV3rg4Fr5ajvVBTaTOy4DTo/8n7mZO6+5244h90Xsm/rVaZunph3r5zWoQN
x/j9UbMB7MnD9fi1DlSxdHWHqtRmNanqWDjKz3POQStJ5z6S9VBDAbdhOvK7tE3P
purxgilTpcBkU6LTi5f+bElXGYFjTrZ7s59w5SJHbROvtpKFwFkeljJUr4sDlGXT
nQQ+ffhQzqxZtiinXTAP1Ya6pjpakkA9bq9W3W5WSRcxtQF79DgmRJNXakKlBycM
C92YMbnUG2YPN7bveeDOox4gGR17I1iyhKn6NJvJ6REhLBmNDMCQs73IzdAHHTZV
2IvsftJdmjIKGtM6TtoJDjuPmH7dMkzCUGIue7jxEtwXaI/+nv+BWt4li2rfrYBc
H5zozz644R+T9ZggWhZhk8brOR0xL6JUd6tfGkZDAaef77t8NlgSBkNgnWCZgq2H
UFUk7vjtmnqtUiK0JONbMT1i17lWxGur7DZfvlXTNZtYuLd8sUbXkS7YKsExY0V+
wsepbPpIXVLZtYmgpNh+1zyAPcTVu450PjWkdRZI1nU/9/+67rz9nuYJ5zkNKqlR
Cn/eeGFrDDH85xJfHRsPaXJayTMTxS7Hc5jQ44RMzMuwwhHaRXNj8ZZjuJhDoiQP
Ftziqd4sTM2cqvJtAbuJ79Rwj2N4vkGf1AmMHOL/luWZNkyW3WkfRJaXO7wTajXo
l448WkLq2+yEwlFqryADYpC0fqH55NTrbBuFJIU8lDXHJvgSBYua1X9LxVfTKpms
X0flKZZ9SBx9eoR9uDXOYikxHEN3ajIELi3WUT/d6tBQG5y5HKAkw+ejQ7aPapSS
hT1xp5hlbLqQbmFzajpmGjaPgSO0kdjXp3rB3ZtIRPDxh7CaS/eHo7TK0MBjOhY+
405xvns2F2Yzca7DOGxoAhw1hdT0PSsWaS51swt550pKmtvpqh5BIJdehJl37RBb
Vpc0jYIX/vPK6Iq/iSpDsbpeoTKyepnC7spVWxen4S86SjOfxZMH99O4bj3/6uvU
9Y+/INNseMhuxbMpAGYa/a+0saVI+9E6lvAbUe0gFB/ooSepe+nXyUcLXNuJXQoB
kfr9XlmlU6Mka+7jSBk5vQVNP2X0xjSDLqNn0lsTM4H066hnguc2OIFQPAz/YQTa
CptAhJuM9dVn8zSmNCmljufJGClOax6KNm4n/DiLZn6ZGHJ3GHf15tE55Rr7JBY7
e/4YR2oDvVF8PJeoAuXsNNMYtPAjz1f4pa++USnHk0SdNrgiMq1WZlX2JdqRNYVt
9bCttVMf1E9wZuglSLisHkpHamYLtx7T9N/QHdHxopgSnI8r9URPw9OruWf10akO
Of97lAc5NWvXxDhycyqt3YzPNaj3EMogdO2oVn1cKffepYgIACoFXZHxXNscTH08
RQ9UtVdGp9eWKxRXFq3//boY9EGjd7i2cZFlIoosBKqjZb6aFgiXpVEDZLmTvA1e
rcarEw3tEJSMA2FU6ljONAo21XyMDC7eobMy/ClwkmG1yvCpZx7tzRX0Xsa4sB/q
8BdbndkVypRZihrjf3M7KeRnkTpsjYubq1bWnUBdfCv6IbACpYKfo4WB5QrKZy5h
ORwwxkGxFvQFbTb7tb9u7d7RK1TxhkUkU1jTxO0xB1pM1VWcbnHzUs8EoD5vQept
pLl/hQ0fbowjlw6V9UdbCDBDrCb9yedD8D23Im7Yq/5iPqw1ggumdp+HUxEzjBoU
Vk44udM0zbM9XUsiIm1rKf2dYin9Wz+EnF+9SwJgN+fPhE12Dl3VBafvKqkTbM0o
SkZ0nLFfU5xaO3lHLzvAJ4hcLCGKnEwB5n5iZbfOMWsE1cMdg1kTixnef9FD/Mnq
sG/GsZg9IwNl4qDW6tUg3iVGdRgxd2IlqXN8Pmk++EkkVDuU6i+qUjXXuMKv6glS
dDOA1w8sLSCxtn4gYjPVLE+vr5PQHfBd7cJGCW08P8dWWRh7bNiG4dq2QVDz98+1
Liiv3w/w/SDB66jm6bcjDcCogzugylHqkg4SK3qfhpmk+8q4bPiXvF0RVAAZONKN
dgCbJ188WzcuF9Ctslwd9bVAArw3MzxWF9u2kDMQiSFiLOOp0Ibo8961R8SzpOjL
SVN2EmvFFjWHV9x9R7QlAeWi/+PuJ4wlO4oOjWqAc24Cgk1AIm231yM+HMNh9tU8
+IcjXPJNq8Pu2uUaGrSvVuCSQa+dRR2et3C2xed1yFSMDCwzHAaQeW/4hN5TzEbW
7s8ev1sCHOmgx1+w1RiDytcCcy4dxWvsYEDt//Gt6lUhDJj3j914rSiKVLuCQ0kd
cVesVPF8fuf7GU08PZAKg+yRawOy91PFT6Ka9X1vHojs3uuBO0FuqpeYlfu6mE2e
ZoPY8z2RAt/zc95ebfVKXx3aJjE2u2yUVOz2pCQKCPdCcbEmYulXc83ZQ91S/7wM
WfhmvhudN9AlAmfefdJ3KTSyo07i78AfzTdMlbKxFijQW8kvw7UsYr9UG48AWWS/
IoAjEz9Eb5mXjGVLf0hTNLOYK/onjPtVaED39gzntFvYCgniIqD2/gVXmMAcTLWP
iPEW4OQcC9Gg41hUO/Z3fKJ0m/pLYfQ2eP+YOYYFS1r3RU5qHZCDh5sfpIaZY0nx
MXWtYAbSQmOhqGFUZOMstXU+zroHsmOjdkSn3zw8BZklMWGyoZEXWoAqohOdxzn5
LOAzHY6FpRyDF8/9E5VRJQJlyNADrImWHmGrlP5AhJvFkZNT6mwKInDAFORyKt9l
vmJ7JVEgpXhncOlJJ9Muadfmknzb4jqMScOWjpGs82QJWRfLQMnBJkaDGyhanU1R
PvKh8iafkQhx7OG4qLV3KQtNzS9pIfmSK0QaUPMxclKNJ+V5x0cuzxl/vmQJ/WLe
ZbX/CX1INwYzS3ziAD4km1Krct/rB1keke0mg15e1kSja7uMuSdZiQ8EJPFEeG96
RIKoN2Oz3cQtaeLI38eJrLsqkuNQc6zzpQItDDqzPnI2pIUvDMISVurNzciZIMRP
XIK8yqgIjU5qo3oaLj2fbbpdsr9d7QnXF0U0MrxseaR4RKFRd30Hf4lkZlI30cpy
0Xfrlgo684Pz30ePnUTEANxYb0vD96m7XWzr2VHupni+SSsWFUxIEu70SBK9tiEN
YyxePNWVi21jPGxLAY4onk0AwMdgXtu14l1WjGkKmdxVQmut+iRwUP61fYHZ1qOO
MwT8WrLfqKB0LAmgv738pbySWhVI8jGxBHE7/fm3VCqET9Z5eq2oXEfeTJS3IhIk
t6H3RIUxciulK5Up7CYXhGuJWxmrcDMOhpFaJf5KdR7fdukgblJMICTEr4DGniii
SYU5nh0DcQMf2jSqxAEFmJ6xWg+jOMSzdxUdrGXw+zz2fYey/Ys73tREhFu3uULN
lcAMz24FAIo3atkEAccKxY0Z1t4W9oEvcQ5SnFatxxzPRqq9VWdFRdcXYR2je3WK
808CgbUf4jrvcscuIuxq4UoWtTSExAwR2CvIPNC6wSBrXeXQvqun5cW/cxZ6o999
DNhs1yoB98LfyiYn18a11hTMvPyHkzC1qxPC3Y3ulgQZjGpEZ9IhGTd4gbB0N1xb
NxAcOMyspCNQfEkpEnOWr+Nji0GLXPo8RSV7bWVx8Z7wcMFYVwJc1f7I4+x6GvjT
vDSYI1bAykDFSRJYO0scJLf1N70IM4yJ6LMZ0r/Jd96c5rgCyUbuAEx6Nrqo5dAo
NcFV6ei//D79sJoaHAC6hh3YRIRBfg7JCz9BxVW4sWWfi5AE9ydKWGZwrJzZis2J
hlQFYCzB4lAZdBiHY1DZBSu1ozguD4BAFvL1orK2XJceYhjTDaBuxLwgiaUX6xdh
VnOX2ywD5GRe4pbvBYW3/OHc208sVaes7VMKrf2DheHXIsz6QQtq9pcqcsmY/h8N
LSHQGkHxMR9WkzWToMqC4jcqVDxgL4KcV9Pn+4AOO4Tb08XPgzOjRftCt5NvKMsI
pQQ4f8e1UpVsLxFdRSrEz1pty/3DsF7b7og7E92zzAAArC0o6rpdxPnNzopcwm9n
RgI/ctPBGjgaKFm8YOjXfis6yv8foN79/cuWJeau9ps470KRIgM7pSgy16uul+3Z
b/n8RnwVGpQnvH3ep+tsDAqEJtndqYT5eaotIwE2owxTMZ05wPJtK0eoPpApYbH7
a9eEpcsWJJ36oGlO8vsOpTjBFoOS9rlr1+TTom5Z5UH5nI8AmGLiL+ijvb9MhXBA
whIlezSqLQojRvFtVvJ7lY7nCi8+BveSqYV5FXlgtN/xKoKY4dNqQ+YsRphOwKn+
U6fXCZTHTyRrks3ZTSM0wFuraEAEV9i1czTeT9ZfaloxdLdujKFIhebUqft+N3rB
Qk/tlYIt8Yjk9cIG9itgYdUwKpxXqgTC1WxvVKIVkXQl0SvVCTg9ex6WL+g5PRPl
R3BkM6mBbwiPBF95KX6fLeaxWMPoVf7K82L4XvYbdBtH2Wwe6V3fBD+yy/uFoXg1
APYFGDNPRAU+PMRJXXgz18TiVPjjE2TP/Y/Dfjw9/6ApC91dIufKL1PQvxjNAYO7
Ie1AP5o16RLfW0fzNhMVOa8vR3HNUUJrehjG8gD0fEWJ9K1Lc7CKSF/axlmeR0Vy
VABTGj8WjkF0g3Wi6oExSTxmlsb/iAZ741IGFQcyY4Bs3yo/K1ykfcpb5K4YwQmP
qkcFFx3sqrpyX0RUeBwzhcEyNcDTkyfSoWYeHeiu5yh32OeEa9UzY8zSzDddR/5t
1x+NhhLqHmQAiSBSODe+pTBTFLybw9aqCHV3KRedGjb0+MxjjrlxO+R35DtCjQaC
DXOwH/EvXBuvrO1uoOnwtJoES2Cp+bq3bNo3+keU5gl8+hF9HOQUVZ0WNt6CgHZa
LD69gettefQA9H9cqRTiG96k0/yLH+Hz5I8W+iISQqamGRLQpawNBwopH2QjiU98
Eh7L3NODxbDO60uOELJDL4HxQZblYaHLWQgv6qbJniJ+V/Sm1Rpw0/KcefGbdPMC
NdMCJ/j+Mjn9XEvkU8MJoBnXgqo65h/Q1RRPxtsIHynaNPsvbjzWMjxol+XEIlhK
rGzzPXwN1EZIxcNZsZN6mncey1b6XYrujLWR6iyMgaMS5+ZSNn2tSVvX7uQomJLM
+xiMMCQKZlxH+JPDVwi8lXEA1jSdoE9hauzJfKbma1nJYn58z4Q+lWhoGSB759uq
2vH+u+VbFK+yoOPT0zHvRX1nVMciGE1SnUFCPfbCYFBrg8eRiPOZTnRcPrz4dR4M
W+3wrfwuvitjeLpUnvu2vKJmiz+IqXkuxM/2LTdpMwF2isW/gAmkwlvAIqQlBPIv
NYtiuWx2p0j8K32NxpyuPBrcVeLPLg9A7fmsJS8YM+ysfuUh2CehAsyz2Q83yJhb
rWKfQSS839u9INOYcBadX0ZPXUaYvk5+7VFDMX6R1os1ohHZucYyiXb8dOoOUqAO
+DhTyLs4IcEw9p2dsycz2ZJaPi/3s32YziqriulYraH+bPypnpW7MX+XqFhlJZhb
K9KLSwVfv8OL1ExWzE0ZAGPxlI5HXwOJqnQWVoAx3fZIicm2uKwlwsv4RmtXt2Xp
Fc6qmhTgppf3pMOU2GQwn/CH4W626lxug26oN+X62MUYuVERPv0WYVF5viEOpB7z
J9LdlCB+JLx2GlUDKhwRgCsBjmw9BQDbHnShtmDgPSRjyvJ5PVqr52c4KT2vBw7r
UgG13o3+1o4xBIlldSuCwXg9B22eaUyqultS9tl3+qOH7ylmG0fgef9esm/M783K
ZZBw6NfdBWDC19+6lWqBhSaQHeEubzF0tsauIeWQfdo1RkmUB2bcV1IW0BM9C5LT
QQik5LpdOr2WYre9yUeyqa5Bynmf8FqbqRd7vqZj3c6s49ddkAz7ZndU8BgM9tbr
mVwaylPS4NcsUgIxsgxd9VmLkxx2mvTXRSl+S2B1MISMCYLQFtDvwtlCd8gwxqUc
rZpYAqLfRSASCUs7/Tj2xY+eIKhXKFDHQGG5qsr4Vcr9hOEdhiPn+5EjRSmYvsgL
qA8RBW3ZrEE33YK/a/CnllUJK1NL2PE490wYO4X6uXhYT9DcAd7snEIFtE7yrI9Z
t6/BHo9OlwpLZBEIzae5cEmkPRNdtsvuzYemYTq+wjfCALHBIPoaiYH9lPJpxXr4
Wgo7yG3nrxR2en8oiAdxsvKfaRqBrFop1lHfYiUhRuQ+RoXQAJdTMbnjjl55+tbL
t4FeDUpQgd2COpWH2SzHjiGmCr3P38uzNQoP+qE2rSU3P172bHU9+qRVfOr+a9hA
AvZiOQUTfFUYETBN/eicjVGrJpKRKkPXirgSNvfaf3S6lPd1a5jXB149366VV14W
vcFY3iPLdG+aDJcQxaVgZAGci789BByr6exI8bctJ0xIV4Y02pU3eQ5dxq5RvNbb
rUKyB5pv5ThObBc+QhuWW7oOJ/0T7Y95hp80f54rWflq5eqfIW24UK3NDlFWanFZ
Taixljh+J3bv8oeiFB1kufyRE2vtVGP89EKp6oNRWzMxjtKGMXkJKPk8w3H4wrz7
9vcvB4qWdfqCy7lztiUBtrKsKEIKvHWSAphz+pXqifdFdBtIAMVR8A43sPRcEZ+m
mSgt6osqgbW04EIoO30CbraOTLY6i+T/tGaMjZ90J1mKI660255U+vpopIZ7JZ0v
uzvUsG24luBEXgPuVe0GuY4F91R4qGMOD1LqYlJPxlHu66+XMAmJQchTteUkx8qJ
LJVPMiB1KUVG2YdKivVEoWF0e1w5TfWIYX9rZOnSuRpLcBpPpDX1tQKPdmdd8WCa
pRIFgc77Ua1IGcJr+bdesC3JTUiuTBhAmnXOaGLSfF1n42TFcxDRReowhSLQDqYv
vSwROuWLfF46OxoRQYx9tim0WBiP1x2AXAFHrDBoY2gplbNm5jqQ9KUI5cXy6WQZ
SWK5p/CNErvRp/j0kt4NJAK2s9TYBf3JseKVTM6OrRUW/sJ6GMmASannlrQ9WvpU
lUlfujCwVKkQT96G2DbwhJBc0bFPF9f3NkwRRilH4kD7p7sfY13qF6m2JTYVB2y9
mpiMchXjz56Xumg1McNiN5zAG/otfkdRP2WOzY49b747pM0PxBWESURUYsvxEcjQ
CA5sAyrHJcXRvmCQFrRXYekeK7bwkRPBTOpud+2zAzTGnN1K5YQLV20MOz6AMVZT
tOiqKwcwz8AN5+LR+f2DmvnBadTO23hs1SPUQClTcDXR9a817ngHsLNMVx1woYwk
18LjHj1YyFb0YcPEAuQU4MPZ/xsn3jdWxEFynUSR9CCK4YBEu1rXF33DuCJ6nI50
2k796XMXWTJHurqry0Qk2uHkXjrqdnkriPwHypbzeUKaks311FkAUKr9qzVR+VWB
JusxHSzwpdq6XXig+7cSK5Qh4FF8eFQY3dEq84hwZ2ccAdgttv8A31WJZkFjZnsC
QWEWsithztdNsSr/9sUUW8u2jtGr6O7GebVGUrLcK0woqX4qdefXxhwwffGDji9Y
mzQd0G3MPzlFvx93pLhEX6OfrhFABe//jYC5toBd0iF6f1pOcEdf4A+YetCmnHRD
O+s4Lx/T9rq+QFWdj/XQYgSswojBXoPzLYokkDrj3ZhyGBasXJiPEX34OWN51zXk
4p423fb1iiiSCVwNYVbJ9IJ17zpDQ99WrR1SO8uq3tCA5wbR2vG9g+X2MrAJmz0Z
y4Eb2cK/jCHLIyeRYJ6aljfMPG5HoTYgrlKLLwClS+KOf6gNqC0jXQ6g97fB/cGP
lYqHnwqGGZF+b8Wx8eyPqv7T420WToIEipBJYt4BNB8NmRuT7RDluillrUFpu3w6
N3to45jG6Bz62svJVleg04o/bOn1nC68YAeynhlJ2Rw5dMrJtOSxzktYWgmBap1v
dIc3AHwG0Zxic2XYyf6yOTNUNyEchom+yqel9R82CLLk3xLabyDBhK+hQgr1/k38
HakHh5or75fG2tg+u7l5obvwW1+0+9L+qo/3JmWYWc7wa4xwqqgSeHi6sD3IoGqW
idf5wDQYkmA5XIBbiIPGtZqTJwbhzo/LdLA5G+1yYH5YdJQWuCw0J2GNRF/BCnrl
vWAbwHlzezUqJ9/h2XyjSL2jrfN18ZI64ozR7/IiK1Xuw1WwsZrgZRKtIjiPbfFV
fvt1x+UWYoFX3oaQi7kOmAqLwB6H7pjlgAqjzwdiTCD6DXPT2xt0Hti48UW68Msg
B50Rds4LQgvfBAMl5KQBenxz51Wj3yxQ3lamPtpVsjt/hftwhNEm35P96lkjVP80
Pq/RcYfgwTngbZV7a/w5Luo/B+/+sWbOXuiCRKocfBG9LyNxLL1RZzfaDWrr3axl
1CWYucE6SRJAHixTNUfdAGXvd0fvI4UyYNTqssWYdLiudsiQr64Ido8ByCMC1vtE
QDmi67WtiFLthS4PsdzHV3NVApqJ1mol9aq1OizHANj+Z4i66Mla07GbJRY6mkfx
iM3jRN0M1R+T7sqLL60+mJmbz72b76kDi468gyFmSYSNvgEPLknwXz/0fwckOScR
VSuZfFdcmAyBgjDuelfTAhttPcpP2FPmCDUbL0K6fXy30R3/qHOmiUARgOeoRzTU
EBkFnWBLEdo9pEW21X+fl1xhOvcQaMdWDNX711yuGERmprp9UNIuAdUfSA/iczbb
Af/YGh8ldQ3iq/U6pY69shHL/rajP1bLqV8ei64cL4xA2Bzizl1HTeG5deL4a3K3
TBm5hFp4awyXy4NdDPwFCWJ/JqbDxDRfTCoBCUR/0Zs7wmpTV87Yp+UzKWSqZVez
qCXbeuNjReoSydCm8VoYVX5kHffZ2DwgjklAj1wsFB2xHseiBr1D5dyGQAft9hM+
6hIPvyxSJ108mZA045UtWjRh8h1qkvlrwKJafX7yMHXlsoH6wBlhn3GPm2MZFH9M
aEmllkxCsTkZvd/a5WUyIyUuyHxU47CYqBE9kvgkVGtTcG9XUtNJlbrucdR89QKA
sNMUB2cSOkz3/VlNIAtZnON+4Hs3A/2nylXVVXZwPq3x5iOEQyua8rJTwvwhipuF
LCPP4elFRjbUbVtO9D8tRHabEiOeGtppkFcaNhsTZEbE/R4gRCJydRpIxc7k6fcl
KTeXSrPlKABadnae0sQyXvy/FmSwuB8H3dGhalM+AdxNKu0HL7dGANRC68WUtePd
hV2AuMHDkhQ/TN6LthAAL0lkuVGy7wK37i34EvL9ghMGAHyiXrTiMjaSuXaIEHvp
BTq5SJHTb8Ey9vm505ZhtQnMNqAb3QycX8pIDoiwO+btMuWkacU5WFsNzAK+bftN
5gCj1A3UyCYKQtprwYX88ojDibv4wbEJ95kgdRbBcY/4u6hJSr1swEjdrWE1qbom
kEd43Zn2gMvOAjNY/CjbMHeAIBt8vzhFVm1MYzIViZaDT56+CWQ9KIMZAyZfyBdU
BqPU+wAjo/e93NPKUGh8A9ySmq2FlZ9bo8suujBy94quG/j8jmPhAqS5A9yAPLyR
niTXX48JvtMsIqsDb3K8aDIsRxSOBFCWUWDKCbxcJBd9WXePXfIVZwG6YrlnA9Xu
g+D9YBlnjTFJL8uYXHBIFeripx0mo1qseZ3wPsHzw0xd5rQYeq6wRrdCMnv/2GoE
TS5Ak1fYgWOb0zN2r7zgp0U2+yiwUnY/9etJijSfFlwtIN6EVt4KTFhad7CUutxg
pT0WItnZ8iMgJ4fxlZJiLGijYxtVPCf6YLmv5q0djhNX3pHlxkLNTjggHLpatiDu
FsQVZQi8vjJc5yUkXZG20E4BV4iVDUrTW5dwXR6dXktOj9zp0G2D7yR8TuMTZ9/x
kv66eci3X+NPhD30QY6FPwOEpZ+j0Lrlbi33Cfo6Vx4=
`pragma protect end_protected
