// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PVblBakbEuGxFoSuFvTzuPtVmyrpDa/b+jYi/mOCg73dZ0gSPHWG1gkK8wG7tc1W
ZeQbp4x9EPVJ1WmzGUhfH6ZPk3M6RWW2o+g9bLqgPO6KRLStcJEZxkrOBvlK0iJP
CBckXlHeRRcd6rQuiAU1Ctg+sy101952xh6jY/Q3dLA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26688)
DxQJ4CXBhoPDp7dfHb2wxsv9N14LUxk7iuRd3Iug0MHOefIQjnhNbJ4ZdIKBIdRP
7B4xYpcHxaLOHPgvnOA2IOgSJXvoolq5TLcZaKp9Me4M3T2Vp3KJsPHMKe2hgy94
bBqOvfx0fdiynin/UrKbqgyUhndtCrnDxFeO8rWpJ9FHbaU17TFqtTEtA0BNK4vH
ayeNSdDERFvvUpj49lbfaPWnsHaSq00qxuLQZ0ihC1TsQOwccDba4lw6M0pkxdEU
8RGBO8AME4bLeBvd12z7S1UR55/uuL4bMyYdnQ2uj+Jy7mj2Raixu5k1qJFzIcyI
fOP5ZmKhzfX/6SuMCdBewXXJz3YCVRE6A3nDjsYDeQIfWqnbxZeAzxYZoUiiG+dv
JMziuONiyK5rsoxjl5Mk7BTviXkmzPxpjIhUMZ50H80uLO9ZfZa8SFx/OycMHvuS
k+KLtWUtty2GfnrKLQdi9B9ozXiNVgkXjbdtHo6usq0/VlIIaWRc79J74MeLgjqU
wplsjPrc6vdNHKnQ9TDJS6V0O1Xi3lGfBt8xNYYPnSzaLBDSKZGSSzK6p8bJ4i8Q
qas7tCxrb21FZvrP6P5oIyQdJcvH34DDbQAZoWFEDItg61MTgX3It+fsJuJbaO2k
5YBZRYlNApmEYUxgKmF2qIzeKWIKTWKh0ggx9jeKxgTgDWgITWDdPMa68yIJQMqK
5kho6KYvB1VxevHyBxUxOdpYXnsDuDACOkCEpIyvgp20Qn075JKxVGtixRCzDgNy
vWFpcqBVotDf/8afIbeWnKJ0s9O+qMm4uKAFDCY+iOTWiz9xq5sxGkT/YYgpeYfU
TioLpDijHu69oZYj+U2foSRKQZoE1XfVQGgYAsc6q12b5bgelVlYFiEZzOToreVn
xV3H9PheKhknBSgxkfSqKfgTVjPHFmGBG8Hi4h6mw2CEZyKZTmqIZxRIdzNYTGXb
L4+6QDLvweMj/L2qKwacN1LuSHVM3uSPMaepOxi9geCQGE/LfpuaLrvausFSb8HN
p8XxyBFppJJGqIoj5r/OZD1Q5sYnlps1u84ptWLM2OA/YwsUlWX52v0l1+gfGPcg
NJ8yLkwDq19NlYmWRDOkNZVdNyk6ecUqojTBRqWwZcsTfICaEf7OHkLz5VqVsiYM
aYl84FIp6N60IdK3dfVNudIp8S0iz7emM5Mcs98oEbFOQZpXTT+jDDgGvCkr8cl3
lu/avzAqHNYWax2AEZnwDak4XcIJl/XhR/6eTqcS0U6DWReePhuBOIO/avbgpbtZ
EyPV8KWShAUmIVxkhYi8RPqEkf6JedpXSEtDQvK9XML9K64EF6ybVC5gD8gggEbd
1gXiaLhTjd7cR3+9EwMlNzXYlwTLKjFJiKHL22t1LaQu3p9iENEO2TwYnBRDmP+X
UGlJiJL85AghxvRyX7Rfuy9KKXAk3uGzGUlfVjOnCClnq0mvgufpfSr6oOZZzH9r
V2JEsj6TWsK6t1GJE5jpJkmO1E/9IUxd5GJBUIrfdBluAaI1R/2ohvzHD/MLW+kK
qrUlUljuMQ2l3attexo1f1S5FsN68X+nvtlPT2jNat1tZXkmUj36PW8AN2M/Po71
9hZJPTfeU5QuJQ30v0J23I3bHeNKj7xgO28N41ZCKa03H0bssLGKakguTvJIr4hv
RSAPbaAwaE7ii/fAwxdwq+dyWnoVcZpN9+HAhksWUk3Znbpv6clfx9XScXTLbG0V
lIjnhklHT/mLwScGyuLir1x3ueed/Ls7Vrz7evojY0cuuqpSji71VH6DluCsZI+m
mKiwkbvCYIFCwGkMfPlgxxqF7J8KPu3YM5/DKfcQXV+XDzfKrtc3ZyQRzeJUFsPL
ugTZn87Z5nzE/NcXFCK6p5NVaj3Q40HsLiDqyXSUE27sVPrQzuaZuRdecWSYZhpm
C2xGtUixLUmCCCm2MJ5sb4wF96d5ZUP4sxSu8lr7/rQPsVdw0yd2iS94b3eDQjuU
Wxz5r+6i4eP9Q+CuZt8sBKaVSjzL25qm+XPcrnbtJE8V9/MY1Izy2jb4BfxeFxbC
UrxdHT4pCBwt1bNQo5/XlyQ0KI6YFodjgnu8b9Ba26wVEkxW4IVJipJ6n/KSgeUP
Vtxdbt6OPytdXQMXh4CJNCAuGwEEvCr9dXE/79qdl4nfpzvNBiuLnMdDQtyr6qJ/
JPbQFEpOpNP7v07V0tpMz+kz8qC3db7gwl4b3+b5bEKsUxNI8doPnwXMy1k2Lf8W
J/8OaDyJPjsBpdb/oI2GsNBYSnpsJMrdR1r/AlZIab0PCQ5Ku6vM/SxuNDp6vDR5
AAxIj/xiBUKVMWHEKwsaVwptHxV4CtwojUgt3ejcQpLs01OaVyh+DBNqpG6cLZX2
Jcs1MyjiQ50ulbjSwl25e1C1rr6Jw797Zc8IpedOHl3X84NiONe9x3ryCj9cEPAR
biISSgWr85fr8DYN6P0+YNm+6VGKKA2DMTP9ZUAjgnSNz7O2dOiDZfK0dR4iE0TK
EW8hYeJOedyVM5+muB7rBc06/21gEBsit+0J9nhZWqUCdK0o+tP2353DWDsyRSe2
/W0CXJA0Ktd8YbsbEZiE8f4DjGjNnFn1PkEOsCpIxjOqUYuxR2BeRGGUKv4MSz2x
4ceA0MAuJhtQh4EzlEsP5KUDULCVh1w/wCSJcNrjO2r7JN2fqbzXX7HFEihcw/w7
FeJujD6zGXN/RviZSLSYEjsrzdKivT3bXnEGvJN7gJOKefyhDae2D9au7ZxwNmOK
sUSa1xYaj6hhNns62gfrU08yiMITBPh/haptGGp582iYZglpcrCj4tjUi77oMBfr
ld+E6STsna9rRSGZ89Qr2jTXYlCyU/0WVAoC7kDjo2diEbZijSaoC3UEvsvV+H3/
LIREtpdC1A3eK3npH4hJsAIf+lBwr79+/9bQzJRTTbIlQ9YwlSOcQIGu6dNgPIo4
UXayBIXnESFTL7vkGNrmhp4tQy6R9vLZgUK3DDHbzjmV8LFtbwy45FSvPZps83+7
ET+/Er6toK7ipjnYdPVBEwyuOaB8bQ6MGygSxOafXyv95bRMUG+ommgH3Zn89Buo
pIcLJDUz6YmxQvd77U2GGfqT+Pgi19FoqSFLlziRGr0N3tS+6y3Ht1jJDsA7ONDf
iVlt1RwI+RftgNmwTNDZ35Use9yivoZnOz/xRMKdhNo2FnbELcfMB6LQW1hh1P/Z
BHGMFF4hv/PbyiVGAzuT4TXWiGUJRZGVORmNv4xWbcYJUwD/6rJikNJICWXFfbC8
auisK46QFCLL5zbQ/2rKArhqdQ8YOm+VWz3mTU+YMeRedw18BKtRt53Nsbu0hoCQ
ikaP4By9vE1X9vQsdU1OJEDE9xTCh7hqquqSpzzIK2EKGyFWcRdYxZdBgb1xnfJi
97WTd+gD+Ejj14mlAO3fGKVDzwukQ6EcKV8crcvwTlAMYPUFTdR1eyiR8Su+ac/Z
0El7DnmXRzy/cMmVnZ3Awtjs9nm6V6I333wukxfx+8BbsSY1vKg9I9EwpxlXDgDJ
+Z9Z4BE2QA8yWXbKfqU7QVQHoSwc9wpEI3EI92vRAhi6jl1kvtNGkqoIEt84xDru
P3s9wHjD4fBwLoRmDnd3iGcMk6vLb0uxn3JwsDYSJExH8YE6U5UXlrMdrII+1ttz
CyvdAbkB83ml3Z8hLXES4o0sLfATN1bB3tLYr/7CnG3pk94A+XlyLqg3RvpH9wWF
vs3lCjaW9Zl0442AQRBKjqQvrfNcQrCI9x7C7iqYGwNtAXTApEW+uyNSymF+gBon
wSX9lFzWHl2sXYd8FT1bSbXjCAUShp8krLxwBMFa0dM3tJNOyNGnQWUFZCLTPXjA
z2RjNxbabZlFYZgH7TF/OY/U+CyhRhXBte4NX9DE71Kwrym5WK8pQSk9S4Paf7VP
tNR1xW/QROsBuPtrD+qbRJwvOXsWDY91vuWrQq+xj/SMfSDfyDaLemc3vF+ewsJS
SNreZunwqiH21GBp/+TsmIXvUPbkEfb9GHrRx2e6GsrUm2F9bltX6mGRPzGzohMs
H+LEbMo50UOmdJtYKjr9pyJeIOzI3Lx3V1a+Qi+XwT0DvIApS7g/qjlKkFeBKR23
oBdg+Ji1l1eD74eroc4+fMgPzqJhvbsct/d9gvPMu71GUTDOqMwavXSJHWOBO9l2
uxhw3WHRAHf2qEQYtaYoeXzGpsTpO3XWUMP5P9PniW7EgKoveJKbO35v5jL+jroZ
WKr75FuZzVXCZuXI5nwFRsKcHQi33XApsGJYaFjQoCcyZbeVOVi7dKE5BCFlQ7yz
F+RBmjfxa67ho4ycaIcHpm2y1c+27pcj6V7eu3OLA/nClesp+VDrw/wjKWQamnd3
E9AZSQQgTI8RAwP1ouKRtQ7pcT/mUOgidh4NUXMsc1fRwaclHHaRe8mpDe5pjf/7
BKjzmjh86f7QVrcq+bB5WisLuG1UHz0vGm4Ulu2rT824UXZAXjqFVczkb8gBJ6iC
u9bRXu3dOt5vME1bWeLUL2bbpFjBVIHpkQxdsnUxYGrXJYb8QeBCBIeMYSf7F99/
BsnEGf/HSv+wSeU05io4uKYeluasGaIaguy252JK4CFEGFK9t+FzptXsLL6gR1Y3
U8eSPsFd6Ks+lzOZbcx+draBC22F3J9yX4XfEWzscdzsybflmzKwqWDmGVRO9ag3
cXWin6d7pJyRxs+82mU339timxgzU9uUQ5Ukb4N6x4z2QSIs1HXhsPqdjag1OY3U
XHXlRANvmCpHr7t4YubSaDc3gQO5bGNjf4/oOlpZAbo/RLSZVPSN+NhOvk18xSr9
ksosOBlDwcVOdBLb1xp90TLlkFjitmo2LBG546T7f+Gm9DtE1+g0ZwWGGNCXgKYj
hVdWI9+ZdsQ0ZcE14Bacr7vq7mGCXchpc6cOFaFRkCTd+4z0t8nAfE3z/IjqNuZ9
Q1Etk46Co3VX+d6TD9iHB8+ZavnpLH4UImvSr52I/OoVbchJLRBtaL2fDThrfUb6
9QxTHLHz62Je6k49jLLR2dOCNYgZSZef5/XO5M1l7pmqkdjhjd3lENh5w8W1VEE/
1bYZjK0NSWX9vnvwDyMIsOG4vOZkXUd2dI16Vixf19Ecc9JrETo+GA2hLqddZHZQ
VdpftoeomFQesMUACXFxbdw4/LHjm2ljMI9DdghCe021PDd61xIh33OoG/XItP1u
xoaN/MnoVLUbMEu0OlEXGdGzYNp8VjOSVp0lC9g+7YKkHG1y2zM9fhDqf5ml9VPj
Icx/OwTpd9MJDj6+zTSnQNz6760KxBXHM9Sz8v+6MtWnTpq+W9XgJLjojBcBiiLl
uz246rtGBdFzmv9BAp87KhVNQzCaPzIdmlJPEjx95F7SAeMWKwtkx21YN7YEAaPE
f2Qw/lHsBQNhZ6AeBXHeQzmwnUo9+L31zZ1jmfqXXJIlBV09CVxK0QCjgstRRPI9
uXkYXQLgSr7p1esv9iIXHfpj6liNr09Qe0pJWx0PUpeCT0pF7zoIwChu3m/x2kX8
4o6ezmuB/z05dHm/1HcOdUL/2n2+Cft/ntJWso/WCmUjvMHogjS2BYNmWHb/+cyT
uZ2ioNeQmYqQZOxXVkVVHqrGIMrWx3gjxUDg3cWKYNKbXiDGw58As3SSObVSNvU4
+lWMT95gk3KDTcc8u2F0h62jQIS3OHXIN3rYGoLljffRfm2sWLndZt1CklQ7GAfC
D+4Wz5oEuLeYqrpxoV/BtKnMBcqu2DAtZht/o6RTuMOlC1PejVWas0WM27JfMJdb
lAuLLrZpxYf4CtkzY6rV4WfXRL91PlNfE569PVoZRb2tOBNlJ+oa8JWGXj66wZUI
r+TwEZru9DvKZS8EMAW6ef8XrwQKvO/+TcICie1P4T1SdcEAQCQnrsRAqDhlHj3n
VmAypc7OUbcOVvK91nLAfsh2QPduuDtSwAdhPa4VwqzufhlckDQaeGPMFnfGFV/6
5Gt0TV3ag52ztjxtnWp9xLE1bOK8yjpkrHPVkwIEcnCCJW/TCf8AdJF5QywAMQ3Q
rW5hZkYg75AnT2+mYbR0Ncd++e7woV8fY7ePdeEUlI4Y4oeDDtXrSiqmysY3Y3zm
OJli/qRh7AewufNX0KeNtf4Yxl9RYsDSPYNORGH8DsqMU/MkYu1ERx2JL3YNlpcc
hz6NOZ9pH2zMAaH6E/Lx4U8PgpHlid5gllhS4+13wGKluy/iF3zIGmGdU5iOC90q
SZLVPYk8n0ITtF5RZFvP7lfQnWbOxolEYzuR0toJj17UI1Ydf9UanbsTvaHcO2kD
V/JZtHGA8d8mxrjJp9tqvx8r5tCXxn6vXIa3Kyy/YTKZrQa/71yiaImPWJC6Mwk6
jaP3aUF8w6GOit/XimvZ+qteivU6RUWXzjyxhFbc4m85VJB6RiY+LMNpjpsK8hJy
ZLeg6GyHFZ3qbv3Nn3Vsw2E6nC1kN+jyIutSvu5yHvCU7b4H5uQ93WfCcj96E2Tg
j55qrN9Jtvw6pcjNIxSI5C73sVOi555UZ5k1OCMS/Ar80iy8G8S6JrlEFYkPmfWw
jY5oZ2PBVpFiFx1wR+px5FAJwzAslN0nCjI85/jPEIt1bJ9hoD9lhZX2BHGZirOh
3h/6Z54PCLv/Zb38Yw9GYEyA9maHCp0CtpvUUG2OxWQd1+sH4kSfBuxkaSjOVHou
Nel56trBoONYk6LBEYvReRLKnq8XdT2Hh4Pu4nmEavJI+fB24AJ9d24VUXgJttmx
DfRI4LHZVckQEjS5vJq1OqbkEhOmzHcB8U25m90Zgsq819EUHUYzKXVODzo4lZI7
i4NxrmHw2og+3E6qK11kKxt4QWVziXYMpOWpcEzwRksU+BdZ/v99glIHwGNzI2GW
jQfHPZFRZrv/BYRT1Mp1DUAaP6mL3rgf/+IBLdGxTeCVj2oHdHP2VJqZJbCXFk6c
B1gZixK0h8NDijk//xEm1sj2Z09oqo5QLPRAKfTdpqjLOmIP1i7pbJnTPvK8tGDE
Q8Mt/Uk11mL3M8sVJaz1J6jKVqg+nGQeetpSVE4DLB8CkoL6RPaM+BHHnrufTNVy
X8OxdlAuYBrosElQge2/RWN6NgzUVY19VvaI4tC/qF/mfPzAksLMoI7jCGVxVqZP
lPjIHVPsZ9uH7XigPEnGMGiFZV08U5O21MRicPnxQqosriHdWcK3lnR1l3nDKOzN
Iv24+8CSij/hsutKNS+xhiSIcaP7eAOHQQee2CicMTejNVYGBbDhV3/yPtoF5jXP
ymsUNnBSj+yaBAZdIpcEwInTuOr6XZGcwSI7B4sEGn1gdKlo3Wv0iAKHXFWalo1N
BSMmo/oZiVUzXFXW70KG9gAp25TIRs4Rzqb2NFHg4GcPevhNTdbIpwlIYfFLEFK9
9ukIbDKnvoneWJ9q2Ho7W3pz4TX1oVEIHSd0HPmNPPfFcCKu2qoCwwb3FDtRUjZy
n/72Mj0zgNUUPorwMoXpm6YyXBOLF6kGhF2Bku2yAogF0xZUTxhqPdWLLUA3Z6Ir
3ewwFSL6ZhkqnBb2t5AtaPLe4ss/FoQrNYtCDk4MdKpfwnYkD1EJs+f6uFU4C955
vLh499vNqzm0wWAymj2GEAA3cw+8xlw9u8t5NMWEqxs18YG60oq7pgi0LcPzwCSj
J17ZaBNCYJx/We1a+zampZouoI5VtAcaMUtnINoBAeXSXIbkN1J9+n5CcHycK4va
HoxQX572/jIuvl03nHvGdgNuGheASVVu3RDUKjpf1FY4LJxXsbDQC7nvB8PLSvcc
IOMwJ5wzogE5Ug9oNwupjPvHOqLSuRhcWIl6wzPyO2BHQG2MhlygQG2rLbMg97V4
eyGBoMcgnOsRuIt19vnXu9zcKCGOpJiippFdH0NYYRqGX0ZW4yGgMZ/nkPZ7uWlq
r9TDSC3OyE8x03ZxMOwrWH9EVmip9pFygnkjd2635H1ANcBQ+UsvZ2RfLdYcmxy+
9fE6G/UafPzJfQzYwYdzNx+XcXg1sBH5UtOv21LhBVLZGUN+wJVEZaoJ7WzTZCSS
plyKERu6FsnZEQEq+fQSoS9fui9l88hAZRP+UopYnMZo3Hv7X9v/uNm+sUWPnUrk
6hTPptrOWMnZ2ZXvjpQ92/Rx6TqmU/Z39rue+NhXD80xd8FRkDtvimjqVLjjDgWw
nLltiovqWYa2Lh3/EIhzuWq/qy80p3dL8K3c1w5bqrs37iHtD98y+TOP/ikZz4a0
U+8rmNtH9zUeb+SHwyN1ARSs/tLQ0/zD586NSBH7T1nqx4fsTacoqydrblJ7dTuv
1hjXJ3V1OADKUicXASBqOkVtHDtDm5s9BIvPY35YiVxiTHj/aBIkZO44pK9FA2go
GbYRFNip/18kmepJit3SGoyo5T9lsCqFna6V/0lgdfEjbz4gewGaHFjJsANzMUOv
FIEK/9iFZi8z8xrHv7b1cF9unPvbXglmdAizDSxAyqqrOiYT69EqIb5ldItC4wom
k5x3QN4io9Or5PNVohqRviMct+MkTWCkkrIG0aN4MGQYRTBMyANh8mmi5RjvElat
alezsRxVww7IcXGqNoC/58EU4F4ulJ4XnG7MZbCbfxBxZYRfOA5+21MGZE99qIFP
vFfP0yqA3S9m0DMBOG97XRtyICi+jg4l5opax4ixry01mSmt0JCibcRKFDDoAH6P
HF41OIigUTjZi8z+1yECWttqhrCHEgNPRAS8KSffb/9dyTL2Nb01ULIRF5O+o5IU
jaZKaWQ1C6bQh/zpl3oZDGSNp6IzJoI/XBLTd4r7mJCFuDOlJW48AdxzKG1puxkr
KomUk7bMbNc9qY6GKeKg9sMH1TjoX3hxF6J/0XRbsT3FfrQNz3Q7abjs1rC3eu6k
pQn/pHHlApxIaJXVVG/aAUuQ6GrKdUet5uLtw57DN5zroLAu8ynGgO1fb0LQ0YX1
3mRdA18D0fAz35E2LuL09OaTAIBgwtIh+jN6mD0YpV977yq3HRnnfAfD8ODWlpqP
7DQKuWZCh100a6vsBartHOauxsAZ7xrRvyIRjfcK63cvOWw7aLjL+kECJbQ8s1rV
04RAwJfJDd6gtjmy9PkUEeZyQXGgO4KFqohkS1PTBxXHNSaU3pmUoLAhfkcCuz04
a+RuU+q8o5Wjzy8PXxVEUNV9se2uQ06tKyE8KzQ4rKgw+yLYmUWJv80kPVb5Uyxp
eijlNgvkEvA4E948rzI2uDBkmmZDan7VHBco0EkC9+vF9sVi+FGYp+doSdzdTf6B
Z6j1lcNNUqGOAmsjOLg9kbYyrXgLfbRTb39m0DtjRL73MsZ710hSYuoWLWfO74IE
rOd4TkWORJ50A9vOJ3vQNX6jTgy0L+XyTMFVT8GAfqY+lJG84ZNFNpJubb2Osg3P
xcr66b3VEMWSWspzHSGV2Jbgb+Gxy3Ij6wx5rjJrBd3yPqFSfYoITvYl3LjvmT0b
WGCMuaB+1iq4x4pNGhpBhEZHVmf1feiMv7HoVZzZkj+x/NCItyn88ebQcPmnQdee
hCWig5G1grDbvhMIOP9Kdz4HP0Mgow/70fdemzFQ/EoRJ2fRLr7RVquGm9x1L+pS
nTQvosCZX7RCjuOX9vnGiEHtBMk4Nzwjk3jrteplENk3y/MXTGxk7eTstmez4obk
cMWB2SBdL7VwT964oYNmM+rdc83bKXenprqRoEobe10nEiEuby/W8yHFFZF2/AJb
ssGSi1wUAUizA0BVRA8Jsk18rDT7gx2v1KIEumR/1PXFdLeSp8jLqzT1j0yOmg+P
N2ISf2uthAyGg7OIMwFg3YgqUMJKtSVAAP5FdtI060GKuKbk6JCpdyKFFvaKwyGG
ET6x9MThGRIiR/K+acQvZJmnZ9s3/3bsEkjaS7h8oCrFT+Gp/F5yq0B8Ijgjxkp3
vc0uN347deLknVFjYiARVk7x5heYWZuQ8x0a0GIsnw2bRuqD63b1zaUsoFsapqA1
BcFpDMvIgvB60K9Sl9TYxrM+YOCWBFxJwlHQZveEWOMacAedIhtpJuj0WxxxQ8ma
MlaciaS0REhTHPFYzBO3uzvls9+sFs+nozcgSlflmbUQGIloA6q5ErCzhNlZUYho
SE4ja456KN3cZI7G94nbtrP+hju9+eTYhJkE0DyHSRgTnVXIWQ7UJB5Pd9W1FGCe
F3Xi2YsfjWQZ6u9YD3+iYf0iuZa+bUo+OctI67BHh2K0qvRwqYKHyoLDPjHHowpy
YfSrxdROGowLLaSt+b6c3mTcl5kXYLg8+P8h3BAj8DqtWWccoWeRxmXhpFPZWxp6
6105XRIJn9f8ipj7zCyU9lpRoGiZNdL8OxkJ/QnrsuONbmu/4ZZJIK1btePRC/5b
h590oVTgLcRhUJrFIDxMBjcDAgsnggPsKl1dotAZZd+89FLWk7akTtYFbc3erdLL
epK5v5oglTf0h1BHObvM918vglvDPUqgNpr+FOTL2s0Zlr6jyrpvCj2Jbd9zTLG8
o114etCqZCb0DsL/n30Oep3irtDJ372iRp03bDV6B2J8mvzfoEZwog9HIwMH5O+U
9R1JACcS064I7G8JZxw2QVE73RkBoJzem840XEhjubwe5O/goK9LozESJl+pnkZ+
8zsQMTRSjLHs1u0Ss34+kfE2XKINrA9gw2zR0B6fCDpcEAeEgAC9r+9SxRD4kpWK
hClvkKm4DIgL031ojywaGpauWGc4d/K6WQccFpasDIRqESbInyqZPoy1ZKZ7RFAD
od+v43cwHP4myUN/SrugzKtwIgtUcyZQ55CsiuHFaiWBtA/Hmcu9HXUdORDtfN6j
M0gOn9NIyMWMGNdkzlA1XBIliI6S5R3Ila1z7EXmeWSmXObfdbSjUhi/wvuBfHFT
EZkhpftjTL2JDsJ0klVv/ITs3nMAqmVK4/AXm6pWCRlCXxTDVzljq/zoghbPoEZY
vKGjx1HGajSUdfycGNuNhZeaAEOLF5N591Cb78tXeFD0BaC6fxrK9PYJM8XuMpGU
xSs7Vd2g6qTEqAUu9XnXitGEhprqV5xgyVpLVeNsw4WQ1Yv4v/au9stcECKfCOIJ
CgYrVDrjJx3aZax3PRYAWTZedRwL4Rl8eBcoy1oP9U/UFupIifxtEChP/PEIok84
OcucBKPWNLyw9d9EDTZRdXwHDe3kG/7P4LpPTlTcrmNlqIHfnP4NCJ5GcjokrSh7
fuIK9k4sRvf2UahPFKjDkihTlcllB9nfbAFLG8PltgpCY9PD/97eYvdyP0X9+FR7
McBjGKT4nuo8uoflT/6vB+FOH0uy019PQGnxJFw2kVhDu+DJpecXCl9NKcFiokFV
NXD+jRxYNMXUPQE8bZvKmjeJC+O0LJT6gKque1U7ZkKSUwlW3ihp0qBUxPuVSjxC
sE9S4UyiABLTrOxpmiEuJjA/57skKZY8ebmZOUHZTLwAnkp879J4tGIf/2WfJzJ5
dtkKYNMsNTwtY/GR7XJZcnhajuHZIWbX3+GdVzfdc8KcOWCFztB7i/s2NIe98ZR+
brprB/QH5O7SaY4IVO30dNQM7GbhYJ4J8fWcojjG0fJktIz82k+VWt4e0SJvfkN9
GQGr728stVNzXrWRv+Bmns29lP8GErYQOLkbxNvyVnaNwnVqF2RpJghs4ocWLQd3
mtkOYocJxlBLwaAbxoTE//k5fG/cphy/hUhExazCIRCy5SiIkLOnXlqbDdj7j0bN
ZQVcVsx7vzRv+UOE5H0UfoitTm1bOm4REg7ntX1GGhVcdrI+FNcGkLeIr7G9JTjA
hezWMOg2LgRD+8J2z4GaKycO44KLP6E2r7lI/ao6FZcyZ5D3pRxE/QP566suxR4p
U4F27alpASA9tcqrMp5HTvGr4QkxS01TX48zd1vdhRQs4Qzq+QezrUiTUODxg16y
AhsAVzIS31Nt5V8QEm8VuHP2MEaGTaQmTjmpAwyQ3ex3u9lpaxkUR8ES86+oHUeZ
U7k0it+i+QTUVgADfzuHqImC4RTWMGnsbhZC2TEQcBkGRdNEp4Z//RkvF3us26cA
xEKYu0jvJG80SZs4RDlTzKZEv1ZK10LBJ7gndelV46p9XQQrnqVHTNiZ0VJP5M2R
n1Vxb+GxWqXPhJkcdSQNvY//X7+cGguecIBh7U+XV23N9HFACG2Td8uJb2wXeuH/
8c2S0E81tO8Nq0xOmPDHLazFM29wLnsgGDL5bIrZdlN957mT0GIxAHYYasgLvfts
quFDgu2bDryBM8dK1ealt7J4ZB7TDH83djKGJixOH7l8/1e9dOGKFsX6nM4p4gLd
3BjvD+XGbUSCN8WxHzwkI8A6iNT4em/gZpQaw6bwkk+3UU9/lUPpvF+guge2l+aN
mij+srw+lnd2x1GdVOBrdd6O9hPZUbnQlMsH7VktEIKvjcMxkyTSPJf0T3pS780I
c0b/EZzUbIcUUpt1beZRoH96ZEUPxs6nxfRW9KDO5a1tGDRWAQfWFCRg6i2368d+
jINNHHiY6Q0VtzvCiEwzSoNii2DcT/fRJuppxUxyo207WpI1Loe56Husn1HcypH1
YGD4mWnTf0G5a39g7uPnk7yiQ76Eavewsedy6ubTA7NpWY1PPxBDKGU5AvJTD8Ii
VdZcOUE5aZh7KIEVZkfO9TTgD173EnhF+kw6bdmAxBWEWSsr14NWx236GmT3SC9a
DAeN79yJuhfjTtQVHwdPLh08YT+M29p03c67UdSLjqLp/oUg+neTySOMzm7aQ38W
1FKiD4R/lNLogj83xZXW8aChdVkuKaDHHNwbxJ2mZH/KMTkk4NXnXa8lFmlCLhE1
IDa7SKe5h6nIZVLZC9UDnTjU3AOMm2pnct3QXQOF2wRv9zqyt8LxFcUCArgH8MDL
3tsVjSp7B020h7iTUUPDwXM+ZEGQqzxVoFQFrBiNsepwSVw+DDDtaQjCAga+eZfG
6DWoqiO31FSET27dt3YK94ExZOP17D3mpt1lMk6XiT3fIdiRpXsKLl2jYEF/IQ5m
xGmyXsxtuhmFi6v1OAR8lRn8it0wKvswPImHJJzg75r5t15gfH3Lkh/I47fWrKSo
2CnNZ89oEdAKwpGz6tlg/M/Tou2GnEiuEu28TeHXz41ga54DPD+KbMO5IRZkmLuA
PN40Iim7sDzyKYNLrX6wLB7pKcIqvp5iKSBujS8bhqLYSYJJvWBmHr7fckazf+ZM
S3ict0ojjadZMskr7ZQSoHcuEZoMWMUiuoWF0NrPHbA7f1oRS37xIglmwEhvUE63
zq7HL6E0rWdxZnME85J3wzEqlFPL2cl45gEx7E9kneTmLW9SDLTulpgXXQIbAoI9
B80NJwBs6eAKxUlJE+J738F0tUYZizy/N5IKUnxunKTAV05fIgKi+lB7Rd61xkZc
qJOrzTfB5HYOPgI6J1q3jI/zgQzUTuso14fmapFLGfS/67cFUcpJw1rCpM2CJoNU
0kYYJ83Q+LLc3OK8v4OLFBITJqwBcI7bf5Yafe544HPg/S6YNVOpg1zn7EpE3JnU
YVxLDvyl+rbhERCDYeLr0jgThDIJqnFrZQGGWcUQTFnaXeDxuwLQugYl2a/aNtOL
Jvhtcx3KPVczFXx3rGflW64S3e9husvdV79C7s8Ttb4h29/XXUBt6QD909yhbz8c
Fb7cgHOwK5Kr2xgWQ1Mph38xvxViZcKnUtIhyxHH2EEcZaFSFlZWB5FJhWvsvZrI
UtHdZqOUL9EigzHp3xab6EdEEwNXrggyN6n+I9SSL9QQBpMzKd2dGDh/hPM0NQU6
pZWOu9ROuzhqmW01PdEOvB4lxdMbpGRb/B0dDl2NuqTQvnH/3rZ+ZIiEC8zRv4Tq
XvVql4uSrKEdQmw7fV1eG49gbFEKVEfD7wia6v0Ts8OsWMIKSSFboO+9o5n5EeIp
s/qaduaZEESczD+iLL5rhF0ZVQcelvyyArXnY+09Ejn3ctlSfMTzNtJtE95fDKsy
P8eztiPNVHzkuLGHBPn7IwQwwq5WZGzTrhu1rD6qjwGR7T1Bnb6unyL01PZSQBqB
vJE7RoAxp9ekuaKg6RF30LMHGuR0SPY2Uq520JiYCAMQXNhcJwORojQm5fA0c9AS
5chRKT3AM4gb6XoXmmErmOdmW8iFypjm5f/j9FJTNItbU9dLh+z9raGExcIv16IJ
PnMcU2tAISzkpQHX2xQ6hSgWOS7GGw+94IwTXyudSicuCCJ140UK8Hs5Bre0nIK9
hwjVE6Nmr80qsJl229X42+dhYWSIX6Z19IG/jRXHzOlo+cqvXgrxKNby61d+pDow
OqOgS68aGqbbosHZ8ZdK7HDSvj1a4jNOL4IbcGybvmlbtYn82UdUt3m4eOB8Y2Lj
z5+UtuLrLP2qPjtPdKohn3VCQEEdeFcbuLedT4r2PLDjwV9mwxYjitvvb1oNUlVJ
MUwK6/kwBWiQg4nhx3WFvQ8KiFDUDPMzb0dLmUzBXWtUxs/0MtX1QvUJrJWWZ5io
sh6/j4rl8shzYuIymcu9Li3i3O9Pck+RwJHxX9oC/YdGFy+N3M7HIy+QdPf7qgHS
Z+KJNP50iusfVH1epQQFMnfzao5ij+EEo6TtZt5Y0Cj9zdEcAA2mA8K1c4OeItKv
izKsc2DxbhSasNVzBc9jXekOxFUGGMt8gCTXRpqz93CfMZjxhPVA3MZIfSrJv4HW
3f9XzNLH5qBn6BVgLUhpsrsTlscJeYRCrNmO5zGSjf+58HqP6dyyZiqH3CB4Llno
6vQW4vHvwVd3BiWd0hzhMzFvZum9Xko4qd2dOr6BNbwnbN9tBSUX7C/bYNEmDVZY
yey25324vJDF9lJomQjeYVOwxc2tczvBikHK/Q4UWjs4C0/kSN4rLKRuDw/FHDYc
yTKIS/vGSKYtE8nFz4r+fzMWhRMrCFpZI3uD5wIRHvFwSgE5cosNNkImUvN0ZT+4
PwXXGg3fgXaQnj6l/Fji9ZF/ctXyUHrkqSbGNsMNV/p8+1bqAFrndZwk8iIe0S+w
WRgf3n7EZCWGHQzb1l9uazXrck4MNqxdse7OAwUVm6gIAh7MgFi9UAqFFOHO29D+
RtlJbvxzusVc/hYvaxxdEkKwVmY+cDQ06FmR+n1Ot+do3xdplZDtxsU5kbiA/L+K
prp5/5VTkiD9sqSjbqTnYzRnEKVCGPu59NtcBLnhdhSzOWuC4lP6QJPUEIL+YLUv
2QhZKV+mRfCOFJDwwDxBgud2mu+bnst6KFej8Gg6yvpHjl1wKP/OAINA0l69/4JT
EGyLAqN75aV9WE7fRB8ds1UYukaNOQuH4DZmLZnUzki0YaBL1EfWnO9eDQCLnNFz
CWnq9XvVV91vnc62zS98p7fyK9QU+JumPASsEZ1wH9INtGjYJlDfqwv6izT+Dn8z
68krLTMhurrzONJghKd972rzMq7xUN6POKlS65a9R+kzyDoCfIltLgzTVwhX049+
JGuotBnT0HWDxOolYYkolOgaG0cej1C+NBGHMxLGt2JmBthssDugCPGZOeV9OrbV
5fLm7sEvPbfBPtjZ21zWmEOw8s0ntzpLFDARDinB+He07WWLae0idQs6QgaK78Yv
18xhA2H/0IeSwnfAqKoee8cngR4eBcpITZXPt310USSzg/oV7HuwV0BXdXXnqPiq
IfZrkQ+UZuP4pKlxdhjOUkKqrNzjImcEvxWng3hvkl7KFW2HrRHOStC0PXkQLqX+
7lYn3lSY7mDD5BCDgKK38cKPYvrryC3MgrPIFhHnwiN9dQelbS3rrl1+GH/lV4Ee
H+TvDbNvfs1l+rxllAyRcdvM7uX5VOjuwhNIyj8xBSKvDT2HsY1J/jyC7veFVwU+
0apOKavRTS0auz+iRaL2Fi4HoTGSyPZ8+hex8lQaOBya/kl75H5LKnVi2EXQ9Ydl
jPrWSjAEhkIHUsopsCxT7iRzSO67KfDWsbyFNE+lHkQtMUSi6vrCNUBJjLz2IWoQ
DvheqaVaDxIKzCAUKgxUy52E67P4eXgYn1nzJ0Ndnhlc+2ZJr4GnU5Moq27Vd2jL
EI6OxxrpSEUMYYowKRXoy+e5n2RsJw+z79AT5o4V/Ftwk14IwIHXcYMmSNct834A
qonza3ZiBT4dAudIDqVfAko1f2sXa6UpMZuYxC1tpCKYHHc5xmX+II6I9JCNpoxE
D4ZVAhCbJTBa2GikFQkJ6STJFxWB0jyhjFy2WUBGypYA5MWxomowsp/OBGXuQFo+
S3jMjaG/nY2ez4WABSYnemVDZxQLJ6KtNLo/oJfvx44r0g5rvyjuUQS1SiyOROpj
hxIcYT+8D/DhtcjvsiRWs6POmuNwgxiOAl42DJgJA/JtLx2bXRa1hW2cF36MGkYN
W/tg6zg5ZEstuyhapIa7AzUhgwe1ZED1ROjAFyooaE1fbsh0A7mzExaGCafzxkxn
l5TmMEvxzeX15nkYVjdqTmYaJkYWrUbx4NDgA+Hxi9cGQX6AxnHi5yI554ofZOax
mPioDW2zKNPzAAkWlGxgwCoDkUuF37P+9zGiXJ3ntXUjPhfgbDCOaBBMKg6meOO5
h953ptNt/vq12YMo+A85v15xJIUg1eeilO1xd0Q9mS6j2ySvuWYR+SnEec/kfXuG
8BSbVTVeIH3NXtI6PhmYQh711i5zyGzw/EXBVZdz/Jx9OuuKQY2jdUmZsCgnLHn+
c2MXro+fjCepSyKIhSoG5CdU5nmfI3wnjRX4Gma9uNNkbOEObwYUyfxMVnrTBkFP
nFlc5cB+A8IAqiISP44zz76uh7xF8BPPm+Wriw4Q68asDgSU4512KWPVUDS+vKXB
auf/sE1KJ9Fa407S/0FGpNbi+C4UiDOd+scOiLDsSDUHq/YKVpV9oU4qAMA6xliR
6TBXDLoCu2bX3bznOm3JzWnKkP+z7mi5FWd0NWnbOFr9/19zhcm4GcSNuQi8qhbi
1qPEXrWuiT3xDY2LpnIySdNWcLlR1eITN73Ny9gsT5mFytmW/ol5/85QtOHIngh9
KZzYqpyg9sc4M+G8CoVt0GOq0SWrXBCeOSy4x+huCmOMvCcOU+xCtHMZ9SCsJ3js
X7H9mfZrRjU9PTJWYOdHEHd5w/ULyP9I58lGxVJJClD4tX4qIRLjmV6OBH/Ym+RG
l0P/3n2zY+XutJ9sFoB0R64fn6jU+DMMNVoZx9Dcp4KQx2DacjAxGyh2anCKWaWD
ofrdtl72DPJyN2BS3bnxMHK5ATEj8IwsIoQ72Ii05lOxYSkUFOTNkF2lmkzshopb
V2dasRlgZ4+JrX37O7nND5dRl/LNVbAgms5bNG0y6lCW6LjOkkS2J3kPEV+/TuEr
eGg2jBse8OZhcwlmBKcOMb5tLHWS6sTCibJ3olrwdhlbOCa1D8P6Wr3JMVspNLbA
ksglhd4vTqCQUS1+BkECANz/CFOkn/nn/Ua8oGD77o7gU4ziaZgXKKVUq4+LL1Dq
0XZoo8AbXXJ77s9S7dvMrQ9IL2QikiDuYtKrN/s7cVfgDRqG3oMOLDKkAD9U748L
Ui/2nIW3p/V0d3X5qO1YZyoB0pJcvP08fz7qxbA1YTOU8fFk0pXKyTNr7KOiDdmG
ah5vYPa1C4oLdK1PKjns1hYLl2uoixkNVmNT2/agOXnp0YWsrn0JxNv55JPdTmfv
uHivSuapwbR1xktrFRY/9VtlA/l4CVzC1tV8BQfs1Q94drhXlKu5PXFPPWKWuOuE
qzOTdGE4Jx/rbNXVPjRr6XKlURvQ3Psh8aucma4l+8lb6U1DR+tLSMi2JaVoTJlJ
MK4VrGG4fMzGfabZ4tjgE/KFIeeQfObnSnOvtP1N2HtYEY2FfC7FcTyGdKXGkB+v
PFAQm1LkCsOzVqv4GvRyNA4VOwsM3uUCjYyiL/BUbu1moOCMcVqztg0kdtpqs4aM
Z2AHBY1o5jYsNQbdSqZuGQfQzhUbpL9NiTZB8YU/r2RBs8Zx1DBkjhVT102lxG+m
6NprIbAyBI8EJUtO5AY+xS0wvvp0FNEFYqYexfW3uMxYCozUDnnz/Rk6Fkk1G41g
YSLeiKcp8TdSAiqeF3Q5w6yD8MWfYN4jQt5SQyjrsZaV6FuYwTv5CkI951bKmCv1
8FKchsmdvj5bSOVnLI5Puv1Gg120ODbOqpD5b3H+w5zY71zhRcaTzneXwGYEJ+Ti
xkFh3VJBjQEkF5nXe5kVrS74k7GhWUP/VnR5myXHc8Dl05VQcYZcezbxbvFF81rR
LnuQAVzGjL6JhXuGVJyuIf4ugQbwNSE/q4Wde/7NGLxqXI8snncUM5g4+wRPs+h5
X5Sn21twx3QlzVAMUsdUeuMAgbPhhgQnbcGaeEyUz+273kagKE49UMx3vFiUTXBN
mGlJFQXdGjugUycRmj8Vs4gDIIc1VjJEEKQleEhy9IYH2/nnWSmFO9APrdoeRi+t
DDz23RghRMfw5mgF1lZ0bPFE3z+xvgUbhyyj8iBaFvtuu12UzihRIzNm06X7T8sn
yDbWxR+FnFNW6bKSjmC4zslYEq0EzbbMlu5Il0OBBFfJP8icN7U3jwCiTONR8YRg
bxfKVkDipUlFJ7MEP79MW8YO5o5A1WJ+zNOV6RNmiV6iRoWTbYli3TQ8J//SkAC3
FYyyHWJTSSeuClE54bZZsYqT9BQggnhKZWIduBXajjj8Kt+jBRzV747AC4k2Q4WT
pvWuRE9X7uPzYqPMbStJJAdIPP52e+o1XnkmMQN92KgmGNgz/31FgpjyI45WQydV
6TRGhZBVDopIlNyFYRMZm3f+taeypwD5mQo8MqHmfWbjVLa0drSULdqMcZwhOmmo
kqt1Nc8D8RxTDp1qFYdtnE3aS4nWzNN7SqYVTFIcK7kgaMrAgC5dgtbUnxhGzG8e
+MnmNdJFCrLuFZmVxWHCyjYyzFQTkBlJhuV8heOjr0duXSvUL+Xib7lF+IkhCG2S
7joZDy687ndBuOmpW9rKaak70tMyIepRWiP539z3ahVLMnqk9ulp3Y5vwubk74pi
94GFVCMwT4whRErIkb6wxxia2Ggt9+ExoO9FPJdTnr5hLCJBnEBkzFGHIPWT1++d
P9p1fuTfTCkH+3KcjBSQJcvzQVAXea4yPxwAm+dXaKxBJ/4dWmrXeVaMnRgLNH4C
lF9XO6EOSI0Q3rE2erG+2gIJE5bQOrUPMmbhOh6Ow4t7RQlb69Lf0rb2I7wHW/3G
c23kEIrAs94yyDxqRTsu+8Pp7HnS83Xj8lZ30Dz0txERMar9oILctl5BAk330rNQ
akwVlrE3OosKsmXw+n/O/+OzQpEQpWkVL5gNliVGKICx32cznh3Yhitt29+ZQX0A
bZ4nwSOGFcJ+7a94TB3P0eeBDBacBIWaJDZszrTD1BaWI0SnrfxI7Q6RBHuXQKfU
lYlabhxP7QfVD0uaBUAng0Kka7NGk0tf/GSR4MoR0GwjzuqBGT5sLdaFGLnzmPIH
vo6EDwkF8OZ2+XKfQpD+3YhoSrsRhPbOzwzFZQVUxkrcEt6rEafQ3oTFgX/iN9L0
JEGc0jWpwlCFiAYLrOpF29Pgcf7+C94iGexI0b53OVvo/+Zscl0JxlGQLX7J7SwF
x145mWI9vpKukA/Cs/3moRw/2v9zoxPMg2ls4MMVY2pDBEkZVoY8Bn5x7sFVnfT4
nAbFI9fumdTRO1DdTa5Kyy0s+dA9xqJQ2yeAChPIyHzb6AY3JJbDnc5cZcCl9f5H
jqVzxOU26ks4g7jpdfhrEKScxpwCq2bLCjD+M0rSO2ArtHkdIf/UMFCtlcFsitdV
C0gPOjXk+9a66EY23jjZg9fGWSbP30PLuR0yOfGHXSWpUOIYU1uEr2D6cHwzAJZw
690hZ5Ln1tBFXG1CfXbUBw2X8u1+HYrEnAg/7ZZruH+DfUKaw8U2BrND7PwmCDVp
K2nasXc6SjgI0sP3WOshOCd+loZBU3wbvH8y36kf/CaLeadz6vyRaBMKGN58Hf4X
1kFFnqJIz734PScGJtRIhiQzXFNUdgOwSSBQ0RdLm7wzNG3X1wxnh92X1yKpWy97
sUO18Ad0Lccgo/9CHROsW+/h+aD5+mvcYHgcTd00eucpTnjXRM1ILewKEg0BgLK4
2ALqqpN+hbenR0Jn43H7xGzXhjw4jnsqe7l/7AwlaNBfHGYBV3yY7cxDDp6aD9qf
73L1QBunkKIcskz5HXUi6JJQ1P29WG0uizhNW2f8kr4kZdxE18r0SdqEI29w1cAd
DmLmGVcDIQfmkxdC/nLg9eBpuZZpgLaU4nurMJirC3edvQCv62cQhU5xtP9HXQ+9
JGXQcaaLz1OJvTnRSxZl1cUosvhqFos69OicYM1fh5mPbbd0W/R0FadOE1Ypty5T
vl154i0R2QAMMd0HLqn6Aq801jbG4zF1rRpCC4J0/pL13cHznUMHTueKHxjyIEkg
FzZrB/qNLSeKAMoFXmqYodIeOIrYBQDxjks6F9Qge9zpnWNrRZ3O+kGwdfqPK4Jh
UIKEeI4WfrIHNHVYFWAc2EA9Z6hVfSAa6D7Hu0DhwFC4aftgy/NTelvrlZaGQDKh
A9RlRjwpEvyWBnF0c4+jtTsTbK1MhDmvSSI04guqJoLQ8ZoVXNG1K98WbrMZe4o3
1Tn9Mj4g1BiRfl5SV7trCuPfAcK6QDJxxcXMN9rd/iVNjYLOIu0oqQ1mgvVo921V
FiHtyMAZLDf9dyjs70amczvNxmSu2Kk5xsl3xQjhKFmOHgYV9cNsZs7GE8N59+wJ
E2fUUqZSVweCte+I8tyH5GzOkE5yxT0qwR48iqlM0sOAmIDVb+OvKsXYdbZ9zEZx
6iFvAihRNsSAiogyMZp/wPK8CR+1uArNoQBWHalV1hYzEm3w3Qdv4Qbcrgnivs/L
ogY3HysuJZts9ITG+0zcaSV6Okz+vG7UJdbf+Pn6QobAflbkVOWKMZV+ZNbJDFkz
6TPDZbaeAtTscuosPgOiqXzPdUA2bzoAgWSycdQNy66Uuz5l7p5aFUPtWqEIZ+vt
/XkkYlKeUHLsscJBR/yICMRPoMVGibSHYFICzRrl1YGoUDDA3EdGbmLPRTOuLs+M
S+6Sm0533DXH16JHpw/P7aY4H3ABmykCnZ9hqFbc1BWGgmiYNObrzu9r/66GFqNJ
LPGZdLIr48d/kwoiUM5GFHLaqJQzYDrglWmBwd0+Ppgxfz7yYH/BYvbaJNo+rYeC
YwCU8shxCRd3LTaIUBp4IOr6a+v4Rfox6Mcro5gYu3hGzC1SZWBmPVTI/BmdmsI/
7aj6N+i8FjFcY8EVu935ERES5LRKSQ0ZB6HdmgrOwcLeZhA3Lz7C3jYEH7C5Eh1K
oddARpZ9PRkI/jI22SDpN1UfBwRTejL+95abbBSdTZC5/Vh2/D94kzYn23ra7P4R
xjH4PfQXY5Fc7mxGClujbPWoocQLkZhe92aRihLKu+x+8kJQUijkODY4WuY5qqAn
AN35o/jHu5225Y37LRZ8HOM59iZm6+5Yhq7pC60vIz4jfGLFKcwfRcLeSWWgQMbf
NS1yJDea7n0FDzQ1QEs3wFjUAXUrL9BWDsB4bhXSkcVOSvM9GF4fMNFDZoyVXsJj
FhkKr6qeG6ynC8kJR0PRaQIBPXhd+r8bnrX1CUAv8XTPcIhZuEeGfi6SDbJy9kkL
z3use1awLNpL3XADTH/djY0lNfaLB3aJbo2i3L5YTS8a2yIOgsFNEr0sBeuQQDhA
wiEbM46TK365SO4ZFwCIrdjSCXKnqhDo8RrU75fRlHv9TZkstTmR1AesGCjHBsnl
7S1G5wm+ERI5wt641UWuBS0SjT85C7mQkUt9BhFAvIZ4g9ftUxpfT6MD7BewjDK6
k/N24hJTzCBZwQbkS4Hw4mG7BbS4e8i/ObpqXF0dGD+hu8AwUrHoX6syFlYPEwm5
y5eMlsHV4QXv+OIDTayzcn1aHJ71r61HZnixu1OaECcyzcVx3LNOpuMCulVOnUq5
ey/+tk1ocNkbETHgJFjzLYvxF2DHg1BqBQCoHciBgViJltjfoQHgbXvxpwMCwrf3
wuq2OsPpx49yQbwbzTf+32Uqpg0b9aAhroNhbENEIBkiEZFf11flnYnl0VinEGab
qrXOxRULC1HW9OI1oGCMANzmJjYaORACb9Qy8lMfr8Cv1PPFq6OKcNuD8bl7bTQ0
A3rif3oxVvQ2a9xYlNOdY9zCc40C0ASMAz1ZWVQ5kOckSgTkErUOTvwoytSQhgLA
KSX981AUwvjys+6EC1F+rCRX4z5wdu8FrBylEwoT3OKhMyCzbq0bXbfnUlbnKIIs
Er+uAoGkrhuwyJUR8jp1VXTlHCcRHaXyh6xHyWzKtDoFBOauZnoiCSGr0oymV/7B
oiFe8OvrrK9agUldXolZnsn59rwqdoEjFsOqjWBqdpw8h1+T1WRvLWHlVvXGiSde
RWTmuncfuwIv1IhBWsmAKrdRIqj+gpl3tHzlHZr0i5d2YB9AEi0FtiTyB88Dn658
l7tPWqqonqfzwJIZJCAG7nCGjwf/c8veuEOM+cXtbegn0CLxF7FipBMd2EVcd1N8
9F9Xwc7/c868halUwpoimRJGu2Txfd4/GX1rB8h28yKns0wJ1TPPQspfeJnqGFok
oJHd63G1+kpLVtIR1fFVx8zpKOjG/U/Mqj2HlgvW5hQ6xOatufy9PxPDDhHdl6Vr
7zFqg4HLT+AXq6yIQ6V9ifzhXN6DoVvkPnMXq0RLcAtYAQMhN/AI9KCLI6fQyAGD
qUrUnd4BONPks5hogjtCKan3R49ZGcaT85b+35bRvuxwprcmEhOui2a/6TTB1ihN
if6ohA800r9rFWGK8F2kzAcaIW8PmRRB6RwJ4eg/CUifMAQSErGhXMmHQCarYdyh
+SaPV+Nl8d7/pNHB6Yy7YgpWcgH2UAeFYs7Xi3yxT8YoOLreIycTTAJHBScyLbvD
bvXLZiYr5MSJQj4T+Fyn9h+1TYUaOmdIATI6TUcEiHoP7JysnXhY2OkW7ybUYqKk
ab/yghRto1cBZ8q0R7VP2a7iprUccmI/y11s6MR2iIjndNGGU6DrPvX4JUAq5Ayb
O021Z72l2WsBSxqiJsPT3wDhCN9d1ccqME8gwNV+kwwMZSDdWVYzZX31zVgvETr+
ETb46E5bIR7Tn/Xnz/8wYW9vnQOqasYLQKBwCaYdY7HOyZF9/pH8Yy6JiRD7pdTF
JE18q6tISnXps6oNPqwLVdtZ0kAez+f8JaxXyLWxki08ZuNF6M2YaRO1ynGMfEJF
F6lsD/abWrPV6noLkyideS9r87J4P3i1DlycLiBZyJI2NUG+5mq4Up9gkflioChS
izBL8d4Gak+sNIG9PSejAQhSiNfztwioc3r+egE2YRtG3+++MronLwac9t/fswiK
WiBlVUttjlPDAboZd2RrA4IAcrDBLo9/CcT+gBs9RfDVg3awAYg0ikDtyVF64og9
BiF41caEiBye9xxvPjMIT11ibPTCXw6o0V5e2ExZX9bV3Y6biHQb8Tp++i7wjdyi
ECQ97T9Cp2R+djiT0lOS9OCTWv7G2nLwd+vJFy/Q//XXHuVONwD/4qSfBl2JTIiO
t5h8griHxiFkQlBNCS8jKTA04crA80LUDRAhKiSmBSLPQlROHziZH3AxyOxzHQyQ
iIFInQNU/yjf6LbeLi5bWHeRSSfCVkrMf0GxtbgDC6T+W66rm2XX+j+FDqMoXUyP
hgtISl8XVZhbqONbypNkc66rKGlkr5B1mDUuUd3YpTxyrFwCsuqA+/S5iQohgFzi
M8hp58MM4Ymgu3A3aBUx+ZZYJGBLpQaYlqgUfUKuY8FO9ASbmtn0jT2G2436J9aV
JPZ50K/cbm1mDVN6jWfBNnFdDrrOSpfpLwl8SkEMcXAD3OsncCug2SJgQkpTy4lm
PcgDdeXloqcrP8Hj3HflF29IByDFYFj2ZtX486lCEcbCvXfztGU3iExuGprmnvQK
1tiLOsgEAydfCjAxhRYRjJds2wr3myukyd9YLfxkcorlXmNOTL3M5FUNo5HxBWNG
cm+qe5FUJryGj0nuXizBrs1TngmWdxAy0fu1PwhssirGklDcnb/38xsZEG4BVeEJ
DbcGBbsnU+d1oqHY2OlSYmSBsaYXCgiDDQqmTYKnRtnE5ZjtyAW6Gubs4oMAby+8
ezrfaD/Uhg1DfhHh5w8btFme8KB5c543celAFjIlWW0XA0cj3jqBB+01XGvkcweO
mT1++B4bP2l9EXFI1ZFFdP2SUH/OcR2JZHMdOv2n/B2tWpnJCFS2dOIunyxJk+Qt
GmuhkQBi4NfvQ5g4RDP1K/4gJjJ9JbPsDnAHPly5LG57U6bMEbO9fkS6SWRGGm7B
osEg3+CYqIlTPeaSY3Za0c6o9zflEAJ8LrmuLMmO3STPpsS1IvmjcDQ7Qnr2nrzW
gPQj3vIQIcNTicmscAGZy8ANNYLsLgmQ7sJfXZjQ4BPXLIYYQiCT4Tbs36HD3q7J
sb/zRX17Itb4Mpz6cJbef8bqXOinERnWlPPbAvlh0LF/kyhXdjEnl0aXHJkDHrwe
xRPvcfR8/Hp0uHVgWFJVRuW3xblprMWf+IYSkM9zru6YXAZpZC8ycYex8eaZLB+9
jrerXTI+xxrft+tgxCSlSjDg5yD8BEUhiclBDYTUDzPz1w3cr+0Yodg8g50iVLd9
k/h8cnAM1EIGN+u7Ib+48jFrxrbDMplOfFVhDK/2dP1m0qxxgjeBX8xQDppIR0iT
ygNQpZCVuWHToMKD2MTOBQH5NUqshQXMFVIy8lJxTWV3VRgqMFhxSNDXMKRBm73q
+S3eLSbCXpdipyH9EUF85omcD4QKVuthUq1fp95j1VURbmfAaavQyn9PTnxSa1L9
9OMgeqduW5kiWbldCyFmN6QF9/cpbYa8o+o7QOIStxUGN7Y0BRvxWNjNV9mBlCoe
m377iYtK5uTHsBsBc49YlNunZstrinks0yvuvKEvPmQbc1ZL1UQAGLPYnr2VtByo
VVfHGRBjO5VLfxSlcZqkd8MLdrWT04f+Tm4zmO6CjSp8lEmVYWcMBnzZJ21+YZRV
XdVtHg/Z5BuQDyTxdm0YHLkrYse2VUUOiTgSNCbqjPzvFH+gkRZj5DNuUy/8+fdP
MwIW6fNIfyRlX4O7lfPm69LjxZ8ykQLZokprvzDczo5ywsVQPiBNeD0bp9ObtZVp
GIZ+nw8Xaxu9GmvNdlKUcq735Yogd4DmldItmqpu+Km4S9cJOU1KuNxhtpgGm8lq
GzDR0vuxqB25u1GDfBeVkAPbjKoeFi0KSWVIuuPNjF/eCYODi+G5wEAg+mL6r1o6
7rwIwVJujw2Lx8Qfg2WhlSEv5Mf316doJLhA9GYbCYpsKXA3FYtBTAHOy4+IDaMe
HVE93RGKuJTf5/NJdXQePASd+hbAKIjhSj0PeqOZOT63vgxDg1JKh3cOnKRogVRo
Aq4c3xkdeMSCa0ESYqyl1FtnSga6oCnoQEvPF8rdWIzZcr0VKP7fJ8gGOV8cKyUa
MW10VNVsT1jWgkXjgG5lCVd2VSxKatwjA1jdbGEZexk2MDzHTkdMT52uSMxcqh3e
mC7XfPC43sHOAYyGKGj2pvil5KM2Pa+Ui5hx+adGmzbU/qXPa4BhDY2tOW2cm+b0
jp8qCkY0WElVTZQPWUZikI2DpLtVvqqQm3EBIqEWtIdx2qrSSLjPz9bckCS+WMBy
2IC12u/dhryhlOH0cyjO8gsIDsTUZ/DyDMts64YQbZKVK/jUKmI0lp9KhJcbc0O+
GWJA8adNrwL2lO8c/EcsbhTn5tTvGPBTgeFOnHHDSFQ7Q9Dcfb54oDznoEk6xtXs
l2bcdWGm71h3C05izofUwu89rd+8OJ3wnGUwc170w6XBmiQQLx8U6crv0gGXjVxI
V2cYNE7QZPbZrt7Lyav1qS2We8X2PY6gbJCcfwGs4jsAmByt3Wm9To/DTX91qyYB
6im97ag3+g7u9yxeT2vfa/WC5IhX3+UPWjc2aNGRc/ZfT2/wLNa+/iYbicKumwN7
Pg8oOndG9nFVwQZzNkvw+BPv0rjWV8r5x0ywt7V35CrbRSfkFGFrIq3DHlh7n2yF
wxM9IEh7efCpPqc9U0QkWF02nIWwTnBixTBQuXgxriD8IRE8erLCrGw6HvEAdM8S
M8WGqeiet8QZwpOqKJpz4Roqc+zQQJhJF4OxGgNp+yhr1psvGSfi5WoHgC9oLm9w
04KfSbK+lRxc9db7otvzZ78daiUmwkFcQunoQCJTb6GyECGALLUkFEn8Pgtr60EO
wV7i8oqEfaACGCxw1xKKP5Zm/0Mwv0jcTLpV22FIom3Y8d/mXLabr+pSc9Lvjvoi
GkiJbIs2NXdOi4SVjZm1pCF6845OG/OxVIxHrBviXntfZ7WtpM5raCSiuJWj5w1Z
j3PDQsa9fy2VIkfu3/2JnrTqENEK0cHVpuj/QOMyfpg9coTz3DPqM0LL47gi+UAy
ATgeHYMXsk3ez8KboSV+hBmCZLh5czdqufVqgVzbKAdESOlUoxRLxewbcfE2bJ+2
ul7VNbXU8e3EZk5N/KBnsFEpk/XcJuvvd2m/l/LMtpSaq5oMzbHxpI2bXlXlIAtm
QNgfCoYDzOkMtE7jakNp9aPOwJJ4lgm+r7yMXSAeIJ5L/5gTzrM9KPO7GItk+rAD
dgkDYS2fXvjfA0qKwlq8d8eIfGLIkvQMaOL1G6G4MRNvo3HwNiuHDpLn6zaOOwZ3
hUYgNqXZI56RSGVeeoWVed8ezq5kXqj9urMOur8W0GGBKo2/eGlqWvTQExZeYoLz
vS4bgcKePdI9np+T+KDNMkbUgmWbubvfK8GX7ZTKALv8q6UEG6FIlC3sPfixotXX
SfdBLjMB/hqV7hnSJGaURw5180FBY9zn4SWGhKNnAg1dBdcTLMdNkVadhFWQZlgr
nhBIaiZ9Sdhrf4OSFcfq/WFDcHdca5m1LdqurYbnFkJBI/VqtAW1sfwhl/M9GnPk
4U/0X96V+jsc/LX+0hBKFjEFj7uzE3CzJXWZZ8pw2PICfnGbDCaAHT9QtgB9wTpN
qFfcqDHQl+2NDCDWudFHx1y/xayM5zDUvUq53EYP3Q0WCx1P7ffADGmBZcMzZzww
7Hqyz/R2D2OlO6BmgiqjMTKBBn4bH+KZQGe5CNafof9x84qceL+Ilb5ypnANTXyq
MuuDv/BResIetIxDZIJsBHkaCEyhxgUaf5hc4x9kXMdMcyOFCHC+qJrA7VUlfmP0
3jqBG0UJtfo4eN8JQb2hrQH7720KyBAdSZMOOFeNaCGf2FcFW0QmIHhYFRD2BEqZ
rK+Hq00M6iCzAroVEfeUt7lvtfSJUUL6MmSbXsXf/HZMqkcKwJrLSjVHFGyojtk/
MlREaUMOCJntmjL8xY42DmPZcSqTk7fvOveFXX/gf3qHKjR3ZbBF0Q9E7WOp4a2W
sgK8W9A+RE4M2R98ciFDizqRPhv3fzOupl7B4/SeWNRZopLksabcvkGfX45cwBUO
/mU1vKlNbTPr9JEJNMPgNuMfeElVkrgGNOQz01OqtpqJkcolEseD6Rti9BX4Z8U7
Q+X3k1WkYn2fjXSGRsFoNHfNLVN3YnEoWD4r1WLsd3afeDzdGjFcRWeV7PW+YocT
cKAPKZs98Vjtz1jxHLVdenmnA+/UWvkculvRx4BJ3XnDt+e6HKjKi2/gX7uXh1qz
4/Wgg18iC8J2QBSlg4LU+S7L83/eSvFCldP4pnvH9CYYZI+IYhQEENM70lrKo/Wh
4XUPtUGbLkA0iOeYdL9dD6BWEVBb51nVvU9ZMrM/ufyXVSCSRMwZbPc7rCKp//LQ
NWMf8h5KbpE6SNtr0z8JPuMo2gKKu9rdxMfn/T80BEbITkLK3GJvlsdjYhcrfAb5
CLgL0zwcgqWYaaoCy1pm9PN/kHAkq0gjzYZAfn/tn7SpkImbSv9XaRggVTqQZPU6
+hmD3sk2ujaj4+tDgB4JWe9LvOMDWUDJLkDfU9t8SPFXYsyH4Z8KBsAQ9X/4IprS
EcI/I5R0QxUfX+88Idv8W0lysWq8cl1RPrR7qKgntn+nuDx/hWXzDCZbfwA7qkEg
CBwfOEH262BwJNjjea/JkYQ3daSh4L6MPjaHPX7+mOIxNIzygwC/GOH9+598/oJm
edptwxoT5lfcxRzqP3ntJ8P/oYKaIq99dW7azDnQorBrHIg1I2fC/QnbQsFBr2MU
YIA5w/sHSAFs3I7yk8ClIipFMxtMiMMi59QvN09SHt3TCYTOlDwOthH1mWax4K83
YP4JCfrT8tAhpAWH/TpyoXphOY+pJgIZY2/6a0bkUkUReEtC778keoddpUtnFY9b
W0WPldetLfZrNNsSCj8hFd60AOHgAy6On4nWzeIlbY8UlO6xmNkkAm+8u8Tn5aCR
gaq40HZtvntXgg/Th5+uaO8kfH2R8r4nJ1bYqA3SYhpjuU3uQgYzzdO9/L8kIYR6
ClQhVyG46PJfzEDzZXTcfNnb2b2gwVo0aNHABrPmyyh0lQhPhcsS3ZG/j0HNwVq/
GLKNrM58jqXOHkf67V6VNDyJA6jRzIk9Ne55AZT50TNnv8JECqJRBqerF9gVFMe5
ob6xfx2s3jh2hiYb27wucUgf3Cn9KnkZFybBemqTsVIr6KveV+NvXpSQHzktRvy4
8pII8P+B+cAWFoiUeCe0n5biIrb/FuwxDh1QarfQuLetHah5IottfyZFI03Jb91/
b0e6N/NcHjDX1zneLFVkCGpWxEtpFaCGsly2auWBycdlXaFEVBTvGRhoDZ5jStMM
BA46R/QEqcHCd7qKcucbsBWixPhwEZ5wu2E4vJDO7+tOrTZsQMGo/PHLp71FSAyC
5rcO6Jpb+XB79ySj7cy4XmRV95E6EO8mSj7iAwljX5AhfxPDDj5pJlCiedM4Syib
0kRRiauQg9/zLuszfmZPFzbD+SJgXnQ644LuHpwrjDGgYtAaonCxP/IYcx+YqGhf
tVFZLAM/WtioBH1rNrfyARUjCns+WenIfeMXEzbd2Z9LyhapTKgiJk31JwwLwcqK
BNmk0We78WuRrVNpwSISDeTpB56uHvv8NqMYO05NonEDQ+JuP8Jw+waQlWijypLE
yHNUu3xh3ytsY5wYzh6559xUSzUV81tGpDnLW8T208Zcod3Y1mQgiDZEMTolUSMg
Jzdy36e0I+Pf3Wfct/8N+mipxT2yK06lBlEUG4HFB+HA6THCi2piS9fNNeLj/oPC
rPO/UPZ2mOjvvlL7w7yAc4OTkCTGPepBMENUecSxs+YRdD15Lx/4ax41kKE6JBgx
xExuT+jNAYsCRJ+I47Lj8W0cZqL8W2K6+/LGFkG83wx6ygj8qtirJVVk5cE+3EL/
+TcOiqJqqZg1wyK5tS3gJB9PbE6F7FWAxH83hitekg9Pp76E4rLwh/EUmxWDlc0r
Jt9+wWlL0aG8ZPedhKlJqeDR6nhFF/F40n3kiARvN/SZqjj4Nfa/8YuKDGXmfyEt
OSeEsK7/dMLjF1cn5d+6ehkD9hphXcEoNKcKsTp/+ATU8FAllypPO93mZGg5sj9I
dQ3SVyYmyLatFIFg2uiqYmpr3SqW4TWkx30BDT3KYEHCDsUaXRqO+hD4I5wVw3bV
cwvH8ytuj3IJljTE8i0IScwBA1EgHydZfZpe0IwRdHQGObrxCxraMR8j7mCjgYS6
Du/fnsuCfsDnHr6i1JU7LoShKfBWplYrihUzqZmu/y/XIY1aXdKPdW1JIPqzO0JP
XvC6zp02IkW7s/BYqmfRrZAqDHXxwlDLugWsAE/hWm2LKfxBCg0Tzul7y0tk/c64
sUosMG/m9vUG4fopPn4Fpz7GBxl9+kyxi1QkzTqKvEnij0M74U3ljqWymH1SYNTD
Oo5YG2uRHj8P9LH+hGSiCUDnzV3xLbTZAZBQNLNoIMD4DcWBOo3pFeBARWZTj9HL
yqErtp6Hs414xNWr6VVTWonXHS2/p6rIzlU2coBljotSZWd5lS8TqIjgpVIn0drL
isAqz9AjucnLGYiJmeP0uTIS5+2XajsIarvLU6RPl1iwRvVwDxj3D/s6JqMvMaLz
GF+RYk3faBLMvRfZoQaoFF/d5yUgkK7sh605isKyWHhssYIVUkmX4AGnLiwrXxBa
SxW6oPHtksgq1t7cXrJDljzrxsYv2g6lNCAcd9MMG06R6w5lA5MNt37LbX4ikYbJ
2R1LsXyRtZ8Wvq+Xu20cCvQfLxN4y1M/utlrbSkovNUUPXjQzY7IC4BViaQ/XjC1
NkSzc0U38aRkRSdErfAlGmD9DJDc3lJ5CIZuSNfrkHRL8i/vMh9ABNJOn6ARz+6n
2FH75Aq6y/BCS3TNynjVvk3glorrYOQvBUWHh5FMmRvFJ+7tOpYofK2pq4hnW12w
E75sI1tkaZLQ3KhwJ6b61TF9yIFmPq8zZr906UjCH7GTnsrgvNs1kd86ZhFWLyhb
F+LhodtUxc/3Zl8EkHYX5QDw/58ep7/S6N8mctvScP+jsN57lOX8O4haWLASnTdW
E3FayxAf1mce36FSi/sjI5NhSen2r/DQDhyJmJrlzP2t9SCpupmol7OP4PMkPRsC
VTzFyJguTmaWL1p21Ktg7idCn+fQoSURm+0u2GKP4nRGTtD6rUQz8ioBliGJSW6r
OJ6h+6Su8JA5OOD9A7GnBiPTcHZCS33wzeMroW5qDoBgC5WT0kRdEqpXSbGfRgnm
hpUIvVT+NXxmKPYlZXt2l3KzmM4pZcAR8J/iWWZbO0TZ66E2jgtbILfi+5Np+6k+
+qBgvUo4jPgMRkYK9v7hkNsP4sw8+U+QTnF7+5+TsxQgknETUhEmrA6VpTB8+RVS
MMD1r4ik6VOKTMbY7eitD3D3q+6HnU9ep7ktX530XX9pMO3zCtZoLw/FgmtORLr+
VCig+4/cWJ4+RWqhI86qeAizGk8vNgSICXH6CrJnVJ4ey5xiDcbx6DITbhuvjfDu
8IPx2HwACnQr1vTjnbs9tQz2YdnAgQCz1L8q7+XKmcmkhk1HURNKTuuHNTKBrvL9
iIImO4C8AxxvFhPHrZS87Y4maOiVBIpMbXmtecpmjA2WVWtkAHf5p1rZPBeISvUM
ScyOFv6i2vFr7MWw+lGpWxoobWf0kykj/t4lJIZrOIa6a7OHqZS9go6Rc9G9ais4
rAJBUZOgme8J+VozLJE3pdG8p+FExfIn9R4H4eRSTYPMkepfPr7qPIp1fhNwAM13
hR+oUrg/7AimeM8UPo5YLSqeeyriKGbylWm9A1e5JY66CcmjfGvHQfWSvNjVRmAQ
j9HQ402zfKhw61riYp61Jc7qvXrQbYwicwieEOD/BZGdO1rLdT/tvcXjhU6lL1La
+qYS3Hykz1+gDjAQjoN9tlxKOyOYyN0JwHAhLUH4is9KSIMNWrrGZZwn0GdrxA5p
OnC25V90cf48740yTXkcGRykzMuoyjkj198vRkZGSULbR5O8ZGp73Co+xkXfr6lg
VAAeE29jZrC5q72n/iKbXXcTAdueT53NGXQhiOvTOdHo0hhXzAPypRkdl9DfQmfa
jACEw25NdKsk7opybomW9FKv36SKEJ5o0AgsrvwVPlkvKs9evTa2feS5/XNUe8a+
1q82m7WlS3WTw6GzUCMPOxDkl35wKVHY/mi2WX8OC87hDAODs3bXDdRZpvvl13Uk
rX/tZu81jHQGvWruySIKtz8lp4ADbsln3r5+BKal+GJxZZK49N2/L1PtFC5tSheQ
Q9Aiz4ipVOfb1C+XcWpo7HloP7h4gYIH1VN2zzTjRj6enwJRuxq9hibSR/VfRXkA
Fj8+KN8tNUu4bY7X3rgTdJp/9R6fN/oUfM6NjYo655CiSx/3jhVTCmxE8oj35c7K
M6oLFpekQ9/VrmxGJutNHra3RmgtKfA9cK89c+isFijY74tQH1u8yoeb327yd+Fn
NiT7AUDDh9YDx7QehrhodGNP9CX9Bj7bXjL3D/frGlxz9xPXk1IC8DifGsj4Li3Z
ul/fIjf5eplNfanz+IS6m2m/RXTisQ3r8RzA7yn5+JSi3lVSLj1Hfw6l4TQGTOQj
j/4EoPHczlAASVg63Xm5v46CSmqFqLva2ckfJVGNLktxljGc9f7B9PvGkVelZYC8
6Ebe/oa/yc1I5kcyLAfEoLVXDIuQlz2XkylSzQJ97fYn8k8kPCFcPElb1N09qu1K
8KijIZlYPiTVBYtrUpSwC9+833WKk+w4YluqboI104iDjgAdqHbPTwD1XX/wBbd/
1GJsAGbILcLaz6ZSAek6+0xqx17H4/LMSav8qBawB1Zo6PCOLYffP7Szu+/XVovP
UHbse9sn8aCogMg3BUMXGb8Y7gdw0iclIWRVUCWWNXdzAa6wf8JWj41hT1ps21xv
e8UU3VMrP6XYywneL48dIECjm5rI8WMBWqR7OCgSok0dwXOrvIx94Uz2ALug+peR
6ijy4CONOU08Tvf3I+FwUiakTm43//7m6/b/DLF2jiFCxOGSCDhqXZ7ffCEJe3HR
X1XLde9FL1H6nm678/LqVwgriH6MoF1a+3ojhNVPQkG/mAKq08gR0397zk4mScrC
jArJiaSA/2/6yMhQ0w38dyluXSCqyVCMu1tV7uCZht+ckERszJl88E6XyKmkZ0qm
NSG+tlKw5IlNveRWBrgp4Pa9YRMrUE7I/lmBppIx6pAvjp9s3XPVK/RKHDlvsL6o
S2UPEQUD6gZV/os4nLe00Wx9HMW/stvTjEAOVLiWdzW7waKztebxC3AbZ6eAqRXw
BEciq31HyM5oqRUyr2u8SgtWdnNuCpTmK2XXT6y8Q0e9JA1ChkuOVYMibJlhtP6w
5X6uLjTvoNCbvtydqjZWyc7yK5S5UFD4ebgIgo6EJr87twEDbEEZDp0kmhGDkXiE
y54Rc3ZHt9vgWRdXf9nnN2CG8rIWs0LzftjaBDcx24QtWuwRAJ4VV+mdb7W3T0nJ
mQPvKDiZxm1XiVXhgnh9RliOe+Or7qC0g9cwAk3AZwzvD2ZCq0s6eZxstn4sN9RS
UqE7h8R+zEngMGQxDmCWxgFGz+g7wK9jcB9EAokDC50LN1uX6plnbFd4YLsFmt6l
yV9oc39W7thdUay21eZBDXwzFvylbpctT7tvnEyj0JMteE+l6RVnt3sPCmDOqmx1
X2Y+JohA+R2EISgWvFIN+ltOAiLwgifnxEeUFWc5ZT8HESfK9MtP6Gktmw9qYgHA
LpDN6XfnWtdI4qwrCmG0VGg7M4drz3Xum/N+W/jd2URUEtHzVfyUTQRnLDHxhw5T
+z7nICnVMQJABQ2i2V6IhzMvX/w95PslUpUTfIs8tueidv3Yg/vrlS21u79vwD8E
QIi39sR3FfrIDeFtAztviJ47XULRnSM7UYkuxnEGPxJDSZU3A0q9RusUA8LwyOWH
3g0N1ckAkJhimlF+EdW1x0cPZv8xi0QCsmhg1wjvuOwj2nZBvQZJPbKI3MfizOwh
DWoZ6P8Ta8ccUBFXHOHEug0bbSXhhjm0gUwYsGkXQHz7WR6ZYBBXq+b/Sqn195JF
RKxW+rsq4u7FjxHKZknEpt+l8z8D/XvnIKxlobck8+7tcpbYpi9ps4KgNVTHbok1
gCE1MFpijTXfPjfq4IgXIMZDQozfpDooS5nNleO9Qs8tE5uMqUp/RT7W6sqXVd4l
xerRcdQSUbUSJe3+0MCHKsPA/MVhDHnK6KNVWHMTaUDviKvGflzHjqHOLHFVsZVY
xgiZS/9A9XgP/Jwh05y8yxmd4MKDk6j3cqXGfv3zfKucoF2upZYHkA/DhsI8ONHc
10tGubjs/SUeZpHy3kQqDqhFXdN0VeG8oVUV60H9dFfVbtQlOIPKKVkutS4P532e
pfIFf5B2lg772UUZYzNOPH53MH+mj1a1q6r5QLWq6Yu1DGtvgvOad/aQRXV6Mhef
CHTu/hykHTFZTRTrXFYWV7J+2kFZAmu4wnIJfldv4HdYLGYEDxXhFQemlNEX6lo6
kzRytlGMDotauLKaIfjU1I4wfbWNbmvTdV9NXY1SRJqDtLj+abvyeaZR+/QrQnqg
WKrv5L0pWqjplyhFp8sOg4NAzl23gtWd1IXpn9Vz372KMha5fdzTgw5V+EBJZP4/
pGyxBLoMQzsS2lfV/UBnmWbPo+VfaMQxxHdyId2Xi0lPQGzuwr1cWMheNJtR6w19
60+QZG7ohn7GK4sclF6RtASRPMEnmgToxeFdnsDjQ6uDMlIPrSRZzKiiBfHuKfo4
30XT8fr4W0fXzMbwZPRZpt/RL5LvKVWdKTINTPVOvNly8GBTPRJTNIDgUJl9Hof3
LNNVeXFmMPN2xyWDfn5bn2NJVumDWLLamU9JHaBoSe/qqP+cgoLMnQvZbSCOJm4E
kHK2c/9YA54uq7fxz+0FoPoz7v04oytF+g5bfL65ZdZkM2hc2Azs0I1uPg87hhPU
VRI++oGXoxHoINRNdO15vWKO7pUYFwADtsqMjN6T+F5e9jr1+EFQmo3u4xmF0Lak
A9mBMKFcVKNTg1RW5TmNjU5JzFAi+JtoIMyCPQn8Hnc/UKG9oKZ82zv+buKrJa0B
wP1PedSNseur0wHVvY0gA/eJU8+CBQnWgmJdwySCLlX+wdj1XY6E5AMVrxP9gWro
k1yMIYK/QuFK8X3r8mBK/qa/A5wVBiKVEHUNrqQwWoT1vKWGOEfTCs9X/T7mlLnL
k0L0J3JdSuG0o4/fTnAWI1H6wmF6cWpipEwXLaNFZjxcrR9InS+7e5DwWRkJ216C
yFDtmi82NZ6QyMWuSy+q7d1BgHEFKBAUOJM4yKeLIdj7B7WQCCYMlClQiJy76xpF
HTHScjj+HzCo0DvBES/dICkZGxa9Ca16DeFGYnTnMPKS3rBREju4KXfwhFpXZQTn
ljgDj7SYcAavOjAnLy7/IAf3JlrAExM8jGhvXDNBgi1iUO2DLVIEqcLr/2KW5Esk
CxeTL07bP4OvyQerx9WQ/p5wkqh8kojVst4BFsMG+gYvemRLR2YLhyHKNj4e7yuR
o0llIAoSjb5wWEFa79IeGAO23gElObBuugXRlSa8RgCifQCRAdcKOc6ynXh6XH7k
gXtA+RWoZYJXqrMzi/7YlF5mT0dXg1ZA0m+eEI6Ab7tGcGeS6gpdRxU7zf1hPIbf
UdD6yHJ6DguWKq5+7MIQjkbC7SpxOIapOuOW6BjBojArPAhlfji8ZNHuhjnewV03
2VQC6OeuFu0pghgd0REYOLieBY9YzDNz2CnSEVtXDhCqm1WEnQ7aWt90wVrImrlF
VUkmiIJYNaS7gn+0y8GZv5qeEmnFTeUWQl2MiCqqFVRxCrk+N/GtTrw25wvH5+Qv
72yxqHdS0RIauBAH3pAqxL/rmlxR79FFItruuLwijveACY872r089+8UqvuuC05J
FWohLxiyK8tS8ke4rV2GXA+6NEM1wd/22hq1mf34qzC7xrCvHfIBW+zLIUflL6eD
vsPab9UYY433z985VrMC+ABZz34FpYfJQu40kOrWGdAJLePWYx85jbME9iF2kSL3
EsoRxr1qQ2tQUIP047wmFpig9TmC3QqpIpu5fmm1geXhqMQmrkQdRXrqYypLqPlc
y+Ce2bNw/Em0FHOJ6j3Jbc99a1JrBRMQfPL/69lgu/TpBGkJFX6g3k+qxiEMgjgO
JPsvssNS3xSGOkVFV7dE4m+veDFS02nkCYcsKcjuTHIf6bGwCzQW5e+uiJJJhpcC
u1qRuND0dYG8kbprUXs46ko4KQDJsD8IYPTGAXqJo5uBOe12agtS45v1xLVYwfwD
`pragma protect end_protected
