// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
rDYI3i+PtpgIxQexcYtfQAQkESqE5/wL9pKDogGa9G6e5jyhZUDTcpG8qph+9O78sBp8DbFy6tm0
1RvC9L2DlD1e+7aa/GAh0poJjoj3dB5QBkEgc+0gWpVJSRGHp0COhxV0/QRH+NLBRfNyzvh1puuB
2KK2eS80oAZd57Ksz0R/UXjQGneKxUnuUFBzfknyzgZfHG5wrvOV1TnVTk0V39DSgvC0RcGzzInN
shVE0SUW8XaHiBadoLUosG7qzy/pA28V1ix2GMjzJ8zCDc6zpbhNdD4y+t/IBtx8kqzPJY8t18LN
5+sWcUl13GRxSJbSAKFl0sVuQCD1Jy0RxfbYFQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
sT4X79ZCvvn9awNQnV+YBdia97lLeUUcRVWfyzEdhVs3cZpxOaIyBOCigVvD21RwSlMw9YJ5k5Jo
2Zip17+6X8Pqt7gGy3WlBzfHMdZu5A9wBxtPcTPSfeZCwz0QlkD8nb2nqfaOT+Ljuhse5rNqCHXq
p6QAWDZdvporPkHvHT8TU1joDQmi76Wd8J+AM8xrK6oTri0Y1NQjyTvkBcIinYKmFucJIver8b0o
KMyDMCvexdlA7ntjk3gDxX7uOgQtbQhYbfvS+P+O8x2dRuqtkledLWMUALyaUwsu6jYl6BZvtv6i
6CHL6PVRlvRcmLQrmHHd6vhJfUptLMn1e4pmlrOQ78oZQ927JAdf/v6u/ABkAJA05Vzbr5nNNyXy
gRjeR0Rd1JjIbbe4LEzkTKCI1v5eKhvbswJNXzbUq463G6Wj3B9K/qbluulvqvudVwcNyTDoO+hi
QLsY794L5Ir0lPRVXf5+WaR5wk8VPVZwC+AHgw4roopeMKKHZJflZfsMkL7g3CoDaQvqFP2l1CAO
u4W/PLNdrOOeFQuMdLzVAq9JuQaJu3wdH7nXYthn6TJIhK9V1ayTKRoL2+xv1QaFCE3OaQ6y/eEy
1aZCc9U7wnH0d9FkpvooHkLL7zmGGs4CvsTPLxsThwDDsH5S5OdRKLlFzIphTd8dsR3Z0HBb6iKo
eymQDXhDNwNZg1QYG/UKoDFLH+xsz6EXJGsJ8AfzPOQSHDIzetrTCNF70CezssovlNyijhRL5i7L
defjRpCjAGjIQiM33qnnPWdlbOZtqz130ww6O91go8yxVMcLii3Zl4briIPDSyOz4NkBx84hGmXR
Cl2x4faLTXMF6rZ0DAswXiiDaNFpGgBZ2hvpdcTYhcjm7P8lx82wjCeGtmNIQJjCKf7oBSPsd6jK
pDnlSeBzAnKzXIIPwrz/8QA1bpXieXbd2cCLi6xvWr+lSlgFLwVN6Y0gVUgoCItPX5OLuqNrzP36
PEKGO+St2aAksku43WO3aSbfUtVqkhNZqnb8G2cgZpfj67CVkVxR5UwCDgpxu9b4tHtg6a68s9fI
dkx9o8v6Oj2NTDjhXP0GNONpNUpkublaf73fqRW0lCVd2THxHUTNxxbAxzt+qgcWvobutzEakvX0
+l5mhQaLtFCt1CJ+IOPoIXtoMjEkiDn78lL6vx78sw6g+XCus3oumcMd1ir3qCCSE28o8E19Wcii
dKkK0ZB26Q//5S2WnW0K5Y++WK7nM/MCqT5gbnWg+YqW+yM5+wE5orx4pHazqka4garRNPmQMdUx
myjVr0n7mimTmbDp6ZuYHCLDVCNH5cdsmdaXa2Y9VGv4Sr2ohps6HsDxNYqj0bB9ojSKpneNLOjH
DfsARuBkV6O57ta7PiKImKMoKNepS+oyNcgzLRVrpMQqzS9Pj7r4Zi/rRINq0YGvx7I6106HGXEJ
42eFzQ8oMA0zjwm+6zyeD/Kn6+O/aVgBZkmpXJoJUitGf6o9uMmjG6pIU7X7zJdemZ6JIHqu8LFq
sfoUWQCJ6avBfAr9Fwfc5tgJIAYFaJN3V93OVE9vbY/g0E72ptlUHQwpa/VUuBUztfmVjWOdf2Nx
4G2dTDarOtKfruCn35VIZsFn8MDofCyMjVGLxcrQTf+XWWRzOw5k7e4jnzIsHGQSdmE6WaxaC4t5
a/0GkXjkbTnBKLE0JrigFXAd59hN4FvXjPKFGoFK0zvcAlYJrRq3Q6E9w8rUUqv0NZN75e/q8wZx
Q0C7DBE9M9UdG74oAmHia80j/W3qGF8mmX/hRZXN/n2gqkoItRl3JPF1CwiNjZzq8kMpeCOZwa6p
xcKdJV5SW3VkHAqGo8UDiuUR+NiYRxFGs56bGZ3DNKLxWoGov3oJvVuYJ3GXCz176GOtlD8QkRQ/
x1MAU5s5h+C4v3E1X8IoW5MkEV7R4rVIPSYCwDfBqfuXPXL+1gfMC6DZV9YEmtdQ04qL8RAUMFNP
dZ4ArVBMghN6TPJtqsLO5n4byLLS87P1QoI6XR65b7NS2U5os/FTBcYvroDV5iFKsX+j3saUI74A
IC3/TT3ipcW7uHKlj58R5FxlDuOAgAzcqyFplQFE5ua4KvYqNKqG7B3cfoCv5189/+HcOCRcCoV6
lMDhNtCr5ItWP6JPy1T3k87IZE8zYR9yXEs+bzheYfaRvAwrG39IgbRP6ejAHiUcrPCfLPyvU5ZD
YFLIoN8bCOni5UO8SClgTOoSo6wuDkZZuWwEPB+09sfOviQIrlXpu5VUMhtm280Br7M4sAkvtknZ
/YIqU8WNeXyfh3GgZNH1H9uXR3/eLWqzWJGckiJqNhPkzQ7sMxhwWfrvYIWYiOpab1urwv5vFV+Y
gJPhq0vXtD0e7+Pz2o4GGXCZaRjrF5CHw2vzk/vg2Ipd6GmC+qR6Cvy1uvki2/R1loNZ/JWtBMbT
kdVrdvfKovQZzKyFNJtNv1c+Ox7XzaRue4yEy7g/bSidy/pkFFbwky9GRO6cG72vLtfKgS166xaM
d7smUZlSLDzCdxxINkBPGopGiG+GC4GSuWoBnofwOhGKRPB280hLRywgtzp3GZqYqPfqRukFy4FF
DJ7ZIme1IgYqJl4MkLMLwK4q+uaQzcQsYNXWG6PbYV255S5YQvUzzPEQ8GnpsZL2s8GKzKc+QmUy
VqGHtBz0x8ZRI5BWSNEngUSJpzrtlD31GQrXVF4XZFbdBY77281R4wN9c+W9PKOLeV4EIH3LhhIc
Y4wTZ8Ti+SFaJfm4sxtHl/a/1KuvfVzUliOVq2rcP8YqCZG6tWXw5sZTp3pDbWRU3EKUC88GqM4A
WIakQQZivnwKXJ2GUoCl7YmgVuJAFzvPlUrHsGrbKQjCN+Kj2aZXeR4LjBY9yfuCV9xBeXTY4wAY
i/DNwVXb/c4G5orfRZIoGBZuI3ftoHuJTtGpq/zx7B+LZVyJV5X6Zsz90o+4HnK6XhVxZgs5rT52
3a01PI7CY8R/hTmCDX1F3aFI/Ymuh2zub11dLG/fPQH1rxWcRBovgiB5fcqmNkMLhjWsEoA4hNum
2LpJ4e/vDQGA+MUlIvYNl40jngtZzEVWe5TYwgK7eeESMMrrlptnf7mKpXWL3h7V++7l1HwHCc6I
cO/mdHI+P2twOJ8wVsW2Ps4adXH+GlvcTxzmw/ZjpHlLeTTYNadzNqKf5+cf4ctGoOKqPLulpi/4
Ul21fWXzEaDTYTMuCkfKDUGdUBNVU0T6WhllkonomI83enjxsSpAzcz6z5ZjJOHJ3W2rsMJXQwfT
np60Rkk7m98PTQDCqESZ+zVbsif159kmDpGMKIaTeKk7C7o0qsh01qTSTSvwZOc4zWkTPFakMp9M
Eg13ecyvtlMmktPufuiqYW83Fv46p4QStLPNSQI2ADlLHiZtEfFY4HVRTBudK4TpLJ1h7v0GKsyR
FF5B/vXN6l8Q2YYQ38YN+xx3PTavFWUw0gLngV3c9dwASVTb26FdBJ5QAOLNVNZ9eyjOYjzOIv1C
w9FMXzRszpE1K816lTNgekJF2WO54GexmwWSRCjgDIQzCJWHy3euvRB23CcV1vjQtX4FJ7ghitwQ
Bn+Uw6kgfsW0GQEWDvuDuNgVjTfCKfAahgRryjxnsa6yQBGpx8FIZYK4CxWfYJb6OhE/G4DMI2N3
Doe4f6JjNoOnvJlraJb3OzzEqYGTQ9FQp97TxgJICr0intxuZ3W16s1pNT3icAR3nQXPmYFdur00
cv311zWFe1Soxfgu7/9mKi/kN249scVyRfJxLiJ/REeHFr8D5Ebyo7H3AvwCfETz9muMM/QA5ICp
BMYUe+vNhg7xkDRH0lhwwhO13Ju9ce0PVO9k+N/RKrAaXaINJLRY32+rWrU1hmR+RUr4taJJWB+H
yJL54psfJ5xAYzWYwgqibwD2QwR547e2hsHzpwdtg2HS2owhl9Zp+9J+QlDznhxRVMxp9UBwYlPe
3hr7vQHcdsfNS5NPGgUtSLghxO5UjVS4JF/YTufK3PQTjdeIf43UfjLlXT5KOKV9cKl+hAqRJggl
DSKW27O4DzdCoIYHURLbBr/PkPu8JghE6LGUFbBHmvfv1+IUjW5bzK5i3ahQ+/EtZeJUReOb9KDf
nZaf2YV9KZgIYomBE7J8+bzGFCC4KpkpQsS5RUsLCERhMK4NgTU+owaodA2wUNQDjV2qLit7g1VH
qhnkny2A7V0b3xjcclmCkSAgoVlWXkm85Nh5oqxH+qDujh3YgA9lmk9VyMPCZr+gjaFvKXaFXYZC
VJUnqhYGGu04kDUcf38DzflhEvig0Dhy6VLLRA50yK7V4vr6M58z3ZEW0FT8GetSAuHo/ehGjDkC
GTLfLV4zPDR8z6q4FEbR01j2bpwhLWvsYpps4MFNudZN0dgJNkDRejaKumzNVs7+RfaWiAxcC/GH
68pTbsxeP08tmmvqqP0lZL3ru+wlDwNznWWDzjG9V2frUcviD7fdnS9GqDWSWTRr3OI8FzG+whD9
Sf1O7zqZcEwQUiTsfWx/tKnTfdxoix8bFVgZNhN3mxtDNkV0BbjjzIK2IythDt4oY52o+5YNF+yb
ceJ08zbniIp9gaSCcbGI9SdLOtd7o5ouh+lOok53NSdkuemsPw/Ily8SLxZVWx0thLeXLWcNR2e+
8Uq35sEjDfnicqbfWSwPfzrWTHHCIJvEM7nHlYRw11i8mW1/FHwcJZQLcyIm9W1HQYUG+dpOPyyb
fxMJACsq1x1yN8LB2P2xq1e99ckszivrg0Y/1u9Zi9s2oFmjSpRuctBtuTWrVZovG3WutrBc0/lr
zxfSTkz6SN/mkUfqpKkLNAPGMs2+bLgAa7fZNJc2fnkTkrl9lxXM9ktX9xd1ZIPHZsQDEbXEcgde
PiUTiDey3qd55uTv9RAM5MANWaKs5ZgDwK4I8mVaI1DSqEuvGNjOQrnCVeBZNhVFIYsfn/DhKvbN
rHF77o6x/Fg+lmlJcQe7lD8L4l/IHIGgpP4FZgQA2iqX+XP51s22MwCSwJsx16K14GTIlf6LnAeN
8QMNLDnOxNhhAFEJvQzqeWBVr409TVHD3WOJicX9/uO35zzBKGwrfkQSKoo+LV3k5vwDDKQt5FBC
5gAE6wtLJBGuBA0fZPhzEwPB0MqvflEpqd0R4TPLtvxeHCmMmNzEa6+MSNZdiZfPy8d/u78wWB0I
h9CKzNdUJvnUUcx2fnENtGbblEwdLxHJIerism29CepxtAgYJ4xYi1LbHYviwjHyRny1Y5ZblV54
9wfvK0+himkz9aoX+4FsUnv+9TJ5JYNZaYuUjyQ3aj7mzoTAZ6y+ktQasTA18tGyTctU/yfCung5
WmP1RSfxqAGCdMjZo59l2ALnpuYlH/oaTFgSxrRDPgEBV+epUs8mCUhMEdLcyav2FHhIDF1/XmvO
dZ1MubQ3XU23CL1n4dqnDFu0twCzOqsuH3o+1+p+wEYdSVqODQvNohwT8+y0VSdW+KvHwbPJbtsX
Nvsjr/TBdsVzTy7JfUG25bOi3Kg5Ss6+1yyZ1r7GEsYF/gP/T9KpltEXQF/wlmPuD36CGRsQ1CA5
p6CjXeDYzmNlqNPu83z0F9gK4u7iAHPSrJMRwVnVuwx57hyM3P6tc14/jknFmLMhmg7OG5BmqWA9
QA2/5tK8E7+ZYveD2Wx5BvrvyiYw9pLmIHwIB3N5F/91+5vJRwVztVIUsMAu5aXxpX3arPouiRuC
s/1oPc3lfThsaePJm5Elg1KxAjkeXUoOLuwauP+OGsYBGcbG8Xu7fL/nETMW4VLqjjgJx285bd4F
Jds/50ZbHLwPjjbkj8AejyzI0MHmOEfNnxJWfEynYxikmgj5PJiSWVT3O1ZLYbiMX5chgVFGKU5x
XIk/Q1ttfQ6Pp75X+xVvksSkAXD/pnZ7ZT0KwFXjFgY11wNx1z/ujCPDyrTkyJ5qpV+jq6ypKFu9
Sb+8yMc36hutYIrvvrdcgM4JXQxJzajENe1swZ9hTRomxcbB2XTWzLek0ysR+q/5GWAohkxy+Nqb
WTLYVa5hGt8jPfcVKrTa70iWAKMOdCfpg6sCTaxlT9YEmINGd78u4SIG8nlvf86YYZSw41wVBK0D
N611JV4uQkyLMLAFbM5HdpxPHSHmzLVSa2IkSDfr6blYq1/j136Ytj75k0bGTU1UsG6LglL0mlEg
/SUEXFdlSRK9ANifzH9pSejkO9vp65RY/LOn+b71CEOy9EVOn3dySBVstIRyPj9GUkO/TPB9xdHX
/P1ccwAdSiwll2wF7C2CwOT1E7uWvrUKDmvlPOCUNgc0DkG0tvyZ+FTWml3bENDc6n5spioE2/Rk
vrIS3j9Wf6GLKUilk6KexvR0FW3B0ZyPGX0mdDcdSqU0/7pg1Lq8VMIY6lbzeogZbUJUJ+fAkAHj
OoHVIz5OgnQQstg10KSoGnSbbWs0We9ZBW+2G7WNzdrxGvvo7zGFVq81z3NJiROR53LkRCHJG49M
Ok0C7UcWSmKWnLrBHU1THOZ0UbDKm3Hw9x0DLEqiScbRi7jBAeorv5YxJfUYYGMBrTGvHgtxOGWA
13MhZjocUzJ6p5jhaEGabIQFiTTK8INky/lEC6DUCwRE+l5iATbFzzD/cVpXWOiRrx4+3nIfG9F0
T7o65qVpWVZ1yaKAoXeBWK4XscZXoajDT9c3iS2015idPbjki9C4Os8DlFNSDhqgF6vbPsbdjJil
5JqFWPGHyTd1YI5eroDoeUp2kr6cI0k0eqPYW4BN1QZgAoZvSlK8chFqoVzJC4NwmOfKnrWLAouG
lsLOiTyBIQh8WTdt8wkwBi0Yd5HS4Wbw1LSPWmbK/pzjI3F9E5ih4OPuE9TxhbO2ZR2dOjGgWsvs
RJBK+UuloerhN5UWBL/jJPEUNg+pkoF/cDw7m747oTcsOhmqdAX4en7csuiTM/txLd07k+BuNI9y
UepTUgOo0lj+jxEkPWdXK9B1NaiHEcCqbrPqdBNzH26FO6ns6arf6K6jHISIeTlCQ1BGwE6mIkGr
3g7eK2NkAC4ap3kj2Tv0iAexTgK2XL/DhIs8nco2R8nmkS3hACbeoBTOYFPQZOgMG+4sPK7pyZ2t
co+g2qNpKOXepvTSCf/Rwsn4pEQ5mOO2A3oV5meZ2f0qfgfBOoUPKKoHujDqUth2xQR8vRJaLJlJ
rguwDUXkoZZHOcPLZcWNN8Qg5gHobenkS3JM6pWZ6xhcb0LotCc/J0rsylpFRtTvreUxEytwSV2A
vs5PmkBd5qLo9tixs5J8VhxVcTeZCf3a+nfiErZaTUKsUbJrRT0kcz2qnAWVIk6iSjv/fq0SQPtJ
5cw2MB4G2E1tlIz5HNad5xljdaFw8aOHSFmgo96q8c2jL0cto9w2UxBcgwh9M0VJE+rGRudhQFdU
7h+zxmhUKLpoGkirvhtxKdyXJcXjD2kMmawGrTWMCe2iC2kb46Ul2Qw/SsAKXjL2ZS9JIWXFR5hc
DYV0fKZnyGxxMFpqdkv+pIM89z0kFWoN7C9uHkH1LTQ646pSZUV9XLAJukRmVtgVAxzs9wNWP+oQ
6cYHBUWkNmH5vhEASmfTzYOBs5UIl7rCe9/cK9zJt5ymuKi6OuJWGuzXueO63/8KEyMDIfKUXCmR
a3rkFb930srFFvo45u1QvYE4pqDSS6Kz0RKy+I7vQm5zFTIsgTNC42Di6lmDFcBndxO8yL97LpgX
NRRMJdLBts2TrTvzgjZs5+5xPAhlrjphsLcEVtarms0nixPfJs4NUWQtRSQB+N+k/rsxnIcnSIWs
ZSIc6hprlrxO9V3WV0HLdnWa89PIiIW0wdwoGcHfiTw7Mu28466Afy7xg1ypha8esR7o3vRIP8G2
s1sNvcir5imNNfayR881jUSMKRpBSos3XCWwUZ/kHbVSSeIyPRuo0+Uqn2wAVga/qJrnMRFMEr6A
tNpNBb23a/g33akvD2G5u6rHJjl6tNCpFWrw+jL4HgmRJyC8nPHd7S+Qt5gBUY52bKpE6Qh+LGI/
TOD1fqfi1qdhD6AQpEF8VRWyZ5jP5qSGGfe8kQvl+7ecIjx5Q8cxHmiVeiZY0h0SKY6wqz9oyY93
7E0w/XoZP6H3nN4QVyDwaoh0bAsGV+wG3/GV1ucRwBC26GMOXuP/UvitpTfTi+zpAfzYxdNG6y68
JXnGcRZYfxMWittrLB9JCM7ruNHdyCaOZBcr/tByTUp0gHbB3WtS1987iS1+uxAKwBr56qr5PsTZ
HPYP+6OKFa8mYbdEvY8dPqJj2V+SOi790OIR+YgzHQ1pvpYZlBx6X5P5WZbeDbHbXiZDegnnjxPs
VYQtNkXRdh9Bz5egFTvEUIZebje67M+FHeD6Q08S9pORNo4ce9I4ocmQdEcVP995H8ddq5Nxp/kZ
RtDkUpvQ8LHbcagatdJppzWZnmIA+wp8vOJrnJruS60onsV4hFgKIlfUfjfEeqoeiMc0bjAGH3YZ
i2CI3baGF2lQUG/4kFngxkHdli+DkMOP9ZQyo6esq9M6QqXJw4BEuPIUtDmY1QGc1+rDGv5Jjn6C
L5EDkPBLz9EYnBx0KGvoQWKfhVuaWnPMxpWq05pwwJOv5tkZbT2h+mNyhZWm9BLjQ9SGNSXGmZpb
c6UQLHq0iaHAWqR6SZ/GXtKamqQjsMfetzmhDzKL75nSOQf0rmE0q72YK1uP89j4DHbVWcb+ayc9
GG73oMRlLdJhbV4zXc8EZm4dYO/wUoneZOs4U7YI6xmr7PaZuTezpELzFYBWkbP9wBhvXD24qsUY
Dcv0UvSWEd+a1QAujtL1+yKA6Hew1eTxky2ch5Pzb5tlkglAQffULjmFJ+7OsfnZTjV19pDgsIzh
Ri7WfsVh46rxhRuNGHuMwhyd6Pt1np1XAdDSbtuoJw5wkat3FNVFskQ8Nc7RToh6Pl/M1R4CENrC
uXeOaHYrtjzI0Oy7veH/qHxg1HwuBLPxiPwUd5Kgk6bKo6QkoRLdAu0v4/7RUJ5ZUa0wNB/NOEZg
hJ36i+QcRIRnkCXrk26HM+BJDfWyJx+h83ZYx0oX0veRvQc38b7NntdHA58ObU1kmp0Fw3iE2xF0
bJgj1X0o/raT0bCwMuw+QzjdAIC6j/qa3jwUTLN0a1KBELkIXnUTvR5GkoN3m5ULqSLBZMbvkOPI
qbMuKbgpkQZVnBO3sVolvNjKhHaKaHgU9hgbceU2llj7l6EHqJHhUnrHMRt4JyIbmlE80RaMQWZN
o5O4/0H3fSuAzvLWwJrrGvpce0q9T9YoD3i3OvUm3jsxcQ4fa+CE5txXkTiYu8qB6mhXIx1FKzzM
JR5RL8oQ9bpjWNn3JwBdLYogy11jIWPiSS9jsnaGr7fbyKJ/qF4an99Ihveg123mqgkAYCrdRa7b
ygF7SSZkTPXyG7Nhixbh8QxTJrkPHlANeWLwOMoZ1LKqGZ3AT1BG9SLfz9nlkuIRbqaXVOdN9WaL
rRrRj1tfSXLWXfN4xyw16i+IN/LYEDz4iBmDmYcokog6sVLqPfRY9yuk4POaz4l77PKII1xAGuQU
p7XOZxcJxswpg8JDHWN9ZOkrd+W/BI7IfAnQ539eXZhUe0aUKLCCS6L9IIr2rTDpjFOZjjMWlond
oVrlwzbtiGvHe9iX3TtxzHQUu/Mz+E4K4DMAVRCBknFFO1W2yWQZ3gtsQUH1/AhO+k+oiUTQ1atT
P4pJgwsfSFSJpb59rAlQsHk1tH0fWuTP2vta1hxLWYFocVuCHj/6bU1JahF+bX81weiVUdhnAijK
+NMS9N4T9D9YZAvt8jB4ZPSfb5Cr4m0c3Jtrzn4OB4gXUh1jjLIvrL+bmAjCngaKKCpIzwjnrpue
1OWw99Dx8764JTuZyEyB8vS/uFgEmh09m/W/Nva4uwpv9OQbeckbT+Cd0dNowlHzdkBUO6ljWk1Z
SOGFKuEQP6GgDiyTW+VRyYQ/Ep0RDTjH6KpFzDW2N8EmDiHNQJlceseTtUf102FdSOVxeI6qCYPs
94xi96JHM6/fLP6xcxNDxNks7NHfedbsr13BwdMN+F8NoSI5smbDVt3BMkl9WbPhJ1y3cGNSdcys
UnNYCM61hNyoZbzQlnQ6AFVC1+jPYSD4guXmd7CXZ/xg64MQx+CiqJsOS9/bmhDbN0M324yd4qv6
l7yuZGxI+HlFgyYNijYWLK4gZq6xGU+Zhakla3MBszeNBSOSZym9GHGPuC0ch4J1bQMVlKPKf2pX
BPAIT7df7cnKrqxq4IAOiGRk60msSlIekXqgl4sDx2Z7PklROUweI4qVINAu2rASgX4Ph8vpi7Xz
VpwgUWIKGFKLFZsBLcHC5cq74sRjxoVKTiXjtOeb5vglC1LDWMmURdyVve/Bknganl8fpIjTlE+Z
5NwqfcnL3JXVGwLdnvoaMDPKJUgtKFkyOvqw/jS/9uGbUwibO3lN90vpsYInMBUx0EiN3n9jy9r6
KhYVgdQjBkBjr60ap7Tn/HCCGUtyox3388yvm1HFHAHqaMjg+9aiGUc4EHRKbueg+FWyzisOrWTt
HYvtwytkqoTmXv6fYwvORZ/bP+2SslbaI9jyeP999pbQu4TEWip+Tbct6YJixcqfyZagQ2Xtfs2H
dwS3tbfJZezhGON7DVoXO0wwP1DBOmbdDLdjlMnpmUdySsStJpAs/ALGGSMke2kPiW2715px+vzL
CvqFGrp9W/MUMXbF2oFvucVORA7MypPY8uhY/9EMpWrgMQepGfEUxwy4ooEOPI0tI18HYQPPbbTA
Z0bogCgoN93ufysiPHqB45osKnqoIl/7YdnsboIfEk5BNQ2RRbKWc05IDS4410PLhCG2hkd//rCD
n3zEbiBpk35tHpoiCtu6ymW0MHpJ2F4mfgBqFDqkW5tLCy8WRo5SmxU+mTs2eq42A9pXGsDs2hIR
wd6gMlARt8V4RuY5NLBfPimAeezIaUmA23XNAQCz64heLhJyJZ9FP8qLrzZDqV8+A7Io8RVsAQc8
H1B/k8qPHHJSEVDYZV268YgI5iSi8VqzUtPKymiKZh4Cc+ErAuk0SL9Lnv24S/76zHaOmyK4xH3F
nHuPQVhEzF/kMfP1m47ZNTwc8D7bypfvW0p/OhNAkKj+8ThosYNJXlVOw1pIkSmyRn6jtjrBLmNb
wB61llJiUOHep2ZtJhSzuqu8q+OQGab30eM6iQQeFxn3hf6qdea/FTGjXnEAH+FLRsIIXovNoVwA
bRnJlWKOgUyZrg98lt3e7j/GkMvw7e+t5KInO2JQLsookbyAZ8r1dkVeMmhoYjv0nLLSYe2vBMJb
H9fp7hQNB3u8LEXdk/hapKmgObdFdkoycUcDWCsPKWwUolQ3+CjvNVYCmY6x0fszAvB188Kdhcrt
OQjubPx4nhLi/cCZj9RlTLme/dW373UY+sDK6HHT5NGBtGCffIMx1OUNZSoqTb9NhNkld3oZWFw7
5wTaKPHnfYxEmxj0upp37DwFDgrsWsakc4XF1TzIIS24Lv9XdARb64i78xzvhp6srvrL6F2P8zEb
0ZsPzbDdgf1F1EE7DYQaYS+/CTB/fjTEec5t/I/1FeS9jPLyiOofmG3ChgCQAFGdpkW/OE/USLBz
N0YzM9QxRMR+obHAhmSvaIs6IjkQLjgRkZTqnjcceIx+IaTK8pmQtD/rS472x0qpAarbDINAtcGP
BfGBytENG5LA8J+WwCMORolLmIMx+0CNpt50ApVA/Zbf8cKom76JlX9wIxXr+NxMnsBQmLPFVqsM
7UTK1s+lFBpy4KvWkdqBSQVSTjbixo0BD2eQXu+kmvIK1GD/244yskjyF+rVv+S9791F8RapTm0U
H8TIMuh4ZCQETpGlmGfOosm9bCmFA6p4U5wv33SFWNgFf3Lu20SBZ3FN2epr
`pragma protect end_protected
