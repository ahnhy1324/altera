library verilog;
use verilog.vl_types.all;
entity clk1hz_vlg_check_tst is
    port(
        clk1            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end clk1hz_vlg_check_tst;
