��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O�k}.Ż���"�����x�u!
�*�*����K�f��\ �<��nFɚ��f�.&V3�t�_z����RZ �UP'���I"���U�ϓЯK�݁/�G�5��#
/���R�|�1{���_����,$Gn���G�M�J]^e��Zd~;Rb��N>@���O:G��o�)��A�ڄN����z=$��TD|d�c")��8��|�N��BK��K<J�a��$������ D��r�>��#�V��dZ|8}�<SN�����Y�{F;y.H�"42�Z`��]b���Dk ���X0Н���	Ԛ�z È�hQ�)F�|X� G�c������Erh�T���.~��z򳥣�w�?��P��!�h�L�%��ׁ΋����+X!4>q��.��_���͠�@�?�?�'b�-��-�m#
�-n��k�h�{1��?�w�K�ZH;y����2)D�U1�l�$���"3ix?S��͢��4����3-d���σ��H/Q{�⪲O�C��F^0�4�j����Z��,�R�M�{�}f��{\����_��d��y�� A�3st��%���Rr�IMs�� ���#t��C�`'������MSI��=��E���)���E�7���>=���c��sv��$�Uqͳ��������R��cV�\%�#�e�u7p(���� ��ڡO]�z[��޸"��7(���#�d�@Xj�L�q�O ���}D��ѯ�uV)���Le/����;��cf{p�+(m�v<���0�L�N<L���Y�r�2�p:Lw,Z���(;..u0+]�Z���K�S��h��V�$���o!�ʂ������� 0X��"߷EV~7M)&�e�T���.���N��\�T�FJy��u���H]ԩ�����S,�ܰ���9�6�����TT����̠��Wq@6c��9��	�ß�:�D���aB+H�-�"���b�V�j衼�!�����@��0��J�D<�>���_Ɠ�ˋ�<bfn�s}��JcA�n곟X�<��G�d��#��h!��<����aW]��_��?��D�K��yRl�V�eR�� ������&��v�R��8��hYy�2n�^�3u>�.�D�Z�ڵ���OMO�#N���1ݵ.P���3������<�t��d�Q)�l��r6��
í1��ֲ�;pOh�J��������:��5ȯܒ����j���
I�f7�ߤ�kD�4�S�WDN *�oMk^�-C��u@����l�C"�6+��i���!�N�d|�LC"�`Ik�I��߀@*��o�|\�`�
��w��y����A��n��<d�!�L��!�`�n��gG��ǚ{���^�M���mD�r@�	�HP�y�H�=���h��Z?c�C�9���;ay�X��}c�<vN�O{��a��i��~Qs���mJL� �������ڔg=51EL*��:�P����J��f�]-_K �@�e�=:�ǌ�{�������A���")\5qx�E&z9_�V�ݾ��O2D�4x~s���&�J@�; 1wzY�v�n�Ҋ�%�A�?�7�݅JÏr�$����ŝ���#>Ɏ�ߣ݊���Eq�GC�%�+"݌Yb��k ����Ȝ;B��y<���dJ�ۿ�!@�_�l��CZ4�?G'֒l��AQ�PEUf?!l��b��!�Φ�h�JG��[�<���Yj��x㑮}�'e�0/�`�M˸9�F�5#Ä�:f�Xrp<�['��+!�tFf�O=pr��3���B�W&`�*;J���&��!��fA�6����l,�]0�>�RJ��Ә���qi�C�Q�
����S�<���_h�=kY�2���>k7�f7�|����4c�7���3%�󬀉g�o��R�.?��|��n�ioHR[�����gz�H+�O�d�y�ȏ���kc��gD"�hņ���7�R�S��x��Z��<>wG!���,+z��m28k#'�|^�y�U�K��ᝎ�]����%�/j���p�t�,�k��X��g =�?��xue\���6U�o�U����P�pB����T�}�G �oN	���H.	�q۱��p�Q��R�p���el�lq��DA�����ڍeM"ߞ��,Z��X
c���������Z�zh�X��R�8�;�R��e �0��=y�	k��v��M��z��$B�'���ėp��j 7��Fۀ���};��s�$M��Mɿ�dZ����Y�3�״��Z0��Re��a��d����#�����郄�{����P��S�G���6��� �"b!=� "a�G*�#��9�<g߫Y-�B�z���x�T�"T�_|EY�~�y/T(�{��-��i��8~�M��\��P���B�³�	���_��y3�g�6��x����23���1���ۦ���z	�lHM_���<c�v�X�����緖�4#	S��P�@��C�mf�(��Y/�ִ��q��P�n���J.k&$�<����k�
H��:F2˰"��hh�� t^����Z�ea�
�H�2^�+�ː��,y6���͎4�l�io�����"�	�74��4���O���x�D�5���À9�T��ᮬGP�fe���7D���IP�о~�]��A ��$
��~�".��*��9�WV�CPlu��@<�t���/Y�t�-�`;�%� ����;�3�7U,��鄑^���<�u&��-iyZ��<nwx��53����%�ME�R�������-����n�0�a�n��0.���Ļx�je�

4�J[`O�x��L�Uʮ�����qW�ְͱ>,�S �enw=���:�a^\��i�K�ވlCVI�d���Y���Ԫ {�M�6@�9�Q�XޙIT,�|'	�׏�Ȍ���g\i����SO�|�t��1����Q���\"�I,��0Ơ�Fi!��������J!��ƛ�sC;Lժ�Z�%����	�z�ĩ��@k�"�e'9�S�L3L��h�%^Ej���oYl�� .�K�.�b���)B����(G)ϖ�g�SM�C�
���y�����8&��7��l0]	d�6B8�/�55_q8��L�n��O	��S�+`O�T�/U�vPf��T�UE{"�P�l"(n�L[���� �dʼ]�?�5�aS1�
� �A���2e8��/a�^W���9���u����P���]�^D�Ï
�������#�S��Lk�[RR�x>b-2_}"��nHG$�7&[1:BoCB����;��Wt��!���2��!�az�NԽ*꙾����D�½?�����[���1
�A�������2�8�����%�J�����|��5����U�z�O>L߿i��Z���0��|�4��+�k�aȃ�?���+b��n��x�ɚl����?Vid.]Z��W��1䫖�a��wm�(]��4q��p	myr��8��Cl>��I:^��g��}�>qO�F�l�6Y���3M�2?����'�}ٲ"j��>��=�a�9=`�Z�8I���v+|��"s�LO�Q����UeQќ4M����*R��_T�s���>�g��a�s�غ;�9Y+����v����ӯN��7v��$��"�(�������f�#�T�l�*-�E�V�FcW{�>�w����c��Ӈ���6�1	��2j
�gK��iC�	�9!�n^+��YF+��>�35V�|���{eƺ,"�0-�2��=ЇI���!�*��(Q�ewna%�;I�7���jDh��J��i���=���P�s����#}Xޏk�]��F����>v�2�/����̐d�m���,��E+����|�$���ڵ7?,$v���M�d(�8ݵ�UD�Ɏ���T�TJ
g|SF|.-���^1�������XO����u�D�#Z��v�I�P�B�*��#﨏��-O*6,�ʠ'�O���rRf��w�-NQ���	��qМVy>��RWs���HD��&�������rܦT_�L�7��87؈˦��p3�#|�9UL�'%�	���E+�7�Bw=��G�%�����cq�LV���-����K��>?P�n�5b�� �	�Į�en:	t4꽇_(���\!2�Ũp8/�wσ��������9!��P�S�,� ���9��ޜ0��b'#5��.���}ϳ�T�{��頌kw]\�झTc�S�2�vA��K)4����z��p�/��\���PYaᣪp�M���u ����p�*�t��/ koE�Hj]��+>���A�S����D$o�M�J9z��V<�;�����bT�祸�d~O�E��޹�{g��Fe��n��
+�=�9(���Je��~�}ʍ;P����@�݋7��G ᒼ5���� ���F���$W�o�V�8Y~`�,��H#)�pϚ�G|��*�"�Xp;�dD8�-����@�}+!�>�1,���u]2؞���8O�_<�#r{g�²���Ou�t��#:{�,y�:�� H�{�%j/�L�J�1��vw�f��.=w`��⨉��m�:�H�9
�s�}��qp1h�Kn!�R����m���C��&�WT�H����6(p��X�Ec�rܹa= �kizm��H�D/6*����"S���А�R��f��m���4xbM~(�T���/Abm�j���B�b���Ơf�"`$h!E��8�m_Yo\���悒-KC�Ug��W�Ъq�a��k<��������U􆡀�ό�Oݑʉ 2�XD�.:�$�vLe��A�7@Z<Fr�b��^�~QԢ�47���� ��T�o}�c�����L,������L���$���L�~9#-�ꑿ���|���f���\$U��*�?N�[��l_9a��=82�P���_.�eZJ�.���sg�Q�$�8����j�����|�ScI����o���/uj�?;ͤR>Ekw(-��ƶ���)8��nD��ݫ9�ݤ��v��<��+�.�!��gI)��K�ǡ�I�8xݖi�v��"�Z<'��1"����;��=&JZ���3w*����t8z��*����U�;��y��e{Tb!���+d>��<@� �`>B����`{�m{��q`�	�e5��߄�g�b(~7@�g�w���C����8�|���f�B�Ҭ���K��B�$Ng��c,[�ڑ1M�g����6+���]q\G{P��*(l�uR���)r4���k�=��$_
d	FfP/����1�t'���`@+1ԘS��w���_(a�pD���E�
�6;r2��#�����eE|$ɺF�s[��vP��_@gY�8����/�{5q�#�\�=J�����Lbb��u��ई����O"�F;����+0y6��ɅX����9�<,��K�:���&�5.�m惼W��q4�o\�����P�$1�}Q�n?�1ػ0��Z�˙����	���Lt�;Q�HDD̕�(�-F���U6?G��'��R�K�A��v�}5�t4֌��c��)�nQ
�);N���ޢ\��Cxө	��r;�x��`*�sŌ�f=�|������%�RDb�����_t\<��E�k����\2��iP,�`���-�q�9�C�x��Ǖ�p3ա)v���`O�G�H�D�-"�$~ ��߁M���O�h�*� zo8"� �u^��YO�'�D]چR? ����Y,!_�����2��?5��?T�(0��#��S�y�#�j���5-�#�:����m��"��$��T�Z����/x�H}��,Z左���1��w��e�a%��^t����+�}�����{q�w�f!=���o���r�FeN�&*�V�,ë�5{@�S�iO	�F�9V�n�#����F5V_z�ڊS����w ����^k=�ͫ�N��%�lwF���-b,>�ީ2�p��P2/S*F�l�o�����`05 hnX�i����b��u��ù`�e�v�f M��H@��h��ơ�	�UK��t9�"uŌD�_<}MR����,�+�m���q��U�?���*��T�(�Z���M�$�{�J2�^2݀;��C� �㕈:8��6��Xq0�\B�p��վ}
`'>�ߺ�����/��;�j,��H����� <��0�=�陣N�!��1'��x�M@��~�Q�c��~�-`\�KV/��z�^���2[���Fr������A]wK�G�<����p�§�"�J�RC��V�I4�jH�>����U�d�� �l+=,R�g^4���gs�_r�bwIP���Ċ h��.Ē�J�\��=]��D���"�%y�q���`��`��KpnF���ìv�ޣ�V�ą��O�Σ�����H����u,^j�z�؁���9�L�S�a]t�����g�J}f�A[�9&f�F�p͏ij:n�d�%]��͇�x��E�������S�0j�j���ג'!��K�X�̏����{�Tgg������cQ��qA��*{�ٕ��V���sG��̍@�h��z�}E���|��9�r�lo%Y��+d�l�J��&���2-'���cMT� :=�	�W� g�Ov����������h�5g�4]���ɭD�W�܁�ƹgs��Zc��]��Vq0�fu@6LoEJ?0t�ޅ$J>niI��Jj)�཈k����] �@�X�1�Vͳ{M�(�w�t�?����<0�~$?k�}d����/���k4���H�Uiw�]"�r]���Q��s�:v}H�,&Yp���� %a��4*6&��^	�d�٫�����]��6]�M3�*U�8���H�q��9������}���df���y-%�/gP�MǴ-V��������v��^G3����h-e=d��mp�B/�r{cx�W��y΂쮅������%���5�ݓ򳐲�N�Õ��������X�˻��i���}����*(�������;�� �h����ڃ�\k��7��`l���Wvv�4�����e��҂�w�ïRy�9���/h.�F� �k�l�xP���Ј~Q���a�2��
l�>{����_q��W�p�-�heܨ%��H��&i)��Y��N/��<��=����T;G琓��ǺN8~��*~'���Z�q��E�BJ�h?t ��j�Z�ѯz!�o��*|�7��y\9�~�(�p)G����W�ë=�$Y�����}%��_F�֢�8�]9���QM@�g���϶'����P����~fJK%�n� ��^:݃y2�	�J�+�efr�]BTVW\LV��l������M���fd�p�s!)�k�w"׺B�y�2�R���o���l�)�.d�mDNh= �;~�3~�o41��Ď��f�kmbf|,���Y�?�Q]+6TC� G�����H��V�|�3��*f���K-%��5X�����^����C5�ڣ��sW8m\�Y��~�ڎr��<i_RMLb\�*�Bs0�'�T�G᎛Yy����vH�=��0r����H!O��֯
����>�j��7Be]뺇�!1��<��B{`�U�#���gsa9��iP�����K�lne�Y����U܀앑��é���ɸ����qDУl�N�� �����R��<<, q-��:~X�h�b}��K����0@Y|(���� ,�P�8]\5q�0Y��$BCj��V{��'����lq��4�P>�K+xk2�*�d�8F�;��nnI���S`��e@��^������yL�w�7A���.K�3$gյ���[$�?`��$�
ǤHDb��r���Y�7fk��M�$I�ƺm����%��my�@O��"+M�z�T�<rZ�U_7񷏴�-.�}�*����ɸL���?
3q
���S�."�ߟ��A<&�$�pa�F�b�24��5��u��n9:[�x��u�(�)�~%����nm�����eX��ӊ9eX^�N����X��m-}��<����c���B��杼j���w��XRy=<�8�K��hI|������`r6@�K���t=
CO���֜�KL� ����pa�E���R'�qÎ�JE��.J݋��n����g0G��@}ͪӜٺ7S䛄�73hCO
�1��i���޿/�4c���ԙ�&e9#׫�`��q�\�y2�h�V�5/g*��F�N_y�@��T��9�&�C�������ڹR;�hv�f��u�=�?tH��h݊+S�%ф���t�*ʺA:�9�L�f�O����N�c;�J�v��x4�^�=:(m�&������!7��O�K?���L3/����p�%$�`���"�:G,l�L�S��U%=*+�K���ɰsr����8��¤��/�ɋQ1�D+w�IX����ߗ݃?,4�W�?�L	1���6׽	�K�����sXDҁ~�2�ã����⃩U�z�m�(:�p[l�lx���\$���sc��X|�E�	2F	A��{S/0�D�Ue�_��v`3raY{7���r%�HPp�����(�.��Q�&o�B�~�����s�+�p���Ay�*g8ql������r�mSM���0��@�j+N��\�kt�BRr?�ǖ
�"�V�T�6]#[W��"��ө���,��$TP|%�N����_5��q:,�!��¯�JCɸ��m)�$M�����m ������3��K�Y�C��,Vz��!�'�N��߯�D'Ƹ-�H�<J�Kh}��P�YV;��`���E@��wǇI���cKG�t��$y�WNK���HL��WQ�HW�,�{z���l�L�҃�����Ui~�l�Ϛ��&�1�%��b��8L�%�8��y6��7�C���χUa�����V T��c�+O�,Df&�
&Њ|tϾܰ�*�����ٹy�}���]I�D�<�A ��ނ:,8ӻ�6E���}'�L����<Ax]}-4��L�7��I�DO��o�f�oX����������LQ$�]{ʿ�N�� ��5�>proϑ"��H%vHDb�	�������ݢ�VO��D���$b���U�م�Avu��~x��:s`&8����T��M��tծ�C�/�n����1c�P����2��ϵ����6�������၇�%���f�P�c�Z�j�J*0��ÍK���B7������(Z�?� -��Fm�)��܍��λ��:�<�������^}ۇ��|>�7(u8�o�y��5]�y�DO;
ZrS���9���M�vhv]�C��!~=��x�#%ḯ�X@�"�pDIj�[���(S_�ZY4T�Pbl;� 9�th��鑭��@រ)�Mo��E��a~�XO�L����]�K���\���ir���zen�
q��Xrf�n�/��-X#�����3I%KI�᫴C�	l���w���^v]_����Z�5A% ��9̊��sn��D�D�E�����t��:>��Ri�b�֤iɑ?�ӏ��S�QZ���!A�ΝT묦HH]�z���N�'��Ɔ`YAߕB]�QY]ai�!�?�4��h`�����* nҊQ�EAau�DA0�����!|08찾����[���Q*ߌ7��R530�Yhv$,�p��wب��-�����S��bv� �$b�/!�c��	-���ԄZv&�U�%XՉ�8�chg�gp*���f�x����3V���X4����LY��cX���'���@�+���x�Gdp����?�Z�Š��Q�׮��&"�hk�CE��S���m�'��1ٍ�b��f5/=��#��<۟v"�5��S�b#?׵x>B���l��J"v�WuNcf �$O,�?sw�U7��Vy��_��Dm8��?�ʳ�򾃲��8}t@��yZ%N!�5�w�����u�ɻ@�P�Rҹ�.�!8�d5�*��(��cs7]sĜ]��{��҂U9��s���J&�R���Ԅ�~�2���
���%�gk�;����� ���Z��.�S�0hY8���2����*�U�3GG�vb�A��߫3�__�%l*K���EB����(�QT�4p�M�`.��k8>7����]�������d'��<��t�'�ZeB��3}U�~�@�v��*�^�0Z�����SN��v9�#����rI�ZlI^��x�~�TS���?�#�_ӎ�p�.�_�
�W���r�_S8s\�T���P�8�x rxB�+h�P��K/j���{e�n��Ǫ�U��0d䈲r�T�e����_#N�S���;`�-�)�c�O��>�mۓ��l�àᵳ�-�� ̢�B�vy��sTHi�`�%�ӆ�.S�"�P$�E��]�����-\��6%���ə�lD��l�F��@�Q��Ҹ����o�3�F��V;�XF\���	i�D��Z�����\���m2:=�B��9����'K4��!��ј���OR�ظ�do[x�|~Ro*�
R��D���.�7!�8�]!���MD�B��iM�:�y�2��\7.n�KJò���%�sC��B��>N@�)'�YF��"�h��s���U���PW�Ƭn��n�P�LUrH���LJ?�%��R�:.�5۵;�E��&�g-o�#�	���ӆ����w�v���l��@���&%y,�����������w��Ƈ0���M�ɑ�����쮪��~��n�4���P��hv>&�� ��V_�"=�=�K�#��w��h�3��,��nF	�E�7s�B�[Ĭ��|8<��|	�&����
�m�'HluX�A�n�n����Y����p�Y�0��`��$g��&�`a���˝�́B-@z�=κ|�b~�S��X��66�S�E�V�T����� щ12��!���ܒ�w�Hhpk��@���L�4������ʦ��0��HŶS� �vT�a�"���II@���fD>�<�Q��?{aFq�PW�� �gڼ�ȵ�H=|�:�%���4ZR��"+ɟt�లU��3�o���bBE��Ґ��@l܂����@w�6��)|�M贻��̎�%ڽKp �'��-���l���hsw9�V���j��/��g�n�l[���ްm�t�.$Y� �<)$�����h؇��/0�`?��?�w��A�>��픧���'���AGܨ)9ݬY'k���� ���X�`�1�t�)���Y2��r ��A�K���5S�tr���Z7�1>|N������u������$�PL4�����r�>�j��Z��/Mv��Ӗ%�@�8?��n��a�*!��e���C�N�4����#tA���C������/7��u)�w���wU�
l��u���:?I����2l� >�^k�A�,����'��+4ltX]�hp�ۅ7���Ʂ>�t���Z��
�P�U��7�붜�E�����h_Y�l��}2�U1�B�O�W��~L�.G�Axܴ�#�<��'[�g,D��,�O�N�|7�S@�W'$C�t)K�$�j!S���[؎����
H�gZeQ�N�s@�(j{B�w^I~j��s~dy�Ȥ_}�����_7 u"�"7[�G���`Բ�l�6WL��zϱ�+�&)m8֍�@�kڮ���k�0O���/����&��z�)4�邷K�>u�"&��J�����Q�Z�����0}���:)�s����kv.!�T����q�(���x.'��WPnq�"[��0��u�eKa�N�>�9�K@'��1Q���;q�Ad;�'��&�I�W�!�֏d��1T�l�b�zVc��O�g�%5;�YPf�i�\s	$��J����c>�>����2�`�O��5b8Vj���@J`�^}��5�nsWǪL!0�=<\�,����S@އB�~u�g��'�Dpg�]���V�����j�߹W�̂�S?8�h��� ��n"H�U�ʉ��U%�����>"\K:@!@w�ы��Í�'���]�a�Z*� �w�*�LؓxY���!�A�����*�n\���%��j��2��MU�k��'Mw\v��c�LlmS�3����B�҇�|�������N�ƒpx���葩����v-=��Ng6c�sP�X�985g���o�`��Jua�㊦ތ(��@���s(l����E��E��x����l�r�����s����}�,��?p`۪�q�-	�ܻW��g�#ˉ�����8l�m/�w�&�Nt����>�~�T��꣼FC��O_��Y� ��R�J\��mS�`TT$���b��j�>ݻ̟A����Z����62�}�+xn�*Z�9/7w%�n��J�Phz���T��xOg�$o�n�1%E@�4re��G�b{7��E�+�p�
��sU��� =!�UNP�A�����L��,>����c߹��g�#6�YFL�������މP7�ة��J/�ן��2����^�������&z�����*͙�S����1�<������Cw.�����+�w!6�������R-mD$�8,Pc��0Xw�}�d�W��=��_�	�+�"nM�&<\��y:V�_��ʕe	t�����RX�~[�5$�m�@~���0űmR�tzXҳq�T��Qd�ux��,�
5�4�n���`�x�REfK�����,ӈ%M����Ʋ�Zb��.���|���+I�ܷ.5B/�̟���1��@#�khZ��"�i1e�+O�[AE&`��z��US�ݱ[�^Vh��X+�t��J���ٰ���)v4q�ʑ��J�m�ZYV�����f㴫�kŚ����y�SMU𶎶�3�)��bW�v��w�$���>�����;�JiL�9��dR��v�,���zoOԞ�c�I���_H��Js���=O��|Ɩ�i��gb�^��'���.�����^�NZ2� ��Y0K�Ѫ�%���ppD���eH�D��p���I
6�n*�����s�dw�_M5���BL��S�C�����n�q��5o���<dR���Q�i�-��O��M��C��Ͱ��)��I��Mgc�tƱ~m�qu�xn�0Ok��^�a;{8�:��BnE-���E��N�V�P	�&#~�CT���T�u,�1)��~�ξ�P�
<s�+_��[I���^	+�[8���x�-���MB�=�g�m>a�z�d5�"���n���"Fz#��L4��ly�7��E��އ�j/��|Br/'۪o�]�K@N�"�e7�|Q-�M�����{[>�|{�Z�CH,��l�?���엚��0��pv$.r�ٳ��JE0�"Zi���eH#K�#'��ㆇ�_Fk��2���N3҅tw{S��t��Xۃ��|
���GR��@��և�$,}jb�/֩`���g��Sb��J�\&9��<U ���o��QS�[�o�.}L|������9]�]Ů��#����h��=~���k����'k��oCpY���=�8�� ��n�6�i)2g}Nt���A���i�_nNW��_|�	��j\Lv)�IyVN?��r�ik����9��M�7T���c��������d'Q��-��%\�q��|A�js5�&=��y�W�F~�o���C��|JS�U�Z~�<������id�9"�B�崋�t�F8�j78Z���h�h�
�I�#2�z�I]-�x�-�(���<y����l��xҡ1����͏[.j������^8v��=�Ŧ_IW3C�w64D��k���_��I��5��/k^����Iݺ�~kyB����l�;��P��I���v~��LH$g�3�0����Z<*������O˓��h$��+�lѳ�0��Qz`r�>���8TM��h��o���y6�$����N�AŢ�I=��u��Ɋ.�$��-^돸G���#Mp��2@+2N��tݏ���O�����w&N� ��,�Ҭ��
�Ks$z۬��8�d_L�.WzB?��������=j�Eڇ��+���u4�� � G�M #R��"�I�����+#���ך~��4���x���mE퉌�߇VBv�p*�R�f�,��*��g�5@���C�5��H�2G��<@�-�,�Q��G�/��\�֙.IPz�y�R��P�ܸ�hm`Z��r����[�^��u�"fj)K���p�yf�o�9��X�6���U F�<�uB-�,B�{ۋS+�����chYOz���vA�0��R'0��c��	=��f�p��A+�%;�"��Uy�l
5�c����mg=G�	��`��y��cQ��u|�@?;<�Kn�&�VwݭEm�~���]�,�z����UYY`�Ӡ-~�2��j�9{�:>�'��0&ٱ��%zF<[�}�Hx����&Q��R�h���c�sjO$Fv)�#X#]�vç�9�?�NK��T��A��ޝ=_�+a�1�|�=k��@,�q�M�u��`�E}ĥnt�e�BVѐ.�ok��i�l�ͤ'�{���T|l��ak�1]�����U&��Z��i�x/#���7;˃ZA���'�7m�Ky�WkڎT/��o�K�2W�F1l�m��^52�(�x�����.])d�Q�cNڰnI}	l�q��;�+���3��u6�/�x"��d`ع��|#�1�7��* ]o��@�j]�`ZWE�5�Y�0%!����V����Z HP''B�e�A�}�o�?k��)�%��� ���

��5p�����*r	�u�1���/�9�5[�D]���N�*k"K�z���H9��>���%�����l�|-�<����r<=�tZ3X�L��k�0��$�^tB�dp���:a�?/���|9u(��ȵ�y�Aϒ�rݒ�gi��i�\d`��b�
��OΞ<��ł&CwY�`]��� ���n0un����(��ݢ�֭�K�5��/�X8�u��Yn�%�q�Ft2r�zG6�5�$��{�}�ci�j�Ǽ5N��{�𭍟~4ii�B�5i	l��@����OE�<��������7
L8�HG)=)>����w���J�2G6��0Z���B�Æ�+�{˵��:��m�څqd���H��'���k��� ���i�Ԑ�%����f��~q�m�	>y>Z%z���t@<�|��!��(	BWy��Ȩ�Q~����.�u�fW�6��d����e���ݰ�N�#�[N0�/l0�\k	٬���� �+x��O���,���MCh"���on)dT�ë`z���s*�;����M�5ś��s��[����<�1���o��$	�,�v�'�q����ıO����������3�Vqig	�D�G����Bz�'�Uj2(�'��W��[��Ƒ�MGF�&L���<-b��h!(��|�3���yż�]c������+Nu���o|Q���,��%��{:��1p��"!���F�P�wӸ�k�4����;vK���j��P�es�}S1���dl��$2;`��Y�.O���;J�0p���^ٻ��f*�6��}������8�D"S�ؒY9�/�/e���_�M�<JD�^��X��;�h��0!�=��,�7Hg���>L��L��$��.p��1�%�IQ�v6W?��9�/iI�`�;��R�T�F3R��e{��l%��tvXv�C��z<LH4����]N���˯�2I�vd$EY���&�u�<��ޓ������0��%#듔�<�# ��I.����r7P���\�v�{�� �/��L��
�+���H�=��ʢ-�7JE��쬂���H�٢ے�Xh��n�DJD��)D�"���p$f��k�V,:�����\��>�^p!��]�)cZ3]b#�d�AJ�,\�wɓ�x �&����L��{�A����J��Xu�k��b�$I��y=�+T&��IN�v[����?�';s��)��p����و�@
<�F4�,����M.?������߷��L�,��@x;���T6�v�w��G�Ņ�AJT�]|r�I�2��"JO#R�(��f�ZTTE��j�Z�'.zOG}7��nܪ���	�,�A�ǰ�	��� j,�x!�y��[7 �iIY�РTw���Ά_�¬6	��B	
)�	����,{f�ʫ�xG5��;��V�y�uT�@h&��2ȲzWAVJ��t�2,��'�6RGOB��
�CnU�(�pQ�D�^������R�aq'����Uڴh����#�8tea�:����.�;����E��0B�"���z�Ÿ"Z�������~�y;��_�B��\��F$U���6�@:��-p�.m�Ӣ� ��QE%�Sz�,��B3�V%��O�͠@;/����Uv�U�?����zjaB
�����w>���%���i&��8�YϤ"����0����/K&Q���tZlO���V�p^�vL&Ô}�~��
N��'�p���/s��B_��-�H������1#,�6���؝��ov��c���Dw�{����z�@��&���@:ɓn'/ѧ.�����.J.��$��D��ʹ���-^J��~����Ns3�9i�O#��
n)q,���~rТ�R!����'��TԄ{���8Ⱥ�Y�=�+�#5�&ڭ�K_�o�����duvA�Wg�R�~��ڠ��,]��ρ�����zO8n{A�4a��B"CC_�j����݇=���H�w�jY�}G�x$#�.v�����e�����j�$$�U�������lE�O8����iU���;&T�U�F96�fc�p��sI�ć�P'����呮���t/�ܺ�<�����p�T�8�Љ�t��r�t��;� �iM������2�伪C��O�]�p�qƙ%"�~EF���Th�,�K��{�y�0k�Ve8�*y� 3�0"�	9�B�@}�*@�)���\ҵ�Y��]�so|n(GG~!�����H�䎐��~Un�h��ձR�V���;D�E���3�fޖ8����K?�:`��;¶������/@���<]��)��
ɓͣE�0Qj��o_�*\t˥IO�Ki曅`B�[����3<P�.���]�TDɥG����\{H5���kd�C��w_�R���@��7ʜjP�qׂ����W:�8e��` ��>����Y�c}'�ػ�%��O�iշ����ǰ;M	�ԧ�������d|�z��w�96��_��Ph�hĎ�\�#𓚱�4�	n@��f��$m�#�b��=�]�y)�����Y��Yg?6\�����p/�PN�)y�o"��Z�P��_�K�bO�-Ɋ?���I3�NlS��qā�8qz���kK%�5� �W�o�39�1�!*
���ўXӧs�b�$7f�A2>{L4�}v��҅|qO����3,,���;��e�U�3�}݀���׮�$�+��WZ���:eη`R�=���MV�!Qv	ů�@�_������/0jef��Wv���V�k��U��>Z�ڜ���'`p[��o'pɘ,�=x�H�D��k1��fy�5�ҝ�ł�'���%}|�E wh���x	v�[8ݢ�ϹG�����M�9,F�R�В�7�c����e�9J����xB���0�iDf�pq����A�'8k3"���Ј��Y>&�d�ю˴Ԁi�g'���`�@��MI��.���`�SJ}Z4DH=��$U��`��3{��d��a�^,�_��)ԡ 1E(k���(��o_�-mԔ�l�(JU���A4��-|��f�R�Y��~�*�'���1�p����Snqf 0	z� ��/�r�P���1;S?�XFmW��δ���_cq=D�� ��4ޯiQ���p��`_(��k1۽]��~w�-�����[r@C�[�T��W����%[md�H3�_�ӦqoAI�}��n�S4��"#��4�RD�#�i�g��U���D��eX�[w��aQ*,	�1^Eve4;�.�JҐ
��G�?� �ֱQ�[��琄�;��X kw�(b�5�j�"�N7�_�Q&,n�3��?\7:��֎�w?�-8}����n���/�H+�<�A�"p�I�����>�M���Z�Y�V����>��Ή������]sjy���d�����[�wz8���YC���Ҩn�����L��Qdb3k_��*Y]�'�)ԗ��nS��(�����4��)<�RW�"5�t<�gb�����kf�@C�/�Q{lu�*� \�r��
g�T�Rg��c�<>��Y�W,���gIa��ef��y��g#�_��b����ޒ����Z�Z��q�dG����;�\󔛿|�pd��)l���LE'tgZ�OV,-��3��3��]�י�&r�i�Ĭ��m�E��
��G=��6 �h�u?��M�C�t����mG5������=/�Y�x��$|��i��Z��d{���{�"8q��I�:��^"D�(�62���Fb��r�(!+@�*ZE!A�I�R�X]��E�)J坎�Β��>:�"��x����l�໦���=�+1�CP爿V=-g\��#�o�ψ�Y��~Q�������5��݄m��-�$��4�u�a���*\��8&�
*�7�Ru��hjݕ�.��&5�?��~c|��5(2��V��1I�#�C=��� H�aݩ̽Ruz<���5���0�eׂP�(Pe��e�% �Թ�W;�}m_+#k��ox^���G��N!�b��-����N5ٶX<2�b#P�(�7 r�w� �k��}+GҸ��(��y�b� m]��i3ˤ���g!�_1����MOG*u<�ZD��~gQ�+/_cn�q�[9��Q�]IS�`7���t1;����c�L���]�DF�,�I��A.ި�v	��h�.	���s�bC��'h��=��k�<$��z2X���!��'�1oʿ咅]� jE �ĒD����A���z�-��ѯ3���E��C�mF[�;�r�!�W3Z@y����4��DlN�����9�0;�N_a�`�\S��^,^��<��HX��t�蠌�ưz�}=P���2]�;�l�V~����?���ǧ���B����Q�-��.���* �� Ǯ�<����F���Ӌ��~����+���/�R)$U��Փ�Z��;���?O6
���CX��b��
�
�?||����^O�8��ic�y��d�tUX�˷~e�R@_��H���E: h���4���h�zޯqDV��I�,�	RQ�W	����2�ڪ?g�[gLQ�,qڟ/���a����}��m�F������(��E������!�`ʘ�{�δ���3u�@�V��$�� :�.Ln��B��(��EF9M�a�p����O�d��#^�c�A�=��Th�::|'݅MɄ��j��2�1D��@:bc�QGkSz�e�#&M�j��am�N�a���\���G�3��BB��$q�	۳34��O� � �#���B��LA*�ܶt���2>e���Y�����0���YDF���B�+��ooc|�%m�H:�����#���� �/��r��aq��z���|d�Fa¼0=D����1^��f:Ν����A#��H!	tIyY�G9���Xz^�y���~�9�=kI��Qp�&��'�ޞ��q ��J��X0t[|��:K�>
zB��ڗ;;��J�IrHF��:����,�7Z��!��c!`��-�B������9�)ky�����>ْ/�r��#����0m�����6ObR��ʣ�}ԬdKďi�`��z����1�0�4U)�ǈ�L�b>�St�.��DW�ڦ�$�,IF7fh/e�s�9���Obk�-]�����t���&�x�\��P����.ڵ�2ݠ���Sڂ܃�:�����_�.�M0G��j�0��1ح�VTU�`�7�pOp+��Q�+W�B
�ޟ�� �� ᝂk��s_P�{�������9��R�ZDzYσ(Z�r��ʘ���ͨUgE���ߙ`y^�t��m�
}Y��,�8��Y!��Ȃ�{^{-�y1�5�/�h8�9J�6
1��bE�v�~�ܚ�[Q>��5���j��4��Z�%�"V��A%��JF�:�X��=J��cEAeϙ%��t�~�a��ֶ}�u�(}�v=G��_��܄�o����h�5�5���S��hk(� J�_�K�B��0��g��PԘ1+o`�-È�嚸��9MAr�Z�����)�h�s[jO�[pl����j���`L;��c�'�Wn��&1������B#8�����-��Q	p��#�1�>�ɵ��˱�\>��1 �ɼ����R&�t�pA�tHDDJ��m�
�H��cY�20<G��[�,�y�����Vm.����=��vD-_�wtE-�`r��V�sC��3��q�W������&��!,$���ѽf�I�D�$hf-=�8$�)�]_?j�u��:M���CϤPͯ8;��\pM�>�U�	v�w(z;�+UV�	H�ҹ!,R���;i��+Vm�}Ī$ �QB��*๓�R�e?����C�H	>Sb6�c�O"�&-9T�i�/V)�^kذf��Am�=x@��dsz��M��H�ᾂu*�p�Ɖ��JCFv���EP5Ȱ���׮�B\����_^�:�+����U0�? ��s�V�_�Q���J��_OG����Ѷ+�����]?0CN+��O��O����%�DM�H!o��9rB��ShZ�Gڽ�+�x�L�J��O5�C?�����B��щ14K��9f����6׾r+�cN1��0����B���K�)4S��ZVUm+NY��gU��+1��-���&G�,�e*��c \�Q�]��k������.D\���͙�!�Wh:�>�*����ᣩb����)�������o��*A�nKR�:J�2;�iF���vz�:��pn�y���d�7������P֓��޾��������[mČ�]�S����?���b䌼���1j(5�^K�;`t�GO������5�=Zh�ռ*��q1�ַM����(,3�q�\ϩ:`?6�G1��=�5ǵ��X�E��@��]�@Ve�@=�So���Yà��p���wiY��d)��'@�2,]�^ +<�:������?��2A*5_��}+��2Ȋv���?���Y�X�8<�tF����b�:��P$e�ʙ��ǡ���6���)�Q���Y��zE
Q���@F�I�P�&4�s���d����,)	��Lv���d�M��r�[cQX�|`��H~������Ӹh��޶ȑZ�5I�55Ƅ�5�V�\g��d��д�^��1���BɊ�d4��S�5�'�r=+JH4�-u*�^&�'yKe�^��d);�Qj�M���
J���u�K���ews;'��mDm��
�RPC/�U�;�W�n*_�M��[��!�����,��oB��~ʭ���~Α��u��{sT�N��Wz�9�������z��B��J��NX�2���f�)Q��1�@<A@Jib#r�1��S �`T�t��G�@�X��/�n>��^�{�r�K'!Q������{�v7��e��[����� ~��_�eߴ!N��9{K��q������
��<��0�
��3)���4L�6�P�HB�X@┘i)4�lӂGٖw�p��*�����>A>9��N�Pni~�V&�c��)�Ϙ�xs����dﾆ��MMR�]�`=Q��.h�7;�^3r
���W.����k�}ﹴ��13��L�_�:�#j�O�Yʟ����ͯq���O@�~��ym���_~rx�� �&���PW�/ãi���l�U�B[�j�K��U�a��a^[y���c�����˘�:���:��9�n"5&𦧱�Ȇ�]���y��S���G�.q����' ��$��W�K����b�Vȧ~gB�chSv��/�ˆ�����X�-� #;��o<���6����&u���r��\.�H~7j˂?�T1�x$��K͕�eK�"#�b��K�m29;�zy�pzJtn�l`�ۿ/�j�.��|X[ 
܇�>Dp%(�U$�`�F~��ܲ���R&zR{i�>4�����PlR�*����,3F*G%�
����
I}�z;�{�U*��4�2����	�a�ZB�M� %��I��?�ƥ��|S_�,��� QY8�K�c%D S�9^77=�;O�>��B��`�8�X�G�^����#0b�Vs���ۃ��_[E�wۄ���`]�0fL�HlStԴs@2�v	��6Pi��^�I�+B��ga���h�ajɺ�Sm�Z��1��m�&����ȿ#.�`�ԅx�"#��
s����u
ϘYwl6[�|���)���2$�`>�G C�Bsh\T�fl!#�'P�<�p����l��ij~<9�����{@E����igbE���]���^Ƿ�w��9�:_���n�������uJ�xM�Þ_���KHA���w ���`)��/f��ڨ<㡉��'��h��D\�J�m���;�[��
{`Y�h��C$D5���ɛ�F�g��(c~��ڄ�=�'lj��^t�v�9p�H�T�L,Ή��xǗw*N%��s�1,��Ÿ[<IC�H�Yᶰ"�#gij[|U�\�ی/�iGi[� ��dq���W���+#_�#�A1� xf�7N�w%�� '&��i#E�P,����T5��e}c#@pV�
���A�!;�So�:�P}�1��=ϼm�7W�����q�#gWd��{�G����W���R�Q��!
������iҗ�~NZ��	��Ǳsa�X+�/�+Yf@���h�g���G7�O]�54���.��Q�V�9y�7*@/���g�BuG�E��$ �n\��>�)>���2[l�O;�)���E1��#�B�cUF����8�y$tR��9I�����zd����Nh�R���(V�$�>72���u7�
�^�^f3���S�� �30P/���O��;��X@�/��9,;���Z4�d�mKf�>���u��3L��ƕ1��n7]����<��:�,��1�8f��( S֙;��F���˘Hi�v;�(�A�'ױ�%�#<lZ/!�v>e�7B-�J�%%o2̦cx+�Eoֺ�aٱ^�'F�qx�W_-��Y�!���`F.T� ��p�G�Q��q]FD��ݶ�P ���yF?� ;����S��Պ�7L��[�i���#�D�)n���W/\�2'x欼&����l�6:'^��|�%HvY����ޢ!P�����R�6r���7�Ա�k��Y�)�[?8��,u�O!��}ݑ����{���g�h��F�9cX��m�[]������>�̯N�����Si,�F#��+Ia֟��������xi��&�ǪX/M�W`��$~vJ�������K����!���:=�-^�ܡ͔;R9X�>��	�O�G��_�4v�;�1�W�O.���Yϳv}ϰ���.��q�j.� z�]VP�������c:�V��Q��z
s���� z���/Q-��&y��V��J7���_�� �#�Si�x�_�Ţ���Cѡ�}��[����I�Lqߘ��	�2�����F�k`�H��M���T��VE��
�ڭ*r�VKߥ����}�!9X�D,(���+��Ћo�\��$EG֕LEu�s��ygQ���އ�H���	�������{@),�H�R4���C
G0�'��OV�捱�M�#��T#�|%��d�Eu�)q/2����-�+v��[`*�Ƿ� ���f�ɦ�����}M�m�S��[��0��Z�Q'��|*ػֵlX��2��>��X����7i�tg��n(���.�QG�H���$�7y�y�
��>��x�PW�b���7<Z��p���5-DT�n�^I���k>M���9��w[�ú�v�?���@�O��{_6�2�f��:`c6�a�>\��K�6��$ĥx.Z��[�g#��;<�p��(�i݅����~��ǌ�� �C��C\���:ڴ�
��'�(�;�V�Ywk�m�u� ��#&XكF�
���X�g�x%�А����	z�q���la��>��
"*�*�'@��e���(�3�����F`�{/�U�����
�QW�3��*`�D����x�3�5�W(#+�Q!�䢰V��'�}6悲����N���:���I4�=_�Eʹ��B��E��P�v����OXc�HG$���k��DeP��E�Պ�棉���9C��e��-�r{°L>���k[E�[Fh���Q�m|rN@}�q�O�V@l �����s#��$�ް5��ɧM�O�Pej�w��U4V��~��3�5�O>�, y��8�(���pe���J�"uc0�(���|�Z?��A��co�&iTo%�>��H��v������D��Ӌ���5�R��T.��
�#Ps�ST�2��ri�^�k������EO[}P�h�W�m��B�84����iݢ$оai�By=wN�N��g�G.Z�Qf�L@o��8�e����*��h��V~�^�R�օ�yC)�茵eA�2
������.9[QD)��M,�Z�m/�>4�J�����3��9�;�1��7�H��h~�´<�Fw�0��1诽�5>��$~��F��L�e�6��*���A���K^W5b%'>�w��`��烠)�-��뭐IgodNݮG����;@ҶN�S�����;,υ{F��E�I�E#�2�bUJִY(N����
c:����׌�~'�r6��Q Y��(Ͷܵ�f6L�'�0 ��0�� �d,s$`�����MHo��Crx+W�o�D�,�&�/ [I�QN������!7�n'������b��g�e/ۢ�V�<��0�W;;��c?%N�Z��ii��;N�mm����ץ<�/<q1��ܟ��Uʜ�p�Ӳ�Z5vp�p �~� �O-�RV&'g�&���*�[*��/(A��a弅
+�\T����NIxm���+��e\9�h1��N(r�R�n&�������$]����
��I�{a�15��as�0�`�fn;��H$	��������>��F��ÿ�Kb�YP� |+Oq���H��<��HI��g����S��H�#v:S���VZ��]ԑ����K���4��c�U�>nH*%o��h�=� h[s�M���c_H,m}GxaI8\������|���:
T�߮ǎ�B��*;�Gn�)M����O���R�(g��bF)��͞��g�[�&4�ѭ�Sw	F�$��&dz�Z*�Z�z�עpv^�+M�6��f� �Mm�O�>�Oj�j���M5�ȸ�%9/>�{��O�7lϹB���9��{�;�R�x?Siء�?�0bNG�9ey#�l_�s��5�t�r�lG�e7j�uxR���:?mZ�VD�M�`,6m�W1�o���t\�Ͽ��io���P�Xx��_cT��P<�����ȼ1���>�^*�0���@ڱ�������A�2s�;��$5��M��	�]C�Y��v\~ި\���)���ʷO��VWFV����A�_�R�jJ�+����`�gв��������r�X�*�����%!�G_�*)��8��e_�#�Q)�O���-����}�D ���PͪO����*�'��]�!�J�p*�u@�sf�P�(�:�������s�
��Y�
��:��qMa�t�6�����B��j!w0����Q�����"����+ﰮ�)�Y����{qfKپp��D;��L
-���6b���/7��z�9>���"�4���gD��E��:����M�W>�C�����ڞ,��\����\���?�v[��v�6�~u�G	��~���p����>�د�c825w���o�!Ku����K�2)��s4\�Oʻ�)�"#G��" 	;b��E#g�� I�%5+�{gУ#e�dr� "���s@bCo,���mꍅ�OJ&�-u$ �-�1������/��nI^�������U�<6�7I��|�Y,LD�=U��7q_����Gw�h�e���>��2M �Nd�`��j�v3ޣ�+�F!t�k�?���+���5^"wR��߿�&���s���R����ș��:�8��j�d/C�	"!ȵC���B"!Q�,Ζ �i{�x㩬	�>��_7��<��B\&
Ț_0� �����D����s�k9���%q�|w)G>���N��ع�|\�}m�=�Ґ��8�7�?l|G}V�}�3q[O��3���^��B��p-J��pժc���U��
�q}���0n���������B��X���k@,Հ����wB2�Z����L�*ѥ����]��'"-(����x�.�ڮ��RH���o�$���N�\ �HK�����L�x`�8����󬠾.-�'�����@��r�/*�pYљ�M�ܖ�@�G����R�,@��O��Um���)�xR5�!�؉�4�@)�+rDn�Ҟo_G_�X`��n����3@�#�}X:U���8H��+�]����Q���y���̢�Y�:Ә偠5W�F�<-�܌�Ѕʦ���,y+=.: �@|�6[�����z�w��*��1uA����?�*����"[�')�5���.. ���\��j3rIf��>�����$x)��4��\ R\VD���N�C&N��}�����(g+�g��֔����+.I4����õQ���wV�i��ָIgi�dՎCV�E��	����h�E�d�U�q�n�W9�v]Z��l�\z�@�:������IO2�ق6�%Q����$V����B���PS5�����_tS6ߙ������0S��^��7ޭ�-�����)�'c�hί�Xh<X�֬㇞��k�"J���Q�U\�5] O�0D�I��7�22w��$,�Z�h���J)��!5�n���0Coǹ�s�&K�
�Z<�S����q���9�<�(����
�o��YR`�Wn�2�����[6E��3��9��,f�j�-~����$*%��j�����m��,���g
(ުA��O��rWq�����+��ψ�8�~7"�u]3�}n��9���������5��2И;�/��?�D�^�t��17�T:�Ŷc�T��7��{a ����&4��Qu�z�����`�,�����@/�r��B����E�v~��0�Z�>�o���_��0�7�)n�u��2�U�:��r���@(�����R�Src�&��&ݚǗ�Qv�z�,�Qjeq�~�T��؇�"�He�x!�[�s�1�Բ�ӄE�}M��M2��{�\m��5��п+|ڲ��.�����b5Q��L�6I��O��Hʝ2R�7�/`�jٚ_y';�)��'J���OY�;��}� ���KN�����W��p�������)0�w7g��Ly�k����}����;S�?�#oSe8�����"@��L�<[��:��SO��+T��Ż�o:����-J��chw/F5~���2$�ϩ�Q*q-�]wCĺ�Xq���R\��I$��%ߨ��zn碎�?�:G����oj��^.�|'��
�#+/��񂻮���I���h�������"xw� p��w;T.�6�ﬤ(�;kW��z�MX)=걚BfQ���T��d�2�K�OO��Nr��{d1���C�G�%�������� �F��M�2���U�	ZR�fW}�����1�˲93vn��G�$�����!�SI�8|@�xk2�.�R��O"4Ɉ�:��Т�Av�t��k:����jy[+@ہ��1��Ԉ˵��̴Ѻn��������h�b������R�կ���>�-����§��x�W�|��uR�=�(>�.G�������챱g��utJԦŐ��=��$�/\��ck�����d��ە[�19�y�F0��"���d,x3�g.h��p!zs��V����D�qt���^�Q��7���f%��=�Ǭ�!���}|���)�wJ��������[j�tځ��4��ݙ�e� ��<V��5�B5FoW���0/f	���r�워���� ���z9�b�����S�C��?_��W\
Nx��E���r���B%��ΑLڀ���2�P�[
��s�����ܤI�ci�+�u]Ǜ��rBa`���k��Z�c�<)h����:�۝	YXn&�|�.�����v�80�A¸DV�7<]pu�Nn"|��a*6J#�kHM�͵b�e��ijFl��s*��v�O�	��F�7�ʠ��/d�0�����li���?������Fd˺Cb� ����+ֺJ�|KӄhcYf�3��_�f4���r�9ru�-�`������M�:,R٨�#!���c�b�R�@G4���e0|>���n��ώ�gd�z�H@��,�������f\[�F�h��g{۠�8R����`=[�!<�^���[տ�7���S��5v�1���I������M�}F�eXb��P�_��<[,�!g��V�� �>;(kJ�a��� ����3�b�V4�4ؼ�|7��I@P�c
B�>f��_�[��a���P��8S�����Y��y��I�uC�4�V�I���UJ��e�L���Ҋ)j礭�u07�V�w�����FM�AK�~4� �����T!}����ݰ�I�A�IXH�K�$e�����H$�9��{a�rcqܗ�����_���W�:���>G�#��'�5��s�q4 �����Z�)�A8�:X�>�n�a�� ݡ���k,\��(�-���m0�����8����Z9�<�"��jr�A,����;~�aLuHT�y��k���ɩ���B��ɐ��0U��sR��������5��v��|n���-���S�����L ?q3�f lR��+��~�[!a�sM�)�s%����}�2W)�����2����M|���������۟~��muL'��*'�����	,��Ł?c�Z8{7�)D��z��)0!�A�E���)�m�n�v�9���b�)��.R���`���n�E�gR;��ǚ��_���ߌ b�_��Ͳ�/����V
��G��Q����J�{�<���=*4�ʑ�O�_r���i�^)��� �-jF�l �j"3�I�U���0�#V6�ʛ�J�q�pӒ��1 i���j�!���5~��ӈy�]<�O\�*_D^-��s�8� Bɓ�͟�0�u:������E��6����X� �"��� UR�����\:�:C���3f?q���T�^[����C8Ցc3�٦Z`Rc� ~~�����O��3�a&bsD�ޏ��g�ޠ�b4&/	u3�)��X@�OQً����Z{�"��_�����U��j[�_�Vھ�τD�`mM:Db˱�K�I�w�0r����L�tt	!����A+�=Hٚ�S���#.����aZВHt�x���w`�hE�HL��:Ko��o95i;�&�ڡ�v�"i��J!t-E���T�R[�w��$r7��묿��U_M�
��L����aU�A�.R�o<ch:H�R�ʦ��h%`x͛:tC@��s�1����j�����v��r�Pw�%eap�b�Fy�>���͞}��>u.�}���I�����Q\\�!rp�j��,�=�6�ܓ|tU\�	,m�uw�F�3��.����n*�V-��3Q*H���|�`-��qNɢF�-h�	�����K��bL��-%PȠGۑ�9��p�f++�f����C@X���qr)0��oJ�z�>,n��D����2
qa�i�i�[�*z�90�p٪T]��"{,i�o�I��Kg�6s7���Z��P�2��x>����@�9�^�E�l֭�����ޟ��b�}鰽Z����D�"�7���VȬ��]PP]�/US?z��?�W��r��F�wN}�fI��T�4�|j�n[�������7@r����=r��E�n�~J���:^��v�N�/b��U�Ȣ�< �w׆��.���$'&S?�z��:gtM�Hܑ��`������xhekn�	[�Ƚ(|<��1��;�/X�OTr��?`�{[o"�l�9�� �ȭ�'Y���(>��m:^�����Y$��ZU���0�ѿ}8���q`@�yf��ߌ��8s�'I�F��Kv�4��s`�m��=�q�L��WV����_2T9�}1m�b�܎���H����I����I?eO*��Ȕ��f����*X0P�ԡ�/�:��Җ���<��[?@f�OA0�t��%~�'��g��Xi�G�n��x#��7h�Q�=sr|��K�t�K�
ZT�	�Vl����9��$\�Q��DS1�".ꦚm6�\���Ë�]��+opԪ�8-��D�AX1b�������f�\,q�=|�ڸ̮2����X ��Ƥdȿti��(����Y�-�=�s%j#�۫#w��>��0k�D�~��x����Ù�ą|����
QO.�c)P��:�4��W@>�q�����o]*�f���q
a3�b1��]@;x���YA�07��uz����o�Hi}GG�w�3�_D�ɚ�R�'I��QJ;K ����.�U�X4�x2N��8>�����_�VmG�@#��Q'�E��k�{9eҤ6H$��1=�W.��YBk²��Ng�T4 ��.��!�~��P���랞r����-�5����J}/�*Y�ewο�7ר�3Ox���cU�b·��ħ�'���w��VӾf,?{�M)�pF�_�]R:��\T�����
�`"�����hD\-��h��t�2m��5��+��7є") l,��
})C9	T3F�;[�c�aÎ\��a��
�6���ω�慊/��ѹ`���`�(CbX�@16P��_�նGD�.�3%��?�.�U��rW�%b��٭+��m����T3Q{�Z�v���[��<���v�<%�M��p}·��'�(8��S_��Eر�1H��lm�׮eI\t|�7{Q�a�� `l �@��Eɟ�٨~)�F��������+������@#�ɔ�cI,���d���v�Y�������a:�x-x�"h搴l�>����
��(hH���y���Wܔ��%AZ@����ܭE�~�Xڏb�\uʘ��-)fv�ᓒ�Zz:	,�� ��uh���kV�"=�Fǝ�w?�4���ȝ��rzF����_����RR%���0�@�:w��(���u�"�����H���Q|غ���Jz�|v�ta�%.�O�Ǻ�T�!��nu�Y�0���h5[���ۃF7v�a�U^Gw��a�O��_����J�� ���B�!��6ԅ������,$����u�^���ĝ}YJ]�/�����'S�8AS!��3��Xp�AEc�-���Ǫ7K��>���4��O}�2[F���>��^�^FD�#��Y@\��*ds�$eي%M;U���bƗ�k��#C��a~���~�Ⱐ�BU- |�y��pn��� ͣ��"Z��'t����5��%Ʌ������|�29��{���:1��rh��5����������)�����QJ!�!;M3ƭq��TW�:4F�gP��XbBfZ���A)H8��|�5ôx����_\�]����	�G�T�Ai�%�zz���2qF;�4hE����(+4���4e���g����41ܜ���`�ː��S�^�Ĳ��
���n	�&��8���p��J�wlf�SN[	���������� Y�^"�ᯏc�kc�̵�����������s���M<�(���F�s՞ʐ�?����6&sj�6�2B��ڜcf$�zC��~�rhy(X��Dk�X�0�Hbg;��t�kƃ=���8��GZ�!yr5���D��4�k}�7��Y�A'�����w�g!+���N�����-�T��yvE����j.�W?�R�됼��}P�ȭ4?Ֆ���t�nW���{6��^�)mX�	7(Ʌ�޶���9��E���r1��r�՜�r�1SOAE�i��|�[M����A}���s�8G�������E���o��E��"O����s�����>���3~|�> ���~uA]Y��I�Hݘ,�ٟ�!;ڽ=�����������c���٨9���?��?"�S��A搈���7����%N�{P�xrѥy�� ޘf���À�_FE
$q�����ڸ�\��Þ�T[�йm���f|Fm�X��1' 7ɍ�+�:��+,�Ƿ���˷�Uvn]~�&����uI=5���_T�|'�F2�Y� j<%�>��������=��f(������۲�'�H�|�����߱��ď}������Ѡ�((���5�0�:X�{�#�s֧�p�^	.�g(m�9�qb��_YA[�Y�f5N���3|~ �tRrE޳3�󎆏�/1�	}�f4֋6���L�^����rYV)�gmSb+	�ܲ��-�8���{,ٻg>����S;�1�a�ׁ�y�W%��AN��k�I�Qr�N�tF��~@}�d=���?ӥ��]	�ů�9��q�Ė/�g#8F�C���gQ�_�x��;Gx�-��n7h'���e���04������O��[�ywm������%ퟜ�!ܮZlsx�B	L�%��g�{n���ҀA!X?{�\B�g�|�[�R�˵j-j����|8�z��Sm�\��؎��D��،�!z��~�B��Kt�y���j����e�_��o��㮧�`-.�2S���R^��W��
U�@B�V`���;�2�����^j�r)�T�s!�j|_�l<_�oФ�A��;S�[n^B������nQo�B�k�l�����>Rz��	F�3�i�GSrnS���A��|#�o�ܫ}ר�;��3�9̄����{i,����O�m�t��I����b�3O$]��ؘ��b���3X�A*��6
Z�u��������7�D�������#l��й���N}�g���e�tEZR�P�qq�q��R9�)�{��O��x�9���'&�.`�
vg�6��~=}j��j�^&�'Gq��
���X.�>���(���S�`��n��|�]��������i�\mĮf�;�*V��m]�c,&n�`��{�Q.=����ovqh2 ŏ�W�O��D��)�˔�`���ֻfi��������!Q�|.fq��U�"N��8^/7D���\���C���ۇcu���@
+���x���|tF��P4�k�jQ�'�9EF�y�ȳ�)o�I�~��fdt�G��]3�+�kCb7ʌP��A�+�sY�9R�3�&�n�B�(J�R�g���c=�'D�=�Іc/( Wn�k����-����F�X�\`��C�E�,v�0f*�.��*wv�4��n���_dи3�u�!�?�L�l�N�*���'ʌ��tK]���+�~����٨�����"���T��.Y2^�4WE�O5���bH�Q˽����p#%�d�� ��uF��4V�T����O�����������M�O�a�w�7�{��߂�L���_��h�A3Da��Q'M;R����^���v�S�� �1] 5��ӳ'�Sì?�3�A��Ysܖ^�"����U\K-T;iϙh �>�GvmF��<��B���Z '�AC4���Z��{�x������f_��Xa��]�����K��E1���FF`��Z��?v�L5ɶN������I"g�y��@d"͠��#��W��A���ږ]V��`{�@�ϵ.?���L&�%�O�Y��X3���d�dU���7i����w���e�.+B�_��)镉��p��CnpuFj��?��7���ur��� ����R�ٻ�D��(KNd0��<���C6., WB0�u����&Z�(��ꭅ�)M��:x�&#��<�Ѫ�[�`Ď�z�,��-G����ܺ(�����s��f�ROk���㬈�EGӿ��jO��I>ؤt��ZM�p����
�����V�0����RD��;�\|΢�:#6�ϒ����-f��!���G3�x^��W�LDwC�.*YR��\zB�a3O:�OQ�"�z��8��ie��5�ÃA犑�;	�r+��+��b�}��}}9�pL
��[��<NFx����j�,��]����Ws^�F�����}|g�.L쯀��>L6�����fX���+j������hb���MV ����bH�ʹ�F_�v���Bi�_�E7w5kDs�V�nb�_���6�f�9W�w����2��>���d���YG9���1�ci����5UGD�Ac&�$Z3vN�"�A.��0�=� l��}�[E^���8��A�l=r��K����-P/�/G�MQλ�ϳ|]�ϥ?���ZAM�f�����+��>�W�=���J4���$Ɍ�aqy�$��#Ͼ�ƻ(�1Kum�5����ݓ��nRU����Ej�6�Yv�m̙m(A-���7�e� RZ8�:��S���0�lLݙt��"k��4h����z��i �}m��_��^k�����m�*k�g�wӢI��o�j��.�팹>��/V�gY��x�%���'��ܺ�&�ë�0�5]��Lݨ�Y�_����VTdٜ<n�t���t%�#�,�+;��8`����������o���18����׹�a�ho�f���F���i���Bp��"���g��ߨ��uj��A��˧3�˴���v����TÜ*r��_)��1A�ǋ��d��̶h�1�!�׿��?D��E@c�^�̶g�����9[���e�IK�Ǉ����
t�)8IK����Jt4��ن�	�,>]��}�a�v����C߃�
<�ˏ�����åuu=�t�P�	Y�*�Jb5l�9�3�ӛ9����溵:����Ǭ��_9�M9oB}�a�䑆쀑g3��Ez0�02Я[ŝ�v����d߲���T:} ��!ڶ7[6���-ߘ;魠_�P��r�7��7�i�����ND��Q���Mj�Soe�P�f�k,�Y���O�@�V޺F�D�F��K������{����66g�!�W�E��6�d65����M��`�z��E'd9��b��H(Z<�؀�(Hjo*=d�7F~�ق�$Y����y5M˞��F�r|O�e��3KԨI�?����$<�2�.��|M�\���L��c�)-dR���ӅN����N���K��ܹX"� ������:Š��Z�($i�*�Ǆ�!0�'�j�&	c��*������g�퀐��>��rlK�HO��Q^�.JK�Y:����2|��6T�O|����YEԹ�Au�Z/E�ؼ�	����ݤ-�?Obz+��^'3�M:�߶%�֥8��fn�F�[�ڔw����#��*�:x�m�1���+Y��KX@JI�9�6R�dm^�cIy�|�'-��;#Ԗv��g����K\��~oݸ[	�����@��\�y`����Q����DO2�[����N֎�O,���24��(��d������#=���"		R�i)a�l��=���ą� �%~ͫ'���*>\俿c���VeS&�Z�
Y�.
��&r���-%ըU��r�Ab0�_JkbA���5�$7æd՚�/y�{b0;��T*
!����\��\!m锰����C��e�qa�5V�L���$R�|Ws�f��%�	���loL��]=�3ĳM�������=I��tW'xZx��'dmD���mtb,iv_x��܁�-�JȞ��Q�+	8$[�n�h�����;�ä�� 3�j���X��i�2�~Jr�~9������aO��m��]�#"��������b*Վ��t�Ȍy�_K<,]�X�*Sズ!�8� Ģ����^G�ǝ����;����/�C.B�X��ٚB�aPr~�"�3[���^����d=s��!P�����aG��e�,�؂�����_C @XO���1�����;�6S?��aS#I!���h$f����a�OB�W2�����W�����0mE7�>ZU�~x�Z�&aGʪ��5ɥ�)P�l�Ъ�
"_��\AS�å�A
A�gY'�(9����F��U�>ɼ�|�f��HHM�_t�M��9u@A*A=�x߼�yb��~�[➏�FqG��۝<P�AvP�o��Zѡ��̀�� ��vPD.\��/�F[9�	b���J��C�>�Ҽ�߃ի��6�@/_y0opQ���7et�]Ar��� �V�?�R�{Oe x�~��i�˶?�[��v��V��'��I�"�p��Q�ť�#���<*�04�K�˷';*F�XΜ�{�N��6�_�'����kTa�kFu����]���R�Yf��!�?�\��e�x�XS�ԓ)�ۭ�R��R���*�-�Y�:��x`��ElE! ǲ�����K"��V Sd��4�:�o����]���+N����7:�aV-�I
��S뾑a��-�;Z'�D��G�4��7���<T޿%���܍Z�EŸ�?XƲ��H@Ma�ZOru�,Eq�� �7���Y�V�``9��G&���8��ݓ�؏�ϕ��ds���g��N[�6^_����=ei�kc(����6����ŷ��Ȧͪ6-,�%ҐݥZ�����]�!��Ew����:��ʑ���p�9���37"~4����V 
��"�u�h��&�2�!X���`UA�02��jܺ?�}bd]�*�-��F�ė{B�eQ7��j��F��S�P����� �M�.
7�DH��%k�E�j#+k�&�,Sg�d�A#��I��~��QW��򨑆��0�XE�f�$�����}��/uU����3�mi�L_:bҋ\�Q�E��*9���pz�� ��[e�PD��������S�'��e�076?�DщS�7�Ƅ�η����w@w6��Jc`O��[k�m����N��nwuu�?V�3ܷ��1Ag��bc8^P�Zͷ�53E���p��#NXc��>��ĳ,�CRn�L�L�~wx4=�͜�v��Wm����� �HC3�ޮT9��B�>Q�	�!Ur��CӍ��ȅ�]~��֞6��G+�_��U�]f�5�`�vka���* � Ʌ����p��#��*��FLV�,�hU��� 8��e:)r���C�5\c�f�<�DO�5�
-5��fZ2z�m�M�ʗh�i>[�ɖUJJ�V���v���	*�c�M	���7�f�Ξ���߿Q�l��kB�([���3C;ʷ��jM��"n|��`w�Kmx�/�;�c�D�M	&욨:����5���wj�P,��� ZiQ��b�����j(�[J  �Ƙ3Ri"�!�L���#tn	��7B�n�P9�\ܾ�^�½��������@M�|� ��n+���&N�C�xD����>$ߛO�z��/����s�K�n5�¼���ހ���L�����()ٻ���@Q�ѫ�PV8d���k��Q_g�8j=�W"	1�;�QdA�հ8{��+l�9RZ��X�0`"
�Y�jWV�0Ixom�b��L���O23�f\��e[i+�����⩈����n�4���3��e��͋}�j�:TE�+�������Z���Gw�dTT��
�*Ǉ�/�v�jӌ)]���6��uB����:�c�-V3C�ҏ�d���(��jHm��*�M�3e}w���ѷс���T�i���n!-"�)=��ޔm_}P�I���;o�?�U�?7��u����K?�%`�y�U�-J]t�����o2�1��;I�g�|�����C#��%ќ�C�$0��'�W�Vm^�=.h�&�����A)7�xN5���I�5�v,r�&]-���I����<N�F֙�HG�����,��e�[��T6��e�T|�2��(#�Y����D��v�:X��h5Q
MnM��5��[� 1���V��Aq�Z~�m���X��[�=3{G��9f�w�¸�m�~�u�<��)���U�����%�mmM���Y��ٔ�2Q4AW�t��N�~�$�����Շ�w+�x��͢���3�0e��z���U�*-���l=�,ly�1}>�]^�ɐ(�����M�@�0#�'4�u;�U���؍E #Ȕ��p�:�f0O?����т��؂�`TJ��h��4S-�겊�zn�/��9��͎���[*�݀��y�8lk|��������Z[k+�C|f0j��n�&OZZ 5������b��͊�
#���@�v�EJ���^��c�^^�B�GsV�ncbɧ�������������<OZ��OM�m�a���/�B΋����9�3�~��H��Ϯ΁������$�b�Y�t��`	��l���yR������D}���W���q�|5I��Z�Юql�(����v�硲Vb����5�2��QU�Cҷ0��e��ֲ yB���#ӫ��b1�2���l�v:�#sf?�$�\�K60P�.W��;�\qM�z�%�E�2��у��Ұ)T�Ҏ,�w	D�C�N�� ���:�Jͩ:bS��=�-�� m-�9�������K�hx9�O���X"6r	���17�8��)k����j��JRs� �}0���)�ǟ0�{qtq��{�6Z���P��mz�7��R�� �'pٞ�Ao�&���cqg产*X �j(��*�y:��wZb�ż�ʐQ~�`_�`<�z�PT��Y-_�#����3����d/T��$�mp�*����z*�l�;�HY$:9۵܍9V5r�J���$Ch�����>�'���˲�%{���_Ȫ�g�5[y��N����䓨�+Z�r�Y��t>��(ҽ+�;;�����ʀ�1��,B3�0�5֓�n�r��k�"��8>Ӵ7g�)�Z��s7��L��c��_���b��-��G��f{�*���(l��ay��D�n�qb���0��_R��JX9"���>��Ȑ����@d[E�o��C\�O���幪�N�<Y0y0pB�����i}f�Y`����o�d��e���ZR����@�@�R��U�/�Ix��b���Ӭ����@��%!ݾ�|r������+Lp�2�T���H���Na�"��le�Xk��8���"?D�Fɖ�)�,�1j��G��(�_�X��?�a�\=�p/�w���-G��g�����TxxJ����~����R?�u���V#�Ȉ�-_����9V���5�~�v�|\}���iK�����{�j"�@�Ո�4O;ѷN����c��UU���)�ٸjZY>�p;�n�/��L�V�-*8�	���g���?0aTӐ�Q~u[��Qu���i�{�r2�&�g�fS���\S�#e\������GA�g�����cU�o��˫�g��m�W�֦@��fc7'k��Cc̀�J��`P��S����̍Tɩ^��w0Rn'ND�f$��IS Z:�8���N��nfl���S=�x�1��1 Iv�<��'�f���TΈw't����}�ӅYQL�ꂃ2�%�y�Ɨ�,q�[zQ^zyv�U�{^jΣ?B䤜t���M�X���qڐ��L2�r�P��f���\���qO0�����p���X1�>�s����m��e������Z�|_f���ZRә	]����SI��y�"���NG�qo�~���
Fp�Y�C$��{�W �[�>g��L�.٠e��|��o���X{�Ї�;0!��uT\+P��ڰQ��X���X�ïc�pN7Q�����N�r��#x�?uY�O�<�"zlc1�t�R��^c>�ǳ�TFpZj{�#��N����x����i]��g�K�>2PI�z�Pmp%4;�jQ�:���v�X�ݹ1�I�\rs4?�+�e<�~Pd�HJ�e���Ҡ7]��-�Z`+j�>2fǈ]����F�k�ՒDB�s�;t9z��3D�W�m˿��QY?�	�ܫz/#��|�9)���e�e���$W�ݛ`���.�H�$}Z;�*\g~���ј�#�����Y���z(f�E�	0����+a�����I�I(���Ђ�Jq�(�`�Ņ�K_?�'��\ɮ����۽+��g�Z��*s@�v��w.������vͩ%x��f��
�����)3><�����}k��]��Bi���`;@�9ߐ�Zã��F�2�
�z�|�U���/����R8�v�?w�t���p��ÕQ�z1��u�w�1t��_:�6P��)%�T#�Պ ��L�����S=UK��+<9{�#��Vkӗ�w|�%��OV*�gz�R���Vt�ܿθ�B�Z�Jm��`����Q���43�,���ZE!I݊ ^X��[\S5�N�"���=S�g\ov����=�1��h��0a,��
����3^�3��+��0U/�M�L��DߡP�q9�0�%=����s~Tϧ�n.��1C{*�"��e�^\��(r�OU�Ȩ.&wx)
j�ND�ڐ��Sw%�mW�n�D�*FQW�Yo���]�vF[6�˰��S����!�vd9�m�ت��I��\#�QU���ݵ;;%l�:�H���=i
h1h���K}@��/�PV�����t���րӖ,�q����m��DS��>73K
�1��ʢU�9��4ґc$���f��.�e�@0)��a�X�gRca���r0�Y�2KB�%e�r$��O�O~���;"��[� ��z�d(t��fV��R�OK�o�T���ꆫ�5T�)�i|��p�GyWgL7�w/G��q�ٟv�Fe]�
���WBU8���{���
2,!=�\��SIK��:Bea�Z"!~V����"M�ǟ9�f���M�K��|<���0	��̬������ѪV��W��Ɛ����UkO��o�S ��m�\$:c����B��`�+xXW���0C>m�ܭ�"��$c�K7<t�_�湈H���~}sf�)��
ZZm�������ԥgT#��~�ա�^w-����0������W�=�[s@�ߴȔ��}��=�%W��ԼEA_��hڽ�D�bx=v�K�Vg�[Ik.��ڏTX&QdJ��s'���KB�SZݜ�n��K���J�H�Iz18�=�`��ކd�pB�e��3;�Cn3���+��T"�pל����
J�(����ǻ�\PS�1��!���X����8xCٚ#�� s���Dsj���҆35�1HR�e�l{s(��Q?:�fV��5�#��3;�c>]���91��ƿ����e�V8g /W�+0%�ߡ[��`�S.����х��Xy��M����k��OXt�w�|���poI_�:E%�J"t"XY��K�0T�H�P["c=���՝��5����#�W%����gef���KU���g5�әJ 4L�}/�+-����j]C��w� �A�h����"=�`daf^
���
�>�Ƶc�P�K&��UB���L`M�=�2��`�J�=��E�����myF���9�+����ր�c��#��:7YS�5l.�e��dq$�b�c��أ���F�V�~t-�$����Ţ��v ��[O�����@����$���/֋��}X=�y���N�����
e�L��/C[�R���:��&��3�NL��1J�e����������6y�R��w��P �sG�s�4��ޕG��fe���jg7ག���[�֫�ЪR���pL��N	�P�F���s�<A˹�Bǰ=Bϗ���@�d�IL�j[��`��;��`�˱M=D�W&�*�c�J'�K�"��+w�M�0^0�E
��_;6�~�.��#Uu��Л��pCsK�#m���=�A,s�C�5�/���&ӕ�g��HS(�̍��GB^��9��e���ϊ��acO�W*y�'{����^�Ҕ3�{�c�4Z���q�T�����O���x��p�UlsU��0�f���$��
j�sE[��&��?&O^�hǟ~�����v�!�@���~�1N�S+I��6�ls�`wo�r4@��7��K.��(b�������H�o;@q�Yd=H
L����u� -���s��S<h�
T�Ypr3�:␘8������c�8rb���*�Fi��B}��LX��R�C�_v� B�A .�����W�~��%kR�:�f�?^V0�Ng��4p�7�f*c�z�,M]Ƕ₷^���So��+҉�D�B���i��b!̳���r5���m�E�{�"<��B��r��A�����`�X�:�Kа*E@5�
A���G�b�к��4�Fv=���g�X^��a�� X��.w����op���(Ķxv���zC��QϘ#�;Â�oň�5���b�� �6)<��j�G3�/�����=�Mb#=�S)|܈�6��ٓ�K;0�jy|�MSY}l�bC'W]6��I�D[%A���2:+D�%����J�@�4���r����T[�<���f��T�DE�īf`����s��{�fVe�6P���[b��Y�������&�I��=���vU.iy:ɵ%Պ�s�MQ�����w'�{�B#3P:���":M��b����.Ӱ�?�K�@��}f@1Q�>y�×p�#>��b�^�b9H����bͦz�.�D�q���j��!���,��i�h*�S>��Q�(�e�V���a���!G��Z�˟��[ϡ�td��`���c�/���	y�� ��'x�yx|6|�L9���	���{�-ĝ�y`x��Ƿ=l)h�a�Vn�c�/�۷t���ޓJ{��̄kI�@�/V+�:�������<=�5_^S傋?�8k��n���#Dw�@ ���'� 4����
zDC���Tr;���Ui�#O�E�	�H�jA��Y���\�ƧT���R?2�C@�ˬ��.i�dȋV�y+١��Wׄ-�J�ӸGGT?
������W���$s�:H.�>�j�̎j������d�h�]����b�^��y~|�I/jug��&�Ps�_�Z���<�+���!�4���<��v-�*-)>��f9�n�¡$��YZ��B�y@n`� �3������N���d�$ξ<B�'��䍕�.U���w���t���h��dm��N���*UO;lP���ߵ�L$&��-����1��E�ׇd�DM�^S�T���ǆ 3+V���\Z���W�6�� pC\5�|�����>�:ɉV'��G9��.����b����gxƀ��f�Ѱo1z�5���ej�:|�� -�HA2=�)$�-A/�)�P���Bξ8xdI�v��+NS��H�7ą��(vQp��^�@2��$�&|$H����ᔙ\D�pH���Qtg�
�-�5�^�|��R*�,&�e����%�)7��ř��oM�$���LdS�nM�f�����3,�\k��^T>Ȭ;�'�$k)���wi��b�y�<-#�y,iS�t����k�s5�C��R=kg�4*�JU�k����P�Ǽn��z)�X�l�1�
���5��3�:7$�&����OH[F�K�X:3����C0�5���l�V�+`���_粳������ ��vbEEy�6���� S�B����H� ��Բ�u0F�����*���ɑs�1�e���$�o��aP�[kӶ��Y�s�?�C7�'�5�r�E�!�r���Wr�=z�\�m`�D�A�-<QL��_e�\�7מ�['d�P�z�.ۤ͡���+ꉗ� :�D�t4u��;��sD�ʟ+m��;bT09�*)/*�U���ͫ�kf���Y��
9;ky�H��=��vԼf!�瓯���EN�����0;|�V�/e��V���A���Ǫ�f����y�HZÞL{�&Q?V���PD���J?�4ϛ/�Aٙ%n�'��L��\_:�ɬ�c>��#aj�	rvu%RF�_��K�@ℂ�:f;��k$�iUHK��IvEr;eP�b�Z�m0�,�!�����zA���=f�ZV�E0��[W�LÃ-�t�F<��d�"Q5n�9�����w���F�L�"CLH�Ѡ�˭X&�����":�^\�7+<K;Z^_9�����*���*�Em<���3"À��~��@��%���m��Y��ֿZ
\^�*Ӭ��j8�H*�)������a�Yū��\3��3L�c�|����`|��}��88��*lj�����_yC��q�ɞV~�sB���ʃ�� (�������٨H~L6^ f����g��a����{:�@����Xg�{�)S�ݽS���W
�����������-��"@������|�r�c��E�T�
�IY�Qq��_�?�By^��� �a��&s���r���������K������h�r��c<�@�Vh�ڛ�jI���=�G�oZ�Y@��/�aNr��WX*,�ͣ��0Ճ�Z��p�Mw8��2���:���Mr���1����R�g^��.�ԯ�ͷɎ�#q���bj���鏫7�r�y`��&W�i�Z�Z�V[�5+҂��-��z�zd�8���<<��{�0\((3�zyz�zŒː�JI:̤�)����Rq��!�4v�őg�>�<3���D���~cX�=g6LGO12�η�'B���*�Q"����K���H�8���^��"(���<�ze����|��z"��J�^��3LL1���z=�z�J~'�ٱ��y{�EWy9��ְ���@�+��2c(�<l�=�+�j�|�{�x���pz���XSFyI�hR=à[5鍀,gF�-��3�}y�a�)�k�Y��V�I [ʍ3
ys����y|�Z����v��vI�V��+I�w��	`N�t�3�o/�h�d�bp�U[�4J�ݱ�%�
Z����a�3�;Wk�KQ���.*�.�l)Ɗ#�f�X�b;B��R�:��9�p�@M��2�T���b�842pg���e�+9���n�� A��t=-σ�:���b�Fv5���T)6���D!A���C<o�%����h�֚%+E���%��y�,�=g������FHٝm5m�Fi�܍�5�\O<+C�m�D�t*I�1�=�
W�Y� ~�|��.��Rho��E���j��i��A
�zz��ڍ{-���+��rY�G��CG�e���;�^M��d��C���WY���[�P:��(�O��'�>16^�]���o��"&h�K�M�#eO�[�8��痾���LA�ӷK*/�E��}4A��<�Rߣ$3Ҧ�s�q{�V/�"sV��ʷVs�R��>�CR��O�\��g�7��ǥ�]�Z�&hsØ��1gx���@��AM�S�����A��lF"x�~�Cst]�P! >>w`�u8c���P6#��lx���
��M��#��W7]��Y��9,��ŭ�cu�a�0�I��e`5�)���O�w�ƾ����#;�����v\��;f��扴V��F��r��X���y���Z��l����8o]r�9P3�Xl�G&��B�PR����Q���BNkcPP��=C��R%+Н��q�-ty�ͅeܐ�:�ڲ���r�c˭�Z�>��uz�:��.� �6��;)k
���-Ŝ����%�.@�2�>Hoy�
���r�����E���'z�
m�>��C�~�R�a�Zҕ�)�܁�8�;k��A���}��b}��tq��6dHCc�t'�@R��-Ke��m\N�./�:M�B�Z��o3J ��t_�b��[�m��)�
|)��7�L`l.��e�]ħ����x�>c.T�brۀ���y3�O�F�_�����v�%k�3~��#PQ�X��06hI2�i�
�%*�9��]�1,�P)��k�/Zޮ��K`^��s��k�g�A��z_��Y� �
T�1GC���Vw��V�OC��QM�$�'KdE����A�E���|��jé&X=+j����L�	��ȧ@Υ�Ww�4���~��Y���!��R0{�6+�&�)0�g��A��pF������?�M"��X�?Ϋ0[���:�A��k�$:[Xf���˯	��1zl?�:O*�q�u��;����atC���Q�c6F<���o]!J�Կ���&��՜j��x�>Z?p���_�&C* �?�g7᪅�KM6��ͼ�j!��b�V�r	�n�"�4�!�͘۩�'`I�X�~���������@�f���m�?�S1ʋ�z͚�z�Sn'�j��/�$O7�?��&��`�����>K��A���^�����+%y�^u��"=i��'t}*�g�ƙ�,��YhqT�pB�/��)���Vf��H���ߚ����e0���(iF��}Y��Y���SO�}j�UAD"��T��y"��5�����|Q��:M��m�Dj���O���gi�T�����l
��[�*񉞐�TL�+���
�QK�ҏ���N�K�F��2���e���\�D@>d�eD�0oF��z����g������Xm��:�N�vx�G��-�vX��Z��1~��S��E1�^.���z�/Cn�K��OR9�B*��F>�X��f�/i3��Ĺ��.-??K�3�F�A#��g<��)��Tj���������.��ga@z�.8�qj&;Y�2��w	�!��塣C�\���8����F�j{uB���` ��W��ٿ��w�<�RO[\40 [is@�8dL�˓x(S�K��Z2��
#N�Z	r�0�5j3��̓;�6ւ�?F��Yn�TD�#+8��Wy��b��5����60g�>U�;��P�I�%�E˩ukBɼ@�A`�4��
������>dV^�yo���c��lp�z|U:�w	���n�2��IyO�C23=c辧9�s���GN��B;G��r��y5xp�sq3��Bv/A�*�3J������NT��/�F�2���MOZcaHo���5ۄ__�|�l��|�2a>h@�C�=�/�fν�$���c�u����c���
�`�t��q����	~k��3B[>�����˶o��e*��ߪ�H�Rg�9�!ԑD�T���Q�s�qgc�恷�>UE��)/�Ђ0��pR}Z�8'e�j�q-{�z�&ypr��`�L�����]Qh�D�z7G��J�����?�j�. r��nہ�}C�U6����~E�L�
$(��0ح39A���R|�M*�����5��������WT���$C��N2R��v��!��rG��k�O��Q^&EK��S]jc�{ҙʲP�U����\Ռ-�w/@��µƦ�w�n�ͻF�| ���
�!�{�>(�yI���R������G���p'`
͵��z�K
�]��e���k�GĪ�Z�|��X�4@�a�����})
�,��i�\���d���k'�G/�r�~��-Mty�~�9Zy�RZ(-�.�<n��v�U�K�D7@5#�
�)P�!Qd>��Κ�c@���U!}ap{3w#�!�[��c�LW� 'i2Xrj>��/�8�
:��I-y����)�Bf�gT��V�KR�r$*w}e��TA�p���D�"�,>G�-��	��RS5� ��ƚ�!���&�*��G/�5�&�%	T�'�z�K�nI�;A�����)��W��7B 6��S��a���w��ո�u%G;�aU�X�k:N�~��5�r�&RvE��v>LB"�7��*(&���&��7�
zw�&���f	~���V��q���2���=1A�jf��n|$j_Y��L7�F�݁VWf��(����S]{ʫj[C��Ғ@*(�cO0���c��v0���kX��[�׳�n��=l.l����J�\Z���=#IoT�HT����ϥ׋�[ԩrˏ���Tb�RU�8�V��X5�*<T)��cJ�O�4s���nD�瞉X�8[�)tWW���ki�q6Hۜ���G�f=���6�AzGv���Ca,�3��hP�����.U�nú��>�V_�WԘ�-#^�q�ȗ�UN�B��o���bh�k�����Q[�i�=1��|n��?!�!�X�4��Bc9P
Fb��I��8���p|��jh�/����r�(ݙr��p�	M�#J�{�ƌ!����}'��D�t��e�����0��`+�ʛ��&S� �_�`�~[d��n����l��(�&�����ױxF��^���ފ�����r�\t'�*��x�|L����y��I��"X��7��-��6߼�ZÀ�G��
�&{�d���J�!e�ΎD�b�8���DH�2 |6AFxCU�q%F��
Nв�b��yI�hڡ�����'�/���K�T�o7�o�%5QR�v��]OJ:̐���֏=o��>`��`:8�)i�e��A�4��h���y'U���w�ן�:��uZ~�d�d�bQ_g^���*��#�_�aD�]����%��`"������R������7(�[�ƫa�t�?K`c4�#��9ޝ�[BPl��l#=m��仝�u�=�ю���gAm_*�|���'^�^��9��9��f]�O�,6=�ۣ��ەZ�z�)���LO��B�̩�(���+i%F�����2�Lk���uې���V~�o�T����7Fh0s�jP}4&�c'S��{ޤ`/�F��8D�8H"�������f v��07��[�����u�����͕���n�8�RLGi|A��<f�����.u��>t�I��ND���o�	�O�Ec�R^�Z��G��ݰp���FD�Zǧ_J��<� �L�k�9��PC�����u%p�4hWq�8=cBϫ�l��6��s�$ӺcE���e��3� o��I�?��R:kF��XZ����Ebv����ntF��@�^6����o�ȣ��2�D�TQ�*�χ%x&�ZƉոv��AI1� �%"	'�Kٔ;���o)%���'�ۃ�}��&�8������t���P�<(�=s�,�[����2q��d4����K��>�o���U������˶�b��~�[��,���O�NS�3=�&�޿���]ΜN�Y��4��/��8�~eQ�܍��U�]nxp�Lbf~��t�.��2�R|-������óP$xbn�6��hؽ�����G�`�����w��E��œV/�Ѵz� oZM��4Ҍ�jz���A��"k8V��<{aQ����:K*��|��� �	b�>卡䫐z�kB�,*�h���i�ljF�+��'�u�������r�e-/�D�K%=k��,H���ld��5��V��_�	O�_�����Х�a��V��I|S�x Ca.��%��Ty%H�홱p�gl�L�뜯����߫`w�%#�yf-X�B�����`���q�KT�H�땗wk\�����T��M�&��$�P��C���)�i���%��^"��b�X���w`��&��p8�X�����r��	,L�`��b������c�I�@��T���.$0�7B-9C��V�4z�C��YT�����m�����S��=]؆�z�R/F9Pz��4X?��ч6���euϢJ�4�.;	Z��C���e�^�������@�T#W�6����������#�`�P0�0�)�c�̿,�zA/u���_�D���E6[f���6��_�&#�O��3�H�FY�l���Aӝ�zBu<��X~�Q3	ǭ�Cn�v�ÙӁ;Ӛ(�pN�[��
�C0��l����=�f,ؖ �x���Q�T���;�ل��ܲ�r�e��T^f0z4ņw����r���T�������u���Lw�}Y4��ԑ�ƚ�ا��Q�oZ�!Q6C��q1/rz�kU��n3Q�j_�|��H���:�s�\��D�������1.�{���Y��ʱ �Pg"ɇ�aS ��i�ƧUV-�t��;�V_�|M�.�O��	i��D��:���u��Z:Q2`{ ����L< `	{��4҈�t�@$"A��6~����,7�$��� F����38̻[�Hk_T�sJ-O����~8�[��c�,� �Z��5��(n[>�5B���D�Ȉ�ˆ�;\6�<�$o���Z�p.<�髇���q�1���3W�9����f�<��[%s���r	��)�%ӓ�owj��h��\,�l����T4�,���[H�ҚfҼĔI���N�H���c
ڄ#�Qf�E���B{�� �G!��Of�Q��	�-j#���	"'h�n���A軉I@��&֮7M 7W��=�
"�.pb�^j���!��}T�.L�8�c7�6]G�(�@!��Z�*�&k�L��+���3�D��	��"X(�E[��{¹�@Kv$47�W��m�Ԍ��,�/�Q< t�� }�_j��Z�����Uy ��}��_�'~���9F|@����~��[�	�rYf�8�nN���pr�Z��>� ]��#o�������qc�I�k�,"��}GB�Ґh��C/�z���%*�+�U�(�[�{"�����-����on��`t��`���wY��1m�)�_����ɯ�
�8ިHS6@��v�����Z�Q�SI}�{d�J�
 =e��K|F��_&f�X&�s�dx���8/뾛� ��'���4���͠�h�h(��� ��������z���C{�� S��\X�62n�@]k}816D�&t��h/]:�A��H����F���`��s�u_|�[k��t`�0�����r�[G��#�-�d��X^T��Q���XN�*5{�@?��UL[�q}�
��A ߴ�eA�L9R�͓��)]��%]םU����'�(;��Mݤ�[�պ;���-�41�1S���l�K��s�D��?�ŖM��J鐡]c�����!���1�tA)S%�n�6o���?�F�.��N���'���S`��|^�z������=���� ��P�o?��Dyv�9Q�֞�.��(j���@)�YqQ\v��Z���7-sBmܠ��G�2�Ȣ[e,D�3.|��^��ّ�1��p�e��fs��0����	q�B�'�t�<9�A�z�,nL2� ��LV˺`g�;�LB�Xy^ 	JH�W�1���y�Q���f�:ឣ��eU���'��Q�Z	(�#��H5r�:u�%�}P�nBmR���eʤ6
!6�"?�ն(���R�Mf�*w�sԅU���ՠ��X&�]��wGG��=�Ah��y�Laհps4pO��c�ƞ|����ڑ��T�O:ː��(������gF#�Kn��i�����f�}��&J��y���3����*�J��F�(^����Fv�z��ɱ�<t�
M7���k�-C��Op���U94g2��ѐ���l�l�p��IS%�؉ڈĒ ��#O|��QC���J*@�����KV}0�bb�h{t8��ѵ���ۭ����A��^��5��9�+��T��pa;g��L�:�
?����s�+�ۖ�o9NRc����}��m2X��	�< -ѣ��҄q�z񑊃\��@�(Ҿ��U\K�zg����k����,���!��#\~_�%���(K�x���W�,|]�����&p���Q
Y�|\����9��0{{�}�I�p�s ��Kw��`2����>{��ۄnN�� �X��]�Ƿ��?ij�\��+����ܘ�.��=�y�t��Pi����0��c���𽿗��Z����Q�#K@��W_n��-\�� ����ʻΫ��K��_hK5��;��m&��2x�SX�ic�La�ێ�9g9���\�:C�A(5jrR�n^!yP���,G����v�m�O�x�{� 艬i�I��*���t���yP3�]�~I�07~@=�~��*��l��i8�N����ǾO% r᪆w9qH��du!�q��NAKg9��R��򬣊�S��KZ=�N7�z&�qu���Y���ք�±GVm�t�����['�|DUxc���[xq�`���'�)�>�_�(�u�H<B[d^P�0~"e>���v0!���ߴ�E�^?rO`��,t��e���'��b^^�uR#τȘ�s��m��J�:�X �,|6"iH��|���/� '�F����i�|Z�p��E"7S��k&����|�lC�0����.�Y��Z@���F����o}*����_Ϋ�u�3�ƭV�M��ˊЦ~�4Oέ�Tw�5�)�$��������]]r�i��9�7Y�l3~	�[�Bj���!�v����٨�R����7�U�iI�Ģ��� M�CG���%)mJ�k��Ji<d� ��gq��Wl�.BG��>a��t����V�h�����6h.��M�Z�C�������F~C��*B#Uy@��Zl��v�WS֦yt��,��r0�����~/
��{�ZL�� k3���S�_GW����U&�[��F��!v}[R�TX������s�qj=�p��X|9ejf/��ރ�xA�C��kc��ݍ����^�{6RU�V��*��Wű����2����� �������~�������-��z{U�XZ#���v� ��`d�Jź}IP�����J>5@�Hql�OqS��h��[t��+�~����8x������G���B�ڹW��%�� �%i��
9V�n�}g��pr	τ��T6�
F��ly��zwG;�!���;j���y�p�HC�m~�X�_�3W^����(���@�~��� �j��wК'��́�_3�7�ΖZUb���f}ձ?О١$�!qS���Ǔ/�M� ��,)����ʂ��K�T)x!p|@H����ļ+,����`�	�}���4*pF��e�>+�ի��u ����|���Ы(�G��gx���������45�K�\[K��UhPr�����4T}��>�� �[~���g��-�������/?�c�-������dm�#q�#��R���p`X��[1_�m�Pq�i�B��]m���S��IT�>?�!�:3�&tOeHf�˧��M���7+ͅz�`$�+o>�Y�1�y���8��GH�?��5�ꬬ��?1wZA���662���t��5X��<Ӹ�~>̇��t�����:�WEغ���t������i�_@t���YT��nBo��6	k��s]�Q�Ǡ_��M|;�z�3�\��R�]
�j���s�S~�m�(:lr<�*�E�M�q]:�A�N�q�l?�|DU���K?>"�if�-�73��5�VĪ@?�|�ei�:�*%.;��=�"L��>.���>d�����-�:��[���S�~�X��&����9�NS|���~�\�/^� �|=a_�p��(��0ȅ�z�ݟ|��'B�`�F|����r�:���M�!gk�/��ĶMI`���j�t��c�"M�b�~-�%�x#��XZ�Ur����������k}�C!��gG�,��n "R��A���*�3�+�^�)n���g<�>ڬ��o�c�T����ߦ`��)j�x�+^�'��P^�`��>�w�Q���7���_�Y�|M@\2����^C֓�伱�DQ\}�k�č�'RS�J�]��n���'����k��7!I�*w%*V�*�M�H��ٚ)�v�.k��G�~л�P."*s;�hΪ?QPT�{��`�9V�I 6�a������� }ם�i�4�X
�:��b%��"��z!�*{h##��]��m��'��y^�l�OY��0n�<B��f��H�м�,Ζ����ڔ�������������ƥϓ7,;՘�8�Y�?��$�p�ú"�>���!�\O�Ϯ�Z���GV�\���ɻ�Z]��a���W�V�}�����[��շ2�dzL�凜�cR��#�B��A��Ĉ4�������`R��lŬ0b���� �l���7遗���=����5��Om<���c���Ξ4sD�4��8as�Zl��GY�+�-9x<5��EG�9�{�ݬ�|�����7AB���ҧ���iV����3�N8�>��Vu�b��ީ��BV�<8v�J2sd	��ˎ�Wy���u�^����@V��w�}��.l.Q;��+wr��I�:JO���C��Ќ\�����<
d}��p�K�
V��Ҧ�v:��͕���|(S�ڜ�;��f=�a��"}��8�ˠNݭ��7�~Syz��Ђq�:���T�j�j��g�b`��� �U�뼨,��Pۅ�8�����~��0	�6 �{%+b�c11���y���pK+�9"?�\u�?'�)rA�.ΟH�ckP�nߦ�F%.�R΍�3Cg��M��Ķ7þ�SU����ɀF���N�'�s;ĩ	]b�p"x>��Z6����ܮ�[��B6E���H�#S>��Kx�5��8�0��#n�^� ����3�_�������z�Y	"�,\�5+�6:�B��hSR^��!�ۀPLn�渁6���$�'I\)dv���(�;�฽�ŗ�xH���	W��|�SO1v%�)=�pĨo��U'�;G�g��.�u����X���!?YTN���a?�PS%�(�+���~��묭�8��'��GF�M�c�vN¦!�֋�e�B��":��H���˕���Il�o�)���X��Љj`q�ҬG��O�-4â��}\@�bk�33����d��uy���t��I�DA.�,7N�9R���LYY��yS	�@�@SKt��R�m��1Y��G�G���0/�����f}$�q,�*��>p�&�b�����VM��A2��4��3�&��
_6m��?jSֈY]���#S{�5�;)���J��͚�K<��+$�Z��;������\lRM�Xz���C�_�uQ޵*�5��i��������ff�{�?gLWi}�:pA�^SS	FY���B��=�=Hz�h7,�r����;�8��\�޷y�L�T�>�R�����r�3���^J���<�H��Bws��F�gw3	�����&�F�Cm�%T����6��#+u<���o��n��&
���[/�Ԯ����v��y<����#�����&�\�fJ���&12��%4#I
jb��W5c/�O$�������4�>2��a �*���6ϵ�7!�o��|�è�P7i��ov�%�- ����3��I�F���E��_ \m>�`E��b|����1Ko�gr�nی=t�p/����j�-үW�R"���LD��A}��ߦ{����C=@��8���A����J)�z+���=