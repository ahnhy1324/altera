// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
g0ixg+Cd9Xv0tLdLLVjRvhuU1u/Mcak+BEkdiDPAVnKFnE2oRpHWhXhxWm7QJmR9
ICb9l8WbzqQYDO8zdTbBpRDfZVNkAGnSfI8e4ATGBTDeBVHoyL8S9JdfWkaNzTiq
cussDruxp8f84y+dS1Hn4zlB0tuYxa3/pXPrs3Anpek=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8720)
NhiLbLRPJBuMT+JdavCWtqZ4nAthlbcm/NeS5gWySt6x29JdZwXG4m9D4IrBMryO
lrV0B5U+JqfN2ub5603n6i+BR3X2AZA0hJ5qXCTVKtwxV8zw7PtkGU1KiM1VkeMa
t3n9/L9XEs56gPUlUmGn1OphapE86c4M9fzCD2LNnDsWW7bfROdVf36c+66+h9bD
yE7hI9AR2psYtQ685h/PGNIr+rOb72rI0txyQ4SpvatYiKRwS6KjhMT69aPDT2Vm
sLpNss3MrI9R67dSSsuAM4G3Z7Au7nM878G5jtvEg+rPaUCSAfm8/C2glPkgN1Go
GZU1uVCu5jrLF+tiQG9NurIhXCNuAKuMMWLxxeNUerMlme870OVRp7SAJ4uLu0eO
6uv8GoOge3HqTZb5oHbPCOQCBen+ORJRJfcfBArIlLxuWFM2dve29L6ZD14B5EPg
3Kdin3sVWldelP8He6czQOJecGX88f2NbhE4wPGymeD56Q/vm4PUZQ50JoAMbaR/
htSVJRHIW1L3DOMYQWahaGCjANlml+zGaGqYdFv7ZB1nSHbW+h31gFYCKxSVIE8V
XKn4GRBB16cAdE1gZIhTbrReGr+YUf4b8AKSSY1rgkSREZHYIZom3Jonpw5S9tFz
DK7gntyimVU4EMUKl5B0JrT/VUhp4zVJUWbUIWTbf6UVBkOF7YA6hsaCzeQ49jvX
5MwQqO2nyeR4x7cPcgKP30JZNER7tM3yPPRzbHvEvWtX+Prvis4TKfff6RNlvqnE
3c3+4qZkGq2nPJz1bCvHmPwKdVQOPZMm8P4G3a15+p0H2l+IbGMhGLmJanD0wASX
/YB+C8yfmlRTTNxhI/92o+fNAUwfw/3PQVFI6+n7LZsxI+2Fg7RosBkOjaoxuT25
pCawF2upej/9Mi90wLmm72TRtAHQpPRzFORdQHXfpRLeXDQqeov4JYus9aMM3xrM
HqY4CGNvGjhfhPNAyZNi7H8n+phRwbkAd3iREXf6PmDoYmRRV2TnohSBkZwTEUbK
TgqelHuVaS50m46uUHPCi0+if35oSmKJO70PeeAAtEKDow0PpO5b+O1s/1jLbFXY
ExhLCjB6Pd21uAg5bxWRpAMkcQH+4dKdqkXOahO/VuQQQdPU8AHk6G6OaqQ569z8
XHnHF7cTUUhRs6JiDVKyAlZGDf7zisHVVDbae8xkkOeRDxwgVMZ3IkghP2kh6AxM
uW7TMAKMhAomAtYMvNXxVK0sqtiAA8m/KbvYPWgjh37nhvKlC+PFIrdPH7jNap4M
J9Ioxtzx1yuP6+85tSo7Nh8DikFGJfp6qpXV8F9UjTB8Vu6QnFWd/G0RTc80VI4i
eM40ql6pg4umfetRSzPnmHVffj5LvEa4TJcrM/j7uS40a0bcn+plUvwZgOGGbAYJ
+zi9qiV04wEnkYFfROlWiIHp+JBtYqUyzlQZhv3mTFFfOmBDLOq9zB4g2kC29rKn
YR1AvxcPS+MOMlfurcCYQApNPROGBZxCVTz+zBA51PneC4q/GUb1DtWYon/K5ev2
M7pbsHu3+eBK/4AwnWcjOG56Ruk8OPW9e4Kjp7YeswY5ZHng25JN1ecvBtOfZKZV
ApsOUENVRE6oqwDklaH2JBaOp8okwY8huOhoopUROWSxzGwWWwaA82/vKsRsh90N
8hF8MVWqfCKbiEYMlqYIBEv6zGIiybrKFldSG5jnqCpR+C5iKgB8tgabABt07Eme
S/7iR/5Y1FMu71GVofzwGHIgdC07S5gzVLuHMPDafu4cnRqi68ZkTUWdWowg2RLe
WEHZGq5NgQ8UfA3dEezFknM+96xkSKmkK58Mfl6ZoRXalBKEypTpTMlfjrQ10Ifq
FvqnT43weuw7QjHnZkDTGMqeiiHfR8pT9u0eY5DLg4Ob2F8HNgwKTZlQF07KNiUR
t1xSkpHg72QfhKeg1rdv2oEplEX9Rleas6BBd4UMgIdRGdwUpb66+ABA0AHPBvyC
dgekB2AlQCkmkB468eUJFNbRKXdsvfwQ8u0e2RhPMnbLhWr9mrDUsP4e1klhQqwK
5qL7Z2TdN51kxtPVEQB9hjjElzXQTci0bXc+Y4GTDT3lGyt5TGt3c2Rfh+/eWtIx
9cvbNNZBzXPXWMxsxoyqdDiPFQdc982Kgs6R3cN63TSINJs7tduVHJKLSXWyK66D
kBEbP1N63G+AUjFsUpgnnQENsxIzxjKdXHE7EQg6eNPQlrlPzq3j0blZXzx6V3YG
tvVJrvAbh1cd7kwPNBjWRfALUT3BCeakfAS4ULIjvOApNVl3CyDev/A4zt0kNVvR
DWfIKL5YSPy1qktoYFcf98Lw0b6ym8EfrPHkfRYpopwfl86IPH7ggvp7V6cqLIbS
Hz3YZ7bkMzl6Be1jw3edcGVVBfo5HKDuU6b57mxio7/WtQzYMHx0Ucrvi+fdpcSS
C6+00uiGoul23YtDaXlLBfWppgGas3GtCNk66OcgiAwYQ3/nebJ8KvCQeD0DW5RT
z2TC9KP0ODqgrxRdl9wg5i5m6PqdFRkeMRHxaK7ZiNsPY3/R8GTG3fPFfomORWJn
ES788Z9WxeZEVOqfSSPEUovb1Nxl8rRMIqdZD2rNypoAeMoJEK9e7I4n3GnKi6dz
SIm/ZlDzAKAXjAFq4beQhx1u3rBz+b53Vp/1yYqw9rnzquHHxoFomuU5QSPng/C6
O2TNGw+JRFWowDUSbcdfkYekaFHhXPtaMYWLaxsbCw67VOKcPMUmrrwcpbt17zT4
F3dLtyOOrN63gBD4928Mt6ktmeezWtlsJhaka5ILCfaAz2kzasFzifOL4YMWJCbY
dVX0Z22nhfMcPDDeRAyRTm6sSq0VdGo7qbZRm1QgVcGuR/hbY4C2UHJ6OJV3/C4R
CcuKKgnvXdSG80NgWhYrFWsJ3induKCLMbz8YkTF/vF3k9HUtWUB+lxblkCXtFNT
+JeTjQeNzdA2g6tg7Nr/7sH4k8y/oFK3wA36sqJNUKDNVdRel8dzVcp0EcOhTAHs
XAUX6owvjnSddSdXKR7ikA3ZSz1+MbX2TRDeuSyICFzfnNiZXagGEfUvssVNwg2G
rM5erqjg6ZbHq38Rl+QTqYiyTGbm0DowmfJgZbbqDyF9K8iWlQsDoWaSC0SNFLBY
3WM429Xrr+N/h4pkZ8+SNBA1TAZMJe7bS5dpi3SAyRqQ0YF7apZbjF6qqa0cV+sB
W98+9cR9jBg8rYk9Ayny5ZRc5H0E+mA2H7xbREzam0nBbe7sOSpO1HqFbpcwRj1D
e/xTTxd8UgDZNfyCzY2h9DY7gohsdT86nOAPwusk9/Ua4FY5o78fDVMOiVTosERd
jyZd0JsrX41kDKC1465jQk67RSo4WOup/v227+suqnqcjSyETj7QCqv/M92QoqrF
d3CahD7S8IGdWJdojLfs9Vnn3iHdkdlVnc8ZHPnKjNWzuz+3ASfnCR/nDWKnHBnB
IRRI60UxCAN9qLFA1ALK1/OC/zRQPHASaTp1EKoUJlC3VV6IJ3rLaNmECu79aojp
2T9BCeYd49i+ol6pRuFuT5f6aO/Dfn2j66MLqW/hQO22UOQWqsQ2ZtL7yEerD6Ne
4d+nkJGK8ljsotM6lH9DShIrqdob0a/E/F5Ty0Z0cGQCb6FJHSLl5sA10axozqHr
mm/DLysWRsX+0OMHa6CBCkpyBEWBkcLKA0B4JgNUP644+CJjMaQ/bpWbyz8/1CjB
bomQ/fZdla05ZGetNR5YvCtCCw0FgH1ad7FNOEs4pAo0aZQxSHnOG2fdRxgVScgJ
1rj49j1kPqERANHYturczGRgmaEh2D9zPEWPwNgvmbNScB1S0y6hIjaGJj/CZqIm
F60Gk54B0621c8NjB28bRdh3DJBtMS3ORmh2n3ypeaITIYVqBzoaHHb1mIZ3jMSP
vY+QbsMJcLNGFdsMTH/2M2vRGHGk6mN241UimYTAvk+WEsRJqJqPFd6mboECyrqg
uZk1TNLx6lCNAgdarrnlIrGxw43Hv54bbANFRblYkfSu5cCPOmsiXjY9skAiQYJI
QVW3H3omyXyqOpDk8ub1EnAdXvRRJh6R+SgnuwOetLSVTnHkA9tAj6GKkwbUgbJy
csyDFTMTK+D0vD/YGDoTR6v0LiEOs61an1TxCpDgir2tLxAaNy9vr0cEG9oe6nJR
rCPupkychkyHPBCnWq0LcTBovriuWwdggpypT180vKLOhmudTHxtxIuXIdxAS7Ms
lSo6oO4qVpUSxKmVp01OJPI05ze6SSTmqMIZtEgUNX5i725mY7O/ju4QQRMi9Jfk
L/ybBYPxz/U+WpxObIvnXDHfJ/ceOS/qTxTdEplVMXvLYKStllUlIV1653bBP9Md
GgylyXUlTAq/KQS0dAIz+iwpYiyWJtxt5Ku87OfyCFc6MovVVKs30ZiYRaVpd0OZ
Eyv1k03yWA9P/OZ081N8/TwfoYSBHgmMR2yBx4pNjc2FjmZqSXSXeZwetTKopM4V
Tay7t3SyWC3SonmoUXCuXDDQnlLLkR9qzk00fPLH3ytz14E7CdQTa5S0VjHC32ZY
1oQ1SWgXwYCr48hho9ZVH3NMKYpnt6s7rMuepUDxJoQ5+AuvslR2vGhni1z/zHOn
16jwt2Mye5RcHjuHJ6u10BPYPBu7PwntC+YJYCI7MDOXHIzoqdlVgwVEJtiUHabX
5NU+c11UBc1Qb3YisbvxT/7z2LnlVBpxYMWV+kbdVu0rEwa+8o1c3Q29ukilNg4X
o7gqPIMyRTCwVGH6xMXwxzBWoA7THHVCvTa7Dsq3BKfdUIH808vtaTyjlUBo5Kgq
5X6uuYJXkQejZa+4iL9Ipbe6oQaQiPOJ6zOkH9o0jF9L8WTOB16h2vuddMCZPr34
5eZo1zvwnL1AOVHgdevKMdcZB5Ltr3apM6m/mBMpRr/s9xNXcnW6Yzkh4aNFLR4z
c5FV6nwk1dlDP/EjJfecpDcV8VdXlcFc6GYQVG5TEk8hn6mXZ75oxc/5VYlSkqt0
4tGDtWRCTkCEJIShte02ZpeHu2d/S+/I8f+ov9+pLenGXHSKYcaCIZs51uhG7MBu
SIMsGCxGztm+sJm+Xp0H9pSUzth9ss3IRlSi957zEG7PZUyOar4iv9KAlWDREow9
UxqbYXvr3rsVPDTJJ2RTuThAZ38xp7EwrwRctDLGrij60xwC7iF8QTR0rko3iIM8
bFV0IdrCHEJthkzqxvZ8bowPYgZ5ASomNkq97AYV8njCL3JXOzyAh2r1s70zOVbP
TvbtEwgjGQhNhxGJrVIEUmyhMX8LtUiZv7vXCXGazZ0KnBE44MD30tJVlFYDBxCv
M8tnexM1XiiNRHvt69uU5GbUyYLArJKBO6zD8oKXpC2BputnFLSrQGZEtjQlFNlv
halbbcTBUaSTLwmPSiwUK5xPfTnHwfaFDbZ5wDsBXjS11n8AwK+C9IfO6Yb9+zXb
Tu3EYqRL/oDIYLQgekAQGT7arDMw1kdHRGPJ4kq7GxoH63RSvLFCjc8Z4GC32Kjx
12CIC+QJJsXuXa9IfAJWCzalI6WHkdMdjaxWNv9PSpaDjqm08722iNAkKeQJATjZ
Fb2LW8y5dGQ3ykRADJktKGiGBlAnOQ8GEfKPRowICBGiqH8EhT7PaOjqpFcsobo/
1hVIWicx6E6JpfCPtmVSdoRywCl4X0cBmpLU6UrhMigmCTQc5Gy3mWkGCSz69gu6
CIueOtB8YPqRxg97jcbxeoP2wQ1EJPniPbgaHOn3CAeoHxllc7umYjvau4H5UD/w
RBDaklzetVoJPJ1w5lAwFdM9dKWMESYIzaJTkkBEGQ8vbBQulYczF86FTFBbQ15L
wxHncFBV5aa2XdGIZchhYOIzvgmiUq3Qv6hywHsBMulDcvedEefE4guk8s2YmcpS
5iNkMuxuANhZ87XXvbkr3n9AlYpI1qFGqHZyN7KCYkaVV3UTgxMzoLPUAjLzcca+
hYAxizZkdT/z2wdn56fuyngcMPZVXN7Vj+dGLxhwBvfMPP7K1fSoPAw5oTjmO1dj
cUjxrzXKB1uQUQ9wGGWkxGLiWyPlKNk+YY1NCzdaLG81A+AWoGm3pU4fWm2risGy
0n7SYVzzaG/Zk/BrBfZ+DQa20OqrVauNBtI3/jk7FyKvHDTmx4xfT0/ikQbdQekN
y2WympgYz+pX2l83uPxlRkcBDtdUcvp8vHEUAbfuaXeXRxJdnLATr3zXf9hNt+y+
M6+rEPxGyFM7NG0fmt8ENG1UNmcq61BtzvI87uoFL5uHzoToh5hPBxWBnf8728mq
vsjXv3WlAULKuu1IQ53xfZjNKXoy1k2QaDyFXItQIX38hnWV5v3be+nJOY7D1UPX
zkSDmGVjaehUnstY+62tneSpHRtHtWxwHANeN+rG7JKgyudJLIgAX7I/g1hsnRrZ
X15W5ps46Kh7fnjQj7MWzftML/0WDYCpRRj4ChKEGTRrkZcodp4GlSM7SUJdI72G
/8nsLtDV3JMHPqF+7fAx07shSw4OqByChoBK5Ji1ahxHQthEHnZKxtIf/JtNudtA
BynL4aPh37vtcbIb3k2it+yoJwQIBqGf8dTEhINzx5Il2VGo33KY46zKy1iy4Nvk
Y4ZOHERUfqqA4b4m6ZwbXQG7c98PV7bobnSku8Me1HYkmrwdfCCNTkGIgwH+PY26
nBu/M/auvpanTj77lz58P+moeVFm6HD+hYUI8rbB2dk3ki5iu4+V4xy8FL3Hn4dW
m58XMKJK73vPUt2LEcW9MnOi+y/DLnH38/sYOeUIozXmmkUbDBef36X7bmafMKng
DwKWGb5tzFCIjSgslyH49NSO6d4LEOy24ryt6q6AXCFK4AbLL1PZ+xetrGZ4OYs+
QbXSQeI3gsZMLlt9MxtI8Qscl75+onc4k9YSPoFXVZ5Ep23aUSGhKcOBVJGdCVqp
0o7/LN8V5B00wzCUZEaxjT7lRlVZcfBiK+hDexddZ7gZyyuCN9WbLUVeG2GUxrjJ
+6I7io766Np50V7GQ+MB31zNtyaI+c9Pv2IFwb5Ek3QusDKh9PiWA5gNoo1AFIJo
th6KnjKUCY3bs93umzNXsv+NFbNUyfauTgpquZ3Qs58zL3Hr8+adPHZ8eOFG5ACo
MhOlCDjL0SBuru6UhKtFIpV67iqXAs/R4S7p5YbzVDzuEmBLSuzjyb49b9RU7eTQ
K/stR0/JQ52fmDM6EX8882PDwRMLwdxL3i2gyPeAANNuIjsot6KTnRD8Hw8hQ8q/
QPKMn6PeJTc8+bWkvJxLf//f8gVvSbT7kcuz5zhQ13SkgmYkcn9AxwDqADMndF03
SbiV3a+phULs9ooQQVhis9AGpZ3fD4OIs8rT5VvTJ6ozITQJP1eWsg9WitLXBMxW
pLo7Yk6fVauKsWPYqs6/FHPy6ndPOVQWB1YzWIa1HQRuJHYbMM2uyoD9SCBPUD75
v21K/5I04qkR5kK82icpwSGv2qjUXMRKs3EnUq4Jl9SdFboj0833HEkc1jrK8hpb
B57vKJh5bvjehLRdE1jFxSfOwUswkkG4XB93Si4YHreWfstB88MOV8HFToFI8Aiu
LcTR4gCXfkyIIVBAcN+iSCv2qSJJ11d1D5Wh2EL8jiY8lPkJH6pDVp14BtTElfV6
/FcLhpNw5fIFqfma7QrO/o0m4cKYQRmGFKYIEhUMfiO6I7S7NUwZmAsUfoBW0sGH
qDRIWrPetYFRLg1yCjggrNiPrrJGtK3dY0hEhgRSJjWBeNeq5h1OHef5VL8DQCaC
DVYu2tHXZhxi74TEsMB7kmX6YkbyJC70Ja2CYtZtyRMziBRDC9EaLnorBBAz8JnH
doib/P3PpLyti5ApG5VPGIXOAgdr9IKv/C0l+xM0zB3AE8WYqpB7b9fooGtmKSDl
jqSPPGUayatJfQKOAjzU0F1AHvR6JLTsETos2ReAoAfGB0AlM+FK6V/6c1/cxTZj
bUiML1pOXW6O+zt9hIoGEG8sEzPQL+kodYqIBdpd4DE+LHTk9o17GkDsJxFvfIdI
5/7tOG6ELMkYwjX3YEVf6yv+8jJBqdIgzp4oDySSfyssegwuevOXGTB4BTf1vuag
cfq2TdPC3epKJ1qjEuAfY7vIO7SVvfIuSXGHcIfHFMtMq7GW7ilcfOsAp18zs0EB
UeRFk5lD+/S3vkjqivKiKnQv50NUp9vvEycFeHZ/+dwY7Pl5dwLMlP/Px48CH6MC
Jl0uaagl0PXST6XdxKBEznnbmcH16Cj9Cul+NMlOV+Z8dY4knnDAo9EzK2Yfeivj
iD2roX2AjyePHWPaFDnxRsit9T8Rfe/qnptn9ucoRB6QDiS8y68FxXdnRja508Fe
jXcYLB4HMbtf3LXavkPxyOidxfhuPtmTA6dr4xdMRT0OBbFNjhH3Jt1N0yoaNNZN
iAqr7almT5ft/Y5AeJGB/GGUqdb6rTWGM1YIEZ2gRoU0fYxI0DIrpiQJKsdpIV5C
pf053RfbtRzpslSYaokz+3LZDBO9xB6Iqssb1SjlDf8yfhu/+MvJiWcYHr/rk10h
HoHDa+VLhgJ81Ob9psr0rpjovwRfpBIRThoSOJ/Qmp9dic02FzxKtIQUyYzF0gHN
Vn4uicLw930NXFkBcovfxeUJt0hqnNBDQs4b+dKyfO9Jp1EIYxBmxJZiMB06i0Cb
xrgtVoXOWOSL+Gu/pClRxNoW5hTGgvU6Jdof7P6PTIZECFZHKZaq51tPJmJp8TaI
92WAu15mENElOR3/s8HlZtkrhJeHCF77+ZFjADbxIaypXyxK88RpGSP5WcCPvEug
AWIYftsNJGLHfh3QSkqfxBP/j6vTPUQqu1+jNM3a4AZGvHEcLmUvLR7RSvyq/SWC
gQ5dAJZKvhA75sm7pM4SlR5gOmWTmzOZoZF/SF0Q1/km18W3b8xZILO9ehfN01vL
U4aVRr84OXuc19URVtzo1sqeLQMpZYTK0aBETS6ge6dwQpMyOLegl4gw+xA49X5+
GjFXcZsNRlxwgy+MKwhpVqGpxcgVWV1QlJ46vd9RcnPzPdfqombMX1/AG9RgOCmb
ZQuGDQELBYm/emLV3lbkv9TsIdRsEhj9K7Fo5terJcLv29TSew5QMSREJmnqyU5Z
RTc9ABQsnUuhLmADVToeZslrIPJnjhVJE51SKr+KrhdTbZLxLGbn7ao11AutrWDH
nzSgbK7RAWsOtfzgiKopxhpG1/QU4F3txts1J6wOK8qWK8MZbnEcqLH8PlQ9ZRxr
/7v/McbsS5EpNDuurSUgPu0WyM7y7KweeQsA3ozdIGfh9gSuzU8QsfN3xUQVjFXX
JbTHf5WWpNa11u3tTNwlqYEXSqy0+gDrtNNqIg1ud0kV1Y/QHXKIDCSMspFennCo
Vhpnn8d+FzsxBL47FaQlvglYYh4wNOSc+8CJIBt4BJp7bT03PGwy92Zj+2yvOBV2
nYl0usXRpDNeQ2YoK9hTmG+MmzN6mbNGMi6iTPbebQMVNRsGAgQM8om/AZUj/OJ9
bZBcbTz37REssPT/5oiS57mqOX0v3R43kPlKwjXffOpiWZFyssScn+v9Tp2d6KU8
QtZGmPH62y3iMVsrawTJr7bc0C7ihr0QALeOBHwtdsYxBHFiFpIbWHIboF3Uuwyl
miAHtx5UhVGHQtcjS9IbEY561dsAmuXD9YU5rhwJ1fETTVgR3vFDNxO9tmUWihDO
4YNfmKIxKMiFo3xDz/hirQ2LlJCT4ul1E/zyuxgY5SMvO/8nyjSwO6C/xliK6ElD
hZj9KJg3xUoG4DkBmpayt8uuNyB1morNNPGTvv8/0z9652CBBKDftebiYD1/NX35
Cum0fg6zshSeHgasWUZr4N/fX1X6JVn+OuNw3zQXtnS1O/FFlpOLKGqIxogw7BOL
s0JKBp8hfLdEprvAYsbtEcr6Sis7VcxPU5Le+jB9nakzRTIgpWAIzLyMGbqk40t2
hqogcZTwKxDgx9SATAGvR2EI5CU7qLQX/+/PctXNiFp3xBjkNHVWroSKU3eB1zx+
qgV82DJl3Xc8FWaiHN5hVjqsoTLFedvEsHgv8XptDet4a+dacvZbslVBKpKXj03c
Uatv9iYOa5pJ7I1J8yXUGG/U91V9v0TklvBNAfNWeNk+mvSOd5EHthoarWhJdyzc
ciuHuCzRAb6fxUh+Gd8pKvAxljkaEDqMH3VKwvGuwW4YYcStPrQLO1fg01wouDjc
4Ly+fb77pEYDNL0NiurobRWobHaYLjAUMvNHI0sTVMxie8novVl4i36lKFSb0JwD
uUcDUtm/tPzfiVqqrVqL1NJpXs8kEm3f5ySN/hr4sAc4KHUSEL67klOtvBj2dv1p
tBukmzfROU372h/Avmf7vg/d3djkz8QjFbHc4wrJnmHCMXJCuQNSNBPt2uqOnYUG
Bg5sqr6WJ1yxG3lnaBGFZCUiMg+7rmmnMAsPwoPx76KMZdD3RF/oFEWe/s8nJFtU
t/1RB/VE8kyEptDRTI8CtRQ6Q3FoRGYinPC73wk8qweDsKbdwvd9Wn8+BQYh1Y+X
e4dMrv8Vqa2TA1z+DgHKL8NInz37XAIf0MjqgTNaxmJ16kOlhjcI/uDNJvPBZwwB
xYnbc9LP6e8hvW0wRYwz1Dq87Nz736NHVlBzwjw9opWKuTWG4rRN7k8B7CgKNl2a
Zhes1+KMZKRQxD2xf/B0OjAIa9mzRFuhSvpvjEWpWqI2i2Dm+gsxd9J0ml8ZYLX9
CvvSckPJtk6sIGbW8ZjWYXPoPxqDfLo/3tXOdO36Fd/yg15wBBLVU6KLaASjHwCD
2HFhZXLmNJkQKbge54rsHLgtkQ/HEDNRIPwaKLqdC0v6Qk5b/5sF4b54tVnFqTNE
ITxUrrLpEu2wx8ux1xsnJYeYtO1d7MbJGzI+dlmEy4A5KgCWmqjg4NhPEMnt6r8F
5bRY0radkjWgNylKeNhmEjgD15niSaTF5IC1PRY/MDa1WIR+Qk3qeLLZiNs+zrmu
oFHzRYItLgjhdP3F1MhIqbWr6T2Kmzy5KMuYUIL9VFlrX87qPatpDEPXeOfW3+uj
SDJO6355I8dBziBtGFEDcbdqP0TwUkI1yUBZdfW+/Zesp+gvkijdgmlzX5WQdQcM
85RGst6uiQLnLHwrUihxoOvghRzp3RzZSOeBqxSsBrrOfcZ4/SycpbHfojGUCGnm
KdmdUnunxx9MVwZQijGfprTzQKFtNDnE680SO+d8AFTMylCbBhdrCYp93FyryxBy
os86HYip1fGCe/grbcxgXfMvcT1l2xs9pb/Ba2+MYP6eBEXNvndKUHO4B66h2Dy2
JXb37NyYchxakQ3/VQVJSOKSxt1vnM0iC24sn6YDFOsECeQVMT8mW9m5cRMEp/KH
xTCuNyypXPSw37aNiD3zQ1Q798Me5EzQM07YW1VJ/0mthx/IAndVnUeEgvY2D+5+
Q6pG1zBHSKaXCF8lqJhkk+F98f2jOrozUfz9K14tY6Y9l07xsGdhRhf6k1wMKfK2
nkbkuvK8xocJxlydROk2C19DaH1nazUL5komnmuJqPQMHNTjIQLl8i5iIRcugviE
9lW51CEfUfjOy9oKIRmOKNN/za2tFMjKWQuJ0nVJ8Y0wCU5feZ5+pKRoB4s1sDVE
/x1UWNv7LVRC3xzno/4fTXrPX36hih8sj+du6iZFltE=
`pragma protect end_protected
