��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O�k}.Ż���"�����x�u!
�*�*����K�f��\ �<��nFɚ��f�.&V3�t�_z����RZ �UP'���I"���U�ϓЯK�݁/�G�5��#
/���R�|�1{���_����,$Gn���G�M�J]^e��Zd~;Rb��N>@���O:G��Bj�C��SZ �K
geK�ΩLS��¨��
O��r��EYщ�G~)���v��<@��os�U�1a!:����;f���7�J=�|/a�-Ϫ�v�!�Fֳ��B�%D/�Mb�%�,�=0HCЭ�����/���O�
�m�?W��!t�`�E����u�d��~Ԭ����#K��{����5!�R\��b�o,�9F	�#P$ �$�#Ѭ1�N�Wb�ƭ��:Ep8I8�ϧ�5�H�%�ͣ��p�sDT�ZK�����#l���g�6u<Q�|�_� ��
�^�<���{�}�^�p��@�Q�`@k���Mh��E[3�Sz'�rI1��>���o��`��J�"�C�/�~�f=-����n���w��$���o��H����Į��[F��/t�%�����W_��5����\,��r"��x�u��p�����3�b�;�k	U�<v��� ~ͫ�YT���h�{��|�cQ���&�=�����wG��L�i�ZL��Yq`�i����uU�gu�����@vZZy8�):%N(�󏃎p>kxe�5֪���d�%��l�7������n)2�*}�`���*֠�L��n�g���k�-��90u�:=�::c#)w�+UX�K��$�wp��r	��ED��5���!lH/��?:���̂�-��GL8SI�3�����O�Q;��aΣx���� �.��ьnR�2�d���y���sըf5���#�go��C	@���w'���&�u�Mg&(�+�3Ÿ������3{7���:�Nƍ�ks�����;&B��a�!B,�F����J-������ΑOv�H���r���[���iɻ\f�8DG�#��K䖖;��f���<w$1����x;�,7kh��QN�{�	#�
ԋ���3�3����x����Ǉȷ:RS�n�2r�� G16�'���TZg~�~u������W���u;Z���f�j�7y��볱��9dbI��k��/n�)�+`x��T���bE�Q?+�O��!-�f��[��tݴRYM�E�2,��S��ݔ8š�1rk��z�i��`��#8�^�ݜ��,�y\7�|����ض7����&Ʈ�A��i	��(
�nO�7�]�0���5(��Ro����k�|�M8!���2Ow�ȣ�ph��oEP�"Y�Ȱ��m�='���!"�H sz�˦��i"j��$`�m�;E�t8���d	����R��o�X���;I�h�^�,�� ~�s�]��~c�!�s����Py�)J�ď��Y��҈�qh����e�J+	�P��a�sy$�V:�'X�<Q��󠙋}M����
f�x�1GCʰ�FQ��8�M�"O�Hƿ	�D	aꉶz����y.�&W���������ٙ�y�zU8~f�h|U{s~1{&F؂�(�*H�Ӏx±=�ŴgE'��iv�D�����D9%Y39�?g'zh������ARAo�V�6!L���YhwZY�t�(�̹��:΄����ݞlތ�X�&����5�.�P��[������^l����C$k�ǹh�+0�M��p�gI�f�b�9��DN�����DF�����kn����̇�:Z����t}��a<��2���^iW�p��r������(t���B���pen��_�k�Jb����
{nI�ݟoHʦ���k�}%^�F�G�n/z�ɉ�b �iA�O@hQ޽o(��QQe�*c�@�vC�M7�o_��>"r^�T��U���2Q�+~&��]
�T�)^J�x8_�a�.%��$���h�X��B/��,��=�PM�'��C�#^1����E�c�ѱ+�L�����52�P���"G�VҀ���X����tki|Ķk�?�݊W��~'�Bj�r��Ѽ��&�z����'�-'9����dys�J�l���S�}xO��O�9�{�q�;=׹n�4�W���]piv^g_�MQE��mɲ����-�����6�[�v6�^�T#�#��0�1�s��L@���W�����3V6����I�Zn�<Ti5�!��B�E��#�7���Q�׶�8J��d���NB��%NwJkn�UE�?|0K���N����+��bt�V���� �ʠ�T�2]�K�Yr� ���}ff��J�Z�X��:���D�Ο\���.$����+1bN=a���w��z����^��)���^��������{�A+��бW��ױ�
����C�cD*:|�`$�W	�̎�?kh n�������g�r�}��g-���ggⱵMCe��ek;�T�\�]��J�j��+�,2�-��H~>�b�Y��e��Y9yc3�v��2�`C�8�g��x�)m��wm��#�֡a
[�j��^�'{�[�O�E��4���L�����U�yMw��.���� -�P�h:��\�?WN~�/�{��9�~�C�� z���~Z���Sv�bܤ�R6eJ�h�	��^ln���P���L���S�	����OԈ�{A�Cq< �yN3��>�m����qT(�yFS��pt�Zt���]�ؔ�$�*�49�<�`��ت,�n��L�\6���S�5�gY�u͐v�T�-J�u����7�_�x���t�R�/2��0X��I6ަ�苗���2�.+���|	��g����֥H�I	�����s9��?\�Z�f��+%�v�t�ޠ9�Z��7�b�	PQ��!�~�|ó2�H�}}'1��ݰ��oPA쪐zO�qh����C�d�g@�w&W���=ס��f���'�(C�G�Mv��u�rȽ�UpӦ��E^Mp�����y��	@�d�Ł껋m
�0�H��ʙ7+���Nӱz��l��5�1���.��6�o��/��j(J��<k���ݶ���i�]��2�(��"N���������8�y['���ѵ�i��/X8G|F����ŕ8<#w�	�|
�4݈������r��3��Ln��������]"d7���+p���P��^�ǝ�Og���u�q�߁���\���")����,'���Ny�x�˧�S�K������C�d�.7����* nA|L��Ƌل�G�8����d:�c^/�ລ��,2��]}Ij�ᙍI�Q|O��ⰌZS�R�S��F�����4��&��<H���Iy��!pᛄ�+����\���aU@�s]X��?g��87W�v ���G��n9I>'XD�޶�}�4:m7V(��Ѱ���d��M�:2���b�?Q�?CL��Z!����U���,�~K?x��Z/�Z.���	��(���6�?�?X������W��E���)T�X��_�`<�&�V{�w;��퓩���-'���sަ�6\�MYk�7�̾�/>��tF�����yt�֙&1���M���9����[WÝ�U#"�F����6�0�៊�k�:x�ܯP�෩oR'�s�uS���ޠh���	��m��k=6�G��C�sN������1��-%�9Ȋ�-��;y�\8̔� bcޟ��x�"+��*������S=��GH^!�vG�&�zFU7����ŀi�K��Pڹf��G^�ܲ��X>F�ά���ے!Z�UC�7�{�-�����@F��!H=�`{NA9ER��ū���f5��v�����}�;g�[u:h�;�K��.s�/G�!�a����a�jۜ�e�&�ɝ�m�ɷ
��5�D^o��F�$�ˍ�G�JFx2�q��{�$��v:���(�ϦڰL�q=`��A�L��@���{�~u+�šbvi�M)  �i�p:�^�7~����������\�С�	1�0��Y�{���2���.傆~����QL4����H�a��W���-�և��zVє|���NI�d�"W3Y@����CvF�#��~@*)-�G��䘹��1�>��.���!��X6S�i�0�R��Γ�ת���4m7X\�l6�b0[(�5?�t��׻��p�X4i#�j���`!�N<�I���D5tu��]/��碑wa�4�ƽy��}�Z%�Nv�&���E�Cd̶�E��e+��|\a3A �Y��].h��M+��~��R@�-��a22��H��F�`K��C:2�=vp�CЊ�Sb6�+A`�]�]�+�����c����u^P�R��+�GC���)��u�kFߜ(.Uв ���
xl_b�>S]C�K���v�;���J����� ��>5鏾������ȵ��V�V�[���n,�%�-�V~���A�(Ұ}���
_ X���H+}�.ZF=��_w��Q$��R�05aW{�8���ı�VQ����ۇ��&4���Wio�M\Zkvɶ��aZ�\K�̻V`��Ї���(�b��g�D�7�3�0N�]����څ[:����]a�\���v�+P�^���k�_�@�Mk�z_�lY7��`fa��/��5=W�CwCep��ЫV�aX�w!q�8�U�TBJ���^��7uZqDu�k�G�&�:X��(��k���b1�/ԋ�g��m����V��'��&��ܦ!��o��=]t���0/Y�GS6 �2ұ�:��s [��z�^09�(��M���~��.�����4ķڿkB���t&M?��%�V�-�zd��4P�xSI��įiw#S`��|OIL+p���Lz_)%dm���)�6&E4=n��n��:<���$����{�	��.@X	��\�af��S$��St�D�9� ���C��G���<����rn��/�@���C�/���e���`�L��d��!-:���	�%�L����w~S������/.&��@F�tt3Ւ�h��y��ӏ��egY8��Օ>Y�;/f�;�H��x.�����������WY6"~*�9���x�ﭕ��À�~����e�,�l�A�z�	/�.i�a]r����aP��C�>ed{f�K�~[�M-M����h�<� %���;f��gFx�w�9ɫ_Y�Nt���k�D��ln�0�n�Og�_��MOj�Z�d�{���~%+��@#���cV�8��z���b�d|�%�wP|?+���z���[�
��XH������:)�6����ޯH��v �Q�Y�իi�#h�ǧޅ�8ݻAf�
�̉�V3|ՂZ�\�a�I݉L�~AI�k��w�������X���1�?����L�8�������ة�^xqH'�?C���[I�7+
��1*��V!XL�d'����6�C�#?l?���8F����)��%5e��S��3���]�>����(�J��}� �Z�[���Y�
79��v���4�'��W�\�(��L<-��r����-�UD���z�O.�Xꮰ�+A;6��S�x�5��+m� O��d��d�:��W�kt�Y�a��@$�N��������#:��$ب�v���<ʷ1��í�ܤ���Nk�N&$�����L=���1�}����sԓ8'��5��>��}��s�&GRd�az�U��$���v��8r
}_��dA׊v�ls��^XI`e��9�I�=��;��+���J#P�Q�7��Hv�-���h�pJqETN�)-�i����a�2!^���o�I���r�_�3�P��Ź��� �;����3H�@���Q`i���#�[�1��b$'sGd������@[��"�3�G��������N�3�t|X��`�\GbQ=�]�Vc��?�"����CF���KM_�$�!��>���-�:�	S H�>��Y��u�<���Fzߩ4*��2' 3�9�7!�^k��?HV�0��#�,dݦ����ĩ&X�hl`�KU�z��2�����BQ\�0����7L�C��{��tf:�G/���r�D�=����X�EGu@��6jL�޿�i�x�!�7������4����n����m �u����j�#=�m?=,
5�/�*}�@���T��:��ˍz}�k2GM���,���|�wd�4�X%��yn��O-�\��x5:0���LFo{Ӥ뚣�f�Ǡa,�0�9�l���-n�K��z��t0��msx~�� 5�#����'aq��4�!@�0kc�+�i���ȦW��"g0I�2i_������E��h[s�
$D7]��_��1^7�hϠU
��!�|��^�LE{���,�κ�M��^�c�=�Is��G���M�
(���L�Y�W���N�$萱Pո�m,ןR6A�Q�pk��w�,�w�sLw�|@�i���4�\��6�������X>}mu�nƄi�@��/"�+�� �����w�wM�/3mbS�������Ms ʹL[���,��X/X_ B��y����9�W9l<c��� UO��S�zmh!z��o�(��<�<#0V{Z�Vԟ�R9��Ԇ�ö����gش�_�(�N�����o�N�i���c%�|���y����bz&J	<��~���3R��=�?K�g0.��sr�A��d�Y�n�h_���v�q8��(�e?gו����L%�11Zq㑺A^I��t*R��۸(z[}�I�>�P4�� ݾ8ˎ�bD�VX/���=�uo���M�;4\[@�gs(�������x�r_�Vq�xĤ�S�kք��.(m�4{s8F^���_3��B������N[��Z��.8	<��/�%C Y��뗢:��K�z�B�(4��'4������-�2�3]�	�r�� i)�&X�v'��KApN>/�=�g =��%g� Z������о�-����0���L�,���w*���T�4q�l��}��?;/�T$��fV��F𪍒e�5h**So��y��*��<|���柋i�;K���ԋ�:���>����Sֳ'�|{Y֕�b#CS��e�)/x��f2T���[_+\�Y�w���/��U�Ǉp��X.0#�
��w�C����qiZ:9gO�b�)-��1{�5� ��RBӨ�>��H)�P��R��gbI�f)��q4�P�n$�W��J�����\}ԃYY��3�� X)%�r60L��A�����<�\�+��3������w���*���|zWv��P��-B+y��6:E����;|�?�f!��������0w�6�&yw<��'�>lC�����c��MP/7����m;Nd�����#�^5���N�t��"�h��9�*&�n��_- 5��[K�*ºHl�H��l�)Ż5W⊒���F��'�Q�-�!\���s���3��A�f4E*ċ5Ɣ�$���5���$ӹZC�S��S�)�~���$ �͆��E���V4g��%[υ�1�t��	cX��F%�G���45���ۡN�#M����P�����iS�Ԋa���{#������N�ځv��P�N����m�d��'c�՝�� LV= &�5z�B8��)���ufY�֮v�PA�H
�7c��������W�����&0�v��/��	�xVX=+!�.r�^}00���:�m���3A�'��hQks�9�b�L(�i���
�l��z3Q���]{gc�n���I�"{�W�
�Px4wT�ԍl�@��pxtq�P��s��V�:)ͤ�7���,o(gGlC��nƥ��-0VT��#�!D��E�4�5��ˤ�0K���j����]8(��bj�J�99)�n�p����������� m��tV�S��<�I$�aQ�M
��YH]]��̗$@喜��{Ϳ����a�# ��v+�U	YXi��'͓�ۗ���@/e�T�Y~���D�|ۅ�>�8ʂ�\HJ���|�˹�q��W�s���L$3�S���D�m(������Rd�X�Lj�tʕ4�r�J��������y*����CV�Ԙ�M����Γ��U!uK���x��էuA�����^E�	�*<�������VAXj� ���H���?: *�՘bmL�ǛM��<ϋɟ�WB��h)�\�$,>�'%�e��@��l�ij�p,�O�@���;�*b����g��:��6����ZQ$�RKL��^N �!�<!�K̠���I�X��ߴ���l\�H�<l�c�)�ƈDŷ����@�-�ʀb[Bi��+��&�l��?jz�Kzd�Ѭ��Hډ�+�Td�XI5�h��q�%TkX��R�Oy��<�-Β�Oc�G �ˏ��x���Tε������W�%`J��9�"#�-CC��ha]�X�"�u�uE�� �L�j�o�Gv�}��,�H���M����"y�S�:F�.�T-�g���	�j<���� ��2���4��ֲ"#/H���NU^Dᐶ3��@5�+�H?n��-VN����>#��@PaB�c/��{	5x��u�$��\f��������J�cZ����b	�vS�j6��L�bw���K�ª�Z�-�3��"2>��X&-�)��&�F(�:��t��Y�=��j��=�'
� $4��Bz,rP������f߸� 
˜��ҝ���DA���Й�6L $#�����1��?��7vf�һ}TDU��C�F�F�����ʸ�>��r�~����~����HBc�-�q[
Bbt���"�X:|�G٬Vhob$�Q�0Nn�l��{�Mޙ-��mg{�����q9��pmw�V�����{c9
Q�~�uz��: �]J��C��v��j�R�T��{��#|��6����� ���pH�G��J�.|n�P�q����R(1��q���I��B��6�Ul^��>��JN�7�]�U�$y�b�0}��	ߗV	�b����[ڠi�����Ncg���G��
u�p�rs��i�)I������]S�)^W�\��Æ�m#'�Z��<Ȕ���:d�B�l��� 5���[��A���,t�����r��\�U�¸*�""��z=V�s�o��������uO�)�M��MEf:��&��P������+j�}Z;����+��^^t�4v�cb�bփ�V����l�rqC T!��Z��5	�h��{~N]�ae�N_�������f#2f���-mH��/9a���,G�M�7)�����bY��-]R�C�<CfXofn�H�(�Ŵ�:�Z17�Ů��9G(/�b>��j��S�1�U AڲT������ǜ��R�e�W}L�� _��mV�~�,9&�}�8o��L��+��܆"���w�H+�ND������
��^�!�#6����S�|��q� ���	����Y�ӰRT"�4����JM��k}!�v��QQ���+T��D�k{�)V��
����o�K��3�w��:��!Jn��]�wFd{�>.�}�$�E�(٩ӊ�}RS��m���1�	�Cy�MP�+�&Ӱ�:!=�K\�ܝ�@p�0a���9�$N���TԱw�r��-��u�[�N�y��͓�{�C�@�����w������1�=����0>�n, {1ms���h���.2�Cྖ_��vsEB�F'�;��(��w;Ƞí3?�d-nr��׉���e�}�GG@N����)�<�������J��g/�����尪�h�&0�Pm��}��I��<Mt����m��{9�9S^[0��0HM��
~i����հ�J��=p����8�C����G��4���bs;�ΔA���s%23�@;�<��Aę���[��db��~r)�[�)��Ti�6`S�"W�͢:������(B~ǋ�6��T&\y}E#*׀���W��������61�ҵ����6�
���dU^���F�mӵ���y6}������{���y/�ŜF!�C�񁶵I���I���Bl~������;G�}��gY�Z�8E�"?q-�U�dgԃ[�ͨ����4PYl��ɸ�v�5v��)�5/ۑ��,�c#Ur�Œ?*
����jQL��z��9����΀��h3����ܱ��k[��PhM�8p�9��򪄽_�,ޓ�v@4����?�U�����X�A�{b�>�Z�����w�gy�PV�Un��S̒��Ļn=�d�D�6p�'6E��ph7�8��2�b�:Rn��,�X^s
Ĵ���bo=�p%7*^f-yu�3��7*^��OB�ԋZN����|R�6���NNPN����N�g}������<�י����-����{`/���k��<ޅ+z)������trh��׉7)��!���/
k����QTŝX�/�PM6�l'�,H���Bw�B�)����B��p7:�#��1Z%���\�Ú��n{1�(�U5L�7�:m��Z3���m.lU�����ͮ`��¸&��HtgJ�$n���Ƥv��7*Qh�l먇��c�H��'ȘȂ�{8�����>/A�uI��7�uĉԵۈ��r��5�ϑFs�m�k���vd� ����X�lJm(���RW�٫����zæ�^�Y%G��j�����g�w�����z7�l���J��{�Av�г���ut�h��ȮK`c°�n
��{u2�Sc
Q��kR��n����F����ȲPR=\u�\��E�9ݸ�v��4V/�x<��%1����UQC��=��r��U)������ʮo���Je��Ҳ����*f��|���y����t҉�]�C��O48��
��������\�_�zUT�˖ �J�].�Ľ�_LH���+"�tKw�t�b��q"�`L�&4o"����i�喢o��3_ػ�Ԥڈ/���(2ϴJ��2.��"��7y��_��{6SI�{�r�j��~4�/�1rc����5Zŧ��ՙ��/���
z�)����l�q.�*���
����KJn�_�kZN������0�i��np��#[�
�u��=�#��O��ץ�Ȍ� �o��)D�s�(0�Xퟖ,�9+�5��r*��U��cp`�!fۃ��e�����Z�L9�w72x��;:qhe�L�m��Iޡ4͡E�%/��&�19ޞ�5�Nai�&I��?`+�7���MH���1��C��-�i�Ιp��\lk{����ųԍڕ�S�H��|��ۉ|6ˈ�A�rZ��?��U�!�?�}�&{���c^��U���5��|*�&{H�
J�J26w:��z?Ԛ=0�S�;�-�H�U\[���(m����7@!�[��/4P�:�Ƙ�/��a�8��ʿ(g�ha�W��Oǚ��e�Z�vs/�r��|g�p~�¯N����3?�N�����[���V�kGZ�C��5Y
6S��=����m�P�IO��w��A_��5S�c��F ���cA���0��$�ПD��G�r���� ��	q�0Y{�q�뒺�"G,��͕6��J{�n��&4��K�?�OE����6B �x�s ;3O
v��/Lq�{��7A��|uʹ�)ŷ�9�'�L�D��1�ۥ=�P�w��O��-�]�'��`���"2M���җ��D_�Bn|[9�@	��y:�Q�K�j�z��W��,�5B|��U=�ڴ�1��U���Kt#�|%+v�uu�`?"���G��c+��ᄤ33��c�o�X/��xz�u��]�/�l��KB� ���
\ޤ�-��+ �mAhפ.[�ƣ���:��^WW��\�0txV"5j���>1H˂q}'��dT�q2`������Mţ���O�8k��hi��S)�0��v��f�5�
κj(EgD��E�z��o)g�̓_���I�t��	x<q�~� 9R��Cň�y��{~�D~y�5��8�`��@�+Sz���Ih_DhѦ�6�xn{�7*�m�g8�!r�:�1�� ��[$�����=��F� ����($���jJC�GN�4gcD��z��̱t�"u�NTV e��3�������y��%�/��0o�~�����/sc4b��".�S$��e��J�ZJ.W����~Њ��(���^�
!��tyA����S9�L��3�/�p�|��[ŇA�{+?��v/St�S�;����G?�b̦:��l�����\�*�νZ�mhߟ����5Ћ#��-�ݿ��չlS7v&ނ��Y�>�΃6��W��y\Ư�`fə�I(OW��x��m�ѫ��"���|4��8ɮJ���6�7��JD����Һtbؖ]._�L\���k��#/ٍ5TO��[(��hH��O�<�P68����u|�P�t��Mp^-m,R�%�hL"�M.3����d��'�w�	a5��<D�VA���6��D��ǜ��� ��I�;�S�u>/� ���:�b��õ`\��&�b+,��pw����a�3ή䵪���u����ѝ*Xq%�<��HV
)&q��u���U���T�a��}E@*䯲����f���-���=�ߟ��BKX6����|��a7P�~3�^��6�Mi�qh}��Ǘ�������H�5�}��_a����z,�.���M���*5o�<�S'R�\�Ց%���j<����D�8L���;A���go��29���J�,�,�&n1�`�Ƶ]�o2�]+FL�r<�!?��koR	��kh4b/5~Fiux�3�q��#����hJ�������X�)�K=LqpE�x@�V��\��0\3��~�����v����$c{a#�z*9����6��D�:quF�{�aB6I,3�� q"���w����Mn&8 I�ҷ��߇�5�4'�P�Yb��:�$����(�()#�Gn� <t�0a��T��Rk�c�܀/b�Rdf�]h�$��(���bȗ� �jj�Ύ����ĿJ��~�陽W���H	Q�F�`����x�|��2 ��w�A�>�h�0y��;��&k[]������r�ٓ?��B0��hm�aKj�6��m%r�>T��k�9�/(�M`Ήt��YgT���d�b5gp���l�
B���5�QD٠�e����n���hx\۪�w���',��(y�J�ha��U�S:��8�ۥ���p�-�-9���`��U����4�+��O�f,�e"�ɭY��a��� 4n�~~�ZH6x���`����O)���W�t�8$q��{��*e�]	S��aB���N�ۍWM������E�鄋�{��Z�ӧ�bےU�����g�Pq�P ��%��J����__�$�P��� ��[v�)��*HnV#����A:�&;�7u�c� �T4]�^�{���s�R`�L��¹L혩Gc9C���M_u�����
(V�1��#3H+�x�p'��ܑF;F������r�dե�������Pbk�p����'H�[s�rvs�B�V"l�9O��B�(�R��V8���K�x�O����<1-�84�҄O)�i��R�7b�f������G��~�`P��F�'�C�v��cS���L�k@(5�]I�Mq���r@��Ζ���h�1�����v���4^;A��fv.�s��{76�ŰȮ� ��G�0䒔Ĵ�Fb�QPg�LDߥJ�U�(�������C�[	�"La,��/ϒu�؏�L��u}p�ĥ&vW���\u�/�f��oC�
�/�dH{	�'����?�\���4���=���l!}��
�Ɣ��;7E�=ŏ߃D��_^&�r�El�Z3V��T�[K���@�	�T���`�3)r�e@bO����;ab�$K����z8��}CzI{����͘������үRXx�Vd�(ca�ЯQ3Ev1j�L��`�ꡯ��(d��=À�n�f�$q�M�>� ����?/�{E�6ˈ���y��H�H��A��w�����yI�hë)x����ٶ@�JO��.����0,?S0����6�-p}j5�F�#Z��'t����ا,@JDHz�\��,��lB�aA���1e��n�у���Q8W�튈Ɖ���I`���j
.��D��kȑ;u
����b�%����.y��5��]=�����K����da�'�=Oj���U� 
�2RG;�q��[L9W&Eu����ش�?�qd;'�SCN��e����B `%H�;������aU�Z��O�
H+|�E�ٍ%'#C��׉TNݷe�ۄ8�Md:��.+3�	 ��Z5��CB�7۞���k>{0~n�i�}d-��9n��L���)UD��/�ȗ^�=u$X�$"֦�c��x��x�ϻ-)��.*�b�T��٥9�U��n僻���w�.R*��B*��$����#�*ǒ�m
���d"�^pJ�O��MS�&���,M]�w(�f���SƉ����{�A�L|�~j�67t�K9L��eTꅞ��O�NG�x�2k��_�=���a�H#�*֒�J}�1^玄�D���\a{QR�0~���lgG4X�~�ac�{l����h �W���30���5���:.{�&�����H�H���{ r�����,\3��y����:�u_��7�f�?��*���%C{��O���g�l�������Ȕ9T�م�o%İ�"N.T%>ij<e`��� ��r�R�G0(ҁ�.k�-�*x�����F���d�^9�!Rҟ�2���C�Cv��CG���O��X�Ѓ����9�L���j���6��<�����젺���7c�
_=�DD����.Uڔ4���#���5W/��r}��e8<w��:[�I�F����į��0W�oS#)��8Ju�Ku�1�1w��;���R�GH��1w����wx��c�g�6��L~yB��~�Cݮ�޾1�k���iS���O����R�''$�I7�,����?�SX����)�38�6�.F [�h"�n��=��8�4���)yj�X�J�A�
 JV�����M��E�B�g��j���l����Ȋ�H�C	��ݿ��.X��Ÿ���;���������B��r�DFW�؜�Q��k<KTSNx�M���`����`�K×��X��W��c�p����>o�t�k>��	����.��elT W�:~�i^�N�8����C<��LJSL[w�7��Ӈ�M��-���!�ң��dv����A�nA���"�R;�h����R`�Y8!7"����l7��R�v�eJ��Kg��5�4�'�d�B"0�ֲ۰�a{:y���Ka�Q�3>��s�!����r� ?���ed{U�A-Bk�N �h�����˴�1=|{@#�p��B��L���tbv<��cU��'vs�L�s��������$�>�$����Tf/5�"}�Θj�Q�Uɒ�q��`M^��HK��O���,Bi�
��|� 'ד�Z&y���/�$OzE#$�������AN����c�~�ʻ� 0��������`
�$l'M���K�%��,dt;��KH���!,Q�*�p������SŔU��cm���ٹe���	{�	Z. ��gM*Xݦ���)\�	f7"8'~E�H|f@
���@��1��ҳ$���'��FE��}��X�qY��)�!g]�N糕����\�'SC�o_W$#Y�=�y3n��&�b�S���r��;��=	.V}h�=�|t�~�l�
��q5!�m�=�lH���8YId��K7��>�T�&���D�����m�l�|�9:�=њ�m 1L�w��ȥ�Ѹ�B䯐V�P�(l Z��NL�w���{Z�Y���%�^!��A&�Ɇ��8��Z����Fv�d���A���͢�ۙ9y��
�G�i��)��e��=�H��Kwc���~��A������>F��#��nBz�:Ɏ����D�V|(z�<^%k�/F�|1NU�<dNf:67��t ��N��"�~�;��ـ�AjC�T�U�Lݙ�=���/Ih���9�i���,Ku���c0�#,._��f�߸4����#zMÈ%b����������=�`��r~����H=˱&,R!�w�6��k+̈́��_�D���mF�+)�\�jԥoJ�y྄E�R��UW�'��L�'�j�%J�w��Z?)��u�#џP���ނ�|�a���!O8&ml�kAo��Ao	��JuY�U�������!�~i�{c���,�hF�̆vح]��b���D� ���3:���6#�!*�)J�h	c�-������c?�]K�X�x�g���e��� �]�m�T� �T�݁V'�#�:v?tE����9kwz_Ff��kz�9X��qDӲ@z�>]�����L�����_+���s/�×�Ηk�_3ꩺ���ƫ�*�W&c�8Q���m�����ů��j��қL4R�'CLq�h���+hP�_$Zj��j����x����H��&N\�9/��<[��@�G%֥-�ę�L.B�xL�x�K�P�[<�T�q�У�Z��4~mVH�6�;�L���h�������6?)������p��r{��;����!(�^�?+�U��Lm�( #�MuQ����g,�]�:]��a��0I��i�^��������/p�:��Z��e0o���8е���U�fD����X�=�g/n�^y]�{���m�Դ�4ɧ�$r��^�(���^��x�}�	@E�4s�UO|ֳHԀSuC�ľ"�>�a
�AiQN���N��$KY@���5�겲���GuS����%��v���(	��X��v�m���.�0���<+�_pOȮB�����'�&%`���z�����z�F�(�i�U����n�_�G]�N���3T_du�o>�H�~;l�A�����!�";�8V!�%D�e����]�|?@��E����{<;)K����F�>i�Ht����9�U�4���U��py=V�h ���Ω'#�!S)����[u1�YF��d[F�4�{� >�t�	Uܮs1��8��k8�]ϋ��d��@ަ����I5����Tv����w���"]8��w�.��;YY2ٙB	'Q��^vu�4��ʲ?u"3]��z0�~2X:u �:Q�Nvt�|���'>�𫳴��n�'�����P��g�y�%K$��$��gQ̨vk��.u��o���_�����D4�:�C����D)�k�f�76~�y(u�n��o? �Ͼb���l��s�[��N)���S��<KcR6J<�э�^8�9)�$�[�!��&�W�wҞ�?��P��j����C�.i=��^�i
��p�1R���*\���ln�%���@�D���P�G2X����T��4���5I'�G�������XP&:!'BI��4Fd����w�6�q;2�7H�5�Sa��ͦ4C�QUK�����I�����t�S�]Q�|��հ���J����������2����I`"eظ��/47�g���Ae$��i:N��zI���՗Akҋn�;�R��/f\/��j�M�0�G%�(�qU:!-�Q��?�P��/3�a�B:IT(����RiF�콑./����|�w�ʵ�GD�^f�њgI�͟��AE��{�=4�M�dt����!���Gd�Y�F-)",���}��j։��9�
)��a��ꠥ.Js
7*<�k]�P�Z�x��6JІ��	G��S٫��'v�-��O�X�ν��'��A-ī��	�S��,=�XiAꪀ�bx�i�"&�Ή���H0��ʬ��ۣ7�|��M��-ҿƔ�Z����\"'�a�Հ`b�KyG$l9q��.�)φV��ą�}�����KXxA�{'��w�F���`xpഷ9b�WjlC.E�� ȑeE������Q+�<�\R���b��5��'nSA�}�y���k&sSV�~]JF���'�`.�-Q�[����W���M�<>PC���������'Hw�;�``��x�{�(h�1���� B�!DZ�pc�RR����h�>��S){T�$� ̿R��JT��W��.��?{#�D_|) ���u{d���j2�&t�~n�� N�L�����\j�M�k�r����o��RF�6=u�3�_�X����l0�>N��(��+�$*
"`?��t�� �,h�y���M�"�-�7ҥj{Y��f��O]���@�u>�����S�[��v#�հwm���
�(���uvT{�)8��Ī��������KI�B_��F�זּl�`q5��b��-�+���9�*�bg%Y��%�m0-���d�s��j:'$W^DmY���G=�|X1�~���s�~�D�>FwHlR�~���>��	:�qpF	���*�T�"��3�b���##�cB�^Y@j;�s��m�ov�]��͑�B�xQ��ۨ�Bn�?��!������z�E��o%
��1b�b�-z�P��>Ç�5enwG5nv"�T}őW%�-��H�cL-㧁�Mק&����d�W"!����=�%{��l��s�N}���W�K��Sk�ՓMQ����Ž�zӿ:r���9z+�Q�������u��fv�x[}�ˌ����ܿ�#�+qS�ǩE�$AuO͸O��m:�'���<�Ɏ����6+����J�4d�-���_󣔚�� �_:����G-58B	�b3s��cG��<�0���/{;R��W���L�ԣ� �2S�*AdZ�iB�4��G#�t�\��V��j�Z������z�]ϐ�.���Kcsi�!���at^�QI��6K�� �*�}���0���X`�J��}x�?7_B�?��lv]���n�0�~���i8"TUl��I��;˜ݫ�����v�v9f>cc�u�5$�=�L*?(�<5m�/Bk%iw�/�o�7�w��P'/�-ssja޶���?���6��&�;bru#�Z�g ��vv�j�����,�ʖ��
��A��E�:}~u1����[;LN_fȩ�$���{�FN�x4 �dM�]����d�>��fST����(�p���0�V��a>=ar��ysmBz��
ɫ���_nM���c-�5���|^���7!-��o��[0��^�C�|#GH��|�xa,��NOw%$�9�W`$�lS�"�X���|`X�J̌s�e�j��m��+��_]��4��]c.b/( 1&�U�O�<]����z�Ǐc5����zC/[_`��/ڦ1$kOW�Z`�;�W�Ty����SF��\�ި����A����X|`���h�7��T�8��,��el�MF��k��9E�<��:�qD�b���.*t��-���̰>��M�*ó�����6�C����#��������h�7�+E���}-1�7��}�4��\ �c/�P`���fA�����$A�R��F���dm��R��pD�! n5��5힨q��dɝ�I"05�O�Q�59���g�6D|_��y��)y�l輣s�E�~�kMhq��ߍ�Z���V7��lfݐ@ʂt��|�ZЎ�HT��S7�a�ϩX�]z�����CD�� FR�4xC�x%쾯��J��S}��D]x�����\GŌ�c\6���߼R�Zi����f�"|wAi"G���Rs��zxJ�j ���_Ҝ�4����a���]@{ԉ	�g�V*8=�+���>	�=��d�g��a�y�j#�},�y3�؊v�&�`>�'^*�W��[���a-�g����GA^&Ϝ2��,��Za���t�B�'���j
?_�9�7>�rqgֹ.�(�$���>o6ֺ�!����?��/VV��,�yY��U�0t�/�j�#�3i�����Sp�Ĺz�O�����o��po:��kD��`:F%M�&/@��E���9kӋT�:��	�N�V���n��L!����G���L���v=�_���
x���(Zѧ�������P��3s��3ʌ�Q�e��V�'� !�w� ��}&SO�)Z����k�����Å���_v%;:ּjt8��|d�Ko�}��S��o�v�
 NC60��j�2|u���,9�d�$�VA���=|�R���H\ۆ���n�q*����r՚(��$f i���}U�9�,�I<�?�~�'�B�)��-���@�!y�/�Q]���N�p�+�	�-?3ϫ#��塩���#����B�\C����7�#?��kZ��Һ/
�����iiM�#�iw%��罼:cR������^�:8y~${oS��#o��6�O��4�m�V�*���^\�����ᫌ��J��2S��9l	����n�n/f݈氓gR�o����q�"��@H�'}0X���BV��29�C�Aebd��'��ɬ�US'��a�z	�b�+m�,�}��HƐ�xI/8
��M]��D�0��(h�5�n���T��}|H��W����N�F����	7��&O������d�Z%���Q�V���?�JH���F���;/Ĉ�"3г:Y��y���c�d���4!r���IFQîu$v��}n
�b�\d-��by1�� �H+MK����0 ��1h��X��gG3�"��M�D6�9`��(���/�I��2W�)�LkN����N3P��T����` PJ��,��}�轢����Z}��
��� ��Hx�ޗK8ԒӸp����2��\�O��u,W�����<zWAg�0���'���:dޤ:l�g1���R�c	Z\)h�OW K�Y�x�cfˢ�,rQ�Ze4�I��"��6����x���@S�i�3Qo�|�>_�vYfw�� �
��p,�Ler���Θ���p��d��&��6���4L��_Z'��Is�U��/,�a�Eݓ��r����r��2їq��+n��/K���}�#�e�j讜�Y�e�g�\p7�]&��潅�����g^*�"z�!:�Dd_�y�M�Ԕ-	�vǚb�����D�=S�IO���^�����EvQI�7��ta����$���u�~�+��/5ɼ�u��A��P��dU�7ѻ

r�<�/�������n��m?sOd1�q;�Ԏ����ّ��O�.6�HK�G����a�T"X���*Eǯ��x\⬜4�a���41LZ#���*��
R��Wcd9�jD8Վ5eb ��V���uS	{pT�|t9�-��'�8x~鮏7e����Ґ�k�J���kE0T}8_ G�����C|u��d��n��1��������k��1�Dh�
�{��X`į�o(�Їl)o�|��}X�U �o�.����gF-0!�]��lH#�_^~��^��<�֧ld;���������lQ �i�v����Th�H���#ߦh�읧���>�]hJ�<�H�j�F"�L���[���f�4.������#���ʶ�}��38&�p29Cw��	/!���R"��͙�g���X�9��-m~���1?���0*qLb�;)�#zV�fƥ����y��;���M���Ԏ�*	`����|���d����:���>���o���-��Q�y�������#��ǈ����vv��u6�����.���O�3�@�X��k�n��3dt���~�P{̻�5�ܫ�
VΔ~�p�(ẃ��G�	���~�*Zk1R&�v�@H�.o��&���v����'?�ŧZ<��iJ�%·J#�*'@a�;`<�5�ǔ�%��=�9֖W�G�o!���f�l۰4�*�UCo�{�x?w�����(�L`���4��ݷ,����F]C�Mq��&MW���޲I�7�K:�Rx#
id���������Oơ�S9#��%Cb#�hs�����t����� Ͱ�N�����`�emKf����@]5�?�5q�՜��ߙ��l��u��BP���"�='R
��O�Y�1��1��҇�u[�C�"���~�x"E��?*QɌ�X�a�v��,��(���ċ�d?���E7o�Q|���_�[�ʰ3�1��5��U��}9m!Ahs���\�$`�����/��@G���N���#`	��ÄB��V%�yq⇄���ʖ��S�Q��2�vS��%�)Wַ�1��O���[i.�mr;�"�d[��t��Ի���� xj��nX�4Kn�լ���NP�%_�5�d=#O�VP�N1��s��;��\�YK���^?��E�`���d�Y:��>�|�j�U CP{>j���p���BZ�6�F�ޅ=U�;���6� ���D��@uB���޿���E���v�I��{v�t��vJ�~�H쬐~[��,d_'0���1[��zX�i�03�������҈J�(��QB$���Pp�.��bp|����§�^�y�W[�-!�!�Ӽ��NF�"�G5-�#��G���`�1U-�����j:��"���y��V�rQ�i���z��+�L�����FA� �2�ϦIŃDWm� ؍sL�g[d#vNն�����WӔ�|C�o8˯���/�g ��pf�8�k˧�į�-C�i�2� ��ͮ^���lA v�#a$�(�&�3�sZ4�5r�O'���6ȸ�׹3��#gpЩ��4���A2X����%9v�!�?Z��I�\j�US'Q��Z�/Pzܛ#����"�T����_�f�F�9�*f��'ZC��\�Zڋ�n���f)� a��� �Hd�C0}#�9Ф[�1	U�9��L{`��W�,��[�/x�v�2;d(���j#�A� �_���rK�E�{�Y��CG�n�"ʁ���k�ܛG����]��s��l	Y�ʨZt�b�������&FP+��3����z$|�ߙ�d?�8 �>$;�󌡾6w�:-sW�k폯v�Mx����m�o��ü��gI�i#X���"`����N�*T2�E���{�<�<s�:c�@���̄�y|m��X���I�ڄ%[�q�AfN��s���B	��Z�6>Q�`�9��MuHp߄���O�'����S�`P��f�3��܃�d0�0��~���R��DHC��S8�HJP��px�����C�7L۠1�ז��\N�%�u	xf� 6�'�D�Ǯ��D�2�[)�4|ү���O�w�K�yE�%��[���p:�HY�ݩ�������G*���5s�sFM /+J�w�(`j(�
u	9��ҫ��d]�m�,h�3�/��J��Wcz8 ��g�b\�ܥ�ŝ!���6��A����������.����q�7R��ti,�w�pn9�+i�Ȣ�]��Nj`�ߨ����`�t] �^hT9O�K�:8:��b*�s{���y�K���@[�<�˔?j�2�?q0���y�	�+{�j-�<�K�DG��08J�"��"�����7�IXS1�
(C���^ ������q��Tl�<�<��\�m~�\�D3'��q�Ro~]�Xɪsx�A,��v��?ɂ���A,Ɩ�s�f�=/�}i���7=yM����Qu*՚.e`z�Q�хG^ܪ��I�#���}^�"���7�k�L�E%�!��y�W���pst���e�`p/ǜ���@��A;�oqˊ:�� ڌ�J��ٙ�75`?B��[\C�y��9�-p_�^~4�w�uR��0f��>�4WZ�sz�q�X��)y��5,�~����y�X�w���zԬL��>��������S|��ՀY	[=���)��aTm �%j����;�vEf�h:�+=Bk�J����X)����F ��O�½��.�}��B����A�G��)+x�T�	��+c��_Z��*O�!ȫ���<��hl�KK}xY6� �V�"`��Rx�x(x�<��L��Ȣ^?��6�1���E�_Α��+����<�U�q�\o쵢E
�K�YvM♴<�O=e��<G�w��E�ym�� s�B�B]\R�2�'��}Z�^_���Q�ݖ}��RP�c���P+?�^��5t�p-AP�pa�L����3{���n�)}[��i��_7�Ίl�I�Yo��}���j@�F�:����ic�/��"'n7�U�ɀ�&��S�9���ƴ�� �	�M.Ʋ���-˙���&/��-�� �6|
�\v&���[���H �?��ځ���I_�o��*ffcݞ,���S�}����Dέٔo&����y#��\g�WB�Φ�A��� R�<�T��y�;ʴۊZT�B��9n��U����;b'�Z�#q`RE$��PM E�f(Z�a���2%�}A'{?ݑ�vz�Mg����6�� Z��'�
6s�;�͢�.���Vyڔ	<J�-B�"0jrO.w(r,c�|]����y^���% +��+UpLg��:�[��e���i�k�)Mx�*<��=Kx���,y����ӷ�1��M��MAJ�>\i��5G]��I�59*��a�x���x#&�%"o1.S�g�?yڼ��%�V[��8�Z���V!�;\�`��;���)�AT�bJvh�>�~���W~_���x�]�#��j����>�꥚	������*��H�y��`.ő�I�'i�-�9�/�����>�L�!n�q<����Fo� \V-9�dk*��_Ȃ� (u3&��7��\fnA�ӵL��pt=R�et�I���8��&��e���̜��C �R`e�|�ʸOʲi4ǽ�p��[_�sָ��?�̾�A�L=�����C%��x&�.v�)��z�O�Fk�[:�8/����ԠbS�<�s���$��E��_�:czO_9��*�V�!Vdӆ7�N�^e�/m�'�Z�nC���+�ۄ��*�a�����deҜ������V�y�"99o� �z{���i�[�ɍ�kO��-��u&ukqL�
b��b�)Tʹ@����:��RX9Z�+g��[]�OXQ�WP���﹮�RѢA�,�~���jn�ٚ��(�x�f��m� �^�I������E�gS��N�/�Xf��������Pʛ|+�yv�SB��Byӫ"�ç̠@������ɉai��f�Z�DD9F�cj����bz�S����6���������z�
��r�w��{ ���4(9���&B-m���6�}H �T���J=aMqB�2��V�0��۽��j�,������K:!y�:���.Jt-j��-. �DZ�����*p8G�\�l�돱�r�����t��N��w	 빕�P+f���WV�V���ݢ����$ߥp��t���t�Ǽ�}}�����~
~p��J��!K&��ro������T����Z�Va�Kz�" ~�sR�(܍���1�	1�!�i�e�R�����dw�J��6El9%`-���e���$R톬���H�r�j9��a���]���h݁N�� �`4�~���Ԁ��*|��$rw3`���ҡ���A �,�����`^�������w�̄A���͝	#��r�R/��;��M��bp��G	ȍ���L�W�g�-(G�&ɟ-�/U��4\��dE�AY��eŽ�q%�6�9��L���� �UF>��%|�v_`�#%!�����w�LXq	�(X-_Q�}�[p\�B�>�@����e�%��z_���)�I����#��L�Z�q�JZ��T7�Գ��eh(r��0��/�NS%�XP�5��̂�{u�{Mի/ }�ee�9�p☨���3�;U��|_ˀ2�{ƶ�ҋ[�qOHY�os;��j�-aĨ��x��e���5VIw8����D��x�\7�:j�\j�`V,������S��(/��4Wq��>u�kM�#kNd`V)�+��1�X�ʶ�,H2���E�/a��_��$^�A�jy׹_���M�cy��֧�TF�7�ഘ+MP��NW�����8Oi���y[���g�@����*���M��hfw�L2�q��p�����cB�Ѯ��\�w VU	RNk�
	N���V�FPO�Wc�����v�jvd���٨MI~���Ɇ��'�'���Ȗ�i��z/x���1��,�'!mH�ZlOUVR��h٣]5WY���X�L��f������o���ˆlT>0E��4W~�.ԉ�W����{��ĩ����
G_�@�sVҤ@�i�+�sG�X�h0���T.m�x2�]�u�O�
�����H��y�����R�2��OFU��3��Ԟ����m�ލ�<"� S�p�U6�s���01�TL���)�O�3pQ2f]�����������v���)��������r�U6��B�*~~��@$'������"2����/p	I<Y��a��Є�L����^�q��)�W�����M�ƪ���0;�MO��SQ��7��9̝�Q�G��Q4�#�0؜*�/�l�I^�YՅ�A~�DTϏ3wϗQ~$"$O�ǭ�d:m�Jm�Źy�����ܢ4�R+�)dN베Jó�rt�v]Q�l���L^%�9�nA��@��\�"��1H%��8�G4�cF�rA��{��e*�j�t֣x�T!�Y�L��F��C�w��1��DMd�~��J��Nal}�źq.�~d1�)+$12����Z�M�Pn�Zxx�1bsOP{��j�?`��Iq!nkL�[�����-j�� &����B����kw�+���Ed���q�81t�������F�@���q�DӒ�Jw����3�$t�H:\ x�Ѧf��� t�z�)�����˃=�e������+s�LH �IO"OOIMi�-�G�^y���g��JҚt�h*���](���'O��9�K^�S�	{n��w�u��í4槣&@����:Sep�ex�`ߺ-��}S_*@)���t�%�T���#���*q#����f=�&�����
m4�y-a��Ǹ�n6��t��+�>s��7�\�V)��(�p�C����*�uaas��d�߶�-��R1���Y�i9��<�6�u�`���d$6L�~����q�n�&��y�$� Wo�rVN�U������w���\n6�yq��w��l6�ϝ�oaD�e�Q��}��j���fZK`����/���iP��"C~�CbLM6BCP+cv8�:=�0ӻ�qGNc��g��N�?��z��Zݢ���|�" �W1����v��z���1d���������/�jE�B��t7��b��l?
8��?߈x'O��<R��.����jS�L眜�{&F�D�!Z��QEG#�=�}�{�w�#������������/7��x� e���Wa�B.�pS��'�{s.�v��ZL�*h̅N��2���5eja[rOe�s8���&W����r~�)�^������̢@mf!Z�{���_#���\ڸj����H6VZ�{���Ͼg��G̵�ۈ�)׫�a��f�:g���OJ0o&+%]:�F
��c�����1-��g���e#�Fo�+��}@o�8[��\���[��/�E�G�s�}g;H7ؽK���Cf��:��X���C|�F��8n���@�#�dj��^�ĕD�.����	�X��h��4�u��1�]zڽ�򈱻�,��"c�և�8<)x�C�S���L-lϲ��o�3�;��pV�*�xdA�?Cɺ�]��q������fQ�ck��͙��͙���#>DZ_����on�Hx�-��Ҁ:r��*��k�e��v�ӈ��:m�-J}����M;}��������H���o���&)G�'��v��S�&�u�4�U�'��4:6���CGh5G�߬�/�BaԞ 	T1f��3A��O�ܣ��o�㽽�$��� e<�vw����?*���t���r#�ag��ׂ�n��e��P�1�!o|SFxH$"�~���;�)��	y>�2����Nd�`T���>��^�J8 O���a	м]���F��f ����=okY������y��58���T���>��Q���h]�
�yM�􋮷�?��M"�L�[ �Z�Qw|�Q��O���ҾT���!6��i/gkz�7)T�Qc��h7i<��1|��%�|So���fk�]�F"�؍��,�C���C(��]�,Ƣ���֑j�3Axl���<r����9���x�,g��4��H�A�t�0WE$�P�7�r-��l��J8 9���k��ɨK�`�
:%Z��������8*�P~t�����cP�!��~��E�������{��;��F�%�H[x%�;;�;�9ZBK�F�����=9����r"v��Z܇�_���ͥ�w
-{Ⱥ9���Bp/)�z��� �W�h��ym�YN��:3��+��K����X��v<w�d���}��K���!(�L����:��D���G�T>��$W�� ��������"�[~v�%�W�h��8n�&�NC�����W����4)/��A��?��XE�&����2�&���8Yf~����m�����/,9lJ���U�H�p-bQ�M�"���g����'����j.�J�)���z�]�@L�4\�����3�$�r�CHEmJQ|���Oe.�4bh����A���Kffˁ��qi�Ժ�۞�֘L�K*��n�J�b��H��x>����g����APl��4o4�f����-���=����9�ۯ��Wg	��5�6��p�+zz驌�����)4��O����6=V�,�4�c��E�6�$K��ψG��jK	\,�.K�-�~?w����b����x��6Kޕ��o���oRC|�K3�>F] �� ��dx���#�;�،Dq�!�ȴ��8�:���V�{g���Lf����Zy��S҇�| �[O�`���t@���Y�_�����PJ�K�И����>f�w,��2�C�Q�j{i��포�5u��X_�Ly�#���P/V;7�y|�B�)n�ޡ�������D�8��_���U8.}R�� ���AϷ��Dű�/��m��+IE�ohT^�l�C��?�js��þ�^	���N���v�&��-��?We�;%�ސ�6�D���u���'�G�@���y~����4�{�" ��/�5�-MX]6��ǟR;	��e��̏n��R�r�埳Gd�e��@'���y��|V�����x��>�NVA,� �U�u������:"hk�8�/�ǁ�=M2�¾��=TZ��,U�Cg��cr���t�9��F�E}��X���~�V8�զ��}S#�G�z�eJ:���cS/���&oL6�F���d��5�Ⱥ<<�t��%@ㅦ����t�5驔��h������Į�%LR�8�Wi[A����-���4TYK��hk*�&E԰\Ċ���˒�RLn�8�`��������%R�H�<wn��b>��P �{4-�A[��^$�Y��h?�#v�Q�n �g���O�����+�}.�K��Tՠ����H.+�{��F�8���N�U~P�{HBV�0�و�P�����.k5�;mSsB�ެ'��P�i�*?$�_y+�
Y'���hz��HQ?�,<(4��1s����\�ƶL?����F�u�1;�b*�gȋy Z�2E�~��@�؜�"��xD�4��H$�>�S|F�PUrg����ܣjp{4n�3��"��t��-|��5�^�fDĆ��?��� ������=+u�4\�~��A�5ڹJ��8��ο`vj^���(}O�垧(On�F!�+��K"����p�>�1�fRġ�B���)X�Y�$�K-��u�ۆ�3��*PLo��>S$J1��;S°an(�y����hE��h�K�e7��̌�@����	1�*���P�o�27�qd�Ӟ��X��g}�}:~���A�r���T�@�\2�������@��y���)U4̂'�O'!԰�C v�L2���|�3�D}W,�[`�5ؒվ�evZ�[+62ld9�ǔ��q��Φ �@���i�ĚiN���M�Z�v{>9z�
��6�ì*�� �hz�e-�L��3�Te��� $��]@�)��T+��u̬*d˄g�]9KA�c<��Zzz���ר1e�זo�9??K�S+�W9��7��:�%N4�L�	"�2�i���G�eZ���DgB'?W]�4*�[�F*��q�ģ�9R;��,���5�Y���qIL��C/}Ejd=�����#�C:��r��1p��8!��T!�c���`�X/�<����$�_���vb�1I�Ddވ�_̀�������O��D|H�ҟnpb����J�Z_����7g��F�e«N9nA\}l#^g�8s^6ґ�W�lm-TX�}f�8y��$�i��R{�����+;��= 2�Z由c�W��f[�s����ڃSn���E��ᷥ��C�r[P��	���b���j��|y��H�P���9��ەT��B1u�5��6��ܡ=��a�g�x�M�CN�D}�~�'��NTԿ��A~&7ӈ��g�Q�G���	��Bf� ����A�'�mw�����*HO�Z���L��t^��g;���A���`(�I,���-3q��a��_��=��l���k�*n��@� ��Vl3Q�"�WD*���k5=�f�U���8�iN���F~�%��Zl�uwZx����
%@߮����,��eP���H4��	2���>�c�n@��8FN?tv=��mS�?�&	���ɨ�@ ����?����-FZK�ܶ���q�K϶3ѻ	�����(,�t���3�����&U�5�wM��l�,�>��6�s�&ۏd��H��	�m����Q����9��������g���m�xqzAg.`��4���qH����"i�:3(��ŗ�E�@�V-���w.�e�vB�<?OJE�@�_��E�9�#EWwV�8��U��Lp��� �u��j��5�Y�/�/�t;]����'Q�
A�VOM�h+f�T2���a��d�8����ef��k�OS@�a�U�ϙ��D*뺼]�IR��>Ţi�}����[�WːF�(Yx:4+^�\�;�Aӆ��A+rJ^�Q�?��	�P�A����B����)PȷL�y�o����������|����	��ӯ��Ɠ���2om��Ѣ��[z��ðn>A���p� ��]���u�:7��r�'_�p,w=S:@���n�3�w%0/9È�� �����͐����&jb�ȱO�%��71�ij�Fm����is������A/��%�cZ�\)�&�hV��T����G��6�֫ڽ�<�f��N���� ?f4�6^uW�����x���P
��c���A�~q�/g��%Ž<���Fq�cG�i9��P�V�L8��v.B���]l��Xܚ$s�B}�q�գ��
B��Q�]oq}�~�;�I[b]�3�w8Ui����s�; ��!T�L(2��q�2�ɿ�|� ��G�0�h���4h�lJ�����='�!"���ӕٲ�vۑ �˝S�毝��d4�L��LU�O��4�PZ		�<�v�\��r�����˸E�m�_�11+�$}�*��=ݫ���71�&��y��_��r0sє��`��v}�A۰˃׭�VeH��ߺ��bR�q����bT 4��e׭���3��8�>�e�`���>Gxz���(��MQ����SFKߩ�V�o���v�w�Y��ɍ�L17$��u\9 �v8�-�{�1�qf�����_t�m0�ٚFVES�p�81٣C%�&!a���=R�OA�����z;_O�-+�I�,�9���+�63F;��8���|M�AY�0���X�/lq�/ju	��{S.��+�OK��m(?l�#�O�ɔȜ9�K�����'zb�ﰈ�E���\)uI�3�r�����2��t��	lՒu�_��3�+�*��(�$���te�g�HZ�����������_!�%�������̜��:s��N|Z��D4�ne&�1��T��w5��[[N����'��Y}��ļZ!Z&V��,����!����'L��@W��B��U(bu�f#�4��堚�G��t����`�_�2V���I�u����iX��@en��������K'�������������R��Gy�e1���2ڪ�*}����ʂ��2�D���>�;M7UV��d��\���*#��D�` e��z�kK,�uU#����~�qF��@K�
8� K�::�>��d��2x	q*�ڇr���B�ά+�)���f/DjK���e�m����@�)�Fj3/�L�R�oJ?�YU�Ԁ���ќq�Έ�ɦ{�p{s�^�LxMwe$_�^�9:g !�AoM��JP����A�j�m�.A!xVц�ky�o���}j���2����c���֏��MS.�{�ߒ	�wJi1�VT��i�ϒ1�9"�y^��8.���mt������X�c���{�-�dj��A%�_�lJVMpgB%(�lи��h�W4�6�����*R9܈a�!�b,Iy�*��uj{�� �A�~�ٸS"�]��$�5v��:�
%�P��?��v��Q��H��Cڔ��2;D@�L	����U���E�ԙ��7�؅RcÆa�y�<^�BI�I�9�����v��v��D�^��ԋ�M-��<������C��+ɱl���{�����ˠg�co��[:%Zj8*e�E��
�������J;�i	_�%Y��H$�h^:ǳ���n��A�¯#f����y;�'�
!	�F�^3��	�\0(�����A}ƌ�)�^|�G�����I�	��w$1�� � +4� �8ʢ���t�3����6�T5����C�$�}��h��Oxӿhu!��a�����4��aCi)ft�T�
��a�_�ze�����!젎�?������j� O������s�H쒷@h�cã?׫����z�d�(E�lp�G �9˛EH}l�0<�K%^�mz��aty�
�s�J��,�uh�Mu�G������2����E͢��Q��'�� �lX���ݔ#�L��%(���<`��d?% ���iы�^�<T�X���V�J1��p�/�p��O'B���|H����V;d�mK��?}Ƭd�S@�=��SkԀ`�w��G��T���=����n���K��zǠ$���8}���(j��0	f=M�(�M�ZY�FA����ί@d`UE��2�Y,��m@��}X��Iٲ�(c(���@�2��	6�;lk57���k���~�/����)X�j$�<�T��^�n{&V���i����w�[r#G���S�/�����o�|cLW>��3]$�7�˧`�˃6�KK�@�xŞ�ļr�$W�ڮ�n�^!�}��9�%J�O��-�(=�t�Ag����9M%�8s�̜�i�d��@)W����`�
���(y���*!���	�
�̼z����j��Jv(�i�Lg�U���H����� F�q!�hu{c��?���,�f�z���d�w��aM|�����-�,!}��~����_?A��ِ�1�$ٗ,��~fi��ޔs���"�@̈́�Z�7&���� �U�S6�Hhg*��5�ڴ���/����Xa�C��9`�(|����CD42Y���?00���\e,Pv�o��� ��@]��(ւ*���W䅄�&����fW	��ef�N�MR$�^�9?p�Ρ���L����[�1+B]�kOŔ�x��E��
p�zA����s>��(�2OH:��~�?�h��t,��G�5�Nu�������xe����}]KnT
VD��PF�TB}����*����_'Q#�R'X�&�7���;�ŴMw�	X�	��B<��R=�.�
tryʷq>hҲK���٣����Jl�*�G��$<۰Od���AɆI�1���)�v�֏�K�����j���YY�+ȋT�U�D��L���P�I-آ~�m���(N	��h�?�2���jAQ�g�F��҃.X&�<`�t׶@ ��d���i�.n����ڻ�R��Y����D۫ա��z|'A.����]񠔂�b��	t3A���L�i�N/DB.�%S�� �j�v����,��`�>�s�4}q�����=�̌�[��"��ޜ�͒E1�Z�+>�%��!�E.�����������-+|��ݮ�u�7�gͻR�}�=K��<^t�LC�}��{7uMzmݗ�*qm����$��W�K;-}���#�pjk�DA��s�

'!əth\��*��zEUy��t�U���ƣ�M(8�D8,) ��,��x�Q�1b�[�
�v'3?P~P�
&f)D���4"��h��P���8�Ъ�F�v�ca��Y6fx�}E�� ����ק�����"Pob����,f�UUJ���ݡ��Vb:��>_�nEX��6��+k�*=���6���6D*�BJܥ}��mN,ዜhS�9��+�EX;���n��F�����3�!���˩f/�>fw�Gx0I��O���R�Y%�kѢԖ���ۘp8��Ը�Q��7�����KHa1�ed`��CZЗ��5�:�ǘ�����>6N��?3l�Z5����|�OuR�>��ET�n�W����^{�ls������ָ�S-���sm�s�z�5�2?�S� �	�͚�	�[�zI4m�>PI�����:������,Ɋ=e>Я<eQ3_��dp�he���E��c`㔛�u�ʓ�pDeyT��>q���iB�s���P��2��λ`�{�A���׾>��(�|$J�ݙIlZ��&�)��P��x�^���"F�� �	�S΢��ShW1���@����<}��A��v�z�������
�Hg��/���3}���,����;6yЬ�����°��p���������2�"5�g�4�*�� �?x$-��/�b&=�ۦA����;�W���ZXǌ��2�D�%�q%�M`�&�j �:��f�,6��ߒ$��2���o��פR4�2xߴ���2�� :4��eGd�d�@W�'4fdv2��( GF9����ּ88��6'ɀ��|�\"�;͹�tr=Y�X�I;1pi�.�z��׈�Y��fU,RA�z��]��y.�%N�o��̟ô��u�ڻ�X��Q����F��˅q��Pb&�ˍ
��MS����Z�,�a��-��n�X!�8G^ܡ��hz���z�4L)���tl��Aِ���5�s#�d�c�ʹ��y�VvX���f�V��%����n�s�޳�e����rs���u�4������G�ۻ�|7)V�-N�6��B�(�%9�������7K們Z�MP��h%�+���Û��
|���Y�N[Af�te�����q� 
��s��%��$Ǆ�Zo�~0�x#_E��c���6��I��BS��*�=}*E�[Y#�N/��M/�;��N�z�Á��O���V�%��8�d1�ԙ�Jv��d!��6�����n�'J������/�!��!ۼER��Z@�`�/���w�	4׎k��� (�����7Yq��{a�+���4�LJ_���`�f%���j8�����P�Xt�"�k�:!y�4|����C	f&����%+|�m�g?�6=�&Y����~u�tG�e��9�ZU�S��gˢ�cP[+sg>m�{M1/����(?��ػ���$��E�b4��XR�^�?�����������6���:c�T����QH#�J(��d?Nj$�����~��O��N�+�g5:��^�9�'��l`^���[C��z�yE�,�#8��P�4��Y�]�N� E �o������xn�l������ZAv}��2¡~�=��j�`��^=׊�t:�JF���yhg,Y��QQ_f�)���R�d�r|v��yUԪC�H�p���=��woa�ˆ�0�4p��x�tݫς�[��b��:n]�Y���;*��:��h�H�g�R<�k���\���>��1��R�̲K5�@�+�*�&��gP�|��#�Aq-�k��e[�ݿ��8;6,l��E�,����>Ujauz0����ʶ��H�ⶄ�*!8>�Gԓ$��g��Udcݑ��dHj���%@��W�ĆT�R�&/�t�a�7��y,���8� �y�+� p�'�tT�D{w���_횈V�qQÌ�$�D1%*�e�7#9{����]S�l���n��	b�f6��z��G�< �@0j!�4_���������,�&��(A�	�̠�i�:�u��)$�gv�\�lHSf4�d��)�?�s�aB���Sj	g�2����}�T�v3:��\�:�B�ao���a��=t��Cx�^�W�F��au.h�eQ�j�v%�4;�%��8� p(� %�o86/7�&=d��V#2|2�8����A��A�A�t��V�ea�폭���Yc}���t�������-5렆�\��UG6j�Y��jyZ;}6e)�%޹�����S�/�w�̔�HF)w�Bс2[�g���)^����H�BGD��P�sD1	�k�K|a�r�w���^'���@5�ۏ�|���	8�W�m��Y��!cɠ�_/J�NPp�M6��x*�D���T��>�ur��'*
5DP�[�K�%�,��7�+�B{F���Ƶ��ū)o�6y9���?ɴMG�~�2���[E_wNC���.���Ӛ��D�J��3[���?�2�l�#��;���
 ��TY~�aL w����8�>0���G=� �N��:���}W \-�M;�	a��#�>�s�Q���r^|�R����E�"U��br��U$�����D�g�f�_lGG�83���}�.�
"Y�V�ZWP��_�q#'T��B�W���&��E­:���\���ķ�����K�F6�������Z�.��bX�����џ	23u��6�@��c�0�RcibT�\.Dx�+B=���*zl�&^,��������Ѭ�[�ß��#=\�m�Nx��xn���sc�y��~�[�!ُ�?B��dy�}5�|�A�/-��4N�M�|��̋�a�	��Hl��VK�����>����{�g����Ĳ\?�ڇo���vZ"�b�"���4���2'C%�5*|���,=����8���v�ֹN�z Ao4��v15�|u��~��n6�P�SP��]�m���u#�|�X�@�P��\���F����2��&d� �� �}H�������ra�y��KC;�a�C���ab��V?J֩��l��~�!wDh>���\p����G-N#e})�y@|W�Y'��rYk���Z�y��9�յ8fxD�/tIΆ��B�e�^IA�]�52���/Kd�� �� ^G@�x�����a?���Jj�M[^툒��<I�پ���gZ=3J+k�kGS5oy*�${��v�#�<CR�����n�nc�P�DZ�������rq��B<I��,Q&{�
>r��䷦-J� "����=�Mso��A�=+z޶A�~,ց��`z>(�O�f2��)�������<��[�%[K��j�MD�ݦ���{}��;j��vJ@�Ͽ�j��(	8�?R�{�'=ǌ *Hb
�R�"���|ux$�;�*: �#��F̏�6�1�I��o������|�6�P�x�Ѥ8�ΐ!N^���;yn@�)B����GT�����c0����~�lQ� ��ѥ�y�H	,����Ή� ���!�$ۼ^�[���B��L7�����O1���ae^Ujӓ�M���=�*�,;���YIS���Z�Ҽ�-��j��7�c�M�޿�l����a�D��I8��3T9h݁��%Eq�DQ���j��n3i`T�O�Ƽ�����D���@��|�mi�N����g�!B����R�9��_O�a�O/�1�#�#�@|M��z�;�杁�����#H��4oo��bz�f��,���@�3���E�Uj�M�)HiX�ɻl�L�s��.1�޳I�����J5-ٔ"ԭ"�(
U`ʦ"U0ݨ�ߝ-�_�bn0f��~�cV�.��>���1(���2?iM�7 �я� �͖�Z�`��'�L���3ʝX�G��{T�Z����(�-����uA�/N�p��)�)�w%8�H�h]H�)��)��bA���g; �1��� ��R2���B�1�1����8E�G�y�al�sbfO�1�L-z���mڢ����H�}F\k�~Z���y�N�۽�|����8��P|?��>]�1������Wƍ���24 ��fW�!�S	|*�F�y�
d*�����R�O���H��E��O�R�Ѿ�ߑU�H��z�.݂�m�T{�2����A(7 7?���z�nx��m�{h��ؠ���p�!��EY��Zk�5b,B�ج� d�%{{�"��<M�|�D$N���1��q����P�~	��]���=FNሑ<�R�i*�wk�Eg����[�˔0��t��{�Z,N�E3	�0�ݾڍ��],$����i� �Òb�W�WqY`X�`]~��&�C�j�A��f����M���,�G aI��A���V�<�_�"O���䔁\�)h8��[g��}Di��T��0�M�E@�zp�"�؞l����ઃ���J��&��{4b�ի:D*�2P���z��)�H�����w��R6h���}5�_�7L	*ɝ���K�}+���?A�Á�~�<V�e�e�h��xe[E�-;$6w�"�����Ek�]\9����#e��}����4�EfO�c�ϭIz��)�U3��i)�i��U�$��~�'Qq������}ٶC�5����]�ղ�7��8�y/J8���떱g�vN�dp�Mp&��q���\0�~��"�T�S7�x�P��v���b�L�������c꫄��Ry�g�|�3�[3!��˚*�s�6�&�}#���W�Q����&�i?��L���g�>�O"�	d+��M��%�4"S�ƣ�5�.ƫ+Ǘ��U��0���{���"{�}���i�_%�t��׀�1}�F݆��1��I�>uk�� ������h���V��`kO��
��\����.����-��&1�iv�HL7O'�qwZ$	��GGy���x���^���p� �y+W�99�����P��L��[^_J/ׁ�43qZ@Ăg͙���$1�c��ҭ܁���(ː��fc��f�q�;H�;�����O�aL��Ϸ�ѳ����Ps�-%�2ƛ�>�����Hʕ�Dj�=,���m��5тXȕ�#�.��Co�M6�L�#7��ce��k�t�t����z�y�u,`���h�F?6��\a3ɘس��(�@HK�y���`PYX�� �\w��.�̇��sg2�Ec�}��D�I~��p�`�K�(�>��"��v��3HabXIڭ<A%��TT02e��Xm۷y�yb9۪evV���S����ncq^?�,�H�Hq<���3q��Z+�������j�(
��;X�y[E��cMF�'0&�������pΎ��DG�M'?�δ�L(�6q̸����xOjB��<̋Z��5$���G�BS�����h'�X�v'��E���,�L�Ct����J�~��;�r��0��5��3ԯ��J�y^��Fg��z�����22��V�ڍy��D������=Ⱥ9h}G���t�H��U~���
������F]E�{���Pa�R%rx�[�jK�
Wh�h���5���u��+�z'2�[�`�EA�|j$%���]�Jf�7�(��p�%}t��\�{�G�9g��,�"Ϣ#�/��C����:�ϒ���7�"ʒ3Q��*�>�8��+ (e|�AZ[�=ͳ��6*'E�w/��u������&�o#_�Lm���f�2�!Wg�~�Np�fC��!��@f�SI ��T�&�?�&a[-^8�}w�?�I�J��/p�rN�N_5\�5�ƿU��..ӝ��#jKs