// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
qwLKFtXWqhwkictl07CihSjWaNCcVPLHQJ2s7bc++kfUzZOhlIqa9iz/49X2bi0VTc/k/FwbNJm7
iY9hGJupHSZpqLF8BIqVP0yHOjVmru3CAgzalyRwbx8JXJHtBTbbW/yF43nx0F6eM9jxwO/zqcL9
2yfHvMD0z3LyWxiV92sgX7JRcCblHkW+m7m41t8WA1YBzIfKJJ4YN58X70GqxYgueJb6g34wgdm4
751Zdx/mnIh8wAXRDRfujc2ySJQkHWeZuPuZDUWN9GvwgmC2Vx1MFuLNqyf1biGPNUlnSGG7wnuQ
Xwl4HwnNgRESdYsL5Mvo4ard8pZ1wbKkt3WGxg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
nqg/tI9sap4nFHDwOYxpT22fOWZ9xQgfiICEBfeeWNA1xjFkotheg7VootOmEKmCTh8hMAok1pJt
I+n8zWV3XXGuPTiFcGIkmAXoab2OLwX+TU0hpGEAxobcsp9aZ/NymeCn31ctDtRwP2sSfUcVZM5j
d61VyMhUJCkyogJxCzhYdFN6JD7hdHl8hEQlCKJvU85DuJsyOTnWWF01LzAiol3oocRKM5NPrWrd
pnr38KRjJpJVkTAr0IGwPbZwnS58eKPYfE7UBy2IWqazX1d58Hoh+EIqS5GD6isq3JxRU3DFo09b
gQZWGSgUYwB6sAZZSQQreRMwvig9zhbVQ1z7Vna26ZIHWA0hMGoUMyMqLNFv5x5wgQIMkjPu5AWy
w+ZdPCoFlxeFLoAsU0ixlFq4RzlAb/WOdXbLVEEBSuqXmADMk14q+q/u59f33WYvgX8dqYfoy2oF
n5Y8c3Q5pUj5UluStWUQZO74zdm9NZ0thKUkxsgPGfz0Iq9lQyWxMcCR/pT3bfl3NvkfL/3mofbr
ts5NCMECm93hxNaOBqGcZHrLAvlGdeq+R8gxMuNn6BaMVDDaL+IX82+2sMuTkcWJ1i/afkT6dBBb
twAohuaoeNy8/lNPqlKasZ8Shtl8R3Pf7eYI5OtdXlA6tDTPvAI2q7cENael22gN9+QM/hheiTK1
uK9h6fYxPvPPqHL2Vk/jBMTUGus4c1Ym8OQOGi1XpUe9aGb0n+aKp/Cy+mHXMH5BqxFQch5P37eJ
dJ01Z1OtXEiTV+w1vOGyUunbufy2053IMehxEIlqJmEGWvn47xL4BKV4YWCu/4nehT+M14qtaRLP
waD91fx3grJnMbksXzf+tja0QxVyVatvvHpghBSWoEHsDLTapNyGzK9N+Cb2v2YY5iVJkfWB/Aa9
h6b0RPAoDIiKAyj10Lj/GnveqG8YzbomRnmfyLGoNDgnIo4dS9hXGKkJyeZR5sJbJxm0lroD93LN
DgDlmsW7DaX0BgOI5Xss4tSb6nFMprF8Rd9HKq9ZAEgoYtrPzrSKaTVtCt3VQmpnPKMTGYNU64+2
5w1CwcOVHpwE+UAHxehQXc1OHeYHtX7aQQtdBVAi7tZh+M1AeZH2W2H4c9n9I2Ost3Jx1cTXK57U
qbGz6AwRUdiNTmYPUQqVwzrSRaBK2uuUJXShd29E3BU9HN20zzImrpxLZzvgcOH2UbFJ81lW6KRM
Lg8DlhomvHpJItGIssMH+VAC7gFYMbmyr3zRLplqBgUSi2iSyNm+qbqWaRF/HZRGYfEFVpdpEG2j
JvW23j5HWu4gDyd67WQ98g33CP/foXdQiw3zk3fE64ctG9I/riG217cGLPgJR/ysCSWASGvM+UFm
cEibszO+Nfd8vsYYULXKwXx/pDHQ3lsuxpEqixhwlaqFQZ2XdHfduKFXASrY37AUwi1Mow7wohwv
+/xqYtKF1HQPDdYKnR8uJII5vvNUlcec8luyT77/96zdDE8yJdFGEJ5WeW/zETFJLyK8VKNa/y7c
yCz6y6nimenbWXrpPCM5oaSZA/isdjSU3ZetcmipX4xk+nn+sFIo3ToOuXFP/caoVEMOUp2LBRtn
65o0jHXqbF75cp9UoS2Cr7eY7/0a7eWUCTo2P+CYDCkHKfzZGxJW7ZMI2siUP9JQELJUUYnDtYXI
PK8YqODOn+L7v3Yg8cnNmhCJOXmCeNh89Pe2a3erUIcS1WL3mMfz/34s2QyA9Xf0jVDulYLP+mPH
6DUdCsWgkx3mmPht1lj0kMm6UWLH6oNLH2YDgml5u8GOfEB0RyGhROHDMG+3Ve7g9i0G2Ya7YD/N
EMiFryBJo9phobllTQB7L60nG7Tl/LPRQXBJor7HmrCdBOJgYrwgXCi4+JGuzJNFsoGaMTMCacgm
CJeO1y9YzuMTzcaFFJiUrYodmMkmSDdhQXOr+dROTMEbp/OqKQoqdrhQ9fI2vpL1XtycnMI9UQer
LAzZTE+B+dDdZz/9v6P8iUTz5gddBn+irdcNY9RyN8IXR639vodA8SEl0+ZGIm4exYjplhP517HP
3UlXw1CkvA9VYBjaPLUzXFT1F6ws3iuIFVLZUOWVfYJP4J3+awOxGM7geO03TVDPnNvDN7lRt4Fj
lTCiF6czxvNTAlSf3RIxZn+bDmtpmGqRWyVYLV3OvJIf4c9qbYaPQW/mqfOhnW1Eo5Vcyr9MGACI
tx4/XI7hZpBCgpLUBfjvn+ZFfLXxVez2e/nBjo5pUfahpVVdte3OcxJuNmZ5DQD+a3Ypig9JxdNn
gxKkRcYszY3x1SYFB3Ho24hKEjQnImU6jSwJ9dw0KUXlC6KtJoz2kvnx0AXkr7R40AGi7fMhb8yS
eKunn4igbhrCdJ2YBgdQugaSWdcLOWt1dzg6JJmU5r5ers4BjvL53ehIFtfrzbugXc1OvSoq/4Jg
+2DuG2rKUUXXPcRgl87RAhvXt+lubLQMngLqejaKLWYsOhaVAyaEtjw0IT9xfjPOet+la5RiZQXo
dzK/0cv/n4kqq1VofTg/VU9pe0Z+PuOEwdGFNEIxlqFNyvXDzQGJqayY1fxhGqSoavdaUC2Z6Fd6
Wd7iva5g2tv4Guv/3FU+/SJV3QSaW2kyiMWHANneXaIMjE6VNuaApSw45xn2aI8WTZFBtoHJM04D
Om9PFu//pE7bMZldEZcKHN9DhfFDUZodBvE1doRBhMgKOyif8JFkbzKoO8e+EvoBlYRpW8W6eDrl
Y7PmTiHifMLEKlNpe0HUOChjseQNfpu7ATgF26/9ZubELEok7XFaBtzf6Id0Co55knW46ibtwdPR
ezBH1vDikFRiZEkXf9HRoJWE0Pgh7Yy7IihDzMde/AGBDjjb/KSh/Reuv8jafMB/e+DT3wyp7Z2O
d+tE2DUKdJOpLEpLEGLCc4m1QaF0Dyxu7PglCjmGEgHyDs8dqgPWwOu1h+Nl6Q37uFPe8NiCVubw
dp5VMqNxGwEbjHdhUs1tvlpNvKjps8hhA9pZ+Ozx3pj8ZZawe2Wr3H7hC/o8+xaiBTRpSpu7TALK
Bl48vucCQiCCKvMVdFU3Ykh4V/zyOYGaVeKwxJCFgle47h7R/1nbiSY82a6WB8vHLm7AsNWPj11Y
o5o4SyrMEmyJxLQw8q8cLtlbfDvNHHAolXOIKD/25TVcKJ8HaXB/rTQvI9U+6S8pfb2x/HfEtwAI
mio3apoJp7wzw56i7miQS0fC9Sdx6UKEvKDzGJLXF3BiYoiKpf8sKQuEBzBzgpkiIlujbKgw1dfU
C4U04S1UTr5e2xuw7TC7bjlCcDabP1hI6jBncx6Oo0ikxhwhmpscqMCeS6r6lw2fpH6DjepkPTZs
twx+OohLCq4NQ8qt52uirV+kGMpnxkvJpWaH5Z/RJCLOA7/POui1jlVpPpMhfn5Cy0+IXpl2n+Fw
1MbJtDEyxbHAgtERsKV/4U4HwGuSHD22fKYqdgz80v/HU4BoU+6XORbhO+iPHC/WPw+Jf4Ag3+pp
MCvYqGrlv0x+cAT22YEBgg3K3Z8nqqsyBzblee8HY7wf/AKg6Tw3i35jFvsjbbU/+oroscIVrkCN
oEfpfPFVa0He6szdjLbUq7XZ8cGrYOC+q0fX1d+xzXUqqnYjUQScwQknyTeowKK7flFfgKJSwAdr
FtSMG34FKeMI2nWj6M2DJMJGDdaNFAevrM14pX3MuFiLj33vZ6q9AhK11KBYTo+eTgtJ+I3yS3S4
uivLN0Y7qn70FtNA7TgpAwsCffV4I68nK5fiwWm8aD0iD3UQP6O2R71DGo7aBTuYSHb+CgGqAsxp
v6hCIrzG09RdjmfI+C7Rkb91UJqaOnlmfEgWeuPJLcO8J7NKYn+DkRHbm76AYzmkfN8fSyUqkhSQ
0vA2ZNHRHjS+xIRPjltKhJaKF8eGVf49M0a1qeRePatdAm1wLjznfZXzPYL0c+LE7BS3xga1ynIN
enz3rGo93JlH1ccKOvhZpoxwoqOsNqllZMeszrI+XR1UqcgwAgYGoX7nmFKe6Yi5mP7sU9iFY1KZ
ucipeJ6E8K1rli8AZyA74tg+v35uw121BvFCmdGfYXUFgzm+pOxAbGRxfwMGMnzUmpGFneB+2kLC
oz/DcABCf+x0ZCWjtwee2ghCjZvllTCYPzHuHj1i3SvRum8Unfhot5cX2QD32hVnxho4BOwXjksY
hw0eQn/uGJhoGEHPOt+YTld8x/yBQP0ZlIKx/5gQpQ0XFoLMMIsUC7RdPuMxQxkBqeofZWkzAJf8
kCR+T9kk+rGzjKnnlo74jaz9d3mqZ2ujHfzDmY1ujtyt13an5/hFXQF1D8W5hBAxKYGRn1VWj4sK
Z92ITGgoNFM+fkCxTOm6qexaFqyIqygz//Zk8rZyFSxrrZQDDRcZHhqcuZjmDNQ3ovC2ISb3qbAG
v+CSuvaPvM11BF79YEVCjFYB9zXj/2/vIRJ6drh+t+0oq1p3HCmxgci30U8OD0Td6I+J9M/9gGi7
BiXsKLEin1nKymfQJEcQU9HoFLNVhixhSLcFKWClA03kD9E3YBHlkUOv82sq1ZVQri8oFfPCTmCy
hqSyIDt+Si4DKZRnyrQf7b3QHlPAfJPmff4f0GOn7izmSDtT3h5orQTqC1KeR0M2dx4eRDcjv9Zv
D0Vz/rR4msfY9FOPlsYBPkX195Q9E/+DEPe5Kf9vV3tY4ObaydSqxkrcaY65luhEPg09CcKQkqY4
CAMrr9WzW2SsxWQUKES/hOFsSk0vzu1evZwP2hedTpnvXZALUNUi096MCxiY3bE0zZHM1vZf4RFw
sKSIndjE92DLk6+auDF5Hs+avO6P+sNZ5OqSueknlsQxB2Tf38WLEr4ZUliJHQsOWC+Uzmx5A7OQ
NghjmOKlPL0t2oLieTglZBzjvJkriU/G479Eww3dH4p3LaYL6+iYIYQAlAbfCSdCT3JIm2MvPesK
xhIlQ29uRA1YmVZ3ctL+Ch/ervZsM5geQNeMJnmOSozeUu8B6cdwnM4Kg13uFz53+epo+94ElJHb
6U4N2QqrPUtEpLx5nj9bRWfrMbLINpbQblDgsEngH3aFseHmueMg4CJkMHZiVnVNYPFmz5MEBrDo
h0/FdqoeHX+0VGfuCRkJ2KsZSLK7NatK+ofLlYdOMlbpRLwBDe8gzMN9TnsV9cTutl8fKkHlRGw5
2sQneeOmYVMorLiyOaWfxsU8MlQHjtqXqTFd3mUJq7KNyPuTltbZqbN3Rp+gzT2PBIsB36U2Ryzg
o9sna+9oHP9dBlkYRE9ZoFpi2xS3xI7ntFSreX300Gvb8NvvrTH/xlHAAbpIkLRXkOZ2HprzYPGr
1JXs1m1u+H3+Mzui2Iom4ZNnZSCEqv5kDPJ/XoOGIjAfqqVsOH3RenTJywfvGQJzoFAlVYYvBwBo
+sTs40weomsaD92zUuCJJVegcmKJSfPQMuwP7B/c1hFjNfPQNt3tes528TzytOXobW3YngkQLWOo
zsjrRx6DU+QMvkaAbk7NnvZMftSWIfCMIut5ww+KPIHKdmfhayyvg2g3WM9nYjSugtyy5M8WCWJU
y9K6h2EeDY3Nl3LqyiCvLaWiw7bg/TPH1Kt8gnjpMjZGygat4Mm9HAcyZIPMXI2kY6RzdeHXXOoK
QQuXSrVTPYmSri5XnsaztX7jkZFXkQHJzbDsN8w9xiyRMh3sfse6TJdxli0a/+oZ4Gk52skQotBH
TRLoL1chDrNg8lLgifvf0X9G0XPt/LkNoOd6PBIhvRdAwritvMphTJ926c7BDFFwGF8VFdv7ME+I
moZOQAcIu5j9phorhZ86OlhoBWHnJwpDXaNihwqA2+XzPLtr0t3mAVLaWnwMsyojZNlIRyWwr/n1
sNEZsI08C52XvokkIi1N9DVN3YQDgYCHYkcXlsCQUU53MywXrExIC34OeXE0AQFTAVh8hbCAl2VJ
VOXb/r8lDrWXW5wsVtFcjI0iStuaNbTIzTxDw37EI58ywyEuL2zAZb7mpVHx7T56P9XHYHBlPVC3
WSjYGuK/5L8cdApkwfXGup3PyE3tGJQSTsj3PV2QYFj215x5NcJ/YPJfSwEToAR+7hp4PiEGJj5l
rzmXotEwQ0aDn0CP0T8xAjrybO0fmjOyAfeQ1LxnLTJ+RwlGmQHvhLL3MiH+J7jexvywi/snNFV/
rDEDOknwIvG2OsIX4iKM8t4eQFP38vkZ+8niepCJ2vMzcseWAG/1cEEWdp8bDdbQtsNxSeW5DO17
msswT6k18fhEyt5Msix/Fw4rb4QJcyX7jr/mxZJ1WzATB9dc23R2bz/PTCOfo1elpW9gCzsdGIWD
u+fRaq4MkW6m7xktTRGnjvbPWmD4f8dZIQOugGalNFj0hMv5P74GFKtIrZMKlv2VvC9/tAtUcxVa
nboARQNPLu9S8PkKzxydCWz684muPdP9zwPi2A94baisi1X2FmZk00RLF9HLhLDhuujcC+QuUTu0
02kvSs6v5qcPmC192Rf5/+OX4cbCPv3YXRXZ1a74TfU8pCZLd5n41Lxqik5OSvL9qKIeE81+R1Lw
Qfoe9hk/r3Rnu+bsyn+GsNP3puJ0zKFifvxwGNelBJ6Boy+mcF55UBFHRzhrCMDB3fdw/3zpvL7E
1lU9DSxbkA8hCJ6E8O5aq0KU/mGMGPIXVUprTHNYgWYHj5CS+xotcciiiQ5BPqQAhhnXkwpxnnt0
er9yqAUJ79l8Cl644SjRx7ycBfurs4sUSoC5X38rMnO+F2c4u4v9XLbwrp2islHAnWv0lD6Mb5T8
g4alLZAHcfLTTy31as324ZVQZy0RRxSKBp10N+IFSJlBJ4TuYtxZ29WbeRajWOeIZdy1jK2yNmbT
h4sCruo5V3QXTkMieUwEJiFSKQVBKGvgt2IeS0e44+1FduCyVmD1HeXmJqCUTk1MjwRJ73kaCv/e
CCwloyedaLQbC1/WZy+grl6QKB+9h3mfApW0pAbcytCKFcMKbyGO/uIjiSss2zQQtSFur9WgINUu
E8vIBcAfBlSe8UAInHXhp9z5ew9fuhlQWf/Tt9Q1GEO/1xLg2OoxPZZcAbUDQHHVwB7EQkiKYAA+
BlpzO4LcXkPAKULs3zG+H2jt7VQfBQLrnm+1kmodyLeSnbmz8mTqHe4tfW1Q4oUH27XxXuRIUP7Y
4GByj/7G9BBpjSEReAYnxumrIs4/offuWBNU+o23Qq4lN07BBWFwFDtUBSZGUQjtIGeikgGZnL8s
qSZMt5+M9aZzeUt7wVGPvwTxByG4fwtrhB9qLYciIRXzePLyCq/u6gLkVCLBNtuyvMx79Aolqand
ljXDsauMwi/smuC/qH7lmCRcra8+sz7MMDIIZrqyYEbSiRcHu7XiO0WQU0urw/hL3b+7HOvsX5Ny
a8nVVATbmlgFiK0mqe6YWqRZnzINpYN1VzFwVdvQrbFCFUItFrQ20Epzbyh4UJiV4hkISEmnadQS
m3fRJdupiprHnrYT0dJKHEzQx0YgWtBJhAxkY2bKzgSr4v6p05JQTFsenIYcpgiP1iXF+YQKVKJA
ii0HE3+lgvECcTejGFOui+jOlfVPory1K8atlMi51Peh/6K7c//ot+aYEGn8cttIR9pOAl1aQapr
5u2pwOkcMwx+iM1WcWJqLq7KTVC03+v8SpZJHIkojFVrAho6Ef7N6hPvOGUbpZMB7yEqVJlNGlsO
TGDBXiADcksRTbMsRlYPX7oyOF72k2i6HqB+K0SXN6axeirSQelBLCWmMhPdCnCT9YlVbCPIoA2A
TVeR0wYlG4DPDq2lOeg41nb9LU6Mtz3kBSUqyu2WqsDL0D4j6DV23Lypt9XcFvPw8/Sd8uOZCVfO
dQKPu68guuHISXfPREMsJ0G5S1wDxX6NmBoXpX9gAI3Hja+O8K0dj98DxP2X5M+8rTPUrkHTbsKD
Qvskvmg8rgiNQHjNPJ9A910fPd/69J1D1LCpmNh1B3kXkAVSy2zIQQ0L+cikQIKYrap7vyZ0qVFA
kxdMNaYGZqV2u9JQC8W/02x1V8VAWoptt1VJ6ydBs+ehiPGyG8rRlPzd7RNW95cD9hqDYpFlmg/c
H4FtKS3t6DYErx4bWvsEBIfRlw8kBQIIfIF0Qy+LB4VxguO0ePpBafItWXvYvCr0sJ5mL9B4PpHl
3oB0rxW0s0d+C1JnXxdKetGevDRW4i4gy0Y4hkFlgchucAEM5sL8KMtF6BYzZi1/4lTPLHC7kmC0
BwvBJOC1s+ir1gjvX+kSCHOrlAzYM/QHz37Bp/ABpL8XKNfpFyLlv0rPcixbo94ntcpLcj/M8dfz
6uMae6kaFJmoaiPWQV2Wu7MhAt0O76DymHV0ZJNodTPO+W98vaWzDE8ORVNjYhWWnqkfOMPdSF+f
ZE4aAA88Vr6eN/tlBK5ipQY9njwHolq29DcuUtJnwur25kOPhVRXdXsjZ4msuTYklgNMTEId9YRp
SGgUVCnqWS1r/WJDPoe0u226XKJ4WgaDIU+8NBGEh3DS+Gb+FyzT8Ave3clD1tJ8tOiOhMkF2GdP
Bc9JSK/AKMEeaniLoGJzdjii1sKhoarBIFblPHMPjKRDNLJD36JoihSdPvnLo7LiWbHYSr5mH8iF
kFfG8AibbOj3AaFGf7Q4QmpkK+dJBMIZm73D/SnyyyUqf/EIh3xXYd9a5jzbcBsPkviXOXu0dXAc
2eSxBYfWEQv1btQaEjCoLbUUijeoVi+pXUo1nm01/St/4zMG/YdBqTEBWwDjD+x3eCbhQFSSsfZb
ZB1pFjJhUF+foE1yUJLY6M6OHyLD99ZhOfE4DD1AcRzYVCLWhGpNil/PSM/0McjRMxStE4QpQaXr
MeB1mPUY2KLK3zzqxN1Vl3/twdAPMJM9TNPxIneOlqgdDqZOAHvD2PakDKpKyKLXPbIXUQMKPhfv
wvjDIE/bwZN0YgVZe2vofVHD5Ixxpn1oi+d3I/ZhATxcahJBBhMmI+2qXXDx53x0YKQDL4d1OFjU
QZPCkCexQs4rtzdLsUIR3SfLPLJZrrRLJN1hsEfweQool4KG2JQ4yiipyDQyRYdw0uvAeLM198Lz
jQO+mvlvWMl8WjGIqoi9mF7kzK9IE68+D0KBvZHidZAAMW35l0a6DGUP/70quJJCT8qliu60Vy0c
uADUBG8RdSOFMAoEPFt/jrBvj9NLBmJtppCyvRTHi+O4A+Y2LIftRK7S3JsrWV+8UCKkMKLX746r
0uyT/wPhcPA6eziKX2/zbRlapRnJQ34O0bPjwuTaTnveNRiACe8RvcDUXrGWy2V6FLm87y5gGHKS
fvJxogCmUNrKGtA4Bjmo3pN0mvIDZF0zVISBbGeh9kCtHztruTiV2EyWfFl1P59EQ50FNRgxU3Jf
a3J1QbAwvFmbDa3jnj2goEmQc5V00gXXdzSe9FFSSQGdgYohgMTUScPeiJWPinJ0evVx6GO72F/G
r7DhE5q7b/H2nY7/4wBpfZ587I0IJRvcV9AhAzX2ospGZjKF511bxv3U4mDt9UP44GLx5RDZP8bb
vBmUhcrQXovIycLKAIdH3YdKGrH8gpXjytu0gIvPkgUpa92vNsHWrMLc5wzAjTxd5dOGZqmrtUkv
G+xj5b47re1KrvsnCupq5NfjK8ZOrHGpPjPcT1Rjd5v+yalnWJ8BhZ7HAnBaOosJLw/cDJtpEKJA
yyBzizlqzD85Tsng5aVi/4DIxqFzEWZ+9M/ioIe+Oihr2NiecKaTnhHG7CkGbJshGnJfsJkuqvUV
ZenfhhFgiB8jU+laODcA9fo6SjyToRiaZ3Ag+QR/c21hb337zxoXaTrRG3avYxnL1/I1ne9lj4bi
+sce4m0d+Zh7f6Ug/0kg/Bgvp/nJfCdDbtb7bY2YAJ61tYQN0Nx3HUKC10DBNQt/JUh7kovNcJYE
UgQPlEgdksUgeH5yOuof5TTBT6lXAiPaI1saUEVwUtZr41j3XSuw8NM/C/MdR5jizlIPrBRM5ytd
y+OsAM59QKbuqUHNf3hDrJJuxIORClgsgEBQVH8AqU27T1axW5/InkWrd2ox3Vxhrb0IoyFPqzZc
gYhdbkDROikuj+sd4aNqheTfHLCfk8yDxp5IEC1BKa0D08aS2Yq5t3pbxIFF/yG3qhQt0yGw6pfV
o8/wphlCKzX7uJc0dl5EbVnxALVL+KkWcp4XGzS7hddwXre4PRH7B6eTguSSXwtNtQbpt5oY4T4k
mZmb8rx3jyG21agbEO6SRplzk1FHtl3dxUoul2AY4SRN83RuSsxVWefwOW6uXme6GBeC8As/MPFM
ngQASIexANZKlFptcopEKgUPPK6h2HtkpgMW3HLMvKTMPatSefoD9ZVazwaniXsRwHXpZ3EtZ3sb
BoHQuvWGYA38YFThPDRccW0CuUbi8EBxK/IZNBwhFQ3rcRvyehsVD6IJ4hTT6pyor2NygulfU8bG
kOaKAD/hkdSrBNWPXHUOZvC3zRyUEQ0kBHbKdopzMRJPA8vWb28D/MJrmW/DernciUIOW4Ar0CXy
IvVhG64Ohs2ipdAlSG0DtB/PcQnCXLa7V+wxTPAhb2XFwatxSK1gns5W8SNTcJ3PwUDk1B+dMxuL
p0cqvLNaqh4WOytQ+fEG4JrOr2G5qcjHGFIczE3a0OaRKJdIh4ot8n68fNkxDBM9C1LMV3u8laVq
qTk5gsm59Ni9bgCrRGjjEpiJGLuJ9yZNquMDTBqYsNdGXiLcCi1zC8d1sKRi6jL8YU2RREhWO4J/
7jzyDlDJKuuQTGRe/UeQ858cEtnkv/wzeqoomiE7RCmImJs4Uk3gdOIrVKF/C92w4IYA1aG597IC
V+f96r0vVDg3agN/xA3cJ1pvT2d/QwlBshMGfzSyuYqBa4a7cyYxwqGmRJH4B3p5vOL7pp1ZcCD1
5+Ps0H83aP8kBlRuf1k3vHs96Z7ItO/NnZ0nTinbX6CwGsDiFRurlFAs6DXYavGZpOsuv/k0smFL
cusg/2s7qZ5eMvKM4nYgcuY0NdhZCRNJcsjdH606I1M=
`pragma protect end_protected
