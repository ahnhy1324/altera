// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qAf2VDEFPdCh14Y2jzRvZeRMO3SiRDyOHjGM90T+mNL03Nl2f/2JNfOQzCCEjNZS
c/8egE0r/g3PuihPxf8fA+suoqOo2dyJuRjn4fUwTH6JgDTbeZV1zoGqoC+mwlPi
OLDg1RCgWeaxx42rb4LFNw64hxmyOJ/vyAPe+p+k6KY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 86352)
7Et9k4IutV6J+25goDAhSKOjApa/bswmYiEOj7tou5AAEAaQ2No5suVMJU9jSxZR
rYGZP9oi5Z63iYe7QLl1q6nle9H/ZFVQxUJ/rlM15fh0pYoWOQjbxFV4KfZHJIeP
g5xXw58tEmy6XQzLh8/xBib3g8kM3A1AUj2SW8xI+k9CQQ4dwjSQFfJbuOUsaxXs
Xoigu0HsLcBQlEeuNDKxDcPl2Bt0p2JOlKehNjk8aVtHfYxuXXi44TPsjKCxgkdN
qpPWkYR9yNFazIsN3bMdRLNfCBUmFZ5NCygSU2a6B7E78RvD7tAyVDcY597D14Bw
C1MyOSe1HV2QbeuVGe6s8UM5OQxRzbO6X9sBFTS9+oK99QGJ4DKOfvaCmXFx/nb6
ebXzSuJMjPAQagbHJb3vCgWbjY0GxbByCtYDNtOmmLIrJlsSeq28g2LZWl8k0JqN
nc+2nfHxgGS7CMVu55f2zlV/XyfZi6d5ChmHe1EPbqRet1EAf09WKWOq8e1y7/eS
/YdzZxVh8NNAVFvJf256vJW/DSu7LlFXWESv0EvwvnyVVGt3IYJXRrkqQTWaMuyq
5+ptfGPdh6WHXmpgENngXQwul394NJtBK7zgRdLl0JPOMYN6OhHblewvjlTbFOzp
YCxDQ7XrS6Rx9JujsGxvtbKUe7tkE3c+nJY+z3hpZyxwmwHaJ4jl4c1bjeVBTIxY
Qij3U2pTQImSaVTefmWpotuwdqtBbFvw6H7r4ojMMazkOcwJRchlfjm2rkNTT9J4
fSndwU/LTMnyYn2cI78DA2Q9dvIv0qQTuBD6ESFVBf/aPT2DsgUX6oSbY/0Q17ZJ
EpJb/VGurnlgjhxwNzHTYSit64aRJ9zRmg++IiGGRO/h4mTygYSZwP50czQ/qMUs
5cWuASEPjKVmN74lBDF8r2Upvb1jr+EYLORCZzkXkqwClBeTs9jRACWY9jjmFZ9e
5TbjUVgoHs0zEjiTSxH/FSK8FjMLYnayNEkXeUsI+oR7dyKxrxUWtVqE2YQtdlMa
H5H0QdumpjnJ9t2qiJVn9Y574GopRBNOEusKaDCcbNsUfCv+3GlYpOmyUAUPUqFS
gVq1PwTJNi1gq5KPC58IYUU8Lv83SFWnjkY1cqwxZviA3yEjfpA30Ayu5/1G9wSL
qljO0/4/lKRyVu+NWKhHHGJGIBjA7e8A39nN2VsfQYBq7JPhnz18o1r8Re8jHMhZ
ndmMspuZoOx6Vfb/KBYQ2b/hZnMZpth12tWnGh9YFnLFqn1V6C5JPJKIfcTg8tSP
uTU8R2jltpkqiiQb4SLpFunqFo+7PWvrzsJozHzQsNELSVufDOY8AiuVRVPuZXOx
K8BEirKkkLWUv1tKB/iHAWqtDzk92rsdPueFIv6Fv5rsvldMeb4b5Fex1TbJZGzW
CxWGF9XXlNVAWZZyNEaSh4bOfYru8pOZ33M48RT06NgeOJHP9HCTymRhX3iEoi0V
rqEwQcfCxHQWN7ELEV8M4+1hhGsCQCuoRSuK68K4d+IGUFlnTMQJaejr8n/GviJT
mIdGb1fuQkKUAN9OcitOmyfGbJm+pG5hoGpEbk1Qt35l6qqwOV/utJZwYnVa9bf/
Y6FpIaQHPU67T09TaxKElX7gNu4dve4xSNerc8rAFMxVnVYLDvYG6s7ECY3H3SeF
+C7nOiSmzQovEd7+2tN/T4Ar+c4vzOMQ6IWBUMpu/ZkCXsIcWCHhHUHs121A6CVF
yzps8PWy30tQDoTWGYt/TWojOtp8XtyS7iBg1gWPU/fwzh+rr2VYFahKHwbSX+2d
YeAnmSY8vxhWXwqDeB4XyPqfZLPizsrlRr1DvGasN3oI4/jlJZxFCGMW0rr2Yybm
2T51PAmC5uuaLosOcVeQITmICSHMvD9FmhN2/SKEnr2WiL13k6wT7ATHwy+12brW
G+WsXyMV9FGFkCp7IiRDzTSQcfNXZjhwX72zJ6nkzDvArPRTp2ZlTV9Qkj8oGbgB
xTlyPkfHQ/8QGhiozySWIFQuNKJYkd2TTd07B+0cW7YNV1101590Nr3m7f+UEB4n
55L4fSRmhdxp7VEMSsOaZCO1UxdX8dknPMwp+v7nruafsLMjiyNslK/uZu8gANYe
LTIlBy+aj+Tb9/YNFRyI6udIrdXzC+QpAUrxFuWENvMUUcFuv3FnRqVIs3K859hM
HrbOlp6P0lIUpBF6S/GISiYqxeqa9hNZxp/9KMqoTYkhJ0Olh98dtwFVuHR1YbPj
2iNDXC0heiqBZPEbqu5fWJeAkRROBS0hKuGX0jltaoUnyUnJ8eUCtj1k6hotlYcB
VUgYn1G7DTg7BeVABSG8v0P+JeShow6VovDpXgzfSkZEi9F6CX/t0LDi54xCe4eo
Li3nRfl6muW23O4I0SL9RXKhn9YyLNWxAEmcCkJznGXE0TR2Z+QwIwshNNxtntWS
CHLcHcWLR5aKiwN0HEfZyAn942Tc+pnw0e9JIqIgZbLDCL8Hrw8o3CoMvfIe8xGn
DInpDluAe7DQ2epyme6ball7J/anDzpGXW5qkItH60AUAxHiUhfH3NIbihxnFEmQ
zhueCJZu+YaCHldVc5JjWk97uG9xFq9u64XK88tIF6xWLvHLWrJeck4y3aZ1SBRk
EGnsTuXEiHn/0ahKCuxwXxf9BdZGaBJpmxyC8dpg77oqifQvDfe58Drwndu8rx8g
WfVZjQx2xA80+eAMmIcoPB8+m9v7G/b1UKSjn5wnHLebuRazL6avHQvBvQx/JuvS
1RVCk5ZP/MAsStZpYSlmLCcYm7vbiayVQSSR7bzOO0AzjVJCOYo9XxV99Rx3hMg+
6bZm4u2MNwdPhobVP2cbBZ/zBXlI6Evq8p0Hw3xKycOxpmH8jI5E02puQzKIyiWk
eEbW+f5jXdrC+TvSzKcPmrj4vppudW4jdGqpX/+Mh9/chZnSDkioXXaWuJ2zKtrn
qMx5VjPWr7apnfTtjfDQvxmgl0ZkQtaoJH2GnnI6e40cPKKGIiBqzlwBRWx/ABXt
CigXFSw86pBtq1tEDjIwOcTamVbI57shvOpcptV/TSg8DJVHFHdKmoQuXHLZPa7j
rn/Hgu5rkKuuEX7Iq6hj2rVxB3Zj9C+nGvJtSgnad33JlzErUnA+feuswDqnGAfs
aSfGbu5n3K5s9jW6MRCiHY97wNgpLuhpbF1zHvL4wIZvkVz4BP8wUozjxPww62m0
y04OQiYiNa/iPH9xrN+NJmFwATmysh4D/QwN0CmqxQEODAakWRVVVo34CtW2hbgC
mPu0IBZDFuc5jhs6B6HqPl6NfUl2EzmziuQw2TpGGCgca1Ye1xlHhtGdpClHIEn7
Swif8fSmwOfybgrqBgJnuVd50U7Mn4ES0ZFtH1pESE7bh5DOTg1IAqxN7ElAgQ3e
Oc2r3tfhQCXQ1tXf/OAXHnJ1lk0Y/gAwg4tJQkoOs4Ys6t18jrpMaf6Dmg0lo4A4
KeRjgYIC6dfhyqLznOLH8PFZAWw1cNiRCTe8yHLM4rNbYfTux2GvvkDehnwx8OvJ
/cHdhPzEuGnM3kYJcyb7oQYzUsMuOFuYHYAlSFtjMNYria9K5x+xSdzBwTxamQo6
4ItR3+LAWwtGHQJNpw2tO+zvUnqMJNvNxJPrNNGJ+7dYvS4QWbrfSHYSbJYqwmix
Cjp1E+PlnJSxcU3k5gzbGS5Vc7J8safwrLt81CpEElStoGxOD4pkAVbWSVTr2V1q
inyGgyCSa8OtQtrjfEmwkizbPaKbiGU4lUSZLVZLZXaCC/gaFw7FpdWxA8/mJjnq
Y4wPgSxLhZZ58F4gqCCLyyLY34KHajSeahmt0kFeBrOja7XH0Jk+JDUgYeL1Xyr4
y2FYX18GBYCSxfBCRoxQsPwKq678Kiam2Bf/QYfK/5nqJdPiCrXYpbZp6XnqiZm2
zcdmvn9pTiggloGT1yI23zT1FDL+vSlThnOQHZK+o/Mz9s247Lv27YEF0tUbEvAI
SLNHP5lShK04CNqBayHt9FTK2yAZXdCaNUMyh//bFJTscpITqfP8g+fc2nnstZkh
MAdgieJSl8hfxqOXuhwkcqldOPZRmSTgdoZsqXKHKaGN546z11HXc2oW3N6nFdt0
2uUueQzFtIia3RkM2y4YqFUlXjZrB1McR7Ofb4oVPI63Utf5IOn2XGRZ2R2epCmI
AMsgOiZR2o9a+85s5JmD7lvKvpCtDnoL2ABt1aaYQNnOVZ47fh0RWNAqoNRP2kld
Q9nOAHUEtrTh0o1l5/XYTopGgfTlpqnLeEbCl/flFnGdAiRKpG4rC5TA2MIBYQx2
uPsebyXLhteK0OVb1cCinSnR6Ig61mSWVPe8DXqx3bfDw5xEi0nPe1HGYz+lvQFo
l3JT7mE2mMaM8Xdgmarnez4CIX+RY+lKEfn9gwq/Qdejm5QKrcg/45iWiVI7p1SF
ebqZBZ+OFmQUHosaEmyWpMUfww+oaQ4QwvyxC0DK5KkqRZHsZd7BGG5kxztGmzp6
PHQnB9j8R8o3KVGlTZ4kNpI5hOWmg0wE7/igfyEu9+4SSOP+bZFC6Svc/lVV1XUC
hJJZJksqowh30B17Ls+PpcwgWuEj220zEkhVZyRsP5bR/Bf8rsmZBxsld7oEyjSG
TqsC5htPrPZnWdsK0bvCnWp51iBDhMITsPa1NJe0x70DqKXqrAnBrkKHJLldpGYV
uBtX0infOB7oiH8YCIra0QC2lNFj8q/+k+Xmxlzl+krP+AQD+iuWR6uJOJe4JspB
d1bWwrUywvJxcKqR9JldD+9d8CM9eap6csh1y8Is3h/D+OX7G+onINIrzo+U14OA
SJv2VrCEfS2uh5EgaiYGaF7SJX+lEGj5BlFWCVjP+6wpM49nF84zR1sDfvE5IdI0
9NoayqS3S7Act27QsHhe08AEo7tB+Mf0B8F4qNWVR1cZyG/+oYsV9B8QiA/6RRUD
dT/nVc81MDIH/ceMR19pJLB7hg0QakCWgchufoCVzIUQU87iWh69/Fr9fkYZc5Hu
DePXjZVZnic+wuJBrgP/diUePx4IPo+F+MeRenXDEGL21BMtf/UGrjh8bXdrvRAX
nX+0QQ7KNxlSHP0XfiGWxWkNdjEEda6ShsN/HMMBwxNAwE5daTgwQYlHoVX+PtI2
mOWrV7HR4kvORQliB/HWqMZtLT42rojsAFDpS2rlT3pR47jBi40gdXCyusCWc9GV
mdAfw2MRQ6Fgyr8keNwlMradzgwJDBNK3nNooMY9AqlUkjcJIYJPGGpExu8cjr5x
QWVrbJjue979TDKumQmvCHJCEDmdsb0P9XqntBBBu9JD2dpGnOK5vxroFTz7y9UD
FbNZbec7HNvOBkyiPw0P86kfdhEP5wfhhpJUHQLRUtW+wGRyVQtyZyMnOc84B0iS
WcSa7upTRYsvso5FT3YmY5wCjqETapc1CKULbiat/ZN7Jm2bEz12u4gje8iVbN9C
gJNyL1XRH/peM3yha760cWk9wGwWLQ9h2Hp/xH+rzwjxT6d6HNoIogYGAxueWMF1
6nJIM0N5AwFVra+cFFkjqUGMWS2O8fZYHGbJH6+f56ldPoPqUhPZkjrf5swdzB82
/AOOAz/zeNpOdh0/43SqexHnzBM/vke9DLNBxr1Be9+Tz4ROqjxDdyu8XZ4skaVD
r1tUGnKiL+fnBTtW2sSmQEown59CCiFTT4cCpf6msVynUlWMQCB0ShQg708b9uf1
0E9EMh6qy7QqX+GuGubmJC7bbjPFFGPb/jH0h6EBdm/kJaDBlnFH5Elr/sg52ri4
nabVd0qefzxlNTtw3zFFQtA0r0TS0FojX5uVx5OYAVDI4p4HFEbh9s2jTFtKwV5W
fGM8uEhoxws0H28klZoObmEPOCSHqld4aGv417hqc5vr8rg3goXxQUlL27o0vURR
Pkk0lkM9be+wDuFH+cXKi72FBW9RK7MHMB6NqyKKHvx3bq3IRlQg/1mYGCKJ5Z7K
9Y40ZmIkbO8h38Gf77mdICU+JDr5x6ARoFbexdDf97FaTAYceRqwyyjhjmgIyDWd
KYjcmw+/p519SvOT0sWJTXAmhajw78gSBPD/6wtowBgfs6batFoilvj3BQmosgA9
FCC7foNptSAUQWf8KdOl7XwBsV/FXHiNjtP6+unArhx2e5v8rDIv2OpUJiKQy4NY
tfEQXmPIVGvvsQS71s1QqmjX/wS3+o0zAU/kFAoqght4FBwpQTf274dxn5aypjXK
29CsObX5P5X1E1AkFh2AeS85+iCSEbBbBOTK5Pa4G5n0pXvP0NkJKdDD/76jzY2I
bkEEGmc2MkPmcfGZ2RKpag4U5A5vaezBjQfoCQ+T8LpuQHGusK2X05MFssNxS60e
ATOS+y8B/yIPQ/kQkCr6xO5Xo2Zqxf7EgBPUOwDaj15yqOli5ZnhF6jWUgJZXwre
/9nP4VP9o5WluKSWH7JbX8UWskYCsybi32LMiqPjXW9tLmVw/qS7/qws3TWQEBtv
nAcWLUnn5jpcHVun01jljphaHDBHNVdqheIv9/9oy0GLXCIN9vqY5MN+gg+pHcu+
i+aa6IsSaBijaDKX4Ao3Ya5SkYe3sPtVg7IqKuXZORyv1Ij85G+gZwVVdV6V5R+h
KYdr+uI3tuaKoUJ/Xi9B49I//24OHiCPu/S3GJLyL5C9R5INB0GaZHVfDyFlT2sa
K2FE5XYjubD8KzWiaKjaPxpkUqM0Bgz+regeWxwj40t42Bi3HrgcnjM44c4s0HQx
3MoWIOu0CeaqRwRJ+M7Fmw1A3IB5eeIHIDsu42/p7Z2E891Y7elZnPUqm9pruxGj
5/XwaPKuwNTFYBrt2scjv/cga1DOIXw7YiGBvR4lt2f7pV2F+0Peeci1lqH0Gldl
t1cVj3rDQxpQEyMAoObxrK2tQ4Np8Qw5Riz0WWoy2h0RGdjwIp0YvOHoafMx3ohK
H8eIhlxUsaNT2ijZMD2jaIZgh/Jg72WF8co18xQiXC5J4qgA6+C3lIWgTjAd7KMD
GsCF3geu4wXNJz0wvlZMN1jKDvKNAn/Fr02VuoAmcK+UyoOJT88FwtiUPmTC1nwP
4c8a0I7qxJH5g/DJf/JZ86tO8xXQW4uEKz09nmBsZZ75F4beuk9WsdaZwT6C9ngc
hwEhgsW6NQDF6LdjaOtYIr9Nzz891A0sZ4RoDz0VxIZ3yBxz98pohDrFh3lrKGYV
qLuXi81fSzBWmdWPktjaX4AD9V09+aRgiDLE6+SIAii1wxgbso59s211V9i9QXN8
osuswDO6h1MLw5/xH5VsK/XISrwI28M8qGE1htD3mySis21G0hbhcWjqcyfSM1z8
X+33Fq33SwvDDf6WihcgWFCLDIRXoMGuAHtGh9nXpgXpTTX3sDgCO+butiH6ZYMC
ZhgJOTefUbCNXDBejpH8qERWFoWcyyAOTdKVWRD2sDDVmKDY126nV28wLPu6J9Hd
7gHEpU6OA8GqRoAQd0w2IkzWLhrQCZZMoQuDL9pMD7NR34VYViEZSnIE/ayBMgW8
arzrQM/3ncDugITzfLhNlZ1w8tOQiInsXJc/KCxqCFR6/b55skDBLyuB+cDhF3At
TY5ucE4vYlq8O8btIBk72++FNWx6YuJupKUreDKkakp4CYsCpQvIlJFI79DOL172
RHwECapvlaKY6xJMT8leQAjzOz27AQRrp4AjoDk8+haMI5G1vWVsoM+NXpSS9aRT
ERl4dNbwELxUPWZn0KtbRHquxuQhjCerRQFo638x5iL3esOYB4h7RO5iW6qj5u0a
r5l+XWrbXvIRts4q9DcEyD7UxrPf5N1thVWn4a2xoQ+zYYMVD5BIIj0R0XpSpE3L
kEI+7W2v17/dQrddPZQkB+cCI2Zgji2wketWAAbc4jTZY5eCosTozmjN0mTRY7lM
CjiF4vdGN11CV3MvBllYhDht8oO/c36BcX9JEA+/V3aFhCEN74fLSi3YvntNOBNM
DJzqoRzdMcSn+Y2mJjeOtPfzRw23KOkiJPMpBNAdl+KxT7e2mUUcI9B1/kM1Z43n
dtGN91BpLkkSJ4C2YcRTiWKBXVGLP5RK2w12wvDABZ7hp7o6O9uqWYlKdqaCTXzB
H0qZZsVo58sqghez9rwY3aWeW7xRqKQ40e1KhY1qJsFcrJ1jJNYGMmkOvkywze11
6YedcA7TAehD3IdpFYtZpYu+5CzwNFvPNjWdEQklXLDl2ywUajMn7+uq93lkDCVT
ixv06N/NX9eFegpgMnDJESPg9nsce7/JOXo1QXaaL2+Farcphg+Sozyy0uTURvhy
vXu5NL95rzVO7plxpTniMsnza8PLSgrYwt1IJ4a8qizxVIzWVUecYHL/xtuU+IXQ
dKN41slTwZS4siJmjNhBeJoQCE/uaVmg01EZAUi19uDucF2Mk6B102brtOyN3coQ
wA2HfHpgVjHvB0qzC2CDz8Z73xWQZZvFLtI6TKwZ41AESi/apFsU8P039TL3EiQH
vVhQJv01DlVl1OB5a8sBue6i5DI1UN9jyU41vknam8sSjD+NBBt5JGceORfJrtah
dAo4zHrqxHZPQiy1grS067xJrcb2Wle4sQz3JaUMreFwo+KNTAiBUtHB4nFOsQuO
RlhWbXxYQY7/cKaTuiRywfpPv+DIMHF3P5f5xZ+cTyJJVT4kN2eUVUlOGjH9LCTG
ehVFQaW9kCVKIlJaJZ+vLZDYL5YtXWVQ0axjr+4igLkg3pV1/46H01rnDQmBe+8P
34F5YaG5TN/RKR8Kx2qPzfDG9hv5iy90Ye8HYYWbJ+/e0o8nVZBYesuoGPY8wPkc
7zNnLqsh6F+Q98XwqPtk/MWOoH2n/qKP+UJn13nv3lslQ6D4/UIC/TtXjyILhP9P
ZWhulmWedS0+q12MHW71Xtati7AcChuAAG9Pz+dYw8lWB8/t14IUW1RJqXwy59b/
KeV++mr0QfODUKI/huyvPF9PAtAdlYAMlj6GeTeQNlDhXcVb+md/q3bdhF4b4fGV
WGuzZ3BVmyhfPgK/1bbk37TA6zVaxZGdULNU+R2rdednZEVz0xoR4++6rfzxvCAJ
M/3JU2ISx7C777DQfDsYhF/0BwMyZ+7YzAtLf4xKcIq7n2ryLGnN6MZKms4ifGNk
sTOz7wqWD6e/+VQK3/3/qbzv63mO2GD+ZmalTIaHfaJPQ8i508/4mgiWS7lr6HmL
9xpNBZ2XisbU+FiioNWaPPznL8VqwGU985bZfCDIR8sVf6jExtyq8NB17BIJzs7R
gAtOkIPCGSe1K3tZQqv/sDQDqNT4KMSzPkVfvl2pjOlfmrCxfjbDSk/pi0HiYSBy
osvu8uvm8X72sfZRUBJ8PEuEEQ/vIlGVFMM1YqdWIdPWp6KjzVldK+7XdleLea2g
Tg8QKaV5KeWCtmqrUrN7J+SYaTcbODwVIHOHCshWhAYx6LGsj2nR5mvbFeeQ5K5u
OpIhU//WEp9wXDjTHy/FLzNEWYPhT+NAzWwIdVTvHFv1qp+v2Z7laj6yx6bRpVrV
XWMVu+e82oDeyTltGSkaY3FjUlKKsz4/rNFmG2P84TXDHz9gr3+STrDKpPC8oeRo
QxcUG7oyRYh7U8bszS+H/1DzK5yZ9DW4i02Fv7QH7VJU5PtWDgJKA0eYNpQCfkPB
PtnzumLKBQvSMEZLDoaF+p5xwjtcFSvrC/w6qU8iqPs3o2calJwiWy0yn0BYIE/g
kCQEaye2/qjilX6x/Mn6gzB9Nut4MbEeJvbc4sd4jH0VgYVoWav958PCs7TYY1HS
W5Hb+CJtUlkAmrru1FDgcaozWb9Ji9gn23wVx+jbPT997pHzGev/T6DGq6XvCIS/
1Aia+bDi00O0B8D1yNLfO14coAi8VCCdVKHxgdGII19n1a9Wy8TmD/UUp+p8D3xQ
3jgYetYbhB/BIGJqrp9QkxZPKIGIxOc65a4Of3F72PvG5QDKQpqUtHGk8ND2blU/
+I+O4ZVSTA+sK4Fbm2h0pqCMD3drXY+tYdW4py0CtfyvwiFDDLx/2+LRwfNs0vnT
aRLskni9tnZZdPz/TicKyXrcGLCdVpLHvmXGNOJJnA+YUSo50wLtXfMu3WyJEQRO
oV+jSrb317MvNFNN6gl9qe63LQDQsz6i783HpFWu7EWqEbIFEZ/FY591HIpcw5sX
3nSV8YhMpRpFZc7jZw//b+MLQfCeMo/X3P7U2cGTbViUdu1tB+uCs68z2vYF8P35
38J/DziSiBZLKUaPArlvGQwShf1b+9legN8EZ7/ATuNge05Wn9lEwk8NsIG/5DAH
PSb2+0dJdC7GOSvXi/j0r0cBgYVLBLZLs+40WUfKY5K+YIi1bmg48IQLkNOIIXZb
SiROlvTnCqICZWhSr6aDjH6E85gVpIbiYxvFagBp9HFauDeGpM+d8Ivi567UJZn6
nfoaehmbnU9VdWQkVH+IBLJgO1srtqNG+86VVVpCw8AhGqUCGVBGWZfXGbmgWElm
G7R+a1NaGSio02PQae1ivj3TSKz4vKsOM4+bTJbZRw/MNe/08YQTU0qV8TOKHZmD
VZH03nTdHY/6FnhnGgG0TmVdTY3hdeDiGtAmjouNVUXLxkKZqKSDjJN96OtnV4PM
BpKQo94lvzHLi7R7g+2OuXeW0+8xGeLrWATaTuI6NMn0YfBq1kQAK/0RqLXTHtv4
5TV71EjzzK7q8ZGnqOz4qD6fPXsU2dfYAklmon3J2ZFS7qu2dCg0eIekLiaGTAcx
szVvIjx/YlVhdzZ+v/MO8BSewZpb6+imJ7FwuxmQ/uRA4lW+cmfE+S6v9ifGRjd4
TolbUj82DyN6h3239FQ3adbGfRxQK1IA5hxJuV1mCt0uDuM/WSB3cefF7SDds58O
pzr7LBGquv+5V1dYSM34jtxsxLfSzhNxO8d78wxxc/8MnZaY8cHvHCYsRt36ZkUL
NC2rIy32XmweooEpndSh7mS52fmkkKBTefN8k7koYw69gi89jgI/QQMK7PEFLK2d
tbU633jR74hE1YRQbXc2y7xOVeV4eMv7aAdXWsvB2jSsb4/+q4c1oFRwY+niCl0/
808SXhcTADkIwJqMacrceKqLnjXGW62Vh/t5GeQR6DfNWYc580NhMX12DxQVHzp6
5HdMssgt6jc7qaoFgGd6A76xxL1ejcj1nCei5DSMSkSGMLhw71awD5aWHYcbTE+P
3xbV4oRaJl9u0gPuNeSZuBsRqtM7B230ESa7rivX36mG4ZqZxEr7jev2+raThw5l
z/Uwn4+7U7ynhlJX5dmgTXZeb/in5U7OUMwV//ctazcepLNRJeaV7Rr4lxXWuQ5N
KL07furyFDYir1j9cqyYsgx5SUn5ZGWvb3BKQnT0sFD1/MObKLsTscgSNcVjCAhH
TMBSn3G0ZAEnTbHFtxGac6gOSy88ya7jyJeKqjOcCPRi0qFdcCBtYbOab1jEEyej
s0xqf/BkMrH446BCZHwXut4px8182esp+JOG5+oVebAiRa9zMLxwgxg61+ZpoQrO
JdgFzLBblgtE8G7BZyD+NxtLR19iyR/WIpbVqhYwzhyZHHC4NWAzE7MI8w6iaAcC
+C52vU/yGB7cGXJJLAaEOGL4Xzczd7SEQDSmqk9a2MlOgIo/Z7LJeCOtz9xzflPq
Mca/y6ovfCa5CRZdLWCIQ6vcgPbk77sbazh4TEH54/bxZMXEqr0GnubFJQDUoIUN
u6hYlTfAuHaSoZ5uelSNRmiTjNDMpCZKreTDM3GhV8WZNL9RCV4pCa3/5eZ17L+Z
rBB/sHQarG8BdngWqHpZkdTnv5vvxFLMSMsaksnJ00nsrkv3A38VNntjum0slAe+
OmDA/m0ftvfi84TKCJ+4Nt/HNwyrsCexnlpQQi+1dKaepZr4wFuhH4CjiNWesnOO
yESgkkPGXzeJcyZb6Yemx9TYyrfMwRL+6rPrY0zmUjOz6Kb0e6KDAWzDRca1XJFn
fkoPLqMOfjPR2/haIUsKAPYPKeC1ee8Z73H31W4jUX0ePDanViTQtyJ/Ik9Jt5b2
JKDa/ub34DzsWzYkMiFIJvelXSPl0hWUJeNiMSEx+BMI3sSF3X2oO9p86ar+6T/Q
ffJ9mBGgWhyXS/YtdlSGJpAPbIQzXNmx0xeQYStRh6lUxi4wZyZNniW49lSbvql0
s71kMfMDC0L63Ru4ziVPhn8flX2eYNefpNu9xnQyXlWoCIyeRpyQOby/akLdlIXB
VYeYWPKeM5i6dQEIejW+D1hnAi0HFb1k6PZB82lWkonJ+4wD2YugzKZKuYFYtBrn
colr4shDHESf0K35mZBcxbvaLUGmKgflrfM4WzIJz+FIDHq6LhVhPqknynktqonk
V+SIgEwpIGOwt9Bjm4BPhoYh0orGPWUkrIHaxd2HdWwN9FTh4akT47PK01Gps/Jq
7xJZmzhrxrDLMt3kPKV16NiHvOOAJ3erISGJopwlSrH9EH2X/Jw05pYbc+3WejhN
CBWTK/b2SvijDTem4lJxnau9BJfe4mjx3Hp8i02RsAdYQektjAcImI5tlGvC2TPl
7PzZUzI+qz9F6v7X50X4uhqFUC23dzpwnEfhxjUWyu+P04Pqnt5W+8hpSb2WQcUA
7n5m99Mdsk1V3hv7L5qhsjEosNm2h2TrcpS9/PKXZoQgyiiFJO0aq4vBk9wlef46
ZJKm1wLNGLXm9ITjFcLD8+lMPUthrSfTgne62MB+rHqgP3L/QnktJboKE9QSwXU6
MnznjjbjYlu4UZ7NogDt7BRLLN5tvLSLrokRUvHvNUJ+jafF7DEWEiIGNb+VoUbf
I9dHzfTlxS0EwrcOqh+ggHowqN1vajuXE0Oq/mYi0yhTkFkXLQBO8ICZ9deyQvbY
FwYGaggWrBWgrFQ784Tvve3KoFc4/QEvk915wbnA6In1GuBW2mVJ2titLfU16TjF
tTYqthrHR0EycrLQMtdvUkWu4QUlSLtWbAaWudzmaMzhVMMQGdCvDWo0rH0vj3Vl
Dy/qIkBNuDfimPhQrIcaPSfXjtWl9M1eudVO6YKvPZHfbn4DApKW941poN3vNTZq
h0xOurBwvWpeFjfR+8NjBJSZD4XtU0uPy5Fya6dgk/FF3lydl/0HM0H4GM7YxVhy
pARi6vES6OCyhGm8K8euf/J9l/zJTLRDn5iPsn7rlvKfwV9orTq07uW8SJIOdHYo
KBkfk9WsqCMkhIX1gdTmoe3N5jg9aZkZJGCQYio15mw7Ir33NjG/E3maIvka/pPz
iuk+V8UotpinNhMyrkg0dR4L+/LoETtTki/5S3Zs0/oLV+d2z1M2uK1/CUqZpt+s
X0GMryHVMOZ0sb9RdNeMDKfNS9h+FthCgEwzzTERNRpvzs/W+tRno8v8xqMVPsde
IjrJZ9hOKl1Bn7tUW5+tyMU83IDamK6MAkvKVVTq1+BTODxtaPLID4qwIaD4wvHZ
KblywFZOczbBfS1g3m0fUyQQIJKJJEOj2s5o5nwR69EEToeMmnZ73iOfA1vowBfB
BwSv9fFNEj4XAbLAhhShPlzSb3958txLy/vWYMWyKHy/MmAswyrzDoAMhPkKJIRa
UahYVNvoRYT42h8xdklJoFHfD0F+ugaTiGqRhSuwc3HFaPK67QPcmxwKIzVrP/pz
OhuNGdoXlf4PajDoTZy94zhnP4dMD8BPZR21dB/rOisEtnZfAWa1GpnKg2tGHK+v
7YJ7QW0kj+QqXak4//9b7aQbt+W+vwvn2GXeajBYotZUniG+wL79khEkLZnjrCaK
CK3FNLkeuEXUtRfQB+UnS13gSzIcxR2we8Jcd3kS4sE951SIbLeo17OJGebJVt6o
3RbIA99dsq+MLgLoJAJbVFAvOp/rg7/YHzeINJ7tYkzYonpF222KIPvjO3zDxXaf
A89m+CcnypaFRCbKTQNg4fn6bInRp3dQ9XicJFQIWFDaXPmoyZyffFa7a3gqUSQ9
twQnZGn/fsf3QXyv8bQ7YBo+c//Odk6up6xBElHmWJoP27Ton59mVPQiNFPeB/6h
uiT0pLhFvxpMJ06Sr4LQd5W2yNCMXaGUZgGxSrZbBCiK7+2IPsqQ+YeUVJoZtmAy
S6fOq3mpnVjEi5drNX+1m1s7eUU9yZjTwL6SwOmOCuiHzc5gHqKRnLl3gmMC7KzS
GQfZBs8MkwUWuGR+r3Lc2V4Q3v73+FvqORHfTDEvozSo52Y81hS09sK4sdHRkW7H
RByN2QuWmVEUZBNhw/Lb+WTPYRWG+Wp8dVHV5fS0LNJkzbA3uXuqrJUUAGfA7rN5
D9cXBRFIzcw7exInJCIKy/h6y1I5V3ugCLqDspxPwjyUYkkNkXM8P2M4eqpD6hhC
nm7G+w0pxM68YMi/xLudIwID54O7gHFu71qUe0hDtF3jClZG5/t9iwY7gYprL25O
vSmD1/YQuYNJYOppEwnq17zdq8XJe7i3Mpzxd7mAcJhOA/hIpQJthRuD8YOfsLu4
vmn8hgEBX7aN/gv8U46DVPVKk0AZUJTH57D1QY+CAt01Vm56rn0RMARAQIRAcXM7
WQzp7jhKpN9IXRPDQ9eoDE2MZh9UINXIgSs4euqPPKY1M1XxRy+CT0YvTHo2D2XP
SX+n6WVmIxzp/blRjJwhr61m6WBD+qEeaejZguziaT1vNP7hbD6R/kvgIj2QC61x
4xHtRh8Zb7igNQp0JDc0WpPSufpbwewYW2zDTOSzf/Xwr/EsthD9J+NCdDeLliof
5D64qauPX4PaLYiTeGG0s2GKsvW8zEeHYy9pAiSxTybWjFVgdLTIRFBTGf+Z+chg
1zTa4m6p2ITsGxJy//3zMspGyKC5cks940gd+E/tuR+i0CGw1cGnNx5G2taApdrk
WMfbu4o2mGgAsHb3sa8PHyGlwPHdzij91/3Huo3t3VuIPSpCTHIqxT5odyToLXvA
xEN7Zuzs7qtZT4+yBNlx8IG9mkjQM3woNafldrBHeCZowFK8zzdSc9VAqtCjUsY/
KIpeH6twU4xxP0FMT9O2moENSB4Nq4bK7F5PQeBUhS2AoqFYtSel+BmOdTSJQm0p
+2kiUQotcBGnACCjfwRxmdacQgbTOdzrMHl6mSe501NJHo8BzEtnqTtAuS6Y7BpH
2jeAK3oG4yK1uHPkzJ0DAs5a2b7Ou0Gt98MdRfCUsIP+rvbVyLsSgE9XELw96yx6
0FxpcLaoaWGyrqUlQIls/nAvwJsoYvjdSZzxkJVKuFqOSeB1o2Www5yWNdxEg1F7
2R4P04dvPoyAUiXQGKi3aztMVaTgWQQqYilXaRQ0dNH1Afz0aoMVzuBdhi7V8IBs
Am927FFE29UaQlA+4qgNpbfhT87pjloEc5VMrwdth72F7aA8rkCrOeogLqsdRZ6l
F1q+9wwZCYE51iGNsog8pmACQQOov8zCrvnHaMLPca4+tYNjMh4IBVCt8tk4AV5a
83UNblnRLXp77OYkf4UESsXOwsmdgi8nEuHeNdQ2Qkd+30LVdwN/nMRwGhv00si8
gXkMZp871OaZ4zGF0juQLNLdv3G6rxa59VrhZYmSnOPhI0F+Qt0picEf5mt4zxRP
YRBw9lUPVpkIBifD6zCF9JQo6Txkv6fc4sHgLIfI9I7fIQwWehbBtXjLY3M5A9ej
sWbYGyBDfNMSye3pCuvTIRWx0cZoZGiqAKSWlYjJd+KF6xboxafQmQLQArWn5gPt
8RRPPv+UHLbFYvS1lYq2JuVm2fSJY4CpAHr8NcTJLV42dQs7g49Kwubh/vbKmG+h
XZYxa3PU+9nfRWnXEuPCnxDnVMPIg9qeEbCJs6QQgWanrGrF/Pq8d3MLSZfcl4Rn
D0Dk7r+ZavrQFknXIV06jaGSPsBCBjolB2zMxtsQzvNDQ4iCk5sMldiKPIr+EULW
6bhzSUxYCdW/Ra7rBM47vA/3q0TrC2e/G+MOWOnk0uYz0Po0S1b9bD0OCU1mqs09
Rut4eB79tkFmdBkX73yxgnmHt8rY2YliZC6k2rbRYGBSIhDe2PtdL0LBo9M3VUr2
6UG5GK7v8+apDZ5lBfoMH4V+C8hlXNUTsy69KBN03127deBZR+PLsmGq7huMFnrt
P6W16lg8gcZt5FbNbvcqEv+h91Bs+P0/SUJo9Ajk2Zyd0H45Bt6KqVXJI5uTJAwA
kekqDSNZeI05oeUp1sOcom2EyQWWeeJ8kSq7jE9HujJP7Rxjk24yjdAWx7Plb599
1czht5laEGYCVyoPgzLf0X71/e7D7AhfKaf1/waPnq1kEevJeO4KhN1xFE+JG0VM
PSAPTLHTdvYc3FYJbehAIRqPo3PYuWddWrOmujhT0l1CeQVWk1XZcJpEhryIMYt7
SoI1oxdvyFP+upAvtPvT/l2O51NCg0pv+RwBB6DetOTnJ8iBVHjoCeBtioY7Pioq
159Ii8AhY8/lrjatPgr6ZVE+BJxn29DKN2zIBj0/XCrJoALI/gUMEigcGyjiBdBO
XrKJhXHflNzn8s/DyeTyTDgud0GX5Xv7cQCcQngGIqFFL7yCUpuC1yM805kipEzb
QFZR9h/FZuzWrZEq+S3S062IQP4wOqW7pn5zRpaJQEQNDt/rGPrWAECkp4WoHN6w
Mb5KBJRwI3oNUqgMwuaOWtmZAJXwY+z8G+Hb33GwhSVSeXBRvbug0RNcedIH2h1l
XTXR9wRbjls/46nawOlIEqFrt06EcgcLHUE1TcybMqle1inGOQHrhIUimGTrrsUd
BNctavi2S4LcI+xA0+EqZP1PIJFyGrO0EZcfwQqiZXnxP4+cXXiJSaUbRIlZ1niB
13hOgMlwd+Rc+DKqkkNKINXxejkCpMB9TttQ5Cpw6ZzDzS94jukcfrdLyR4xJfsf
F/F0IkLmjSkMeWNdyQ6XvTtKM1yZNysn8ObrosYUb4wxjPt2D7en2QM5Zk5CRK8i
lA5pG0455Fx1iwOAzaxsYU2ek4kgwlhNvFR1DLsQIBHw4Ezj7+7jdI8rgpGFgNyT
mhQtivRCrGDgcdX1spYasW1elCc4u5ClxnaCXMYGZEpmvTMI27sfgPnasTvjAFMO
ZhUw9vihpRaclgOOTYLmw5gXUfpCou+k8e6THzMt1EJn/1N0W6WK8CvxbSjPg+9E
CF1oySwejY8qrxQ6pAZamKE4nF+mMbanoJXrk8orKoNC/6E5zdVP5R53JFxsdFmv
ue+gKk35hRg7Epdb7cnIRewF5hXQ4AQjYe0nSASPH7BYUUZzH2bejAhnZswKen3z
Vmk5fRc9URiHIJkoJwpfnNbM0uZomnFdXioGD5WJQs4W9cImpAtrqcvNjfvl91O5
D6al6c7xx2x0UWVtKbgjr12sV0xDCMqgBOSo+0i6M61pmX07zkSrux6eryR8w3xo
nSk4RUWZZHPbqb8KlCs1ffQgShUuh2bAq90vbDVvI8tnomFeUOW/mQEIMCdE++kV
y453/Lv/RV2m5NZZtpeOyryWnLK8PwZmtuCCihKFtidZk5o39a7wqZoPxyXKkrCb
swVJEnLh4GYMhLr9clMIEaDGKs4ybb3h67/9ksRFqPH2lz/zGHtyawUC+8+6LDpF
pmKNPtltgkqiFBhHIEAw+6IrES0LVI16Ltf+2sfYdYAS0/CfSQpSEzrJ6w1rRJM3
JbkIGCr1++raMERTa3IrEjVB5QYuj6suFd7K27MGv3lOUm7Y88fp6EIeYeuaDkRB
60ZOBmRKcDknFisM5yFNj1YD3EcYtObse7l0U4sxxwZLuNkRyZNsQG0WGIJEfpKI
zIUae8bYuwe5UDfe+1GMAHRCRoxwfd71Ojnn1/5IVuleNyseMwJJZsXnj8SyQ4jV
BEVsbmX5gwRZzNuw+7Ea+KAxEy5eZXgS5pAzmSxL7Nq6EDc+DwYmcL9Ufyr/5I1D
uDqeYsR+u26NDMhx+VUI2Yeen+0Qdo0NzBlenC/Cq6PrQIIRnhj45MzZQO0EBdsE
/iyUMStmyvbqolbx4SIkXHWXZg23O1fd5FkC8aAS4wMb2aaG1j27jkKDXNvoFY/Q
rLVZ4MvHt1MTQewVIahzWSTdJYZL+MUJw3iYasTldSA/Yiwgrv3h2sl80W7KJEz8
vENyO10wb9l/sGRCWX2ECKu8N1669BhU1jYZxOek4IZTf8uih4fMZlQgK0ddaoOP
urUufUDlM8ne7SbjtrJv3H30kBgGi++o0F0wwrhCMLfBVBXCaampgvwV1HzjAi3k
5LTO7wEqkOyz622GRjajUqpDahAHRFRV5UyP7jgbr5mCulxN7HWC9vmzQZBOhRVj
mzN1YbAKtJ6MG3LVGqoNwcX/LXf9PjHTpw7HgASz+33gv3ankpqjC2MVrL1n+QIc
1vnJoTn6VmlHF6toINL+p59nRdEwqbb/DY7IobRvYMatBNuynBOhznFDQBPclT6e
rTJ01EN0GBASC4TTiYe4VCArvQYd5MnoDpl3XDDhzlrtiI6r1eZfkbXE5feJlNAo
TXPFzBGJ98r0CPo9yROYX7M5vlYIptLw8YOerCpIkDWjQF7wwFDKUbNV8SxrCQ8J
9a5lEJM+3JrWI6+QgLChXTyfq+NeX+lt+aoU0nYXQGfZnbf0/Qf1wB/gAKqR41sj
bSA+T8ZL7hKq2oDYR57u7SC7nWUVF1jm5K/t6f8en/QfWSIi1ktuQteJCZwlRo8b
xbXljXRVjBPEscDVBv2PP7eXOAdsF6P3A6z/ILwxaGvUuEWMP3hbNvJLibtvnJ8H
6++VFyMTIhAURnCXWb5jBNl7C++zOYvLAkiWxjuOKrAqtBINUtzVDzhQynsWesp6
UamYznhEOMILS0lwx34SNc3vuoOxx6RG7EM1+gQwBuWvJGXyXtf62YtJ6kcPTCHo
PBR0GKANUUJ0xZ6GpBOeNv6E9gbemtQdG2rBiWGnh1djeiDBLgncAr9XdomceEJW
IeOU858NnpesvE8SANRxk1TRDqs4Avh9wW8+8GE4RLBYFUHQmLZXrYZ0bCQXECN/
R7xw3nOKwRzpz3ylwPyO4JM7E1h5uGFMIbHPdMz6AmTwmY57oCt63LM72t5yHQiI
asSGP5FmKDtkmfQC8w0+FoxN1bN6d7d+gI52j2ayr5w9b/Kl9M2Zc9Fr+MnFZkuQ
b3bLdNU5YJR1wNFeSNs6l7z5xPpyavQNuUbhZ1QX7AjsT6ngapABzDjAnLrTdVaj
yHi+1DB4H3zLcMKluF7qYDoMdJuJ5g71XCdMr2WNhFLQxQ6TrZ/KM/XMspI9CKFq
TTJ+ObTWuXvFajTaN4FyfrG93LyfMtl0BVjfy6PAPcg56dv96HSSDARdtL1jCUgK
bRjG2W7sVLhCfInXIzJoyJLqycsgWQplnY2OCkCbWX4cCc4Kr/ZqnTezmSIB7OKF
kjKN7frou0CvlYw8t+VEFHwHIbwRF9Oep/d9pGylIdJ7nNJh4YzfHbpCbkyKIClS
2l0LvwnpIScNxt3DVLB0lF1JKrxi0++VDAfkD+z2fRpB6qWPk15An5vxD1Yg8DwT
EY7ebyXuCkotvldoKNL74k+NSLIX09qx0xXmVo1lZxhoZyLY51sXxcAMuJkmJZAU
EdS4XnGfFv1+54Xga0g3l51kJwqJO2slFo85loPkchJeETn6HUgIt8AJuxV+Hi8E
cnekgQ1Xke2a62XjeFISfwQ9v9zI0nHSQHdfwRthB+AaNB2sQ+vk5E8aBH1x4BDh
j6jZJdtK8ZKUsfQvPyEmFUUGm6HBDcSl4UNdpd/fGpwEjbuv5E693r6PdPMdmkNb
EQYxK44qPQ+Z7O4jf8YySnxqtxmx+Z8f9l1FilLHvsd94UhaGyQFWEQoqH8MlrOV
9XhKsxoOqha1C/zJWYfWl4mo0t2CMnpD6HBY/q1W2MzYXquTIrH+FSCVdjrNKT3Q
LXdGsabKRHx81ZdobC1IjbCZ1Zi6X7pfaZPZP/kG5Iaan9+M7BIRzgA6vK0RAuwk
Hty/iQ0kG2UDSHVEMKrT7oJDY5zbtr44Cu1pHm5xxRrDcVriOpDRL4ABCByxXg2K
RtfVh1MqzY7YlgKk3KwTNkjdkRZUHPSBW5aCUb6TG4w3euzQHp3WE5x8AUBWdBxp
6Zwm5X497qmLzTwl5nzNwlMqqKde7pmbnZX0iNXKu00+7EnZla+HvFHssiXsR9k7
PuB69CwIOzmjkDxDfY7uUC2Zkt0mB0Hxi88fQnsix1UZTLY7ZIwgKQAQAwtmChFn
l8Ng36hanlgVLIS9mXtiq/C16wr+H9tLKSriCA+ktjGlgrNNps2gMAxKLGCLUCaT
FXhJFevlJmfazLuVnyoH7RHmdIXZmrDL/0Fl+LB2VVdqzgqUHsUA82+IVcsyrwXr
t8dvn5i+ZHDf5mMMSo7OVoNX/yiWYohpP6hy9A4PDxeW/zXzBLZf/HtG9Pxdwtwp
jVoXio3FXSdtJUiTmgNvpfgvHLxUt9Xtm8yajWB01Wcc+Z9V7wgXEWzsCUHZxGPn
BMa/x2urx8rBu2koK8+mxbptFr62wLkVTFzFNgHnYGFcymRnw+P9nHXbBQdXe8Dr
c1NfSfhYuRjyV0wPDuzd1Ky+ZVkcDCMfrKVlW9ZvxC2FpOwQrXnAkjI+xh6G0faN
6KPV/N0D1BA0LB2Ah/G0vbzWEO0/pLT8q2NteYXOrqSYnh0BU1U2DeisXKv9dRqw
51BmsriR2ql7+l0+ksLwlsL0zbf1Duyfq+XBKNf+PWj0kOllcrIy5l7w1LpTj3lC
lUAp9dSmBKqarXn1EjVYdUCH6gWedpHLIM8IXl/ndJMluwnkv+/DswF06W/v7Sc6
0E7cmh1SSXQIkTN4g35/iIIBw5T7upfBZI/2cUzL/+S3Y+3XYMlBxFGCAIRP+tab
5EdKO3EpxuIMQ9+NEtGH7dJv/52FKWTLqtnpP9sWLhCX9bmYNxYA0TlJJgnhKM5B
OrWh72p6PYZWMBsQTVxuOhlS7Dql3c23sisol4+rtsCFummCqFiHdXMQ8KPB00ei
JIEliGHyok5x0s5qYT7c5oQNgeqpp083haYdFrzUOHQSQNokjCm3kp45wT8pPZUK
I362lIE2GnyVmS/WXDCHLOB3ZRXfstgKu7vJT9T/uTih3RfUEzqpxKRVRoz9+tKJ
a/o9/iVEYP+EVmgAXsaZbFheqQZPcna8viYqkwuyJqbIS/yvPrJPiEUPQ/tOp1nQ
KCpxWgo8mL6CVNuVpvp1Lo0dYgP+vWvsgmTMvVtsvdh8chQ3D9ZamTtbRMFhEbow
+BtOLgInjkJBZ1gj9cP9bshhN1qO+TOtqcc8tGTlxM+f5gPXASl/weemv36bmQY5
kK65Y0Qucmw9QVhtD310eNV/RiWTJufxk8EyQWhjtGy7cXmKreyvBm5Ni1ojaX7j
YgScczFP7r6m9DbGyPPHPyE1I8NlWf4ObC10s5JE3dhjZJS320gQkb6uiwWT5wkK
LvHNqF0ajc45bqiKMY+9c2kdUVmyDEN2WSD1bg/BoZDrMRx0mk6ZIiKS22bLnduD
0J8BvrFovSDZL67vSQYpSWIvKzMfiFqwyDOqTTO3Fitw88M6k1fNucWhN9uc1dRI
yX6EWHDP2nqe/FQVi8NfRn1yLoL1+Id5Ch4DEKkU/peTcZcF5IW8LFvrZPAiYog8
gy6VgIdjxgSdt57wuuACdIfPgbCVVU7bvS5Os41dk2XeRm/7GV//+t+BW6K/XODH
vNezUeqF66/pic5Kg1JBp9aPPEHttunxSSj6fQFpGD1bHG1SwkXHl7gUhrkMvZzM
9Wkl+i5r+3el3MQbP74OT/ArJa5nxSdVZvVHq/zWqXmUZRQx3i7lPUbwLvt0Efdg
50+ar/IHHT+Yt0O/sN62xKsBp1esUim+EitnkIcueeue7Juo+5sEP1p8pwb0WBwX
MtxPb4wTBDmM9fqRUTo+deoQYh8KtV227YLuYvr7jxByz+AU4bSNwgEtxaCmlt1N
idFZ5dEdHiS9fRc89PSCb+IGYWmvPfFaSkqBns2xg+OR6QFgDTOr93d7N0P0Ey/o
LCO4bMX/ZARPjxuY2pTJI3c+2lOYX25kO9tEsEJL5DGlfrh42WodSz6d2sug+J11
W6KxOdIezfbgEOVhjQchtgXj2gpdpMxYU4BS73cGvmoW7FrHAMDaoqRzE1GSQpzC
sUut6+lLi5GUbL7Ov85ZhjEHDXJ+sKkwK1vNOAE8HEDvNSRQpx1kFm/z1orad4zX
YkL8woTa1JOCyFAB5lct1XZfU18Dfo34QPqmjIDrsiYpnvcyBb8BZqC0qE7yi20p
y8pV8FetjN7+hepWdtNe2IEhfE/SjKai19g0GpV1S6ymNuiAtH2i6UAMwMpBeNjw
vcMXPuKhzqCJUwASimzYGBrHE7zNKHcGu9FVgFijscYj2kVPAxx1kXlGDJ2fsF0F
pibQjCYjXaUg+zM/6x9xiFekwgMX7NXesMLjjpoWVMvATbxQN/V1sSPWCvRsIdxI
Q3Bqlq9LDSihOdErczLNvZpHE0uO4hrZCIrrI8sNPeIRbB62L4CxzPzgwN2wv9F0
GKRf24S4AweHk5jYXxxYe5viRvYOuRpMrs7pwEL+QrXGHU6ZX6hzmPQbjHMJ3uKw
4il1mah34SgRQQi21IPiBQvQcr8hPY5Tj2wHzjAZ0UmSqmGYWd9oozQqgQNYK2uA
bhVk1kQtuO8VYUOePCx6wphu+havf1EnQYzcXf23zStu0guphyCLYdfuqSuobi8+
3YohmkMi+GAKSXo3eoQJrKBdZnTLJiDoXvDy39sq2PEhbadGIwzFbRD4J7S0FHZu
MmiB5hlst1B0xb+J+4uHNhGGRpX4c+LsmLY4x6lXfZpXvJZLeUcEwWm7ugyFLtXU
O3VQnQv/U8W7AOYvZ+2N6yNRRPN1HCO64l8Zg7Dw1nmczYMU6lKFTYT/twQMwXG/
TpbvYN7+w55cAxT4sNemzzbnoqLcSuB3POmYGxUBtXr/pInnh2izCTr+L00KLxed
NC9UDe0nYj+7Xva9sNpkv94bnpoFpV9oe4grWGK6hn4bPuTYVt2X5IKVflX8V2Td
aigU7EZUUNLyPNSZnrg0nkk2OxEDM/A0BY9iPQTweCjCrtJgn9seeuxkmtPUwBBt
v824STH2MooXirPpnPEyS9989o09ZGVv5bYJFlEynC1v2iNhrTfPP3+D9zxHsiC5
hhpYqLfsGVLNYEv7mQioXbfCN3TlH7fbKKW+aXciKp09ZFb5fkHumhJ6U33dQWfj
8qSfwprK64knld+IT0WOXk7aSW6FLWbl67DB3UQPwOWPRpCKLHhmBrXBPXUtUdYn
va5DcZskJXyzqbN7v1t1dxPcF5aPQGmOqKgBnjbjiZ5x+xu7Uk3Bh+JyCcucUUyn
slyaOqt2aMB4qsrT5YJojR406dR7BXSWujuvkBFyiFYvrYQWxWHQyM8OCAJdDs3Y
hg6DRZfW4NYqZY8oXGA0kB+0rmrr/KeKyhU7OeYWgyo8zqKIfkd7x0/vdrmyXMS1
CD8wLIJl6ruP3BcDA7XfFVS4U76toRcg9StTpcnblry7KvJ6aaoGtm77POXJgJVP
i6GL5QYbVy5ZItpDKHSA9furdWNhQnLRmB8GKuKkIG3i5PNr03Je9To08g/fyvxv
tWIuIMKZcwi1gAR5EChoZ+eJfEVNT/xKeR9wB6onnFDPye0gB6dMttrPtB80ANZ0
26YVcmssWZjynAjnHs3Dgb0/u5vAzhGGzPPMHnFtsA7NyTP+C3HfqRTUuAzFMUwu
aBCGz3uEl9sZIx4ZljtjoDZdZK54kGwG7rixgRq+KVjMDimekyngEZM9c8LEq+Rn
xkVa/ttfJW3SqZkT84aUiyWOqLWv04MSi8YF+IwsONeHTNH83kYWoY0KF5WX8Ivm
BL82q7mvfh0HqjRY4SWJdflg+5nb1AP0HaDBhbm//wzy+oV+OldeHPdwEnq/Fy2l
i24GhDMTcNnRX3vZfXcvurHtKEXWcdFQd7j+se+wSJ6GHY8+uCAIQ5gG5PQO6Nb5
wVo8XAiyRmg/ww8RxuLiTjfnfDOT0ynjfjYUtjCgoWL5J7YvJ15jHuyHvxfEVfh7
oGDtqKqiGzdIJiGS3ubrJN7Ev4GdvXI8vTqFzojCR5NHVxWaOZc8NeiJIuawNc70
JEWtAPw8vlCcbTDxQsbw0hJEW7RLFz+WipZP1Dji8Dda17zLRv3jQ455uoDeXLeq
RYw3c9SKmM+yjlWLkaWCyBmYhH+hJBjQH3ijoqmxeSM/UFGviH0rZEfgEz5wopi2
Nb5fGY006RQZpBYlQyNXjq6Llv1VjWuD09mHH0M7B6DdNhITa+bj+c2CV5FAaaHZ
XAoQXgolDOiUurILGKI0sCdVAm8BMp4b4RLhD05UZK7GARI33EFO84fLy7dJO7IZ
KNnMF9sAXbaDa0aeg7lDyslhEHWiuu5ErFAI/Ak6TK3loXQauL9f0Hdq93o5EOoi
KuwXZqpj+TzRDh8azPLEIeLOe/KM6SZoSMGxaVcWSnldHHyzJquivLuVLoRLVHQJ
1lVN/uDe6OVKRkfI+4noLYcNjEI1M5m7T8ebyDodwmz3l9XMdHCW34WeJswPruM3
8r0kXhbCbVqsAV/ObK+RgwH3ORRDHn/hBHbFEC/AFNaLJuOxwIMUbM3ARx2ujZBZ
CrwDuMxsgfMwosywHeyPqv7jyrGY0gZTqUwdNVoKU9rdtvu/qaYhPd3HHWarAbp8
Anzdgif8x1IpL8gyP5QAfpt32QMWlLht/Ie3zWglvKCN1dPFlhSiNKXRaCvf2Dsu
aphc9FTibri/z6sc1w0RJHpmcbVB5U5d7Yybj6AAznu0bMCKaubDvk6A/JFMYjvr
mzr/Sl3D9wx8CE6y0oGyjVK8zGu7kOI5QVnyynz98GFZQbwA3DJ/fzcwH78DA+gG
QR6Yxp3AFzcg+PsegDF/chFL5+H+8A8p1QDDu0hCWKKuLx3ZWBD+H78tHrZs+QZG
yY06mzxURnn+uogQjWOTWCq6TpWta5KaKRWJNbUrRfyVS6o4f7LXtaH7hGjBjcJY
xOg1KiNxoRxsBdIanCt/s9fIQXwRvslZeKhOLytjHU0x7DK0WTwHB4LDlSkGV88M
9h/9KJ3Ptoa/v5e00LhK+izd5Q9SkWPy6uVKimsFXgqUFragb1x5EsNBZ8CiB65r
C5uQNpvs9pajcXGh5j/3i6PjGzXaaQTxG4J8xnHO33KfhfK0h7KUGfzCUyP3VkPv
13+QIq41Hwt/tt/p92USCkGrWwl4MZfKWRL/il3rJfDnKCpt5PHiNDKcyBmumxBm
mpUsNoN1t5rfaEbUHyoLSGJfonZSqxVAr5jyQeVtXh7i5F53Zy5RZZ/qvhBTQ0BD
z8vMGa2tDMjqXjuGCu6MS6zc6guOoQg5M/cUu4x2A3OV773DgEmPJiKyqbyId9Qr
Lr941TShcHpk6Jas/gfJ9mGqOFqaX/JRYZKJYEEO7gxumKwZYbXkB+Kdjs7+N6kP
DP+2qlP9Ut2iYiQ7cIDX31nKZ8Z8Zec1jMOje+okTJvZ994wl89rT+yLRSRYD1/L
Ch7lklQ5eGL2p6k7RjY00zZ1Aq6K8H5AYYAxzgtwF35v+ndjZCVzkku6J59O5VRy
R7zlPQhvpvuiXlz+T5e84PO651xOjLrho2CwMaNm1D1T0Ehi3kJ1iif5PHAS2nbE
Z/0CJ96sOor/dag/wp9ngblgCmOAHCq5AlW7+zHT7+NYVaopfJmPJZaw6fIF8WtS
gH+OPP6yhxIlmTY2K8hqU5RZ3GLd8eCb2I7wQ76n6vPR1HwpCiNrHgNSQRjvePsQ
m8Lfum7o6osGPA2717XyiaLpeLF282hyvDLzNgQOhAzw802RjgBipi3N+gG61T6s
rDGHcv40KOKoKsb6arf8MfXdTevtB07/tIr93C7jcxgILdOrgE1AwCn9mcu6I09v
8syoKYmbFSNh0eSAhji+bT5rVUXUKTRqjgxvdFnDJL0a5u09ydaNWOs07yTx3ZOs
eHCOhQR0HWCIxZOKZvg//Zf8JUVrhBLNOtyNF3w+MmW7Bcf+MwppAGbVY0X/DH2f
cMJXmnZpeJUBSpjUkOhh+r1stbQfpPZ8rakQQf6EbNHvI2+PclwGGAiZmRjx2hp1
de3Rb9HgIq7s32w4yZw83ANX8PsyPbGi8So4enS/scuYdRCbWpfTKK+brdJt2sMl
tLzax+y5NwYB+9+liz7wTeliZHwRzp03laTAvNlbPpJgQ13S6pMz5dsnbtI4SOFk
paSL8CACWl4Aw9ldVEYQDIjl6ifN+IWQ+aTNnJNd6Noig67uAxoiGTv1Egweb35h
2IJQgLE7RKG1/so6Qq9P8YZzOillaLk4v+tfv7w18iKk/KhL3HIIxe+lhZgksl7u
S4QiWbl5LzN24zZOpBE35yWs1b/+gB52TRzhfQit4iVDE3HYvCyKdGPk+xhORvOv
Q3cHCbrSKSOvfGIS1x40dWGxSc+LAgk2tTK7hdmUE29WjVqYHf8XuiYw128mEyse
Oz5+XdC/ugncTxZ8IfzG+q0330f1+zMIqUaXTcSMy9fUiaANzo6jufyGW5ttnlWX
NAYezM9kNw4wkGL+komLpi7VZsA2U0NzPRSiYlXW55HJf9ofLBi91Bc1iOJf8H6R
ZoGY7FP/xM89Mf/4ONRbN50zDLz2Th13y96xK/FRz/EOaNi6GraayEBgibWKsc4/
aNLV04bsHNFkPNF+a/CVKdTsTRBUA+SJk8f6e2g+GUwg1Uq9xw7DN8453m+226sh
hCJZSnUMvhPIm3pn8kliNBmKtwyl8mpYi9VFKKYcY8bIL9iXO5Q8FrsQjN5WD1uf
C4hc+RBXoig4FHwVDnn7DFcUYHde6DU1si5aLdLN0lK8OLXO774VceuY5kEaqntH
Lau02z/JDVLwQFd1eZ0N9SAoTtMDWjTeXwaYtW/qZbtbkNzl7hzspDud7b8v+ioa
Z0V0PW7r+CLnXX5uPpzxw8280mo+ZU7bQZFlavdC7oFqjWcChGWipe2sfEpC2Gtr
bVzJ9cwXxWqW/D2RKXUR0aUtcmXpz1+ylUk/VZQY1ityDSWKHDWK/nUPgxy6Rj1m
EmjzJyXuxMGnclOzgUMyWH+FW0hpvoik+uw+6RwO87gi518IWrl1YDt1rCoBPic4
c7H+frihp40S9uBEQdTdMPNhI4Z7DxeXPoOO2WlqGCJcGslTrJa76ycY/m6dcIjj
mQnQYQq6QPovRp5vIcuzJLZ9hTkOYzQErMGYSzouR09j24FZECnNQpSGAAJPLeNp
M8j4zsDjbX0YFckoX6QKq2x6PY0mUl4pJgC/4ZgO5e6MEqHtUC4ESX34R4rBGsuD
RHsud6ssG7nBjpPILzFpHhjwj69CRyVvc8cvll+J7MJSOHFuhcB213+6mU9MHp7v
Nc+1QUYOD71lICAPbLGH7DnOtt2MYvBXv/XnZGTpSZhSZG5sSL3oBAdFKrC8kRtn
2IHc109wzUtQOz7TgHVk9xcabhJ87AJaIzphGzr+EFVMEjv0b347Pqd45Ep1HWTv
4W0ns5J9/LaSK/5w01k+1VxxNImXe/lpykBz+JaL6+h63qsg2BnIINwXOIqz+AUz
B8Y/y3bwjVyXhzNWq+btif5KMOt6Aqv4hI/1o/blGxjJ/6Y8GlfV/lr4LGH6K4Hl
jfob08iiEcidgSaS+aNROyOhxYYlAU2PmV6wrFWIGxAWGAqcQ0XEMHYyZ7NBBtlj
hzGoDUjFh0LehhPcknFKdVL6F2nbaB5tXR8enYEHL0+KF0e03WAvvVoNPXGgMsUm
/nWTgTiq3QggYNlZsytRjl5iOKP+8OLExBe4n7v9VaujRWsrPLOv4Vu0zeBqLh6M
389EB5XLg4wBYv4wdhDFEFacC++cyVImybXC/0+ZGoBmId3TGSiwUu5vb2ju4MPi
1CBcsy1wHgHlF6vZMbFJVt9nV/qeh67NTQvlWtzQAMykYn+7QDx27Dx9cR3mbJNi
t9rulbg2GtD73SoPeiUxooV3kHkv5f3R3eSBCKKLMJFD9ELsFQXsxsyNNhL1IJRB
r6bi1NHUrx1NX2iLaYUkTvUWy/pVXl4HeUJmNRnMmGqMQlJ521rYLM70+gb69W4U
zdyU1h1NPh/Ln/AKfEkqJ67vwMN6Cdi37w9+LYH+WGv74RjzZKPVaV08jqCTyYly
tuJO+pH0VwKrXZY5JpirKmGyubp3rm0k8gkinQUVFagTzB2l2dlCYSESMfOIOKG+
xbra9m+GRfFBRzpmUr1R+dLf10+XKX3fjMYX386/BambXyTRkkREhzE9nSWBv85f
gUJXjz5eaDwBTYlbJXzWEXxdatFH8wZ+WruPa7lSWF1Wc19pIYm7XwoOAQd2W/9t
wvkKDZ0ToEu/3Iw+DQ3ERhqsO2C0UkhXLRCRVDNkRh6DwCLypnXrcc/hG8Um7QGs
hBJJ43JF+1uzaepDs1jeiK6UgvaPslZW7Yw7q58yN0/Pj+tEBPorJs7CmitB80Pv
iHXs+KQxog6yP6FthiZcPfuae//zuxwkdZ7Th2J8NxR8Q2gL+ouWHpFIWm1jmeli
9BrdEHodqLPqJeWvlwiudjOnUgzeMzZ3sBs1N6fu3FbMs53fSHeThQO1x8I3uFaJ
VZJPnuWOIZ1p58i+hobK32geDOU+X3EzO8Rij4kpyO/WBzen47OB+WmDw2ctWGlb
saZg98TAV9WKUiJGCm90Z8d8xzldPVGLLoA/B8KHwhxK/rl1v+4PXig4sKJnWidZ
mG1Oj8PCPEQXw9SlHTfChy3fkBNb8m67TAxtDNdUxZjSmlMDr52y+hOjdmqaZveq
CT4MxcdHRRqcP8X/v2cpYacO1TXpmxcmCN4CqaEXkl6IvqMUmoLp88X+axoLFcOw
BycWY1B/PCJXJYhjsDHKe3ynuDvyCPnDRMT10FGxFJxDQbieqcYHWmxEfum8Tu3k
h6Ysx+eLMCtmrL71m/ql6louCQwfsf9Bg1LuwlHot8GuKvoprehhbfys/2oQchHt
BUzQnYf1rZ2FsQhADNlgzQ40SmZw05tG4LH9lkJ1c0IQyMsw/7gwH6BPBdRAVHZ7
2nYh+l/5u2ZiwnJIZpoi31LS0HXoa+88m4vDL5iwJYHgfrwhLi5KuwsEdbEeQQ3k
XFhqRkz/Go6HGbOYA67S28NQxSK4N7dVq79AYy4i4gP70lwePcg6XTzkBIVLgvkE
hDttfqKrv+EFF0nWAFel0V4LQWFUOPD9VYPedQhwGMIqvkw/Xl4y9XXJwKrBrls3
FJOoU1JwpdVhSYid4hQGK+UlEtUA2V/lzSUiLxQKPLKQcyRUCJM1+YeY0LNKn0yv
RoKxOWhKUnpO+sMmV614ap5hO0/w7uqqohCUcwe5714PxBj3lNPtOYLUwMExALxg
p1xwgeE8ruwLioWryQ0FACTnO/XbP9vB/MZNrOHjK1fln2+4Frh5jAiauc45jC2+
hHLGucx71d0ss5W00RHVi4WbyHaAif/M/eUcXM44kKTfkQD78AEx178PAMJ8Lc9x
KGcjriy30lZulbC+UidYEuEJnPaL2T0To/kfq5BLOJr6Eh0LaYhKxEeWlEDZImHT
iESjdwNq81ktKkQ0UUWu8qb8bJBOWS2tVJchCY8/yClhT60eRnLu/ox4UtIri+mB
ogMojYIuvIE9PXPJyuw6kCdVAQlvR35Ad436Pf8LjdiAKxUMt9y0YExPJhvo9FV/
7LgadHJTgfcrhYoEGjMGw3eknc0bWNXsglNspvWAw9eCI0458AyjglZD3iOlJjb0
6y+3c/luhLAzxgeyA5IZMRnVCqaD9rn9jUabpM6qOaflXAZ/wXMXhykeABpHsKJ1
15j6ZTgHUM0cAlM50Np/aJfu75Dv/51H61KXOCfh4BZPb4JqHOhsZoqR1OTDqmOg
HUu/vcTVhv5UmMgIPAcumSLVULpb+Qk0fGN+jRiL+9/dN8jbvLm7+2ucfGCqI1c5
p3RxR0nKmNFixqn8lS0uIajtF1P8Asedn5f4kJopku4D7teVzykxMG6J68NY96Q0
Eam9Yyr+yV5bsd0dk7WzQieV/tn7BxQ3iTBD2LEMNUCvN0OA28nekPXLR5iUXGhl
DyIWklfjfIzqEq+uUcucWKCNVGrXdMOuq5e0Ml5FzpI3ExipUSrgaqT24IsgJFTR
hQXzcm9ZJO3Zk1DCdZFnn21E0Nf9yXOUevXHiVARJcl6J5xSxmmuRaqzkoeDx/V2
wSaWkW39RZAqfNJq4XCTnK9OTgGx+b2mqCVP2G4rwirvg+IPYFI0av5NzQnrgu0F
t+vIQRTv7eQFJcaMM78L95IWqIyUjQPfw3vz1eG5uB0nE552eeI5j0cnb9aYMsyT
c0ygG0IGi308neiGOJW8msdyGisjOwrgNbEYCTQMrEd8t9RQ5yi/eGgkZwqKGmHL
wbgFCPsVXibN0MIkmAqTYcrN3YzajGmtQ5bEC8jD4reoGwuw5QGX9bet4aTljNNt
hGamtgfK+WeuuCMETgQUfe590nZTGKCttsO6ldJcgXjYqP0oI5FF+KK8Sf5iuKTZ
t+6d+uFNZ7R+zUmSdr7IqcruaA4H322STIwS59lWK/mfP6YZ6uXzr4UXi/B194Ro
ywPLkLKgDSgYAAmqjc8lmbwkRxIylU225PvCbIdRPpo1GI+GCDMzn8PiskG98K0x
V7yzkuYWyw2+sjdBcmhqY6m502mlSnM2wQrj5dQV0a+AECxSUZ2BXG63dFB8c0cz
PWPQ0ZWuOdIiXqpWXxcOasNgs/Gk0WaGsH8VPAd5BC0dyTX/9aGJWddd3EPH0mur
7mmY5bmbdKgjsR9WpCMjXujCr0cXk57cP7PK9EV9O0OuFPa9TrOY3qDTazfKcMUr
G9oDvWtmo5RzGL/7ze/FsFityXVIuZpLtypT33WF7q8QY8gGmw+NoXbm1n3yiQ/H
uE06lTxnPUv7d29NJHf7DUoUEbXsrj6h6O1v5ehK5KD8ck4tYt+rjBtjayC3tFVp
hcdmWw3Ws7lyvd6PqZlQXZnpADOnbZX/7T3uSSeDrZr7+O+lX8xPJ3EJr34LlpUg
bFgAmumJABgQoIVlk4WK7ULX100rGjePllN6RvFT7QjgVxi071sjuSOht5DDiS+W
aRgksiqbYo5L3ZnqLQH8hQpiIqI4yl9aTwuCHXWcxKKQrP9dv6XqZZtvQjZhthLc
noLrQuxqk4L4UG7F4dBw3lMJ8HlCm5x6PhWpXYXx4gkD4I+OXuzuIqqCGBv2923l
+HuJnJV2d/RFiUEKGLCLYRJ3CyICk+byeNwhl2LWdStIVN84MnBpke2sNlLPBiTP
kuODbzL39truyRpf7QuLGkpLbAEDW/qK1aV89BnbeKyefHrxXSdx4eX9Z48VuddT
mKdyqoBJQHt9bEGsAfTOBDmiCGUUObuxemOIcDciCA4FzW+tftI4gRya0jHZufuf
lJK2JLFqEIBl2LmvGpCEIpNJHVWKAgscaNiIpXev5FxqLjfDUVYZdTSbfJo309+t
E43j6uk5td2dZMCQnGVlP50w8bdLeITVqdbPqII9fm8UDui0dNNF4EAFsktiGpXz
2iFUzJJ6GyJsrHMTRTYT0sVvKjRFy8Tmnt1fDutDnoxYF+rJ3xNKg/xW4/W0YvO3
l0AChleVYZX3/40aRV60rsm+hkNnn0JKqAlJ154ckOfR2GwnYmOwerVufO0cittB
i1BC41iOsGqr3EQ0Fa24KaD/9hCQnLo6Dxy3ZrzdlMSguqjgGbywkcmLP5W7nNVP
pPr9o/7950HSpVZbmFQJPBzxr0gQKWu9iEcUJkBVJxUxNG9vydh24m6v69sp82MY
lXmeM+SA250H+fuW6d6kpNpb4zupdmtYnTmAbe4+Qv48uTiB1Fk7ErZua3YKW1YM
31A77HSxXf70ViBqfJfGPMPBg73MUAEWDSeMfiPzmfITfgPqKW4aiwQ8Y/3XYOgv
taP7WOridHTkFEngHywtPEyEBTx+cZx45nwswnMQh5itRpbOwRCQb90kjus0I4Dj
a4c8B4twoVGuDHhKHc1y8QK1TiIEkwnVCO1Yyz7OjAhA3soCb8EWkbZxTAjQQXfd
IJHgYTm1VsI50qWQrAjJMKBY4yVt6orGtSXzJzbxvkcGB/siiaWHSOBYMTQRpyNr
it9tLrnFNbw2p/sa9WXg7ikXSxzLqBenB5v8m1YGcqKXxTCPOvua3P2SG54aCgwc
CedsIEJiyBb5XnTJ68op7ih5o0XR6Jcp5cAS69k1Gk8kWros5htjzfShUchQBD+D
59+6ql8xo1Ej5AzofbCeIFRjiq/RSYk2eGAtL5cVRGobeudo3a1YukMQ/lSasZxK
Wp1D/nTzs4YjBPRHR78u9izJxV8bJpxvdww/0wqSnyGtrhCcrq3ttMTrToKC5YTS
S06cfPGm0MG0/3ZFyIXniaHP8wljAZC1u88Med3RTLzd5QLjkxTyaDyW/q8vL8uS
nII0Wv/jymQWoAzaLSLSAKHtWDSLnlSlji/CTP31kLcdfm4BATXUUyAreAOd/S46
RP4XiQtK5g8ZQKxJCr/h5it0Aqn7cJBlCXPEqd+CZDKOfZeu3HubR4mdvtllyHSC
gZ3NKOh/Oe+1kcu+9ggN0NBXv6XhCuoAew+YCfpo9BIW13j/PovQCPuJkwqmSO1c
ZRNSc9YrUExdzZNpXzWefySIfrtgtmP8Nvywi/kbxE2+Fg52nD3f4b/cnpsR19tc
NL9RIW19CdE/P8qjMEUHQBX3UIPtDMWdoeROgQbOCjhT48NUSC/1AXWS9htDkAiZ
lKp0pflgiKEzh7xycYKou2OsOKVyQ1MQwVSRmCAN9WlSrvBu+uUTithFubfsMsqC
QStGkWrIeoosVcM7B/duHVE6GV0CY+34HsBcYnvjEOFgOxpHQCeSeg9vjATPIP1D
YHENmDmazsPbJxO+CYiEuFvZ9gU+4kaxC6p0OfcWeodfx4oRAVOr3w2Zb5IEL4TQ
JzvyBEqJNxdf0mWFOqg/9Om+NbxBAvNhentGXd46QKqT+1W5MZvle+UypDCCl43h
CoCNiBOrfbu3wTO8z6P1nf4oNZUWyICsMztJbyqJrFIy2+0fXC3kn8v41fh8DjVE
qUILWvz5EhMYxegb/9Q3NtujLkCFewUvJymJsWOgWMkyzltFYIEMOPjSMrsHFtCi
WYu8rL3sZpIyksDEgZJsYKzS2ffTCN+wv1NE4s9q3Vot1L0HOEsoV8F4vjemGDNx
TB773JnwlmY/g6N95T4WTkypq34Sb/XR7QXvQTFm9+YIFgnT5ihF9QkcCMfilt5d
e6XsxOQCuOYda0xi6YvOJHRKJmw3GkwO6r0zzLyJaDYr0JFSNPDyvt2fBFlFSKv3
HCYuHcK39c6j642uJ7d0SYslg/cMpsnUTzpdfWyqxGP1bkwb6Pyk/hhnj2lSa6Xw
NR2FziXO6pXWBNs9X79PZ+I3AD5G4XLBmkge51nn3V0H+cy4xkviBBqg7Hwzz4N1
7iIwzbd2LudFZiyUpMH3fTREU0a+jyoKltNwkcz2phxWGHrp80Vhf5u2zAcNi4zq
/h+/FImNUray22jWdxuQczjHE2pabGWU25rupFdCxyHhNncODdLDz4oZVRCploxy
NVzw3k+L8Jf7o6EvV8SH5DCaexmbRbbQnJf9yRVeX8+GHgB0gY6I5v7vsrkdcnF2
fPPMD7st18lcbjFylYS0wZDlLsKvFkLgJymvyPo32kKGfy3h96v85qVwdWZ86qnj
Oi87QQUhCBsgj/nQFpjYn3FXB0T4+NTJ7esA0CskbdU36miHS1rLdlCa9ZBDLSDY
FL58N6cPFSTPDPUz5AUN/Myj+YvI0zLNGWMiAxhvPhEskUQ9DoKnI7kyYvTKEnfo
EyxJnxn6G4hDN1zhuCA2NR2bmXmbo1jlsgiXFSAiTV2jqZe9Qhko9emjTdC8Hgsf
6BIdN9y27bcPOXyOU0LfgBLZYznIIc1u5m3DVKkjEcyiAXFa73vgB9KlMUTUkgfb
dAMmjRMYsAFLbFSz7L8iZN8QNDzGwINeBTaj03OlIPD0UbW/Crypw0I6FZiiS/hR
p05YRTi9FQaR4owHxMCsyK++KVRSesRNvG7Z8DcDBSazVKvlVPw7Z8eHUgMjskKj
Wu8lx7u3KwiB5pkbVeRgv4/T3H2cGpyiKHNynmTewBynURw2neE2SqKqBJZAxW75
AfHCbwse/udonqFsQjYNGWw1ys+zznrUUheyZKbtLLo5ptR/uBQ9Z4sl7Qbfp8XT
bSzIu7SAEn/CjvB6N9xqwG0d/bmxn1dKDAqsOcmkNelarYcw0BlIHLl9EQXrbjBS
EST2GJzmmvcCdTskR6nFRaf7rqZ878kfSVeV7Qfu4CqQJoNfiVvKWwDXQuMwPHCu
qeVi85yLjxOh5VErzE3cZRFw/llfxbssUirpHA6U1H7AKKy9Aafvm6HLFuj0dVBK
UF5Tq63FBda9X+sNpW2e/pjOopXInPyqON27R1iw7EPBI/dpNNLwQpdkbSzGhDU/
nN+SScgMxQqZvprkUuHaaNP075AXNArqG9koEHDHY43WfnCS5n5NgEDO3vMrETXA
4tt7joK1qjNq7vb7yUpyDyPH5HnFnbIJX4U89lHFopKjX9hJGCUgE0Xg0b0EeoqD
uV9nzVqeQsDoRyX2HFftHI9SKuS0ZgBG3ovDFYgwEbonHj1lfGnKSL+J6/jQqJOa
CFdM7UErSuefhyak0TyiMgcqZeE+2nV3euDtxXtPYEt4lKUN8JEGeLAmoW6kNo2Y
qnQIus2IRC7ftaf35TuCi4TMgt8ooVsrtwONdDd40SUhfmyKN5MpXM4/gIn9nhTG
r5UXE51iebowKnX++flaE123RL4H3pc39hWV/v++WbEw3Pxy9rhfdUb34daO812H
FCC+HjJ3bmkJqHiHEjnuzNGqFUn9B3B+XQOqm4GQNd89VmkKghXU1L5GrCLlURmH
qz6h/ZvEHd9fugpJnjCQB/8rhzdUtrGt54bbr4ugLzWVHyDqqHT4R63CuERWRYQB
ILoiu+QyAhEzyuTVHt3/k3vsKLmtJmp201sksrgFA+NvHpvQj98cEc4W5QZ9wotr
KedstLOcmLePFErga2KsoOvNa7k/lW1T000187lmuxlBw8nbRrdbbF+EE/nghQLD
CDsci1qAKzUixuYS1pWOsR+ut7ADZ0BAeDTkIht6ZPA/EyzE7xhyK1AFS2yFNtmR
Kmdwc6MLck/EyKzaay0AVjedWSzWF5vvMeHtmG4yJcNtMTcChyTyng29+mAsTzW7
0Lf/qE9JRJ5xpIU5QUlbTPwlveIjPVxOzBVVkkBY4U3oRFIYXalSHYXb/0SHHXsh
zWxVS/JEQC1NwQWCaXg26sRT1FG6AkHPYd2ZsGomGhLgu4qIF3XdnJD4V/qLzc49
WsqjfSo2Cry24Nc7EGuajuYIYGLcvn2P/y1+fq4dIFyOazoLdSw2GUBmJU1dRBOZ
L/6bF+2hbRuqo9ouWiFA/lZe6A3XDWqp26+gJjuKd9AZ49mZ7qF5tqiQ/eAsaoPZ
qNdZ9CCETiW58Rtt87aJJo+HeTaOFU7MSk7Mab6pBF7P7p2WX+V0t7ppQiodso7q
7JYio2yuLrqmj/5nRDuAeWc7ncf5p7DudOyYPlR2jFNBFwR6P7JpUAObBmw0kFCX
FUobRvh6NkZg41hLS6+ZQj9ZvjJGI3bOc30hFj0cc3UyyNwJHmHiOJvIDRlik7C4
ptYzNwmYRLvNzuKAxY04twT/Q92YaK+XEFoGo9zqKANX4X/1rCCR9VtmZy4VWJJ/
4frsqJ0eBz6lX0PqCokYv7+ByRL/xAvz3zzJpgPWgdX61ME1iv2IT8MD7ex8Lf72
jzAxVUvmxkj7ETA9hk4iJ1K9110rrNKK67nRJGMuIIfAqekzAvqKMnZTun17Zfbc
XV7LBImK2gm5D2VqFn4SWaVPRnOqyTaFjzpNjXwJBwsiUKLpI45oODALH6MtItJs
90fp7iS90JvFtgb8kz8r0sfy4B3in2E6S0YL8gBfeWRFSU/Q42ZkYlvuC7sib9Ve
SB4+8J7/+eK2X3IQyG67rC4fzMlzd2+s/D+kkgMqjfLWE3w3QZBs111v+B6swXnR
gQRZaAzmSjhfu+LpItjqIshkN8e6YDltGZ82CWqtS+fzpwkk0W4E6CyzrreBaFIX
tP/vs27tANA3qJyBopxUYz8TjH+KWxIrPgF3wHC0GDBEFc6QZhAAwJIBam80dGsE
qPFFlHNMalQCBDSZgxvMRTuYXg4lKb+cMMqgzpqppQMGDSp5njlE8pbLAiC7fxiu
25DTfiJVcSkLfyoArWe5NODKlFVdF0djtRsSXyMvaIC9iV5fNUK0Zsv69xHKuBuk
dWH8RmXQNcjekH0s/V/lKRMipgLiYGWdpDslWuRxId+41HWU7oc15k6xTOD0MLqd
mQXfLuZh3+ceMfKO+/ewNYXS0QFC1VMEE/Dmsrg2GFfw9jEMJTUlUHjpZhD6pGUt
52rhVcJZ1F5iLfXYDih6mTsfXHyLwN1vuAtiyLThlzcCH/PbtKmUTxmuCy8AKdpA
4B9rptk4Vq/hA/pB2Br7WkMS0zbn3uZJqNs6qAJzS4zugfyz/n0m/hglPtiBitv6
bo9CZEu9+JudFZccOwgJUFjAIB4xOU2lMQUpyu5Q/1YPy4oUQ7abi+TdHNtFxbt4
wEQaWqzkFs49oD+bxRUHBN2EDZ/X/XCYHCItBxg3G5cRt3XFJUNagTIbKyfJuK5b
cXi7IMi1O1ge/Sn51ugNXrfQSR0PUVJFG7Z/Q72zOsxC75Y/Em5qM/+oahjSTX4S
kCjX2kk41/Yw6NNnFlh0D4nsSv3HlOEKy0nB18xC6r7B+Cpea3gKM31xqr8mhURF
/RcEhgJMwCRApy7d88Vt81uALz6PASEXgONdZyIIJvABpmtEtVr9sZJ8+EDvbpWt
DFKjPCD1AB5DJwkAjJ3ziLceS2QEDuh7Col4LvsOgcaBjkVjIKeUZwXGuCX6DHsI
k3AYvy4D2UbRY1OWyu+Vk/bQJN7MWE+OsaFDkIK+hn/sEa9OxTIgnJUElnrnlPs2
lcWNbe2yKoMaIVzFiiYaoaBN4/WzutRY0HOnr4sY4Gt3x4Ugwg0NfEaXzZPhDLEH
wJiY9A0VQeIb5oCtGllJYeC12Xy7690zjGW3lNTzgTOck2NAC5un/mDPdKMGVEV4
uiLoHAR0BY0M+MDb13u791EPGb8jHTtZsqzcS2fEA5zAJC2fSAxjp/WUXX+FFI0C
zqVqfqlTx3scX0fUKKGy6h8x6/N8didBUCr79FVsuXz0bmsazUcLqphZ6dDp7l7A
EDZeYILuGnVszJ/DOT1cpGtvaJegk+vUQeNztYkTqs1GilNEE233FE/Xp+dxX8d8
20gpbhCXC70abB2aFw1dstmc6YDHI11KTk5rEkdTqgB8eHrx1rJS0f8vtiILgQTm
9Zseuv40oD2nUs0ybfqcZU1/UmhkFTRe3nTLz8IZ7/jnMxpvOgYe2cZ+nzruwZwx
xi4jtg70ZB9IANCRbgxOiEPV7KSkZWtZPpNjuCLPz7wEbcsYZYq7JopiGeVbVwjV
KK6Ys+haM1UG86Cqeb09h8A+bbxun8h96puMSKiyDJqfBHqrDR+GDg0GBq74k1TJ
RrAb7AUdYwk880O+91FndQDvpkGPhz9HY6MHzIa2vOIZ4KWqqn/KmJKRezvorNCp
CbYB7cEBqkjeqMg9+o+HLzgOqTV+++lvP6XtwKOO/kesdyIFx/hiiu9jthhqHsMK
a8PEEdyLDReUgsRcxD6uhIbYFYvrYOCVE84etk1S3spkv0wl1FAQNaS7xA97de+N
H+/zn2SxT4eeFQHwiHKFL6wWI0JYQh2kwX2RSdScE9ME7lSLEwGKoLnMjAGfVMz3
yem47+OAKGczewlsc4xnKqtL4LVFom1PwIOB+cXq058N2Ela5ucMXhTU6ZrzsM85
xteW//0szXWzB669Zl1ZA7HycnrDa9xtjKI2rPYh8/381hZ3fi6YxlAnNweaeszW
uYDBYVVmB6P3o/2YsSwF+glCS17AXtu9cND7Hr7/0COs9uylK/urTaMFExjW917S
mtV0lUrc037pPztBJKJ8NZqkjQ+bAg5wlrNU3RSi6fYIQcWDwEJJHdngQ3pbqyjK
KJx0ZKMVqFuSFt5xuCNmr33IDVgn9dujvtlw6S11vhWxqpWq6On+oQR7TDr0E+Ed
TggTG57zpEV8DyAvc34bGfffEbDWIq0A6XxKRODDLLYp2dF+Xclt9l8qu3VgHFvI
o+qhpnahnBJD7t+juCj5PPz5SdgxpwXuFTQtAFu/JcKvGXSsYF+waTPKo+by/OCG
6pwhs85fJaSnPymj3+Th2ozyyeAhwoxQer903/lXCkDrBlhSkSpuYVew5jSTxgX4
0lDWP2+BYUjCU78mEFn/4YCrDvA6atL84LY7zokktlYZoy9pC0QysPDVGgYgZ1TY
LX+9xHzwCr4H2IAOCF+F+Fa2X6MaFg/iwO/FJEvLwqzv8q0t+vyzcxy3ILikMW+N
fJ25ebRBVJBJc5bal9LOROOYkBVnYbdDnxc+knZlxUhSNy6WesBTLcTAy98bXVSR
ov+5Y6oSk7a3Olzk5jhoh156A+s1R3rkOp1OCDHZgF9GkRXzlJ658JWzxD/Yv87c
Tzu9uZQRw4W2K+Arsxiv5hDu9Lcb+Wbk0IuLu+8zdTh2Q8KJ6frDxhuGF1okJ+Gj
4MAi4K57LyHMQ0rYhxMxWusVh9OCOJpQGnnxSQkBFWsPizZrf4nrkRJvf7evoU+7
XtUtJOn72is/L58XzPXgBClVQUtj3ieD94sTt5UKUM8TxSAwfEdqTv3Ztkhytw+f
fvWC9eI51ychpOp83zOGmXI/JngjEqn02cTfcYydY6fIwzWxIdZgZS1VtOKmkeTt
+MRWsSCS/ub78BUS3Fo3wNJeJBmGnfzC2Lxg8ddUCKI6wMNNJna7EUTI+z3MHEPj
ImRKS2nli6AdU/DynkNzrG5Krm5s32dqNCRTS51DDnyrrVazf69VXsHBlQ+JhEHf
XamcJ0XOZZBOihWkR11HsVYCsjMGNH85dYu/GStPH+1yTo6dyjlcshUvnuvLF9iC
KqdmQCBRjmRtyhvFLf+G4ta45Bft6yk0bCdYv1b5n+08FcfyP7wjgRFH1f6RL0nl
jJNHlwmSS9TkDxHF/enmgrFLltEt6tNVWc7jGbjI0MIuyGJA4URi29mG7ISlyb9O
Zp6aKzdUkxs9i+Z8h7u9mw9yQtaP73jGXVNn+4mp3fy7HSpaPiqJIkg79V88d/gp
LFaLPYUqvN5iduHhHJpU6CxOZRUPtR78N23hQiPBLbvCAeHU6G3AHAmb6ySNRp01
fWg3Tq3svIFlWeXm42FxLDfT0Gw4dt1nWnMZtOFmr4B7NySo4G3lpGr8eVFCXb1p
hjKnIkPRM0RgV0yRS9TIT2Z3fhn2dBiLvRow1IKIrKgR9dgkRIf6e06evSyNe2cT
Ii2xTKTUvQKoRsB3uKwLfQOXa2r7yBoxE4wEqBwWZd1neuu4/lfQyug7VWGD086a
vx30Dtwtd2RxzbQ7+CdKOYfnJHXbBaoDuWbnpapgoM2do/ncGtvSfHTyXpurzjsE
reHjLiWpTMzJjlXMzc8wu3VXTunlRuNh9O6ZbQpMHyTUM6cniUTk8+gA1WocQF6V
C1N2RrJXpIDOjlFtlQnXx3Tsp3830KSDRI6aqwUZunoiAvVga2IonHtIWVetqqT6
xo4617jfqet9fgqvJapZ8npakZwF/odMBuPtYdRukSgzr91EOGK+8MHx1LENm95j
L/d83BYYYUlrWi7rbC1SxJrQIhRlnoMmU5jrpalx6xukZ2yeKb13MXStRyX6NDLw
cV0qkqmXsA00ai9284ye206jSw3f2opLepDgU5D7dAugVsexIHf0wam6xvKrjRBv
/X+50U2gI5YkhOnJk+4FBB6/pu8+vFSUXVPBfx5c2380zPe7MREv3xfkAb+11IjC
t+g+SIIHjZDs21oZLrBA+vlWgVmMLNdsqnKur17xi1VdN/DN0rDlvvSAGccdZ8Ks
1wjFXEMenPARPZeBs9ea/qGL8fmSYqH8ECM5+T9HJKvmuRn9mATQKUj2ZkTLTsFj
ICKrz4fXuUkaLV8elYvwOIas/gnG3fpewxflCJ2O1kGGPlm7sq6YukfGSWWWu12W
XQEq4lSW+DIZ8+8QAb6+9idw6arvHECzoqYjDbqb9k5PYbvFIntBM5Q3/g9eI+jQ
GifB84Iflo8x0GEzcRNeYPqzzpTG2VmeMBVfEbRXrPcIoifzseVlHcaZmHwpOpgt
oSWNH2FAgA5OBRTIOXjjeSH0Kgp4ZTRZM0/5CpH7cr8M/cyE+L4/5uHiqhTAfxco
7w5z50mHX6K7JwqHmrTo5LY1b1yi5odhYeODlW7GGGlb8pLO1Yn0g9eFotkJFZ20
ZuI/honpnSOZOS92R0Xvq6H3gsbalzVYu2CoXFzdglF7h3R96rvw3QwseZH2FTCg
Fsn/TMXPdUkA7KBx3n6mgm/H4YwB1S4fR5GqQ8ngMUluQ6AgohX2g00kRs8LKo9L
AF4id+l7aVLKvATvbZi629S7v/7vAuEnD2rmLSDJpdlf4Cclahweq371V67VFRD0
OZnl2MAsAhFKqOD2UYfXBCslwOm154w82arEBc6PHa3qN4oNDlt7wWmrm6Ia8j8B
DIgZxqdnjE5au6xq/AHov9PZx+q+k8SmCf2r4MjChDVLo5KJR3JKop8fcAnlDgkE
wHXU0qYJ9PZAGduriUba7hN1luedif1fyBuUdMHlKXFFduKwHnZYePCRPbSwybDx
EFJ53EoGwr0H5xrEvJ32ahq79zIpceWdrD+h28IhW0d/AvsaPtrqyXahXIXlkmmb
ThjEkvWVNBNqna2k2doDt7tjMMXcuJvQh8RRox5kG1gva7qZYhzm8pdzoNKhms1l
EWBBtMQWU1hDBC4n7Sq4ZPoDc+pbISNtLxWh1DA2lEMGluId7DDRyqQH9CwdvKsW
VaYWaOaxACGSdaFeeCeVBlqV+E7Uu83c17ELwUoxvYg0EDJI38PUKNd9TSuo2sHi
dWDhbF0v5NdnaOjMyFagKo3jamzNAj6kzqclkYeM0gUs0f82win5CRdvx+t1Yrg3
Rwteodf3w7CHA9ktd+J5JYMOnGi1bBSjmLbXsd9/fI0rCWdSN77tlumDuCTwietP
6YbMGWBY3dDcJ9Ltc5xD5pnFmYa0u24mXUwRtvKG77x5crqS+wl0e5OwuOSeIVSk
bLLbC31fClROv2wV+nV1vUySm/HlFEHhxz3j58HdOvLpWlHy8XWuJ+ed5QebISoC
jXzOhfpH4ipbYSmqpP8c6UVS7ZWX+CK7z9IjfFujgw8X0NaN0nnbup2gMJKg11QS
XNVRaA/4X4X3d9TnFuf12VQRyZ5SAry9fhV8t0L6r9k11hpK40qTXqmc5OYJdwZ/
sb1WbE43Wk9aQYERX2o5SyMZ+N7nSug2eNdRfrVeiqG12PJp1qbYcYarb/L0OjNd
JjGp2294Q3yekJVhTuqoODCRR+JrRft8+dpRL2hd3SKuoP1ctvNw2Kmo0RiZ7m+p
Qv8YqzqD0899N/NbZiXgiKhpNPj+KNQzct0IECmY9IeFH6r86dNw5ikPyJHYaNDu
6neGg/c48QX3RDytuz5zPtgBQf7gI1jeOwtTV5Y48FP98pmlTU63pt5PrVYDk0eF
9IhSk4/r5uRJ+LNxh3/Pl58dHsocbDVxHx6cnqcjcKuXLvZ72PoI3h85tfqHgpaJ
VrlK9FwjOk0UBU9L+43hVQpg2NOMv6vK1Qnr7flAaiv9mSJAe7JaFvoWDSlAWY8A
Vv7XdjD09vltzNUW5hYPCDYDzRSDG/lhq4N/IRqsMvk0TY7s+SS/ljgATTkzPSn2
JdXSYJdCx0JrLiu4TB8G5FKUcVXx7UiUGIz/s9/S+3OgjnpyouC8c3jmUXJC1/Dc
U5zM8IqyTkZYVRRF3wXEyE0QnkqbhDKi+vmL/erOhnGqxJ5fl+xL+0ZqiQxLml12
bTD3b/wKMR0XBgf8vq1RcSE7AurmHeV8+HgxkoYUt3PtjEJ0wsGDymf7Tq25MXHD
dO4g4bkaTOLULhrKwWoKpytL3KwBH7vcDkrHXYEH1WtxgQJ0MJ+nPUu/obWykNZ1
A/HqTXgv6m6gUy1fH0PAfuHzke+Ey/P6YQ5yR4DBmjDFenY9cR8Jy191bVG7HXMg
Qs4xSHIZqCNPSItWK3b8hyCHMt80WavA9VtDqRQeBX8oZ5uLyFZB7TJbVAkJC1rS
n2wePEDIoLLWKFWFtzJUNr11Ifu5hqGwOvEOd2wWGo4e8+pJDMGOf0DMRzJPeuOc
aG/1EKNLDJdxw2pQ95jAOPFp0w/32Bxb4Udu6zEjyW+9hDVQuhqH0/t2JM429316
M6OrujzM/Xe5/pHS+/Q68HJk2haMgSIIVNIFm1z0It/hLTKNO7yuHisPVYeDst86
Pl4bZj3EAGoIbKI9NiJ18yf2k1SFKUtNH0EWlfjyZPljsXaXOHOQUcFPME9HPGfY
h1xiyBziB1zBSOe2YvP6vyo84Xpo+5oBBnikoNE2UsNEDZVkzI+2VYpUvyZxvPOy
L43+lZVJQqnNnrxAFoIi8S1CM1CIhyzN6aybgoeTse0ObahwWDk1bwalot2BX5oU
io9UKkBvVtE2LLb0Upp2YqzCFGEDh/IVBXHL3bjb12jVY4paqek0R9k265zpK4AS
r7rYcUoZ812e8InMl268AqWw0nF6YdJZa49n4hTBQsI48B0UDZOnspY3mYU+o81s
pOUZgEu2hcmcrzYIwOzmZElkpzGcwCLtv5+IEI7LiPfH1yKBIHpy4iz2wjKIZInJ
7Z8P0krEOEdgRUl9UmKkua5sMbdiOcVnJkEKJpVcXEwdjKZ0+Yw1javQUNvfQitP
eFmxWn0kWDQUeQuSjhlPEy5ED3k30tWy7jhHZfhBihchTLOqy7eEYAg7LUH/PD5b
KueODYJhfUDo7kngOJnT4KJvCc3CHjDYICgeMCY5Ntkn85phpidlQzyqIe9fqXe9
Bkz9kSU5Qwi/sGXJW0Lv6D6oWzzuMbXsljtui2ICvDrmNt0nfalNhMEJPIe6SSQC
5irVb/R6orgSVKYPGJ9LdKerZtew9Hb6uSZhjHzHNjTAfoBZivGvju01aFu46Nr1
p6pzIaf9x7YM4mlLfinP4QrVuV8OQXz69Hqt06wRGZ0EYL0WGtkXJBX5GuR71mc6
pTWG+UDV3LQPS5OckvP9fPlMpM8kqmTnii39OTCiqkv+/CRWoDS5d+iNXzg7XMuS
3dnxrBUdxHrggaYDHx6e6luPEGoYE/2VqKGWb7QT8Nu6P2Cc93vc4MfVdFMQ+kng
C8m14vTJ4rWqh0vMoZUQsFhQc125in4xHlU+XGIzsk8/GvbAHs3I8trKMW0cCxo8
Z4AvlqW3wWsPf3NyJTvicGe0o4tu+hKgkG9whZmET4kXqziVzPNBRjN2t3rL/IT6
4JOqCyMrry1HwclPoZPqW0o3SLJN54JmMKyvjdqUGldSjOH58mi0xvm9p9uT4OT3
CcPJQCuDNjytKTH3tPwcUuJn/1TYJ6N3B4Vp0xf2OaTOJgl3YAAERpINCfmsv3rr
VVLaZDeXxWDMimPZo6QCMuajZwrgQObMLc7zZ9dQU9MDeAd0zhq2NHF51iY7vida
9XWTlRy1aJ4hUkZ54aH7Nv95p0NuN1UHEuCIpvxnxA7jmNFhDWNqEJuDryKhkoRw
fwVhW+rzJYNyLFXaLups4v+rlwaQMDRS2TyKBaLVr0M6vL1TAgjri0BVcc6nmn4B
qnvV4nCsjuz00dQXiIQg5Azqw2fHWJaoVW9W7gK4ml9BVtT5GSa3C3xlkqgWT21B
BtuXxDZ/QZ2auMbGEuSeia5U6kBuG+gpSTOgltQVtESJY0h8r4BNJzAdwcKINrZA
9fIESaiZEFBVsR8SwWEFocTCqepjXb5y9DjYqDferxiIyK/+vViHrDF3VSY6vyNP
IaExrdXC7y1x8EeeFF1K2f3IRyO2OLfVETNhTkYgw7xAH1VT571DiniqajAIkpl8
Rt39tmr1Wq0QcynB7UP2s7xW6Jp6fY5+yEoDhg8qHAhjf5qQsDF6qPp6ll5Y1D0q
ulXDgb5fUPvQQ3C0o6fxQnoox9nJ4krCnL/wBSqOHIpm5uBssWBh7LoLZcQsdOkW
FEJgx25UWMQ9/lw6t9bwEWP79HsO7LRffVVayXbQlhReqHFeh+4VMwNzcHES52eA
Clq+Q2Yn1Zhway3/rvci6PQ/Ju2/KJcvbOE6LLKjtdIFTQ1Vho4l7/0P8oE52dIb
so83Z5FeIWJ/HVn4Eu+QIW682Pf2mrvWZ7DiH4iHkcmEys9eOqmST3W3bs/qoWVs
mGRt7Fzs5fxwV3mgIX+o9NtXrT8kDPoDFIFJvjJhs4pux4cA0qLp15PmI1jAoE+e
2e4GDroDV7jK1DEAsgr14AXFqvjbyWh2/7yFKb2sfFTGvG9pBksCKgGd46507jlH
s98zj4mFQpefnqiijA10tfsnCoN40ve26g27rszJNziA5bei2r+33lzBgh7+5OwK
hYEsWP7od0KhirK6u3riN2tfWh+DRwyxdYGKYzCRlMUqBL6jLUKOZYSbN9LQbZpj
52a0CORG4Zf7o1b1cm98O4U1ZExVTMNqYf1kRfpLDyrOY2+RTxgSV03ibLPwhNRg
NOGlw46EQZiA9tvM4GLlnBpHGT0d+O68AJyCEoN9Djwo6LlHcoggSSZ4oSLKI6TH
HdNmje5QtyBC1Livw+wGtITkQHbRC6QOTz183uIMjW2QceXRTLoa9VbgJkHXhsZF
sYf+Blz9mjyCE/AEvMZnIRMilpZ8P19Q9Fa9xTyvXzqIbglg4b+0yxxEU8gxcKiL
csTdS1eudR/ypt+dGXFQxGb3GjCZchyAYyGAsAfRsJEm8SGUrIvIpFGWngRlw1uH
hfJ2vGRE5Zec83snsQDfF9vC0iB+pZmID4xiHm3YSfm9IQaaTtCXzV3BHiNdQiDD
Oh+3kbhlVyXfRzhKe+mKN171RhTqTdRyONgvrOXAFZWHteRenxCI3JL5ETfo1d13
OKvJwwcFfOGBi2tkpGaIgf+qOx4lLH1mDN4RyIBdRIF/lwmaI4zeD816pdDewLHU
Jfu9CP0j0b7k9gHAD88XzVwUfuW1V7jLZsAHlzeqza/LdncS36noyire69Vxx65A
TPeevIiTKn5lBHriM2uaH24CwSBZ4oQ98d53C+55yFRkIAP94np6tv/zXLVFLjZF
qXDAdgRNyqbdzYdNY2bpFM0IOvVBLX68Af6gWNQwDOL/zNRjIMADPFAZuz65LZH5
SmyNEz7tJ5RDKVZgw7wdPgHeTFcfP1YBnAY8ACqKVU3Aq4yVPgQoIv5z6WfBasxC
5rp0Tg9BN1gE5Oi/P51MA3N0b2nuYAYpgSDJwqbq0WseHdH/Z0Xv2P8UzxDw8KXo
fkUaeJZQqnzOHm+Wsaz+fHNAPwUdl91m4BJ4/lhAesPu1fs6J+pxw8o//el1OEcj
1EjlYD+SEJ+uax2z3bTlZ8x9VZ2Pn4bS5/kOEgiE4YmSlZMSly2CY2gtlnjDQX1y
j18IeL4vNPOaqWal2ZjA4YV2VRXfaamQALPEp3PA9QDKLSjJht2agGjekcC1glCN
3WN7es8WAF5yCxeTVxUMnXHfzGLT+79JKQdFJxRtHYvmi+CgWYgvEuM99BdlaIkj
yA9TV2X5Y/fokzC1dTWMWWBw9+fdw0+9w5+IBnR/G4bmQueMsWQI4ZalQLC7gFNU
sYZ6z7BGUxl/Lq7HxbxlGOkeSB3v4AgRnBv4NF0f/RZOqDrcmwoiAebOmQcQlcK0
6GxVB7jBfqWHg7rPO4I/OBU/l1BgqIiJCZzBrEnTX2qcrIXpBCxpt+fOKDLG3JI9
jt8ndvEKrsFHNgjasDqKtNBeoBPZkO7HvFNdVeAdI5/soJw3XUWutCkk2bKLcgVp
ScL4faK+h3b0mkRgzh5XHPhPxYlTW5XVpzXna/gD6wTr0/ifrLGdvCVH6wF7XIon
upQLxL79/7mRQgYn9o3FiXYZXKDu5ho3U+WHn8TOEl17LXTwFQZgTvvTXQ8n6AH/
jHSwkax+GCw/t/6Ts5pNyilzA+EhgHoQYJJIfWodjneTP8VmNk8h5tZ2u9aQStJM
1ryWiwUIHwUVP+VeadS62WwCE/9ub5tV6jkcUaD1KnRK68PT4yic7P5FdEqcqBo+
972Djp6R3CsOyPfELF/PB75RUtcvjizEXX1zARtPpDmEn+Dyv7fKHW8ki7F9Hide
pV2cNkk0IYEfCUOGNfEwCany32l57pW5OJTBXwIhum/JXCjp3qmkzDBpaHQZiqj/
iQTYzVwEtNOyNhzrvuzUXFHYeLp6REPHShGRihY7knHkEHXul8+e1v4AGYuAApn+
xkyiYHwxc5vNf9Ve9VD2Vt2T0lBvGf9uxVMKwbsmqURG9QWh27cvCPjOJoGbfoJT
xa6CAZJfUFfEDREp2bmdAqnOMMJVs4EmJgUlsvbKDKM0OYbZv9Ary8eFC2L+rlnt
PMsjBwJNZdo1LvkDxSn8EttiFpCYtLfTr57EbyZqoYFmfWkQ5V0BRLUh2KE39SfU
tSwrYCPqNJE1QjB6znDQRnqbsBOCjUHJkjZJrH9ydmH++xy+nhonlRk7rlgkBj90
ZjV6l2SKvDtyAGnHqHqYK7EvGzhUIGwp9OLtk574x/dQRuMBBfze8yrcq7eY3Iba
z4+zH88u4ajrFRWN2X5D2Bcg1fnDQQv55BYzKYFVAXZ0tae1Gx8WTd2gK3UWdTEx
o0cjemGNE3nlHVL3KMwyurxtWpTSoP7zg+R2Wn1P7gsUlQe1ZD+ECZ0Mc9K0weRn
Z/X4wz0SAexS1gJgAi972Rmc2SFEwzILty4A0DRipqKTTGWC6FxS4a1NQChkC9rx
64xkp0j14IwgRJWl2LnY9T7NhGKOaHMSy1Oisv8k8NQPKjPy9smEAhVGMJ8DezAC
d+KRKHb/Efk99Fcg07zoy7jTCCcWs04UTLVYJJTi0wExcVGEsdt68gFSc6t4rZG4
8nhF5RlnjKMGH2X6cvhsy5Nzj6WMIteoZVc7b/GkDf6pD2jrYeXAPp+omhTe82od
3rOOBOibsdRpKigE33jD2EU2mlNN4OT88tfWYoUQZBA8u78kEImoSIq7PmWpr/aI
B4EkdXyNLfBzW+7X9julo5C8N+9Y+MWWRPk65Q8g2x/dx8TY6ZuZ/o8J0JBo3r37
QqGY1emDsGfxL4KH6s/gc7DrZ6sMZkBLKDVlJS68h4bT7vUcUzt2hUra88z0Fo0m
UVqXLfV3FmXauJ0OHxsVUc10sh8u5G5PlxWO7jawiyfPl7acXNLVC2c+0x87IOef
1aUo6Pu0rQItDG7ZGJsfBFwJgrE2cz91Z3eY4HZoNEGbbvVJiCNevwFmg1VA4Tom
YEaP6iLe4zXToFVtSZJqdacJ6o9XSHI/C+YzpGjwD+vrrGeaYAf2Hn2tI2yM9zAG
qCnKRTzpTacUoWf69VpTZdGW78CBl7FrjZLMr5xc9DkmDUSUzbt6SK5fQhnllnrF
7BVSM7I5g5J6bbFqTO5E/DIq1knKrfprajwvYKwGnLCg+zW3XcXVZzXJp5r904o3
WalCrarA/V91QixjbqpY3/t4cIuQaM828bZg65I5hXxhxodPBH3SB/B1HQfPPB38
m4oAEEYjjgjwTKlnjgih2RaPcG2cCvaNgH12dXxBAfCpjJ+EJ2ev/MZ+VchZ7YHi
sFsD0y/yCwJbhgDBS2aH0p/FOlXKaG7pTdj3u7xkKeBVIxTWgbF4lxHe7qHhtDxQ
Qh1qirUSTnA9EpmWiea3rsZZY89ukI7l8a2R0aaInmQM1ht6XDnCpwLTsfVYaQz7
YlXwu7EHcUNEwDTLstgQNAsaEWj1sqY9907XFHTmcGGGG2YzxVNA7pFE3XTm7b0L
DMwgmsLMAJ0lGSx5m9bcql56yL5NWy/0is+6y+5gj31KO4Pr85sU4ksAizDCTUBF
JH5J4dpzRglH7Fuyoa/Sso7+Ur94SEescmkQkHR6n/UIGywoXIDCBUld3YtYyUoo
8rmaxnXZ1CgOgadigo6sJ1TwpxV6eTs84+A9Hmq/e5zLhZz/TQyzENAMq7GUIQMb
KDOgLoQoXU5tlxCvlqK6Uvq+lNYuFQGPzw0SCUriidmZiEoOYRcAiY8hYjK45dH+
HQQn73unRzM5G9fpxlAxRzkwJxaFgzNZ0xkuEPXS9kAcSfFk+nPpABoqbHPcWMlu
Yu7+41kjlaS9qYotj4tjhTPVr8H4ItC3I+I2u0ktCnqRMzds6F1+iTnN17IOF9H4
i8rMPz3ZbQvzoh/2gbmeAiLOcZPVi2sr6jFspNzjcsVnmtLkuNhi2tTus1VcjQaH
VFQQCt4KmrTDOiWUCV00wDDeqmQnw7wTr25jzDkE5ikbF1B1qpnBOzq9IxjFv+G1
P9+pg7oLWQvD8MGgkMNN220WHDZfyD2N8ikqT359Wr/vVZzXwlY5kfogir9HR74x
KjMjtZhBLuCCxsl5xUVAQdwvhxrAd3/Vj6xHvBzTiBtEK3EruUHlWmWw31R33jUj
3UFEvwqt0sO/xHYnom33Y/SNClCbKbzxvB76GCovhcXnj5O4CdnQJL8YH+ZNzLw0
geEtNoHREvLULAWQ4UDCNsq28o1Z4Dj2rS3QNDU3iiQGMV77dFkBP/1FdE3sqLQ+
d/PXV1ZAw8daQxQxuHGEKQ5AUinCth4yOpfyDjeG7r0Y6ZSgg2J8mEUfJBlbTnHc
/5RwY6wzt8el3IqEoERSIU7RwqRaAgSGR4ZXzt+oqtuLZy1QCG1jaoYwpPT0wcZj
fOs4Gun7dQW7hyy3+xbopmqK91G3wm6Gv72V+HmH6HcYS377yvXzM5S4cRzOeSoT
z3wOeu/ft8z6Q/POM7p/VHeZdYV93BklGBRpVRFmTe1kcemxYNWhODU+doofPEV4
vHhvSQSbKt53PraIKyvESWAZf9k0BnUz5UJetwR6F034L+x7IwLL5bpcQbXnGfst
xZbrK47NaqrxqaZaA0XvkgAHAoWTBsKm/geISXCH1gxSJC2yvjQpygBjmDZDnSGW
E+vi8ERmaFR4keBzWEkXh+AUrVb75MXFGINxUvz30tkIjsUuzJrFssLDlHjP43ki
4lb6d0E/BoRVimplWAZn7+nErOeijB/FCfN/18TElMk5R5tHj0ZIRV9VyjOwKtzP
KTgQV4/EYje+BQjClojhpQjlFmkoyg34FSbxjVkEUK6KJME7eRuIJWLtdRzF4GlL
J1QWvJGQ8Lt8cOR1cKu0jpWQ4LrByU6EBTn2iB0ohWcstTIIGaI6rGnLPWV3ALps
PWppZGtRWC/02RBvyo/ghCzH6RDZ4XZuGVH6Nu5WaoqI9tIpwHA5YSDOfhcbsoM7
H/LepT5vqEspXg4zFsUs/nWbe425P8tARHDQCi1RJ0p0r4S/J2gdwqw+/pY36zPR
fCpztJwSO21L7C5I66AZnU1KlPjaNgM5NvAiAXHbMTIXEo5Bpb4Wuyw5VCY1l2+0
j/FjbIIozhY26q7VYJUCQbrGQNcxw8pSTSx9+mhnDohMNnrrHYOm/GjU6SzEIiMk
aA44Ow0obntFcfCVfDkorOGMlqQ1a6Xeutc0aE3wJ9hUylgV9cKp7BOPEJ4XXYY+
1cXeHzHmIQiPoQPYs+iW6hj7OjQaKG6BEJv3I0B7Vpj69LdS8m3I4x4XwuO/C72D
rB82MCT0J/WwEq7Xf+qypBD2ufBziygGq1XmBgxVhPkiLfo4WuRIZkJtOQHMV8Yn
Of68FDouF/F20JQZ3hRAdIYOilgzE3PSBZq4LH+rD61c8/fOE6CN212yWqWIiE3Y
NveWD5vNfywLeyVVe3srk+8ht2uQ6GOYZP9Q/stuBOwCxXEVn6ar52cCG6kOWtV+
57a/rwQ+XX8O1i30GOlG51xcrujN3ZQAd61SP4Fyk8ASgm+k3WwMb+eUrazuispe
7z3R9PludoAJWhzbR3+yMFN3TwgViuCtxtfM/Dn5lOLEEdDTfwZ6fOInt3rRoc7G
4zvJqytZiYp18iU/Nl79ALR52NK+VAZz8PDocCMmIO0xC0A3PdQ4NIrVodPJiTbC
GmcJBamZqGI+k0FeikkO4W77QpMmtw1knlgLSo446VAj63AvArP/1qxPurwOX6VG
/URzHsxfhp5C8AWcJTeMjdEPek0UsqazLGynN3t8vnFktVYz1zD5JpsABEXb09mN
fW5xLROiB9cZQsmiF2sbqsnQeo7CvEkcPVpH+Z5It5Wj2ByGueiT67BMCfFn7JIO
ynOi7r9lCi3je0qUPVTmPjSB2X1u2RhKSex4xcROlANAQQsu24E4t7RxPWXXjd3X
7OIyK3zYGYEzO1VcuP8aATtyjk7XeyIvVvy7PLp5DwCHJF0WZBkFbJjpEj56iFgV
FgW0XmipbOBlUxUD26pg70XIlxre72I4ZRsIllF0PWlUT4YNcCzGKESEYQOpupQk
G5qF0quhPElZj304xAGJ+qIaWj8prychAxZT4nR8dAFQhkytZFH9q0MZme3OfWbF
KLPjb8vX5isJQCeRgJDRsPffu36qYoe0o3pwT0BmDmXmGaoO6QrBKxVqJFYcbEVS
B4PEL+FavDOE15ZMb28JRIOlI8GRknn0hQJe+u1RCB2DUhtMk59ZUk1mrScoYjeF
AsbUCOMQuUja2bA3Q29Is4VC/xe7woILK4PyS1catqeshdsGHQY1HkRCNTvwJr4S
w8PCUIRY5f5OP7sP2YI397O8tx8hFKTQnJZspKGPPQtn8CZS0lxEOeHro7HA6PRR
WZvZx/KRirt50FCSGXG9zWQWJtmMPP8ufAxQJ8a9Txax03M5Z+Ob3quy/mo27ajO
79PC8dLEDWCbWQxCLNqxUG8ZruFUQgBBzUJYetib7DLYirHy8sH0jmpaVB1lZvZV
5epLWGSZTVdlLaGTZiDrid5jRiUMg2afHM97AjI7fL+R9V4d2GmOHD5nZvkDsi52
N9DEJt1gYjX4IEQuWTF4SB+C6OTGuKmvhD1lcKIFWz3E+iHWCgme3m9OrjBy3p+N
N/PyB/pFluSs+LTH4Vh+Va16ZTCwKEnAyYhjN/FJBS7QPEScGtpPrmWCblTk1Xt8
HitvtdqAzxlradhGPBh8LWASK4vH7w53N6QYSvO1FWjWXUvdWWjCY1SdIp+5WfXm
pmQBpiQAsl836sKtwT1FNfHUcXUKuhqMB+SB/zR7fTHcy+JfRwx7Y7wp/Xosqit8
KCqT8/n7GNVNUduPELlq2bLfMVFTvWZ1Z2dL7cEB11TBvPdhwQafG+jRde2io0vG
IWN7iNYM1g5zQZqjyIxJlRP4LMjwaF7IMaUA2ZGuvbkdDxUecqCQflaHqMOAk9Xs
gj3tZoYZ4G3HlluyiJHGeS/j1p762ITQD/nlGJTJAaKQTidZJCe36xIyTRrzi+2T
Orx0PK+/BJSL4NVeRkt2ADJYiiDGU8mk8+WZVXZ+7EHHHMGS00apGuUA7Ds5BlTV
heGTJBhuicaBiV6A0h5m8jD9BiAOG99qeEHC9o6TWvjvtWsvmeH1P4kxVi2PelbF
uuptzPz7QWHBde5cEEcVOluvQ4pXesn8oHLTaM7QsT+Ir+rcYX6n9R9ekER0hPww
7SfBOnEOyqRmdc8l9va1EDqX2uMCsJHeknPrFmAdN0KQRXYxNJfyWd60LF9GwzRe
gLjyPx1TMv5D4tH6mvoZqdJgeWk0im+29qPmwpusNldTmIVvljm8GAmGf01h+Cka
qo5CHhT/+T8aRn+ttDO2kQW5XBBUhQxSGFt2GKydOt9muVgic66na4qKAoyjw7NH
Gwd7GE/WiIlGisTSYmvftBvKlipoxGKoe1EZfuf6FCwWiMAC/tbtGuIS5VXdJ4G3
Xy/OZAz5DJz7ilEe+v9733k/JqQDGsqlHQ0kM5yEo+VGSujfn+TGVwq3IqyiJxBV
FTrRxuxK6BCmTNgxEAiPWT/crxLkDmsuCe3w2P1+Ktw1tBULW7gQqC3fA38Qj91x
UOt5HCeWHJi3lduGxtn3Go/L5Nw+cKf2eVytyh4GAepHa55nWX4rQjL0HqhYUcdS
sP02PActZgFNFYAUOhkuluUh1zsXht4gGT8cSBpEGRYRe58lnbafvJY0s940hSPT
0srPJ802cktcY477Fp9ioDXHSqjyC62pWudKxFnPnInnVdVomhSQNa8jFKKDEuTM
zlVd4fgn27HrTumsirGGRSsmzONTASl8fQL8MoIDH6+AckXfy1b2C+dxFsUy+sqZ
CgG7WSTYW5s6LDbtXDg5CcMOHu4vx3cBGEzjGCNVF0PM337B58y1ODKnJUOrKvGc
AhCteDXWZFQjysgs2ojko7AZBjCQsgdNr2+B9UjLHynqTp5EH8AC4gcBSkoRTL6l
jxkjS7amLOUXXNlrWY+xJJaXC4b3p+cH8CQG+k92ocnc5mjbBsE/8w55IOxlcxZr
nJ+dPSOOWFUOxOBeyQiK78636eEcd6dU5NTnPCkUoOuJZ6fHrR+H6ksp+vLNApan
oicJ6yR/RLlZufl83m26L6B9wgA56QhTne2YDYxn87qam5aWEBkLmqMexm2hkn5/
UR681lS/PK7ELTUrRAANEvYEh7oNL3hq39xzsASATrW3mDcwYqLYDjdNMwcICzkJ
btLYzbuNNlYZClINJ76sV94O13Ys3KsTOhTe1b+aA3V5ZAOz0cZaGp3XSOVRLhzR
h1Gu+XGbHUPUI8BhqKjSYzMypeQYSL94nFoSYFNpnzw/yXiqDD1nTKFJ/mz5oh8x
Du6074QUQ2srJx5ov32mUJwtZIBD4Ard44ub24pKsLAPzGxl/p5npHuXQSIn7EXz
SRW0NQiSqRazxC30T9D5e+eZoKpK4N/hbT9HkHPRKv3zg3ATVnubMveWbH1NNOuw
E+grKMLk5A10hQJGqfLTnWMoNMTcUeM36eKk6uINuDszTWzI8GJi47HmIkHleN2I
Sa877qIvvu0us55EnCVnH0xvIShY2EgPnr7E99YAkXFy5n0hz2JYuojh+s9l4xn8
o6I0xZ9udK8ekf8AoTDJOjHE4VYD1nSVBhdcFs/5QhsUpLwA6r6j0fCeTNznKcDS
v817UPgsf6kd60mt83DA9Zv7tP4JXXgw1hL0RdyHIDjQMygTKF0k+29WYocKF5aG
CVCDb9d/NAtw4O8bJq4tnBAe8ofHCAX8b0eP828h0aDfuykVHJlrRqy8lQoR72yY
VOGZe+xNvL8IQv+/DbjrWI77hLn8Ruod/kwkaSD2RFl0IwHPm84jIHyMUO4Id+xb
9YXceApf2cJEm6KFIHANHBSpdwaJqQRinoEVQ3/iLlMpmgteD5d4JIUzn2SfTQHA
+Uqh1m4PE2ArxSsgvFDl0MxbA7bOlDJRhiDo3g0Wx59Myo6N3N9FmqeGx6DJeVd9
0et/dNQB6gXQCelURLPaS9ZDXsNrdzJUpwkQUWv37ni+9uzuUaaRYN1COofdsbHf
AoKazX52NpMwZwi3OYXkPiRUDFmxH13EVkmcwTtiijOz5ocQhzuG6uwWydO9H0JW
gTwtJ5LjrdCWqOle2yuxpANf/jyMDgTtRHayiKl+NM3vFGhG+GfcknOSQTgnI2Y2
PZumNiJjAh/LNm9o+Z33nzxVPbX2COBupzwf03PUHF1JiZJNKDVFiNaY6Flc06f3
If3mpC1V4BLwNZrgPXn67b/qv0X9KPr20at2SdsS8GbupGBXlye9nRgCvJX3NoH9
IoIEJK5NwNj0YHJa5p8dt79ktf6Voq0Gp6bCYCjZ1YBPbGDYPq8fusZij8/3yutK
Xu1zS66x88UZKaXtq79tOMErP6OxdtET3ViltTHu2OhkWhsZ+XIO3dJkFNUA0U8v
Qvdr97+tOUCxFEqn8YqcGlfKPp59lld2GNLfUi8hp4Eu/Rpr0fWFGe8AonH4mibf
zBiZccDVVowZWC+mX2yV8lM72/vTkSd/FyXJ9J4wP3IsYx1+oNXmWDOOLWEJukSq
mISrfa4HW5knh6ph98HoR0+be4IIJ3tVEmkIPHYmmRVWoo3OYEPlFjRAsxjXix1t
XiYahtUEklXqoexrS3wi0FbfxKKvbBcJWpU6+CvlMYqBkk2SzKsSFROv9QNIxSZS
pAqRaHjI1lOuiPxXbsmk693kAJytJZa5r/V62lZ0xd2FHeQUEftTZw52mXo6NWvl
Gp2YTCM9LXWTvupE1OiiAOE/J+ubZcK6PxFJqyvc5GWL0xgwjPhYivwIXaom9oze
1vaVm7XqgTksybp9Ph80ELaxKgmB1h+5KdrT2fuo4D06Yi7ptkBhnxIiYsCImkK8
7SQNy4bsfN4X7rY5/e2LMvuGid5OiCwHjBPsQ4oVXnZ/8T2NsqD1frz178wDekh9
ESTrlImc5maVvS7XAXBWo9woLqoqfstwWXxJ0Q2lLQQbQEPsALnT9X+h9HItU+Tk
90A+nBl63jo34/22HVhSwj/vk+P0ds/WETFvpx3LyQR/nHvy6eytjpVPZaUFBArk
If93u1RtszVZvaontIwrbgAXNG5p3jK2zYeVzDnFxaBCyKCeUTPKuMcyWYyC6Q3f
py4i8VZHHAXtzIjyjjjW41X+O092Zpjqp/48CO49KA0bfKQ59vnB6by28uKAdHl/
UMFtIMlcbl969oHwS8lv8uwLDGwQVY2YIP0XB1MlXeWxSHCHsv1GImZQGUFcABd0
bLSZHCXASNk164y4V6UYVHsgQSDKeD9+E0NEUQl4tCoLy1DeM+35KyDduwgGpKoR
DJntlSnzMIFt/MIUOnIrsaJfB5++AmN2d3u/QMhpNTrwQaH8iG76/8POM+vMxvUR
xBDsfgUDGo9KhzDzuxh/clrp8v/07XmEcDCkOVXsmteL8c5UEY6MAqwMsQZa+Vu3
0/qZrQBlbOlI7oynQxikKw9bUGGidh7bzYu1lun+ktaAM8m0NncJVrjrecf4ZNjN
VOQ0SIJBGsCYyx4NjT7g6enWuOjLW5nb5R7nZuAnjwXu+hurNLvN8b617240VuLP
rWyP3AoUO5SHl2kUzhkeavDoqhQpUB5QrNWYEa5/dU0XzLyVUysThdHqpafPWVvC
h56q0VevbOht7LBBWpC08YdXP4gXf5lKFxPxB5taTs5lRkQK6FxHre44DbuziZWZ
OyG9s/MRuKYj8iz5tmt7s7BlGSgK8RAW8HceJcfHjdhPOHSBNVuOcTHyyBYCOHir
p7pkzbHWq/gdqYPLp91ab3fF113nK3u2bRXmCbdGOqNyICtX3iDmEYITF8kw+tXw
lzVXfo1P3ZK89PFZKuKqUWoBE8uk0f/59IDlI1jHz+z1KzG0gNT2UlthP8VEKsq/
jl843ZlPMDctGkbhTRLtLlabp4TMfBhGZq9ZsLudmwucJFfQ40nYKZt7Vrxuv0wy
gvQ7xpFGJwpZPn9Qff9XYv7kc7lSnr49l3aW4JaFGlhCVVEPOGLNOpWfSSCod5JX
vwRY/jYUHkd00Vc0gQIu1acz/+5jDw7Oxv2aQIPMJrYkYulE6wOZvoOEA9/drbBB
H7sl828RCIc8Nu1V4ym7MHKaoGmWiYO2uVHcwhYr4wcPdH+4yvnCexzJQFILSCOH
+kqsgF1ai62Q2sN3gAkJHv0M7pDvi08kmvfic1b6Jsmr6c2ml7QpLwJiJlx1931I
hiQ6BvIFUbK/EIE2q/6Vvx+cf3VPQ17TpqfYm9GwrUXBDjdQezgZ9veavpwX962P
SyEzaXvr9WW29zFtBmHFg9A7u5AO3yYrsan0EzNuHKaY3TKpUOwswpOEQ+XODKRk
PFwSN0+Ci7E7lHOGdnzjmEjfeXRh8oafqg8ARinVhQBp0KnCMSy3AgOeTgrD7qv9
NYnQVms877pi4sVuK2FK19reb4dRNHH/N8YyGDVj0fbchPuhyJUA5iuwLY4y0gP7
g/WbIpTJBp0kfZ9JVWAGjunf4jss/GVuWFCce/P8tO0Bk+bu494IvyYEaTG+NxVK
AUh7y9RjMeFVVIkkf1BD+oBxeOibx11yPjBzZ0eNesh0b4RVTXozUBqgOiIe4EG0
ZM7WcLGv3pGS53JFVs8KX6HTNfb2Cqc9ui+vLucrq7deZlajST8/JlW1xA52ip5+
MvojvmKjVPpQMxz8cjSiNkytVp2cf8JHn+e8PGARcW0hfRkVflLCs53Oee2quBoZ
4AI7rNMQg7nuhoTcQELUaiuMn/YUIZcThtB5GY0bPJoVIznTn7OnDBxj0QKR1rvt
IkUyg5cvusAfmy9vx6BzsrlUCqw9ZT5Q5V76KkHETXBHIEDbR1kKDYZq+ih9hWVv
CjpocEKIfwscI/qLYptEHFcUS2LPEDlnrdDSmslpXHABrJ+hts31vMTmBI6a60WO
8nEySVk1hTE9+y2Z0/UjMjTgdc/WRdPwx2hls5Sy2fbc4hBPI50chb6XaSGqg0Yg
NYSSyrvmm8LfhNWecWVkpF6EsfxnPgWKjfaIRjIDSRDjqqZmlKZrKsXIrhUOiFqP
q5pK4lhdG3+V8W4P1ymFaS6pmSuzPMnU6wvTS5/1Vb+mszWO0wds/50v89CmCi3s
cC4RU90BEcmM3RipUUJOxEGpYJrQLLlKyzlDCVqihdnJBJfgTNBxGAj/W3JqFPUI
LYXqfSkQIVCReTbFVn6HdL+hmXro/ODsNly48GK+uLdcz4ZAn2k5ZJZMUN5hFqdT
gWA7rlPiPd7jb6LnJ0gS8Njw8eVRuvCBrC4+Ta/s40iInMI4ZGcj85G6XVszIbfP
QO8dOpa9MGUMkQ+wOw6tDeESJ09mXdg4eGLlIl9NarjfIIUWDh2bKNLlEAqeq7/9
BQ/0UuuIbUlwhcdjBgfrnIcvEcat26HzOlivnvj4/oFSraSZtbKZbTSdn4pyR7xJ
/l+58etOnic4Ybbhuy1OLOX0Qg84FDJdk2JfwhtYEAaA7zZ3R2n0ZZQoIOtQr6WB
yRB1IQ3H5yqHrKk+U50GBzbn5GnmqUcrfnPqN1yIunPlpmrRoBIUKIGgXZXppR4z
EKS0ql4EIhuojIjBLAhDMgcErw+6+lsPXVpE7c5sGpFJxI6Qp5JX/kVal0OYfmx0
m6Jfel1k5dhjXC0rdBMGcuib0bfxsbHctNe2VuMvOM0uS5/3CFduYET1cQmyqA+d
Ao6UELjunjf8IiZj0ZAmVCCKAOd7s0K+HMG7FnSspNRXsR6RvQdyZZX+CeAuVYFN
3fiR47i/WJ+26MUjBUZ7XV1Gpp9Rx0sWd3/gF50nPULOhnWs+ISPHRBhA4/elFYW
PeebsTCVVG1cG1d7V7s640uTjfXZ5MR9VhjCCd5zsC5DCEzeYYFMIDByHRnWk7tU
Yc9m4PrEr0dKS1D/+nK9ubI69GQ6SbMH5qVT/LgPN1x2cHK96CzOqNzHIA9dlR1V
0wcjhwLubM57Q6pFs3WMz46WNPwsbw7+ixdrVoV/9rog0rCUoOnJTkqn9Y+LxZ1w
RHw38oJ+l70LqucpJp3qY7bg5UxpjJJvUUlqNQY07x1nPpd7uluMi6hWRI412tg4
t70AkjQbT9gvap0/VY4gFVP5OXToiy13JcLy9o+ILy2qL1qhe+bVKaThEi71V+fc
rwOxXxOjtrZzbsB9giqSAy7ePiaqD5LGM8unka09PLcwGciL0CEJ0Li506HflSH1
3DxP+W4SSlagmDPcTVvamWB8ffD/xVbzC051pKDSWBcBL9b8UaQQE92s6P3KNIS1
c9HiL5qCuTNy928Cyr1MuRz54R/EQmPfsqpvM/lpkiJeEq1M1760+XP+P/A66idO
xGIH5RqFFhEcqNLIT1P8PZpYKaYEJdPc126zHfxoUoQK2a4lObsrEfL8qGgvL+Kv
P3Y//kZZ8t6lwMWejMIwEFOuh9VSkLO/Bd4fMhKCacQ3ZKvb6kidbpSvnBAQUDJ9
OjeRihig8kEdTDMJryBFuqEdu+l+f/aQ9n1mLSF+xJ7Uq3518oqbTycp02AyJAas
VCwbySiucH2Rsu5i/eyaUxzsKQMhLok6fj0Lg+RT5we9cJQjfiAansXJLtt6eLT9
4iaVV/QrprAOoACfNibQiE4Twj/NDSMJxlzTC5/lr+/zL82o9d+JC6XrnqEUJECT
iig+vGS8XDZ757zQGJqq0qdak1XuW2Loco/T19BGuUEH5cRkoAYuv68sTvgJdy8Q
5IXBXNCrzRD84b+FdNTbS+SQkSLIzNF9xlA8juo+5ZawNmF9Wo4EXP0nsbslCWFC
iGN3lMXU7cAmETGBggo1Kr56mjdi9oMleZFhzcdK7aIoD6pvQ1a8sdaW9bp3iZAI
A1VXK8AGoE8/9z0mL7s9zduoMqCXoGgHclTiMso4WjonhudiWazUktWcA2/mk7rg
31UAYAYNp4vrlJr02RKD3NLVuFdofpkOim/wZY0in27oFAjHjlfj9GGh3xQgLs4R
eOJ/FsKgXH2iobYzxphjy2kmTgyDPPh32AgzkoaRJqOpfUQvr7Xf3WSL5tgk68MJ
00aPjs6lRW4e8A9jpK+mg9HrDnQicUkDZa2DpCI6HRdmhP9oGMPsQR03SNIB6qsZ
ay1WlaPdMq3sXEM3/Q+N5xDnJd+hfY7oglunYNlRX86n1nvgdzRTkGTCC6joFxzb
fNzIE3oZ9ncqGn9sRQTpUoKa5j2MbgFAciJJjhS7F24jhVQMPmYdiFZIInL2U8G6
rkQ05XTuPBC5EszoI3zRmy5aksZpUsh8IxeFXbEp/mUeohzmV0Gcwq3zgMksmesb
GYr54pY7UcDOVyGkb2dLyTCvxiuy5T/PFzBbQQEv40oyVd7GJnTUXkPExzBp4Zyb
Rgo4uIt5g7yu1VeqlqQ5lL/8RNfdmr09A0zPc9a7/ScSoiVcIYfc/OsKLUNMIcS8
82iMp7kFzsILDDAwQW/fTLhmCSsOwSV/eREP0FcRJ/j15nXR4B33xhPU1WbUhKXh
eSevwyPEwAbvGYX2RH6O61PW4c14RXMAw38pUMkPcZmBMA/UZS6dRWzKCFutFbkh
eDSiCGnpJ0VaD3/JZIDm9yNRo/EXHivTwpXnCCG3H6irptRxyWbKBW6N2Y3N9VtS
VcubSqduqkqhnoi3yJhYXIkL+1rQnDzNbXaQw1NoQJtRykrwImRbveDdKP36wkOO
Z8kjjC2jQzqMGxtcMAFvtE7n6iJ21G079VbbnKB3/cxdPQ2Lvvmk5q/JtwUHBOrH
d6V+jw0RK8oCUFIDMLyoz1fP43UYGlbDl75TnujP0UnlWx2EN97X5myJXO8Vvodu
jd6Q+zeBOsiadtUApDKit11Bxb+wlPretkifldMS3zwGXqbFf6mg4m8Nu5qRtT7v
iEd6EIJo8kvpgTdTqPKrZnD0NcSHgXtRkW/UbhMD5OUB7vCRDs4qnfU018MlxKbe
2Jdz+q2gRQvIRMqhcf2gypJYBKFVq7eSZhiwrEQDVDxvsPHmOPQxuywCBJgbSjiV
MfbNCKJl+bUR0pEtojVE1pJ3xJUjRNqfN89TBkT3HRTcPusI+Jqd6W3s+qkhdtBI
OuMDG0+RYZHaXji+jVUrOJJOzTHaRhuaZUy1uhssm1UGYo0aaP2+E/M3D0jPVVhL
FWHiboytTAsBmbPAJsxFGEnyaclTDNLUCt0wTGgByLEUKEAI2YJLe6FbBZnBWKxF
b12sTPBUpQ28Unsbkb3dc3eRoy2tSobSzK9w9yOo9WsA2K5IQ3xCy6sctwqfOgq4
LqWsWmhal0JPo6qnd9Rf9dQdHhyJ52SzrsdZxzjBRkZ6wD9SkRlJkpUVONT16i7O
nClBHsqd898KtNdv9zx3EV2GOPWU2P1VFtzTN6xhlMtjouFVhSe8cxtNc8JJBwMg
PVqKOqCnBjv1O6I/ZR87+sLpxvLoz0Sk1SxoU3KJxmUNBIWU0NK+Nhh1BR33I7KC
3IrHcr8XdAoZUdwqQjnEc7bJxTNkXmnV9+Kkm6AfV2eORvt3XBGpTWtZ7n6ZYknn
Kh0s5ula4zpnLg4SkOOSeBFLLnA/O1yOX5pW9KbM9wn1tcWZW9iSpieyysG2CECQ
ZBNynzZgPThxNdQIAkDpF9eE4as1B+yM2+9IxOlGBCUNcyk/RFvY6o6m4w+rGdq/
iVZUq3KTIW8JcsrzSHU3rX5JjYyh6h/kRJ0/hOzcPRSj+isxo+4NZKUssdzHFLVn
ZkiHo7WrroKWh+NUGyqMHhe6ZBfdtKvCVKvuo2YkwdTXNBvx70FVcXzNG5Hx2gDd
KDLX6BNy3r+8KjX3IcsNbGpNzmR+jNiBKkDWyB8U5CsG54/Ilr1C8SFpzTYbqDQ8
NOKzFgK6uYMEBJfa+SWWxwHIx0EowIAWyB5y9oaT6SpE9oNcC1M8gKBh6qgHJEBe
CUeRpR+6HdLv/yiWkmdDboyM4FF9chzAmmKDqip6UMnA8t6g81MmOLV15g8ZzL3d
2uz0c0DssSTKR1PwRfWDWCWu2athGNZJfNdubG4VjN5fkwpt4iFFqeevLvTLIo9v
0ZyeeNsjD2MvdxL06GiwMMjXInLqgrQJ44EmKj7CKtpxSzha9oJOyGhRl3DfVUHN
OhqaEtkF/LYB1tKUltJwf7o6++/1PoiKhq/u4Hky0K7guQrsWMDUGGNEM4tJBuyy
bx16+l8Z+EhwpBZ8QwiKYLeEHP081l0Zh3In3/UIdswvhBMXHppjBiBIOUU69ZxE
PMkzCJQFB3U2lcwjQoI4DtosS8NS9tccalvSsn11W43dkzBzQpaie4gueG2qZ8wH
Afscf/HEa8lbeLnEckpf17GvmgMkGQ1kfIYHi8sWLyXVvQQH3H9+ypgDoro9BDGe
NG3BcKqe7TT9/TAINBZQ5ahwK9IWGen0H5aLCBzNX8WdVwm1OooAzZTASxsWkCjm
z7UG08uoBxz1boFPqWchHgDQIuO/OdRZqW/YFGhxitB0QesvToLHNCcbnk9CkIxg
sMuWPLuzibkjYWHrbY7Ps5Y7CWqF18uASyd2e7R06pRzZU65DIPokHKeCY4zJxY+
Z/pb5J2iAVCIRiZjjOi6XJ9EgTKD3epkKZHOCyRf2wOlDqja8m5UOI9Bbehxs/EM
/jDSlXXraXY342CndcOlvwFwpEGI8BSPagORx4njgsNM1mBoQ62sax5OA4WuP0v1
XOUQddyhbpDPOdvGhfnUeHN0nNM13ekGJMlf+/UzLtCAGct1ixPgLpm3snvJOsXL
G0vfApLHLhGb2SH0zpGwvKk3BTo6mZJW7EY2LHG4RK03OHBF+dQGUA1wi4arEhVV
10wsvU45zfCHTcPWXEghb0xol1MqkGSraw36w24Zx7N20lglPU9G+l2FPqdN2rNC
2w4C/Fabm8Ha/0UG6M4bb8g4MIWwdl0gkRyLdOPXufo6c95Owm39cGRn2PUzTxmY
XusJ0MT15ejX+3iq9wFxXdzgNEGjLCa0VRg7PFNj6ae2pPFlFC8sHxOUMG4KCyQ5
OUaxsKnpnM8VDOzLBudYGkTaqTmxZfCyzEleafVGJSheu1Q/EXROVvJooHG/mIAk
cTVAnd37rtMalQVJFiTVum8wU63ycmvhgpthgLTnNVJ6y1+iPcr3xoYgOxBNaxlk
w87pmL4sL2dEK5HLpJHaGI0F42EuLl7wO4eCYP+QxaGtFOelRSfTWCyLjevTQHBv
mtKwmSQouPRB8MidMnXlM4xUNnvB3fKR5zK4bAlYDBO9CfzaV4oW2Lk/CNW0vsG2
IN1vhEgxhON0N9ecZPUNimO5H1M5f7yT/SJjppPdnFJBw30J6ekS1delwWrd9nwt
OKM1/WM3T6u/dwuDJ8lGlFYNHQDL+sP+DQE7wM/q7cQfDQ854mM2yHoSj8L9CbuJ
SY5e/XywzhwxzvGtDt8hUtpyXfWF/DPSpeQSALot1mLz9FmyVT4UwsC7+1ZOJLn9
CIG/+DR9FgGn+9st8JLI2eYSGV/dFDatWLB19ukfVz7/4o/FDnbL/nBZfQDzTBPl
bI87YSnjApT9Yjw2033EQ/dN+CRObGMgecTuQRK1YGxDy2JjzsiQ0S9sqC9ly+B+
Ac5xo6JemUN7vVTeN9tN8gD4UcIjWliIhxMPIt9gt2lyIoDeDvL/I0vbKKxLPCqI
RP54kxYp0xiEAdlbSW/FSuF4GSC617D/IrZfgsSO7pT+Yd7HLZhOlX1QpnehuSwz
5HY4RA5VWL2lu3LRepWxjqSymBJdg7OObG6T9p5QXlkAyx4+cVY9NpTgDIM+PZ5n
cL+r0kutibQWH0UQGcXv+wKJB2xl5S+esFsMyWd4nmLv18UugKsOGFdWkLWL67zE
BIfp8KeWemcyz1anipHSsPEd3JZVhTAIrb5sq8PgPsXP+A5niPC/IusK+t9VwE9J
aSQ16Tc0AsEEKFhGgfAJOISk0lOEtESG0f45H1rB5Q69u7tfrEpQZogPe69g/Cyi
NtDGAV0FIbKoU9SbqZ2UviDuuVgP4Zc+pLdSuefMnZNRrYAhMXqMuHrVhP6NNdHM
SjiRSArbeuTtnHqv2/ZavXpX/e1xGk/ySWDQal46ZcwxqCXE3i/Sx+bMyesCOiMk
98+2O3ctwhnjVZu5FsZGfOGNaOCNajlp6WRkLV+K1IfHlXhzd7Eh7TI7RciG/+o+
Q4noMqIf+FYJrHbjE503QMnUFbG/fBbkGf4s2oej+KLANTFO/H8VuIBqL5uvplqW
1n4Xm+XiJ54z5aSv91pb4CeXpvk/lk8CDXVZlm1pqZxH78z3fi5pCtVppmiw+OBC
Gp2DpcBsSM4lfvZl5moL8oxFBE8f3FkLwvwgHw+Z2q5PvPQioOOpcis+AbDkw+s1
aQMDOiM7Woask4bsUfGRvr7GoPP9aWF9AE8Kc443Kxl1PgX1ffdzIW4J3biyyt1Y
T2L7xKx3eiHFmzJYkOSjTLNkswtwlGYBj1ey6i85kn8Fx+JdnGJC+E1aftxcUKj7
8bQgiS4OBYPEcCgsnj9bD/mCWao6esAgF/df96qEBADDzC78pkClaUYrj/f/4raJ
slc9NSULqtnBTCRNz9/NcPNrZ1sW1/bb5i2itwTGn22vLK9xwLirHEzrfqUSY2DO
plPiKS3W5GMnRdg7WtngGHBCMe1Cd3i1qBlQ0I+NIUZBXDwmwZV+aXkm18fBhpOh
WfxAsmbmSqPzbwR2ffT4KIhaWY0f3yWM+9r69a31+ujqIilqWRczvxHUmgrjyXSe
sDETH4kzoQg67wDgHRoegVjnwTtampa/LDNTzMtti356ULw+2AgijyN62JvrM5vP
qw1TPJQqQgKkc2pywSZcHYnae9ekFnQTy5tRJtSpXWY2/1Cb7IxMxY1tInT2ROn+
ujNKiLvI3BeeQsdlUxtEeAgTROw+M1EmA07OfERi1xYqwI/rvQieKzo2TYxFFql9
0jOq2S28DlNKA6lD0vJK00A529csOEBAB+gPFWnmXMxuin2EyAoFVJRYSnMkEkZI
A8YHDuGP0RnhK4cz/zLHnLGYotYL3X4024Jzztrh4BJtDd8hWP0r8e1SNfxEipTw
9M7HdS6+5mnZuq90pgZd6X9SpdWbk8CTW8TKFsfvcaDGrjloY7IN0i5i0U3DzZNh
OY6kIhoJ0XdMOBXb7pYcVQMVHAdga3WzX5IhieYMqXIT8yvsPUzaSJ6aX9ZIoFXl
2lbM5BThOnYYieBanr34PdNGwfDsfEJAyQkjSykBy/VqePCs53vLtB1gEoZ8vXwC
BmRfprklH2cgWCVpTnkXq67c03dX0h9oZL5cvcbDWEPYZFW7MGpK40o6bIIjlErF
c186e/QiLwDQQ90QlzydLBcKD8rbT229wDUeO64pDZQYHoBHuF0tZsN8aUUSyf0k
fThh3tiPZMDVoIyjeuYx9MsODuiRDK1e0fnIherqvY86XHYDCCUOi7yqgazXpqfK
+gmuIMM8Z7i0IZYX2O8ipnlaGotcFTkW84aZ6I9/mGL+wYKn2Eg1pZ2DDNJVZ4XK
u9f7mvpcrSiGMEAnjhD0wByZnoSmdWhQoa2z8aqJ4zaqFHKJG2LQ+7KDaJnAKaMq
1/t32O4X75U+cmJnUQ+9nc4Ktk5RGQxGB68wsKP9yKmL7AsjZGpO0H/JcYnmFpqU
fhlsyYOhzl1hyTMAy4biSnj5347QnqS/F4hAZ1087ybJ0bnZOh0ZQqRLK/mthjYe
HwWPDexTbDGftp0tKcbHS/uEhPaQTrrP22fnlRq2b66Yx3K/NexRa+ZSOqfuUxyA
BiU7GcqWEcUHMeMT4vJ6aINLVyC6OBGUZ/SVb5HmrCFDsV4dXarkjxZMxwyUwhvH
uniWWSsEKL+KPtfycPV+q6CBOj5bT0fnlYf6Feku28pWT7mocAseDhSBWwSXHLIl
ARQqxVZRS+ETJIUoFahsNNBOEhoyUCbF5gwhM9iUPRY0oBURLCQwdIfrSXt3Gera
rK4cr33ZZQx3JS7CtIV38GeKMI4iij93ndOGWkIgxXu3PrW4kgWPaolGZNO5XkI/
NEX1Dqd5Cvp2CT8HUiBZZmAuJczrXZFdOuHvexdvS1396Mx1TVPnG1QqNndQu6hY
UG+SQcVA5j/2RCCzwmh+ucLZAXboirvj5RfpNO/m7Ct7CGWG9yqqfe9siEGdqFCi
39gsrp6wDyReijcewRZQpgNGH6HcMiMgBpcIqvuWAnG36baddHQbgmWdPfjL9yfa
Xk1xnqzjSSG+VjK0/iO8jvx/Y0LfRSe9JKwYJHnIyl5Z4RCdA3GLZK/Y6H9pZTo/
6k164kwPv6froPUb7ynzgtjn7ZazKtP5BAdJPNA0oBHbH7oTdWEJLSwrHod5lCM1
7gwBVpEX401c6gEdJfyfPZ10ciMVVaa8ksBhYPRY6LSZQ3CEgQAwUSJJjz3WhXFC
F/6C9X9mD9cvrSKGe5ny/wiVe/4niz+2PtbzVNbEPIKkwZ+/HEDl7dtv/pzMdMdV
vCsxOjeFNO14nOu8OBJGRsc/0ONxbfEHym4T0H3k9+6AWrULpjTlpNlLtVowl1NH
Fv/8zqZGZhFCVG64/4r997xPpNLSEFtnQijEmqjEekGgx9boKOh1yLdtpz6VeclD
I3LMJWiEfd1TyK4lQGeOC0RwRZqjCEiRBfJB3KOtjh+b+9UGjqC3zwq7F2xQO0Jt
9MSpEA/CID+jj9QmRJFHqMvhhhDut12QJHDmZPbcMzK7y6q3smfmFjIs7DdbgpaB
3o268l617shcHwgGXRIEnQefwmLqim+//QQ3RvmQZuUjP1U1Q1iMo+W9GN46Pvgr
Y07iSgrUcwTSiH80+jWEqdnBscdhBfTIzhlu1lDg8ZBbfq9Qx+47YMDZP4HCPFzC
HjKnvk4mJzIgsOsOfMGXLtEd3anbgcqRaxJHYpJETgYZeCy6sEwLclxTvK/nzqfk
5H9hfb5Mxs6kEq7mUUedNszFpdjI3TJI/4eKXJHUuXRJX0ZQrfEU2iyRiomZzhEe
8+009S0J7vdBAZABXFN4vBOkpin5WMf8csoltU9j5EMPqqJx0l27WoGIlheCuYwi
zVo4/ozsGXv1BMqLPji1OqUYo/iwW1qMdz/RXq1WNnJWeOZs7DdTxq4OO8vJCEdH
jlha0v//cOxBRzx0O+V9WyEuSiOonBsoxMgNrMrGmlFOBMeYtvQaLH6rTf03Tm66
3HoZ4q2664q5splphBNVQzc43eNXgFDm2E3P1uwwmnBu2PgfFvJ9QBlIxv7611sm
HS2I9GlGuq7hmjfQbv9QlFax5aPGKrB20M3Q5uKwuSdgJic2qH7Cwt9NJ/hrcfdA
VeppCpnJB3hPTuhXExDXWGDxvtMhVa9FeGk2Sg2OC13+HKrbgGHduX4vx5+4nHoh
McAmoGiqUelzNTeHUchm7Tjk/YzNPtxyahkWPtal/qhAiWGxuZFCthbDULAyzJmZ
8QJU4edmeevhZErTls0SD3XB/JW9r1Zsbx92/c6DeVMV5oWSyqvwRgx4XLMX+IXQ
qi4Jq4mNxi8gMwoi1AURivMSYszfD3OJZFuaajt1x56dTXGWwF1xe7CMxMYmnmlT
ANaWefm6glbyJa9G5QjOmqd8ong8sVLL59wy4wxJQqR9D53Xf8GaAkBOST94QbZG
7fZXDwwCGwGKvpLZL9jimzQSaxeASXqn3oOzLOnhkNzJLQ06tBDZCKhnhmwQ+Y6x
hN7/LVxesbRHz7Ojmu+U5WvB/cw9z25rODSmKOElwzUMxsXxLir7mMMoSxV3I2ew
ahRaED69xekOi4jPEibgAREFo/GIuh3qAl/KjvhSekVZOGezgwhMbVx9urHjhqgJ
dd4KAmeAAebW9PrORM1Z9XutFq+K/vD3QGRJy41jJ601vuadBG49KasW5ygPhIpj
KVn3je8+LH+GVdVWSnw5LUIrqbi7rHFBQj7e/X3o/aZH0q3KxJSmFY0Gs3qR+Tr5
aqvHa/py7KrjV9ELqJBu4IJqiPAcabb+74S+s0hU4pqFrU3Y+jwMi6a5+MxrFMQ+
nKMNnmf3KMYEy+CSDYiAK5HXin+NWBg74CzVgSAi9yI4sQgFD14Wz+/MsNzTml31
Ydgsn6Zi/heC9qDlofcpHLHBsvUjsuBhTk0C34bEh9VilxS22BJt8BrFJZweEH9j
7/K0oG370FuD7QCalfQGQx2DGiHkylM5Qq3xAUBQ5bXJngJYjWSECQEx/rRsgnnr
GQTg0FiwoYKpTNWn6+qfvj9nLHKWudtWuey2dop/dt8PvQosjoe2GVTud8LKTZad
rLgAt3WzLDo+h6o/xRYPOkueEwkPa1C7hFGpBbtFSUABR5TPGZ1v5A3I+Z/kONrz
AqOEnuVq/LDYjORiq0yRYkqTMEnzK5n4sZEMwrFGT0XiHcA9m2SVxosKuhuCtVw8
1U3bzYqEROF3XFMrgQB0HhIhJsNCF+53vRV2dLR2HGkcuu5ULCT27S/9wvsXk+oU
OSLmjuddCTx8uyBzhvO67k+yerrjfGaczsWz0aOBoPPjFrjrbdlbKnfPUBeB3TH9
uKvSj+RktSFIbk1Rf1l/fleDInP64LG0DUFPRjE++bRhTQ6eEY9Wm3Viu5DAAIby
zURwXvEFRBmxb2+8YU3yAS+fvMWzTyBcYxO4hk8Y8I5yVfhjtsnbPaNs0vUs435x
hnX0KMq1SNqD3a9vnNx4dpxfQc/bURXRxh7sAAY3yFYFbQDgBMyVBsfBb4yYkToS
AaIe5wq6VWJZqm9yJO9ZpZ7rMWjHOjzDVdOT2seWquxr4EnzRjvSe5jH4gr04H1k
H2Hdns+aC+Jfvo1JMe6PE0PqbVfYOe+LXZ2XQc2pEZlo56hPguGmZEze7T+P3qvr
BB9C3+V1DntD5wzrCK0Hxl2UNObjKbDYJyBvnmosLtRBtV0SlfqQCPSDUjVw1x+U
PV0Ffm21idFmVOs+aqm3yWDSANL2S6BpSE/Zv2VADvWY7l4UkvybQZMuRK+iiKsN
BWFmItLg141aqFEfdIkjkL7+DujuOXI9lCuOn4yM5h3CNcQNiUSoKlm2K9r2FYhD
OBFfUx+9nyuGahqe+B1UwXiKOpSmONDMDDIqhvSx4ZMJ4SbWXEOUIKQ6Zq/7lc+K
wQpifxNygc3I3lWmN+21sSeIJ/xEVZ2F+ySqWp3UpJ3MnVqac6jvNMmWzEiKfQHo
5kz1Crm6P0AXMWe6qOh6vSGJQW2iN/WIxYhB37fXSe/Nq4aFY6aQDfCWPHKolSce
4HW0QmcAAhhILdX2Rd4TLe4qzBPp0r0HB8RbYwpiojqFXiwnCqJ5QKxyVPcb1waG
5tgNMNNh8yhSajKrmBTQ5+mcdJVtL9X5/9RcDC7SmBF12RINgb6vWEZLH7dg2Ocl
nEJIuZGkL1iLGSZqr3dh6V41Mw/tSavVKOLYK5mFz84/gnXpbqfRIgkf2ewQ98j/
lEV2fHG8NjW+4xHFctMGbhQAY2lT5LC3A5QuvSdBsEptrbsD++LNXIzyakjFba2C
zaMtnjLD5dekGtb0H5TEJaW1f+Ji7+FcrJV/o9LmGdPZOUXk8zf0p8OkxV41v/hT
Rd9onkZVNZVAWucjE9rZvZtyW3iC/w0tzz49gWTlUDu4gvg/N3FAMPwdKhKfRJx7
XDiaQTl8klfgi7bQQ0xqKK/ZlOmS7650YOJDrXSNJ21Yr0Z+Rtx9T+VWcaed7Wu/
yPvdBCGEzDXu18PfnmD+K3G8sLIGyZogKRZTS66qL7GiNNll68fuHSJh+h0FxYmX
dS32h2znVTs7eD3jaQf6C3mT1+8Fd1JiY7f9LSxPe9ricWgFkRmYAHLT1KFENWJq
d9SfcUNcrRta89Xj4nJ/7vdHNNa7y6algSL/SselJ2QxUE4z8Jm/Y5Cp/1geCcix
rJj0QiE/RmrPKcbUE0I2RMnKTUy4+ixsLYMxGO6yzDwd0yb+I9W1j66G6MgZEXaG
XYcfliTdhdcaEHH+letSIumUXROxcR5VgIXZPmWSsOSt2AfKhFee8XpLlJm2skna
baRO8lU88QeFGuGJ351yki/nVsYUcjPImfaX7NgPeQJ7K0iSIjPzOrxcWVFJr+gI
lKZCZiIwwMYvAPmPD1cWa1P2F39cOqHP3YPr45eSfjqv4+zEvucWruAXfx9SvODe
ZnAMn2WGTleDeimw3RQKvgRE7RTloePdlEZEjRnomP/OBYLJHWyPH809xDcZA7cu
OSwmzf/2anxPoTLArts1BkH1Cm4R/lOGUt+euKtb3hkFZ1tEFqGm+zQYby0rVRAd
zw3Zf7K1vOjxNwPmXN5e7IH/GtOW00hM60XytePgD9ub0//KbVn/eMyMxGzU6D6n
p7gOpuYLn76ArHj+a2Nb/KEP90g64cWLKj4UlLdXvcCHVsV6ME7hZCT3kN22VUSN
8zWNidibpm4ZKC0rCTkjhFMp1QCwtgVygqKOVV/jfppSb8rUvjyY97n2SUweL5Tl
lyQHoIK5CNAe8mjAKzrIWa2CqwyVRyMDwTsioHb4p5qLGbmSxFD2Je8SQlXqPbUr
SoIzEn+9eqL1p2b77ncXIMhnA5CnfA/E5tMGX6qG6qtwNTvO10ZuD6CozH4Io4d6
g55c5qgPoAgo+cD07x3++WuwVZVKV6hC8pFe7Y7jH920Jf6ku16OFwwKjk9CRnFh
WYdwfBbjvSIwjmheh1Ig+QGdL0shYMbwP0lToo4apvjdCTLPQwU1S2jan67LvVNj
q2RFve3ZpIkpyS7I+SEnj8uayVuOOw9w1ga/PpfV19xvVrIT5xJz25sKbDIErqm1
0Xe331eB91ZKh+5NYhfL4I/iJBhhRu5vO2iUFRzsenrnpAOvB74mAD2ZAkhIfZZH
M7ljTDI/0pqDL08OHxm3KP0ozRD+2nz4fyAvGLHDGxoeI8LrcFLJOOVyoKhHsWpX
CTZZhwZun3QBqxP7sJBsInUCERInAAmyUk8366dPMnv+disa6APz8D051ro/rdwy
qmRW/MaoXtdI0nDNcbfCD5y8uSxUQNDuqgNsPX4mCxzabA7OD/9MnH5LT+PNLyso
lQsgd/gSOA8TgJvrBrmtaJCsEURCxQnfGmECB7+nnCPICX+ozlPzecxh2WQKJ+VI
bsZA3J38xrJFtHlVdthVttvf0HhnuQpu3LiD/g01qJ4s43UuUIv4T0TvasR6R7iE
a+TATLIOVFoWX7MrRHvbsmsFw2C+ycPiF8Rvv11R/nzJ8sSLLnjX6SEakM2A0bAu
m/lB4XFQsVbgQWq1zU4buzeoIKpdPmnB6T2LHn45hONJfW4oYXeFw2SnG3U6c0bk
YUyQ//9wvrxdSKoYuRih/V76SRL0GR5RRxoztK7x4mm95TjgC88MNTqpPNCCWSKw
/aFcOEdRrc13pZZlW7fjgpo8/1owNmxEPZvausHJilgOeb6mbVlahEKY1imBJxWj
VCVUx9aP+YpivPT6UpDvPFGn/bNWaxhNBZxY4F46WMiw2E4CRsFP8ZYBa/xdvcwV
ybZUXEWAFPIIXJQPgGTvMXei3AYY2zXaATdXRi2Cth3WNaWemTlvHiz9s1yci2t4
6XmGS4zmyW7/huhd86OU6m7okUrdeMinbuD3fDy2yFAnBCDsyRBRz4KgLjBTjcVr
XJY/0W/v6BI0+YOfyBZMYXlmkuLqjv/aFI4YjYe/ucU3h7VTwIWamBo/9O5IKWxF
kO6LX/2n/wDc80BMd/fkBXdkYRikVCkh6A7KtwVoTRvf49nxvDJ7geQRbKplAaZB
+Aynule34V5KSN3yQ/tYSZ7P6tS4fzlJYkKIBJVIFP+iqzpdbXeVhWVtQH5j1mGg
lqC4AuXPqkNru0IJJZ6SyULMSLFRLGcSbFDKRQGVQRT/0rz2mO4T6dtfe2uExqlN
qY2dPnA0JV81fs+O7F3S9LyTo/1xmKjEA0o2MdbTqaKtWbnVBaUbNkGmb62QNS2P
rCjyE79iBlftrprp76jktjCv+sKUtHmJZWr+lzWjtPPVjncoPjie+fqO0Hhj2Uhg
3KCqB6hOrKzgEuvZpixqCPM+AaM0crykXxo099WUXsUwO903eM5j6VAX8IF+bRff
ZqEvkWj1xPAnItZAi7uTwTh5U2mF+utFu6rRCepd16b7DKgt38mkbhe8cpUawVCJ
tDRdgqSOvI87+SOIyv6mwALJZuYR9iiR4RzQYdb5M0me45B9gWfBJwDHpOO6WKLj
qnDFJNBOHDYYwpoJnt1LRjtN576GSKF18kwdLBLB3uN4kINWWe0Ig851ew1kpvvY
lzXJKPmqCej88l3WZCE8khYtUGn1miKMVFa1co8GWTPVLL0junHtnT9IcDtWahV3
1KYHzgw3UNejOZlmJDoAjGp0ajdd/AcOFuI5nPuRRYLf8fAvaTSlt0Cyua3TfSPA
0Nf98pUOBG0nvUsdGhOB8LQodsp1PFvV0oo3GzG1yn1u1p3bC1wdj0Xs3r8jK0wp
MmBxDqKk6B8LUDfk98Uh86Tb62T8oPplwvIxoRQ/NH6g9q+THJ82KY84J+XdIhbC
WCJfbriYv4zB9n1eted5Oon0v2lRVXEdO8dg+SlVlgpmUBOShCSKT3jNXeNVxPNJ
4Gmfi7xt3B5hFXoXZ9LXub3QTnISo98hmpRqYJiZeXTLzwpK7bNXyUAPzZUFlY42
lf1snmhOBe3E+x52zLB2vDfYE4zHK5cAN+n7ywJZgif1N38k2u8qoIhYQ/nzcuy8
8X8whGMtb2AnurzHPIuj7Owuwf1LE2jui+hkrOn1UVNZvRh1aG6Lz35WKGtFOSSo
/UP6gjohEFBXRAvb7eQyNElaZ1SOdcCgI9rhqNQ6hs33RO5zopBhXx8TvVwcprGz
9+Vw2ILew9I8lj/vtaLB9wPAqmZEmLJ5/5DU3N3/rHhUyzT5DiVHttvzTyHTh+n/
xrv7vD53haryRtUOeKK609HQ4bA/ifouBRbmHnyDowmqRf69P56NJEfiXOV6SAvl
4+XtKf+V5vp5E4xszdneRGkWjOUEVKUNa1qJt0PM7cM8YXZ1733sQaQxZumgfPhD
6AV72jIsuppSrZc15U/YDEMKY3SFj+OQfblHlLucsj5gEoBMjHHTitX/hIQKYn+e
BI/iY34VVWVVN5Xjc7M54KorcW6cFErwUAIDlDt3cBjjcVRYE41cC0EnH0RlOfH0
PCsICNGxCGTrhwhdDM2FH5CZ7PHnRF37J6zyih8nKcIegcEGqGmEXQjgn/HyWWaW
/R8CyS9cTvQZyGVhjdc8UVupqnU1R8WSICLMyVRAGt89+JL9YtqqmYIt/hQhoY/9
g2eDOdtUqqKveSrMvEUqqzKSbTer8/SeEryllheduygbhHvBWxoPAUpjU/t8Sqb3
8hul7nJFGdr2yqrDXxcQFsLw4Y4Kg9nu6RPwSIi5OJXm7XYU9ax4Eco59yw3B5Fd
z+4PLwHaY1u9wvuenGqnXKG3ue4HVsOymAEo9gy+xQ+N1t47+1vUEmfrzPiKqNEC
kY8+80iKmo0/8vex2b0JlLKC7IsbzX/I8gQb/STV3ELeX+rwjDyfNsjBiXTSMT/9
7r2OXw04xyD4K3l20vV1uq2XLKrXFgkw3Ae9KVd/meNYPwyS1FeTkRuRZEhNt+oJ
Js0d8RPxrlEy5QUi99ByYHf+wdwgAlQez15f6XPPkxG+g5xEwkyzeFQTwB02022o
F9I3MvplKazSAxJq70YeAeVMVqvBoLBoN3XB5PPF6BCwtjrlwUVeWRHGmeajmt7D
bh7Gu4IpwsAW8mKtTgr5eqmHR15EHucOGVo0M3z1Uy7+11HFk6LZUBAnMNSWzYgK
EVBOQnxVFmvO7jVboH6QxokqKq2Avhfv8JU2w9yf4A94Q9JS/cxBnKylpdvwJ1V7
5AAcqJNhP7LozDjD3bZBJ9BDJ5kShg1AUyl3PgQ/z99rlVMYj9PuPQfRt/YCqsMG
AH4ZAK9V+LQYHOGkpFmHeocmeF2s2It2AOWrKeLbDZ5HIhhP91pc/QpmRol6bWAQ
r02l1U34NrnDmm6dJyRZEGM0QLTSQGpGuup3LvepysSOTovgULYdGLUm1S5e3wON
p4H97Gpmf5ZVsURoUdfELYgD09iQKpa4iPxGZih0dSfp6/l8NEp5Ripc3LjqnFYh
/UYirWvUclhV5Ch6vLjOOuUTxSlK0HsnLzuxISTki36ZGghgIfyntmFcVnp4V6G3
bbBx21ibZD5yRjAdusWwoOPKU4LIWTbreA+yifcSOGO1uTbR8qZXqlRf0VlHvZZu
5PdJVfmcJYLvaFTTiy6R/wfCJ8cK1hhxNX3/OBwH59ZwtILiqgcmXWa+nlU+LUFe
Yu081HWlwnrdVg/0AGR8me436gVet6WCrf4BzJ7N8XgoZq6Tf/Aly5l8852G6Vf0
sOHiUfpMrttEU4BjM0mwXjLMN7UqPhNIojW4D1fGnylCcsFpuQDb0eHsJLvkxSvg
nrDSZBtdeRLRJwKTSER7TjkYtN7oolOo8ncIrdLf8p9E4McLQ20znr9zuTAoVU8s
Qzz0HJlOVbgg8ELiXiKxlJioimoO4stn11DMiUqR3qLLPYGZ9zp8p94PW1GGvDEI
FgzYbw2etEpMSbOK6tU5joH+0+aE4QBAChSz6/iqIjBJ7Jlu1QvY7QOCONspbLn+
gS9tS/TxXvW0qwNZxhgo6laXu4qrkzXXT9OFDz/BVOPi2RQhjBuS8+aI1dScPR5/
A5jHxbASz0yT4mrNibOTjNYsT9cyfOHJN9Zo5QZOx0Kgl1yK/zvLFe0fuyNfMy/J
bqCvtsGNDe1jm3Lt6mJeG3H0bWZvjHYhS0xOnRQNrH/KRk+V+kuJlT2v7pxJp6HH
g7i2qsqn0PWpotgIWR997HFnwMIu9UNaSLhHFy3x+u+6tmKJxW+bzGhvMCoS0yjr
N/j6rXN+tQoLtXQm6OwY9KSE2zQ3k/2DIh0/6CJpXZYua5i2Rwmdnscb5XlbWzSw
FnnXBJxH4+gClg8mD8RBO0Qy+Vo2Mg5llheNTN4C7hY1DY54CYbUDiGPXMX9zGJr
X3xJB0jWZ0PBySzADBqfWGjC5pnML0QJo3qAkFRyThQgX1oNgj2cWzmG+6goml/c
pNTZpg9dJsKuu60p78hZYjagtgjNGVBeSDfakbCuaalJIAZdSoPaDT7rwUqCOLDB
TV9OgmU05XtZxoIRRKDOGssc32KHQnHo8qCzIYklFXBq+gH/D489DOhku4qSpGSt
AtacdUU/HnUaGi4I7iYwySQa87T3dv7oso1oO3D5XuRrXpEw1zl5wtx50wiQQ35t
xBmYULJ5+5YkUMLwIyhdyCjmYm5H3l1qP4viFoY1FyRo/jKLkqcbimHzWqjVbCWb
f9XC2Cet4Svh2Pakg8JvHq/bmPAdspjxHH2c0yzwUNJxOhASjUsG8cFGM1yW1m4C
NJXWTSjhg/i1ZI6H46XFYX6qMXpANHj5Aa+wfI1PGViw5dSEL43arD6Lz6gneXIK
VAHgj54xnaIwobOxBUhmygxom2p+ypxBJ0qOMm/KSW24nt8d0clJBGYggJQJEaA6
j7x+kak1t3d7QdyjMRsBkJHd9TI9C5x4i6XrDCsucoEu7ePVs0txaOw9PsCmv3zY
omVj2SHFJvfy1XKgulIwoQEcYFsW2rsifAUpYvLeyTJJUKX2src6W9u6prDCB8jt
0fRltivXo1PLAg6LybsRq0zS1qZC98Xs0Ar2r+RWnBKBeiLqPlmTdSw/smTud9H2
g/7dIl+mH2ikCVTC4XWmRxwZDrJ/EvMqRmSlgeMbV71GaGp8HIjrZG+O+qr8sIdU
yRunLnE253X+mZqJPMJp6b9x1KUPi3SenmGk1sZcy7bcmVpeUsIL8Y5XuqM4yn9w
za8QO4fT5SEpAlJRUlrQakG62Eb1C6QsFrrroaEZuD21+jqEqjXtgZROdga+lMq4
j0qEnMUi7kfrCghD7fetvXXneMA9H2ngz4bbzki886ya1qb8dZRsHTVt3OVkphHS
h22OIG8S4YluYhZHc4S2T23Q/zgB6tW+qHmGkd67wBy1cC2lz2R/hrM3sDX/JOcB
boEpGIhQkDWp2M9ZLpsQoyesx6Sg4fBiR9EZpgMaipm89BwOv1LC4VmXIuU7VEQy
y1kzcbkSLb6PS2NKifsqj+1V4/mq1pr5kSX5R/lgaLMoJb5EAvAEQqUL3x4/8WUi
5wZIYvFo9Grg4kVxQFXsbiI+rOBmtIcWCPWGSIGQg6+l5i6MlBEB8c4kFV4dx15q
Gj+oFfmz4dpfCeFHKmOqDZcWs3jLsaMqIz8dQWWZDHNSSSkOna7+4LA/2kUBMX5I
lkU2JRTYkGFc8HXy6yyFIiInKPzF8YJ2nx51WMF+PfoM8DwxdMwpvU/V002dA/Pp
y6jOrkswYB9h+d9abyy4ap8cop4Pb9pycA6/5z2ooFKVbH/bjZHTnrCCxdHm0Khx
/JZQ14yuOsxc7R+9h5QfaBX/Fj/VR0CTyKTsHT8xfnJZlldZSY88g8EkGQlirK/k
8HAI8hD1A+KYHAXjWRTNmSwSNDnMduu5fVmnsLNvKW2jMaaE2zHtbODaqem1/58J
xBMsDeF191CATPY4zcjABi2yccBsimx9QWV+zj1xVnZmtUmJLYP7f3PHJECPwfb9
q0YYbL/ndXPCJpJPPi1XzG/pxPC33iKCWWF7U7JLZ+QVsv/EWH0cT2dA26cArvb2
M8mOMfz5VnnuJK6Ni9+ih/M9ITMmz0UY60G7ETFF1GMTrZRmQ1MPo9jxJXAhO6uo
saxFvFR9uJmcB9VHCUUnOUC2p4sUF6H0h7qceNgYkbjTSaJwHKfEhsg5j3qc2USu
Ux1VEe5StTK/fUCl38VggekxCStiZmvL0LRddozuKLAq09K0UCzAOStwC/6U2RI3
+yOWrkKONYalVXBUEqyfDJ57rpPec2mhvcGhb3YBMAQskLtvsXR9wNgvuGgtM0dE
feAdgs3paBLs3qA/RgcsQNGdiDn+MA9EJaBH/umWzebRe+7LF5yB0p6CV6OQZdTG
s6ysmHORkuxnIZqh9j2kR9DVN1Yvgl1ANBhiPYHwJbMlQcrur4W0Q+YheUUutBcd
m0hthNpbonAg10hcJWXm2zSfF3aNdvTAa4CSyfOZHYCZfGZNOFkWRIsLKJqXEvYm
QB6TpAoMl3qFGWqbfjR/G8ufDLkUMfyJiQ6lUxVdy3DlVYXKv2lit0Nzh5ddB3oO
7Qth7XJD0kolTSdNqE/auuU7x8T2x6xWH01WgHUbOmK3tl4Tow4zSvd7HUNQauxD
GCTGChFsNsyr9RJuEaKHX/nsuqIrXhDK2Y+kxIcImWSxvmwnFuQb6j28SX0VTTaV
P+qnkj5D3o6hax1Qnrek5uUsFMXUtemGzDzMNZkC5Pi6/Bitsuhh6HzHUUGWbkpv
2uSofy5ZQdyyI+KguhA8HAgu6Kia1CYBjtsbeny02L4XMC7D2hUBJ30qkiwpFoII
YCVHED4qKrM6d0heR51sL5bTgX5ggdI/JMurSkMG1hUVcxk0bvXPaQ9bLBgM5pbL
9mHzbDa3wwnixuJvJieh2B/t8QggFTEGPP36PmCuPiQ0LmE6GZG/QMQkD1H+zh4f
3ZFxVXTCv56r96HnlzKALiZLqdqjjVZzjppX5zJD4L2xcKiW3tP+kUj89uuImdGV
imebuSiMmF7m3DR46fX6tPyNNvABH432lyoAGtVt9hwh3ZBR1/tqP6gS+O8iL1ws
UkWCRjtk/bo3vKeAacy4qUHj6ps/izPQgYzp74kjgIarWDsVEmswZIFogqaip82y
ELkozU3XhZapOI0exKnD8wB7Q0d0GiTRcq91Y25DI+7YsGNTtaASle+kiRaaEl7s
Axxfq/69vgeGXEQ0uF0G6+t9mg4jNUArhaqnrJhHymCepxEBEKq7xUNEms/P7gRG
DHC/T635TOU8+aLwQMFpq/HankHwFq3lcDfWL5AwvHgYS8dffI/2pCvcVhd8NoPT
/Jzrn6IIjKzz1y0I5P2czSpdRFcsR5BNZAgkXBzjeymdzznDV01AUUAxxw0D1Eey
3UD3mgNfCmduv2NqL3Qij1S5xJUxfSD2YcgzJIXKZn5Sefssl6WkJpfcmsN6cLzi
CJ5GQeO1SOFFURFdM32GjqW+9GbVshJxvMo/x46wyHMMsQI2Q8A4H5M/ujVErW9x
x+Zab5MxL3Rz46ID+Ud/b/cQVZGi+y2SYa2T4rck7Mm5X/FXOblPXuM2SdLXCZI+
wf73rxL/dAv6f797w6aaGZG5vzG6yHU7VW1lhos6jfEypAYLorRgwZTAxH0FKMcF
bg8C1uZNL+MY1CaT4U7YiXfYWQsCAs5z0lHkNASW5hPxoOi0bHncl6i9lV9VB+d8
RiUXpvZMc3PCD4U3AVv0BvaBw1/vxWeWYb8UEdEQIDKBC1fJ9nHfnpCJHk4fgyv1
Ty8564OWoUDhzRdkVKNxQnUKw1abgnuDRXLNVocUGh2ivIIVLJhBcY+uIwGIH3kf
By3OwZ+2A9h1QWCZtlzvRr7InoylWaeGwT4UgR15xummMgzsNCKQbL54UkOqcJp6
cCBrVZz5Cm9FA3juZW5GfWejS+MPlb5X553pKolbVMtNe7d6+K4JrUCUYyZoTq0Y
CXrhM3iHDzzFNvlZbqnjRiV3s078w7CDIprQFN5pwkKtDihbSwBilQGgJAdS2gYH
S6WBafuf+ZKzYVjLV9iSaEH8Ia4+Zdut5lVKWg/bqwUcl1Iizw/F22Q1EoKyNMw2
H41U5+PNyWCV5OtYy0m7xJqN1pzFG7gr6+dV8OhjJdF+nfrUvlhR7LCamL9AAlSK
a4EBapgwtQKge69a3iopHU9mn2O0kg93Y969UtJcKAW0IZ/Evj9IyChWmd1II6Ie
51iXeGqta8XPWWifbGniD/NpBqYNa0z/NygGrqdvgkHHfUw5Z2UpG3Xqzf2HpIkb
VBe2WMr7ueeFOvPeAi5FcjNqUMdiyZeZhi5yERzecDERt3at8Hp1AvHTEhuLkdPJ
K7z1DpkFT7DLgRcf/wSzZB4EBIw33pFcuRDENnpoN7+yzpMg4ruCfmSHvP8cL12x
dIH5/pXq3DZmU2KTEgjTbMfFLij3Pc31pXLbmEiZdXJwC2aRcgKxqOPwGvigi8Ao
ItrBZDGm1yfwneqqwdIaVL2RbIHDnZ24OkJpGPcHmvz1A/2+uJix/3A90o1jiZjr
Oi/GbyfKDIF0iusY0PIRdIMZdB6RDronp1jfYec+OJI6STx0/hnf42NBNW0/74em
6hFpN/YUNvNPcFRbUDUw2JLTO54rpJ8BGNFU24nEy9pyZv8oRLYwGbQfA4eUn7e1
0kJzR2zeEOwSQnN2IN70B9vrpF5Uq24R2DzinHRYKU3Ut3tJ6yCHRT9fQ0nnZ7rr
oPoZo/SJ8goZAzMpHj7M9Sh8AlXzJdp0rQ6UqaJJPyhEyWtjc/TtelEuL5IoS7zh
MvhaM2yHu5iSNt0+nBuV8WuAU3b8R8mSUM1JvksIQYDSuOJtFBXL0Cshv7ena3sZ
n16VXPjuWr99wVB9GGt7sb+VdD5Q0Lf8h++8FEP/j4MaI5h8HbWPHsCZWDdHefbC
MztR7EQRd4OVt5SXw3ak4CRtNxWSFgtngLoUxcb+TnNWUZFKIaarVR6OUfQhUve0
rygsVxi1f0iwnejwrKe6gy70mQ9GuFTyo68sf/03sTV+Xd850MeabTvBurDTiCi5
RdB7a2HhbdIAKGCvAOvNtHu95QkI7d8lUk6ehda7P2APYNoJN6u58Kyc/yl7maUr
Ob7oh6O+bKUMg1W3P+60EYitcPleuI2Q6f4m/i1bxTdWtSHinY63JphTBOYn8VB7
gaXjaj3agl6bXYwcPCML+mj2rmrpmQFHvb6rqUYQ98c4uLAPcF+DdiM9N6CVj73+
tSEh1tef9XMwdE3zT0NAn2qXnM5NCnPUhTvg/ehvs2cZk5MknOwsz7ojupK6OW5i
Bpq+NuXPOQvhqqY1waDiMhGKPMF/Mc0g8KMcrZZKHI18uvAaGW/y4pxiZLKZ+ima
horP/iTMAEOWABznVwGtASChMTMIFF9V8jY6Wxe8KaILC61NvsaqWXcgVR4zmaAq
QiyuRbrBZlbaR4ifWnkCGQ+Df9N8Ncv8wCoewujewlkj189SzhdvG/AQ0U21C0wn
8LjMKomGRDOBhvs8GKtesK5tXBqP1Ovg7Yh65OTX9R9I1RMMCifpxffiygPIu176
uoTatc3UGOyTmX6wlvUiLteIQEksHJ6wpquzvEnMN1GIE+m8jhX053AYKVOxR9+U
ZYlNO2d4lz2Z89oQNgZqhsm/yFublaNRfNLJOMjtvw9odDtLrt7VmIQJrHbcm2nT
FAQ9FKEqkHQbcvIY8xWuoTlFcM1DgIpeB1wwsnoESsMGZh7OD+WAqQbCWRzd+f66
c4mYFdUGVtseSLY+Vu1u4cIGSgPYddC1YQYnv/QJPxboQGJs9kuGdhZmL3/wHXLW
+DnTm+Kh9OuUZdAxWWkOTsJvMhX5qrOfBw1J5GuFaNapImGZszDa+5/r1F4JwIj7
ZDNUZ2Jq2rH3q8EEOPerVmaiGGW/r4+5mMfawux/ct6NWP+jAW3ZNTKyhh7zQewJ
Cxf00gARyhiwtTlwxBFc1GMcGNJSK15n0ldRUeEu8qbRTiSW8oCQhhoHwnZoFuGY
B0f9QltQA81BC3KAgBNaRuQyjfnBlR+rHQRCSpDo01hEJhleHEq63V03VixDYTJD
NpB0ZrnajK/X6O9ULQ8tKuwR5f50QiYItu2zps2AQTS+iJOF+m+vO9a1vh/qdGbH
NUiVYD0bykaEIHVkzf1qUpVsO+WlhHFGJULvMDWyWnl+A809npbfRTueh20oF7/Q
+nEtCV9jkJjdS4eZ/humnVRcXdww53iGfzSU6MN6qZvg2izekIO1ZcFbBdQwJsFJ
+SNGA96WfCXqBHbv9zrLBc+61EFhrjzOOjZXCkvFQ1n1Yj7vGW3LnppxOEO+0Q8z
QhxW+d7WIGF1mJCaFFsjGXvq1d70q4DCZl4tzNXD4P1OEKrVejajaYCiJSr289PC
q/wd2gFNd7XuX8M5Z9Zrlot6dTkXfYQyXtAJp1pYWCLE7Mk0uYAC/nmMAx4+0eDF
rkIlo1U2PXRBcBpstPq+oHCOYDBecB6iMtGwA4Dr7AouIpMOUBODofq3aC6pqRhe
R1GyjWaEaSzvZGhE+ikVyoRvj1VmPpZ+5YiQe+Fpk8PmKoqC2ujn12uZE9uM7SfK
Zn5r7vgCVwUf84eZqmACSxPQki3SWFaJO+gDyQd2RKJfmCByXRWnXVnlwV0fPwN+
rtcWcVFRGfWQCTksjhJ0+RYOR18SFo+hmXwzIJmpeLUA50OKm4QYogMcUErHF8CJ
y23ti3+EAN3grDTMRVAa3HaIJo3AJXjp0lLREChUsRQYtpoj+ZQORwqb22jS15OR
Ip4AyLxhn1CGZ6Mc6zPpedAgFEPMiUTwguvz17SOoZ6SIPaW8CT6fUA9L/t9gqEk
F/S1Okdx11XDKK5MjHh7GTE7F7Kqv+++1JKeNiq7TlzyIaiOxRBf0fynfYA7F/wT
bPGz5F5VIYH9ezyDUaeLQRVigHN+9FCqVyH+bjueDz7zWODqN7i9zp9BqwdPhkOP
iPbBRRfaIiijHNSPBssmKTIYbzrQ2Ft4kyyE0gxSM3s6oImdaiyhOhomkte4+0OW
zKGOfcAgPxhFnnREr42YMpO4gLdPROXhhMqkqmA3K9EfF7LL66lDi18zs2saQ3d3
KoQDPUn/0/uiK+jJPWo6qcP/yqIGKf+BaTfy3vTxpupYxCY0iKHNyYeozqUUhSCK
mKs7pQVY/pLqXNxBvyONpcAPxIuXLixHlnLYaSuF2TbOsaQBJVmV+TF/2cT2qvbP
Vxl07EE48mMTIXe1fRzmnVJLPifcVEk7/47y92WYqirv0126a4mlojEbTudtwYrL
Xt81r1WzlKLRqAU9VYcw7/R4uRD8uVbnQPyXmgj4bgxVJAscCLXqQ0AFYX4QKJZe
oqEArSttwXaAzYbPqDv8ek0Dw/eZ+UYSesKqSPs6MqsvWEVHZ+0fO6AO0eZnlBoF
NoydmntoSnVVvl0simrsxgD5j3qupVw79ltXxKJx3w/KuGurs9ggKH9eL3+l1T0I
JEEa0Pt07z8ZU7R4Jg23P0R5myjzR0Z/z/b1oJMXIOBNNLt0YYIHR1reXexSfv4q
aSG0sE1mrPcC6Y/1Ak4bBnm9Ci8OFJm1trRHJ7ARyla1zR6YsHPuglq3ghfOtz+T
0NhMJLTvGPLjvW8b/jNIXGI/A7NR8oQ00C6lAe+gJsk1IcqtF397VoI8VFxL7ADJ
AArMgZB3l+LzefKfW5LYV8oOASii7XW6sRc79Izdo9zqp4viO9Q2VS5uHoAVYdxl
MM06rsa9dozhZQ7z20AvuKmzoJsSpyKTaUsby/J0hD5WAUtZ6CEjxGuC0QusdPQz
e2WAoaPA2SK5rzHN/ycQhxmr0GAX+oGAtYnj0xcoeDG6PEtFwsCrDTDNi/Qo9he+
D01UtsPrbA7plGGXAY4RqvGR2Oi5qp70PDVEzdjS65NEtjnLxZcgHY+luxt37A7U
fD5n7Hzc7Kc939qlYIM3UERVEXOytL5D6N1cxv2edn8IFmT8nvFm5JiuM09EIAvN
tq8L2+da0GpbjkFXpdfi0eR59O/9WMsCk6nJGxN1JkpmZeA3IdZyqWgnbmv9oZ+G
2ilQG3Jgop6Co+Cu7Cqn0evisvdZ0nvNdJbFP1E8Zvxu0Ml7YjLt2higjPmzSlXQ
YsMDWpI7uelCaL+mWxJ7/2UR8OSWuCTWHbNyfsW/uxas3gSDtFYzFfa8yngS+CKM
siHZzQ7aBlujyYk6HpjTqwMNrVCasOaFXi1MuYgs3DS4rkMqz1TaeRPKMKud6FIw
UnqCkPavwxpnkLhCaz3ABilxvn+Re/S7QnBt/qKH/eVfA8315LJn989TpZotFP/q
Rji3O291yXbiE7GT0k07lPyFRFGlENO6xWcSvIzSUcfSKlHtX13OgCRuwyXnvmT4
XBk/9Y0vZ4UMPcYAG4PO6RKZNYooEuw+le4bIern4lXyY5l2jYeEfLHJ7R+RD9kA
NP22KeL7nqZF7tybO4C21xDGrJyrah/QEgeyBFi6tQClmqZEi42eT7E1MkDxiv8y
amh4i7Q5yxYl3M8OBsuLUmO5LjuD9tMto6H/gQQTafH8t+C/KciLroKY9zk3vwgC
uHIpR98tdjRcTUgGFp8oagYEEBUJjJkBu46MrTpbCZF92h3Q2eRPi/Mf8uVDtf2D
DWXu6gi6JGZKNG+RvEi07HZ18EUrw/jN3Rtl6Bye2mQxTlyflAd9glL6sy/BEMTS
dVInzUEx36pVs8U/MqR1uY+ebTFt9SJQOIAXoEFX5x+lRc+k9ieNPwJWI1Wrjycc
NsRly7Bg8asHrWiusHQ9RYDEfmAsxxP+0j3eoL9e+4ErRiEbrixMBsEkE7RMx9cj
vxTEFb+uUBcVjXS5/5tbBoXCajfZavh9moEF+CcsX9aYAm63euu6fNWlUEPt+y2I
UM06ZxEYazQJiMXPmnXknnEAk7PToUzQQU6oLeUwRKruTeYJMoWxNpTPvhg60qDc
Xad0Bg/DRpHX/psrHsW4aFf4b8jHhStI9/SzNCExeh/5oK78ocO2Rsicc7XNT+WM
m7Vwt5SV2N6vmchH8bj1fKyagym2VZmpte8Xv6MNFn1d11nGACFmBQ7o6QCfA2sD
DX+LqADUI+WyjbGsWN129w9be7T6thd2oSY2zEILE6vF1Gpkn2Y9TL8X4Lgx5M7G
3fqGNsnWEKxg9JqTDCZAQHy1mbjqZljE9SqrM8PuiQbMVi5Ep1ecpqQZy5Tq2/YM
bBucKtRHCcOe4KZmHiOxYpKOUy1ZEGQRJ5k29+VJuT9+mgHbc/zqUJXjFIwnrmI+
C7yApVjzRcf6tiumzJIYKZozTGV5gij2XD2fV+wRWhhJloqHnOa//4JGDIZ98eLr
RDmnNcgqPYUCYx7+5ZB78xj+46it7WshLs/fIacWXSUsUbDswVnfqR/ftPDPl6QL
tL1dp/xhOhQrIni9voG6KYc1/zYnCvMiadeKwESQnZKlM4BC4XbRDsCO+gOsbVbD
CFdVxKI8rMHP9rTnQA5f+LN22pJlI/sZv7eia17DX8YGNmpQYpdQIxgJEAQ59FXd
ciYavnIWaF4aoeB/I9QrcLs0i5siINxREb6oSXy5pddknS+2/j8lbOdfNsAUXr5M
g/mtBOzxN5yEIlnhh+S3FLqJ7DEdPDWP945EvrGo+N32IoM6GiMzIqiADLmzV95+
9KjQXCs+ED54VC22ORDIslt2xXWbJLjMxL2lOWIucsa4LGmpD7GlB9Xagp7vK65B
bz+YM9B38mEnKgRS4Y9+gedFJm7xjfPxC4CJpE/YKgBB+wvwHxvnzCWRjdqwxA25
RRY2I6AC2Efd/B78oYMzphPjWvfp5JZbeE9Zn1dUwAdls29l5xNCBDfKrL+lFSs9
N8LFLd1coCfaLvkRL61j5acXRs8+rX0ZwywnJdcwo7mKuaElzYoCL4WXrV8A/rZt
adF3Za73IOqPg6Yx0N1Ez/DAmc5nurYX1/G5Wz0SzL3WDJcSgQdiM7ZVM/nNMvHf
r4RDxwL8C9OqNJG/7RZzSdI7o6jqSEZ/mBKJhk0jwvOm/m9Y4BDMzGPQoJxpGx+z
8HWiSD16oKGoXs0pjENpVfK0rWZ623UTc9mUzX8pDfvDKOA7hsSsM1j9MZP98iEG
z56gZdwYcP63hnljrFhrzO+BqFn4AR4r+beP30lmBQQGnTw613F2EOxC0e8kn7Op
eN0nrzX14oGYOA35xtUgokahMReWR5q62uH2ErJRKuHWpDqSIeovB8t/cFVq23LQ
5XnBxh7fVccLcyc2U/I4BI7Mt9XttjuauuZtxnpkzptr3AHCcWODKxztEbNeI4UZ
oDA2fsrOxLzMdeDY1yr+d//0KNGAplaesScRHJ4O8J3cxfrIBdZ7SKRcJD1qJ3Vc
7vNaMPSE3mx8F2LybSNe10GNdwu2ZuhQKI1K4GUP6ZxbGnlwOuP0hAaY0i6zSa/L
DwsGQ94gZGldh6tNsaOCg5tviryj5OZg8BHJDKrTWLS7T7YOPmW7RqKkDx9RfWby
NaPB704bOnoFyyGkULv+ZbRDbsdepXXQ1+mfJjHKQ8F7q6wM3SKow9b6b7gbxuER
GDNJai0M6Gsb+Q5+I82YODc+SC3Oah8r732XwZBhsD3D0Z28b5EbXeVwPjAB+82F
YiPGcZ2opTobLygzcpHxNmjIWB81nUTadF3WQZPrbfeWlgJsGJE9gvBK5Ahymszc
k6qRcrbQDUEAq3r8xZAx660ySIJniLMgTYT/t9jRIE9HQjw9rNJlfBDB1I0yO1WA
1m/zI9VWANiSQ/7pcvg4wn+V38JBkOMYW3LYue92yOMM3rtG1ck9andlw4qmks5D
YPOyh4JSIZLVTtSO+umYg2n4afWRFtqHdOlVbbX5eZiVIvQ7imS60An5TJS/udlr
qE9VMVlXvBo+yzai86Q76R/iynCFvUtntTACookRT7SPfZTvxtjASbXIPpeejUuJ
AerYXapzZmiYzO7LbyvrS8lPlBpwEVf6XaphDF5w0K4cwiNlJB3ufrmaBan4kedA
hMunwtqNGYKkXwAjBljBRg+vn5qBZVekgxEbPuTk61OZKz7s4ChxlpOeqt90wXgF
FCe2nzBmZLETwaNrO9cARsksYp+nuw71fiMTqWY0zGBKLgf6NQM1YUj1VFRkJqtx
kj0StCpeaSYO4kLprxlyz2kjxWWsEDLYiHpnGuzF32Pd2iiWGT2ZPGtlvydWaO+u
dNdblw94XN7WfDAQggOIf9+msSCBXxS5n6A7GOSd38K/paVoIRbh6QXPl9D/75pR
sp+1bR3wNi0UJqYR/O7rWaCIspVs5yGoTwZgg0vWP6GV4AdcbBeQSPNToaJFUKuS
nE2Xi5/+L1dWxzlPMwRMncuJftvgnfzUdGrFPu+96/WIssUvOMxoy6PicNLVZzkt
twkrKi9zMf8ZWZ/LNl9zjd7TV4ARUvd9ldzw1xcgGNGqvVPdysiLDqsehq3aZeZP
fq4HJexe6mrOFW1DLM6mqEh0MCIr+zlmIX/uPnHOyhOn5792/aZLrKk128iRUNuV
TaBrie1jBEdOP9nVWVa9cM1UyyVCCJ428P+P087FBVVtr0/Byp4hTFIfvFiWLI6P
l+TsmLEkM/zLviuxytYVxF1z6DKJjtjUdSo2loRxRFP/Tb9MtJDwrzLAKgngdDrU
DtrSoRQr20kplpJKh91qfUs3ltu8aOOpnX/LfTQWWcv5b0q6imuB+xpnI9JFn6I1
2GMolbaFDl9kkNonr6zQTOQATJMyipgAb7QVUTG5w5nNdoHb8q9mQFcLg20UrSnd
A4JL4bPxA6rb85DgaWKzJhL8mi+SKmjij9gEEZCoWp7pmDvs8toSYAoWguBqCvTz
k32LfwPptazJiuT4nE66+lLnMj4sTssMpXieO1EgUuf2Tw6w/6GyV/q1GPJe0M7T
QJ+C9Nx2DMqZH3mxf/0Jsul1kIEPg6QcsLCg+O0354/2mw6UC1ApxDhWwwQqS4tV
x7cUJbrdjpbZvWkKBKRPJ4gu67NF/26SlRa4COyHxR3h1nR7ewm1DDheUfL6hZUu
TiIMtxhrDgtdn290arssD/1/BTLrUKuTAc7gXnsyagqnZ0hi/S9/xIdwl1er1ety
NE45w2dTnFef0XGXNyKLl+hWqcDN9+P7alLCVWymSG7xt37KWe3/zk1yoSX0DQ/N
Br4kOg9xFGfUjMY8zT2WhjD1XacFfjaXS5EOy62IqkranC/QpNdK7o4tJaglpBvo
DKHbH/ILkwJm7JImTqgs+EA07F5tGcyUVacw+S5wnVMqsT+1K9xInoEN8druFEe8
SqJGqTNYBOs7+09DbkbMdCvD3/IYZ/8Sam6tH9EMxfTYHZ3hzmT638n6wBsyC5nt
66zwetSkqbqZtLnhwF22d6pXhJ0dkIpBUEUH4/5h8qC1z/PE/Mr6x7TqJSVNkIKa
7sN9a5HPPamI4sYCPqSnz8o+ApPPptdpC7XKSsVz2woTTn5hE92kM6pAQXQDtFr+
wX36JYaXHKmukZsalBSiQ8svaHIdJDtCxzNw5kMiSwJt8nIpwPmlmRMWHZZTaXAt
uIhsT7KTbogrm317sEuY4KqKX7bPN8ZjrUVQyUCQnegxNyeiUuRjWfkq/zTROUCU
uxsjGamppoD8EQHUBhnbO4/wQbBaM9gbWXPawKj4kvgHBg+K9qzpBkmrzkFTqbSH
ddULSsqsrJi/xkGS7nhGMfpbIKEY40fc9AmGFs824fFn6mCksxYEjzN3ijCZ3Wij
XQpK6lcrPs22ns/SuIO4p1HK2fBFTBTffwBEPFTknVRwBUSkv19oZP/+vBgtPfPa
diU+F/jUoznxqUqoiKdl/kkg9uJGv3mToMoi1xMX1rStbZuwplIz52P0wbWsr5bv
4LJTmessMSw93u3wEUu5E3gy+A9SHK9a7v6t7419MMYLG2lAPB6cPSOigYev9AWr
d+2Cay2APhpIrpSwenCd0wqsbxmrXyzW9qsCDKjoYXAb1773XW3niB4XrdB7DZ9d
DKcoKY4Io6lmyFPID8qgM9twSet9HcluNkb0SNQ2zU+pLNENpay1K03qbsMv9cVt
5FW1qqF5lE3+I5a4CWnd9709WnAM3OnDDySRMpARkBdwJoyb8Q3ao2dPW59e+1vr
cTmTEhjxO6Cu6QejitRsGxQm/oth2W7XKv12OkKBtveU+xUQNDDRYA2BQGdq6k9I
AkMjTlYsv4CoSfyiFcBozE3pIhDnMijQygyqfT/t/Db6kvTcG53OAqFWpsb8Ufzp
uwNqToBGFl7ohHNpIHcwKmS7/phzsL1B1FY6DN8m/8mkINh72y91zzf4isYaPkBh
hgXXZQk2w9araueF/PRfZxHx/gOogKpRK5fluIsmHiQITn3JFmXTEZ+7qKs0S2xe
jJy3jpNTKReM5241UrMWISdXKumIUZqgO+RQ+eFbEx8De9p+U549c8AzMmMc2fEI
nqXV+SBSAYpJydyh5BbaSKLpavBpXS7Q1C0LlWgBVxou1toUJDyz2lC4nWd6rk+N
y8ngBW7aRhukY6Bi7IFebbN12wueYiTnnYjFPuWhFDPsrBJGqbFHd1gAPWfz13lO
m1/2uVu9pwEDl8Z8JSbgoOm0PZ3bov2bXeEXjpRsUuFNEd9h0ukFN0ddBmR2FEpS
NrSwwLP8D9OfeS5lQb2Tc4DULxJMSUk77tssqkAfFajKQ9AOfnQtGlk29Bma7Bz0
9aXVvR4jUn/sYkZqjE9G6oMcRVjOXv2Rcvnyr8Emx8ql2C8Zk3VeVzqQk5PQMKam
qclVV136x4fVHTDlbaoTTJ+FBJioHXrx8ZfWQW7lduPGA0KWo9YmOf+eZei65Hw3
1KZ/Akffr4BtA3HcJyM2PzSS1PIOL3+2GNe7lFItbto9OQc7muCZNLrcN+r4vRwQ
f0H+qlWRat/k4e1Y9Q+lJjz3mHzU16Ome22bfTwXOsaRbBmsyyh7lauwRJdLNcws
/cHxkZ0LVM6KDRW+DADCCvTMjPRAQySPfYZjUOAMzoBKjbJuPwjSGnlZ8qj5hNzU
tuqJ+8QTf+y25AG5jKn4kHrVPoi/JQVNTwnn4tMzyYt8NgU6dPhN1hMWi4fIeGwZ
OFWikwOqpgKr656FmFcDEU8L8M30rCvrWwTC4+QbUDB9cia/vNeQ4SB6FXxRsvwW
nRRWyxjpNh7pC0R0hInxlpOVB8GcWJyLuXC4O44jDkddlzveMwkoamv2XrodALOv
xrTHT27IqRvPVCeenPn3G7Ox8mn5pO/EonxSARYZS1nkTYAJvxyx7dYbE4tjprW+
x9XdCjIr7nDenqZk+ZKNC92tksU5dWtz4SfEMOz59QeqYRueiVu184ER2wJ/6ZBE
FPGj68z9YMShtC3+AB9RlUOYcYMddiAstaPBFwvsA3hKiyoWdPEdZlxIY3h2rg3g
dJNez/MK7/9tQMN5EJubREQig5BmUCUTBHjNon2sygu1vFv7+4tVG3bic9JVoDCj
XOMTA94qRO4Nl7mN9ksaNqS5d6Qpp7V0Ej73f1Isss5KobjnAso0KAaMTPopUmQV
zX1vcn5wmH+EJCtz1nlRxY/cHYolVgF50RqsruO/RrCicNyFW8+jdGpNOyZxLUPQ
wmlH4ciqzdpElVDiDUXHkhku/ZyJUIRFG+yjgRzu9ht/CnOmCYmMUrivDK5tGLn+
By8wHcLjT1QogSM8e5OKVJ4oRDEFqiyFRp7S9PyZ7DR169Yl87UuA78TQGUiyyRf
9nFEI/OwqOJI3PM3JlpMqq1JVG3YNgu7jwKCBD72wshNWH79U1pQuSBPtYe7GPoK
xznIOxLqf+h97oZKRAhMggJ1HkMwp1yswqJPYva3kkFLK6fqblGIiESp197GMQhH
jR104gIDYSG38AayAIPmHaE6nlRDQL7CC492NK6/3XhSnZ/OgF/aWlhXfvCgBCqG
v7CRY3Re4wceEfbvswYbbBNH9irhwME1W/udgMEPg/9iwkBPoGhJP/kIuX5w/uxF
26aJv19l2x2OB1a+cZCN97FUS7cHml33dmgnUzlxj1Th/18QuASKSH6rF/2iCySG
EhwefxY+/qmQYtfcVXmQAJSP8WM6oQUt7shgg7cynZRNSoAeRH2b/T38axKxiFtv
NJXEzRzRIiuPGfMAOPMUz48szxaRrkEuhEp5OarMfVeeR585PWeFDexXtikOQaia
h4laAuWoQvidp6QytLy5pWmIBgimLfz+vD2m2hYMaRA5e39Sp9jP6EgL7k1pUn66
+k9eyNUp3kFm9PsXYiMipWkeq1QLg09r+gpFy4dZhVPh6PJH7o0OAjuJOrzVcK/0
cABNcBfn46bMzZrd4ijeIbGRWq0sV0O4zr1dKk76lT08nD+qhaIe6xSSgB+tYUWT
YG+9z2Zes0IY7ghrM1ZfvKdZYqFAjHDmALX4EAhpNb44KrF+/fwHiZJJfj9JEDJ5
CTIcNJb6gLk0tVyCL4vL9pRxl23mAtnCL1yy8tP8wTbL6oHiutfrpJqYzShaBlZJ
uA5XK0MNrCx5Uj5LSUf/XDg14BW0DVbuRGfVuOYNz5M10YT+6EdzXh2sxoIvZtEA
5tA5IM0bHhaWCctGVF7IQ1zEgxfbnls7/bF+5P9sROctmQtKoQQesLC7TC8ehN+V
brFbRIZoVZdRh4lw7liCowdsiC185wcB3FJ5N9xOqZD9klkCJqSOHOXsxKASc2Ru
JmEiWdodMjAwwvd2Yr+XiitEWqj/jETRaqzht6nGTLIWRpkrkk3xkolyAr+Fr6NZ
G7ZXxxTO9WVAKazdKkc3fTXeZhIl1f7MswITXgWUgLSQo0HrChmSHKFMAVJig2X0
rKA9axRw809ukxWd9YkAGIl9CBI00oE8q4X/dX3Wqlu+JNz6EK1phZOManAXdLUn
4QfG3deTJ/HQrhXNBrEugylBnmJFLPZJERGFe1qC0/EdKN2M/6ffzSAWn3rd1hQo
RC4RGC+vcKY9RR87q737T9y69q4vTMmeMP6hBhzMsAaYSIQPphTCmSSf6hqDsNtz
7XRauiNIi4Nu9t2tLD4XipGQRg92D0SVFAV1xJNWKOyBfhcH+ZkiaVqzYfCsLpsb
7INt1p7k6938cGSw0rGk0zqh7Tlo/eSq+g6XxZggk0noHWbn9bstWWnZZT8uvZT2
lT5dr9M+9c8qX24nFCXI05wVksmN8Yc65nproiBypKrbyJ0xHgX53nU8KgmadmX5
6tUQFpbG3odbajw/Odq3WexiU+a2ylTetNFs8amX58kmH3O79dyuI+F1mGK6wbuP
jjr39KOTZFbrPdrCBe/MEOCIbUXesuEXBl35APu4/o64mNdcqBp3Cv0bzL29RJOP
GT+k7/oOXzbsYyL4Zuw0VLbxbuzSsQGVHmbic0879gp82BEoAb/wrCBBwvUNGzOm
CWj56h7xgOohjnLcQwsJnprIsembZhQ5svVejCULENmlJpj/JH4+YAyQBBuTaoRo
iULAbWs/DCq5Hy1DGuzf/6vsWuOWqhJAPRC6WWUiFjTHd+rE6bOHi1pHdgSAcFzF
kYs/sEIE7TeVXVenmgVPkFh5riH86KLqJ0Y4YFiJN/uIiR95Y/fnJu7xr28BClEM
G8/KZyseIrv4ND7raLJn1CVtxDkULTK+XpNG7psAWkT63n2eTFVJQVsD/VW2RKOo
//WwjGkvEAeUfWfr11FaG/JEdRHfBJz+UHUlOzQlQcwRhUyuT+7bjY9lMUwvkjns
dIEp6PN8yInOV2AJCopfG9JmsqS1phnnZ6sHMelgJIkcPNHob4Qug1HfDjhVjRpp
bbQYNOwPLUV32P9Vc+OHHT+wQIgkTE/m+BzGCNSaR+Bo3mgAeQHRGXWZYTDDJPws
Yez4LdXnrKIFyyS5doCD+VSOpKxu3k+7cwHpLBeh0di83HXshJpPJdYlQfXqmkDa
6dxOXKIdU9nvFrCeOjOkqNxw8yb3XYtNVLcu8AbCsYJ+mKc6qPtyerXWIvA/YEEu
xJ7Gt7I+OQJ7bZTn7xSEGGjVeTybq5LSGN4JCH3V0kPRYSwQz0iyJi2x3rWif/cj
xTEVVqUEhr/flMpAWbQAxWBmOsX97oSiS8y/7sInHxUEuwDngr4Yv8viN2Ty+rkC
P9XjrwzqT55+po0iYyELUEXhGZjP2lmntG2kZd47FXhq5bXrZO7An1i/MSZY8Ed5
O92nkEclErucpV6GpjEb4OrtP0ISTDvvqk9rGyHlvMf1ADthkZwjZcFrXxhR6OJz
wizBlstlOFDrTTaxxDof39xitCnUkj8WYQ5PNXvHvPHgGpiOZbk01Q7FzFfgeahW
z77kaDq5sfX7pnQqxti45ESfikSSjpmkoP9/UHcbYJj/FUzQJtTwxLtevQsg1lkT
7W0CMawKNnw3Emv4iaN1FG3WZLEraI5oL8IgemVpVJyx3u2tbKSl5n+OIJgbaF2o
lTNPMECpSNVEQez2CRTN5qGYeTZRdKPXVk1sC6rInlfhqGZJb5nzlM2Xv61Sho6W
f5bPxdBwaXC0QzCeTt5W24REMC9MHx5mABlsM0p8QVr+umrkrjm9aN3Ldx6WvmCc
FnLc/1BevKNLF6m+VHqk0fexJhE7haLtGrMK0ZixaOfBkevozbOSxs0GzCmPQJUC
b71hmP6WzRfTh0wJE8s9NVQM4V0jH3Gq9JQ0vXgACG0NnxwAXzL0r89sFgsmUkOm
CZEYLwp9lRZuHB0kX5aJR51KbWmSMqzCy5Q91xCWwgzBJR+EgSboqqJSU05ohE2H
R9+5L6GtEV6cT7aCYstHKiB1zgR/q6817CXMS7VVjyee3XkNUAxHr8fyt22v8mTj
b4Paegfl9b4LSlazn3fa3dwN3UBYTLMcHaZdPSZLKtBysd/6J203rVD1p6VAsiUa
AtjemnFyaELXFtJn6t/gmfdu1tzcD2tHvxBMiGcZRzSKSGh6MRnalfFi0ocgUhbg
NVppvD9COCOJDFgeoI3nUAgG3Xa6XhOthxYhYSS2tp9Ne8Z3WGNiWi8hH2p16afg
V2wbZzvy4FMHVYHjpeKojsIJiLpKG2F576TKppn7HtTXrJ4P6ANCWhcG3MHOvr/y
0clxopMOuJn2xmbN6lmdvI5HPoM9nlA6h54GypLE+DG/uGl+fKpeAVyQo2If9i0c
bqXqfYXZG6uDH6n6VF4VgtirAKZU6oYE3nF8aKGk4MLlrAXHzBuG9hJ82S7ksG7R
etsLf7kIbQOfasHf4g95lBtAaLpRYrI7x7rzCfUgsNsrxIjMIH1pkmMtzCq1U61C
+3sk4SPlFjxTM+fQ5bRIpZjKt9yML35P9o8B703iDbDEGQ7hHCvulg8gh3YPD4Ee
4GqZpUEn5k89562fZUzRk3u0npmxUs3PyYwodeL79J3POlzkm3oyQZh3rYNN+3jE
lzy6IGxFJYHg4N0tfDQTZphF9fUACe7WMSWBh/oRhClnlk2s//g+sUb11gFc/9jY
6ZpBLkzrtB7TsFcM4Vf6br4y66+RMhfMLCKuG5sLnQQaxk6lN7obqDQa/NxeEp9b
O0nvXO9anfR9M3vEkK9puT7EcoJJT0REbZWNddrzZxQ5g6FQaa9B3ScU8wFzqJQ/
cLdGICTKPZVwJj0BT7sfr7Fz2psVXH4SDty8/U2UInQ0X9L96UgklHh9wALkVe+H
RpQVlbMc/JgP7Pvm5Q6rV+qh2VZoEToDKxkLz0zSJqs3TJSL+LlZXUTjxUHtTp4h
mIgAojF17bsMp1bI3XDKgfwyzhVeOS3gc4ohQE5tnWlvsL5dHzCgMjGg+kFI7wWD
Lx+A+zUF22y2+xZHv8zWFijIliBPFF5qjnSDOGf/Gu5Mrq0nLtoZm+fmKASDWcOx
x+t5FK6CGaL8eE1JHLzfQMzoMzGorPKGHa4WlEuJ6YIr2i80NbsHLHOp3SnULjXb
boAcsP3Xux5LTBktWDbj+GcKWLPdex1onMwcaWfVKE1XAwoKsqRFLsQ2NH/7YDH+
++pUKr/ZoTpURRNRlb1POf5VxZBvXeB20FeVLlzJ9lyZQf66ziautfKTtx31/sK7
6HKQnr/hgbud4qYVxLc6M0HvxcOTzowKl3cEuaLvhReIdYY9+ow0Zyc3Enf49dZl
ChiqFghPMEaXFeyQv9i1gVNgjEbIjKwqsFyg6Ep1KEb+Kdz+jx9HYxAkK1hL1vIn
rPsbYyRquOS2AYaXmhpn/5CgMya/XNhJ3lsoETYtLQkhj8veMbLGCyDlWlRcqZu3
8m97CrgzBlsmq+JlNtiFW50i0KDghidy3KpbeNmHIvASVHLJqYqX7xlrIVr19XV1
m8Og9FHhgbkkgtJ30OzOQL4jo/oPt0SUHhF9XhBdEzV7kz770LxyFUTqBdks1W7g
4sx4t45qroexwIGJg4D1POdcJqIPtiuzgvfHUdEa2G4Co6FYinnBGChSu2G7G8hz
7vNwCSQzx3nXSW4qocZ5kvb14JRo14qsoZgWpe+DFLOue1J7BiqTEtWSzTc9Lcm0
zJQjMj25FWuKcTmqIx80p582ggf/wVxvggy1ZE/ZOpzF56xPqzMBLl9FcW32cu0h
Lc2nL2+i1bzKWZeStcgMad4e7uOdTS3C+cDv+hz05QKxkqY9VCqRrFWqntj7M0x0
riCnG/h9RtXvViIXm4IyPQ89HhVZfCMTQKuB82l09Xgk87oaULG/T4pzlRDBUUHu
nIXQ0vCXj+CL/IcJHOPQev3uzxVEUqvmCMBdfcBheDVu11IoyaU7owXSJYdtYFnZ
mnZsj4fvRarBBJjj+Xogsa70sxyumDsdSwIRo+/ar/3g6wGJwjv4NT1TYpbxaEMi
s5j2QO+r0W8Xnkqej9/QE/XQXXXCCp+ejXRSLR/oJRSTBBeipKYeJM02+9wMH4lU
1cnhHhLZOUPedHHOeaBMBQHiLfIaPJMGg/nkrPfa+5KCTcf5MLeWWxDt1ljGxA4s
bt1ePra1fNfiBeyEvbJm3Mkiiohx2rNLNNDmaAfrCprdMc2LH7jjNJ+HP1MLbRwy
AIw+wZ6KO2wrwbfNB9VyszBYZEyYsdPMegoKVWXyqWogYTwWkNSy7sZv6ryiilsv
+HLu7QXYX0KpUcsJ99Iy+YoqmxaTkQpPvu0YXvIshIxhNq9e/JkcPUSGPS9t/8BJ
EY/st0ROU2SL9PZG08rLeHCWlwooB/x9DyEkE0Uq6U7BRxCj+FcTBnWP7Bpo3ZLx
0Wp0XLLDr822FoCqObU0np41wUGwt2BGX42mhnDa2UXVRCg679RbXQlvhr+mKED0
/WOFrSk1zNKwcQNFcxw2H21RCQ8DVmEXBbfln+u5vzi+fHq6lO3sJH5gl/nefGca
SFwmaA6tOpEKv+crYsBPY51ELMRkWraTEFU08zoj4+1aJbdRXtKN16HzIiVKQrXr
CXY/0CbJ/B4GyRcVMEq8AYpIqjEbmSjS2LrfAPshWrgvWpkyyZkFz+Y0F/IkqBn3
9aEBjuUnzGqXDAayEKSkIqTMrLuryoy/Ipwfl3QrRDV1dv9e0NisZpdZeSy5Nw/Z
o3mIa34g5tijsmbC3rgPJyx6dfGlhRUx8Xn8hQkOK5MTBqQJj4gToNFiBYF6Mnyz
nURIQWhoaPeXeKUFp8tlHuem4dtGs4ScOMabire6hFh8rmME194WAPWFtifKUqPt
ehICc5FfaVWLPkgEKB4c9DAhL9z5bJ9eakBWhLKNluFf9iq1DV35VoDaQ/lqI+yh
ebDRx06W1JOwZplkd6CsGETadZf3YGpVL4NY25ouKsx+nsPXDvWtmM5/zWiv+RFI
r7QW9rAf39MczWE1npa+050LHSM9PnnHbR72wDAOfn6+1mNe39iNBiKyolA8ztsU
DEPAKK9bMLdKF6Di5QP4SZqHLKw9vstBBHYH1CN5PacFQkJKtW95pospy0RZGbiz
WrrmoTXSqBZBO37MzpEH4udQJyqNo+zqIgx1Tf0KPUa/RYh0Ffzmi4N1hTQ3ZO5J
YuqDgHQO/mbLo+YZqJ/wKixrVM6X4Qyu9RXs4I3oO/qqwruiPQFTfHzDWvOCv3tL
U9PxZxlKVDanOXhS5bq8a4MHLYZ9adB7EhpI5Q6KkDFOf6oyWoFiQ9Ey8A5MigwT
qDmeClILCJ3UdwVvTC7h5FMK5n7ZrgO/mO0w/tkQFQQV4T4SqvqJePPMMUpi0eZP
gdmZCYo73pDuACbNVySFlcSEfhSi77qXK5TpiYpv8mUmppH21ZNH3PZAcnVTvDgA
lTCMx99qu0g5UGo1sIU6jcjTGQhPUxjoyBjFUtcZcQREfbaMtsyRTHsdmLlhNUDd
Mtl3XWcf7aPO6EktQHjq/k+NujeR2afrwRQWoOaSYKCyrTSM4xwKf02i/sKJ3Eyg
b4sBi6ZISfdA1ZR4bEkzk2a4Ovn8JMyzpokL98lQplf1TFdp4MZrUvoVSx8w5EVM
3MW6f5OonKfldqhMFE1f2MF/4rGRYr1aiq9WZrNjugtcYwag1gTL052KECsdKH71
Vis3gCLIwedpQuAs0LFwlH9La7r93rhJttsgBh/VWjrQDcGtBW4YJx2aY2MWzEZr
ofBIBVVqP7Ju4hJHBdFavjOu23X+eYzxKi2LIziQiAv8zzI5bP9ITKPojCjCJBh4
JMgxAdeJIgvww4xCgOZgf+vLU2ezJWFAWx6vUgrcdv/mE1ZN/j3gc+jSh5Uh+pBg
MYnrFndENN+4MHrYx08Cb64NSxBuukXTBNedV6ICD566nqGSN0rQ/QGEzcsa+kZV
j65zz2WsoUFOm/lkgHw/1a1u0h/PtJkF71dio7IeRdKEM2XRrVuPbsQSxR1LRG+c
gYJibfujUesbCIUaLiXdpxnik31IuBFniAEx5hGA99TJjri5vC2Ejz/SXjO1/TYz
p/AZdCjAm+kCCXIRkYl67GizuNT6DUFpCYvQyXy3YQqQh00QPm1sDXHoDkVQ+Rwv
lD+i62fUuXLP0RS1lVLYvozO5KuTjZlgNP8lOwUsVo8w90LaF4oRgHYUEOnKPAHe
GQK4QkekvXiFldUTHLYwtuJIsJSTqLgX0C/5YI8QatOWuA7PU2922358KhxM4ah5
PNeGGNnCHuf877phTU3dUZJo9HQ+56tSlmK6Hr1a8Kg3mqtwtpFL0aWF8BMswlVH
XJP96wKDDr2zQeFcvyXAVxoLuByHU6K8oounWKqEihWEWI1XJv730zqp0kfguk+g
fQiNseffebzxidrELihI8fWIHv+vSMynig9CGkQO1ooyIojOua9pLm67oyn8Jz/n
SATKd6lHrJhvBcAP1+SjzsoKJ+kitSkoDracGrJ2zTzP8z/lLor5FAA7rN80Zenn
kb5k/yj+SzBIGYScaFWUqSLqRZ6bqL1MXy0X8uYcasEBG29WQ+dsDKtqDXRRZnUE
DzmNiPiUzCkOAe7dUdoNcQOJwTYPcVZOjVjT6Uz3upqZuhIHf3EtCUFpoXBpVM2e
FnWaMYqvXSzjAEBLYSdvYG9AmHBAcqNhQZ1bjxmN1YHXMU97HTXMRJyW/hJDGrbf
HDnv76+wUzYWBxFJ53x+CgLeW5Fbwwbjwxdnn8qtsdKXdIsjU7HLPaVysU9gLt8A
F1+4ryUbndks6ih7Zt97vpBe/5Z2z49SV1sYq/sBnr25gMPIHf52tkgDMWURRNm2
NGQw5NEMbSWds+141U9vlToeb8O51zy2rSMZL3xECzDwEsbmCv5z1posvX3x7dVq
mcfWqyAoaOfFxw7F5RR6WwNqCmSrfKKLZW0mfxgTpHZCHjuays4ROJhtzQxCZ/PP
YOrq5NR5PZ5fpo+0uLobkl7/AkHszQ3SUhUoG+l3lFOdpcOwrh0LWSN1XmyZ88ut
/8TnC33MFQSyaWejvwlhdAhAM7TMmlOtJEc/862h8RVu+XCipkcH1CY0MGrW6Fqc
PilS5Mfmjj8SUyxZ1DFGiKKe8tCUf4tBblWNB8eIH86sugqZ7vsoYw/2ZA1bzz44
fzqxVWUU3/CD3dkOaUWJ+VmzRD/ghlQj0FvG6qTtapB8rInHD0bmYGlC465b0nVv
OXSyb7SllrCFJPjOYweWLr2OnClJEdr6HGDabpTWMLRR4uYPsCGEW1mVJmuUkWQQ
ZR56ClicyeSyW4zVxPbcDVKf4h7cAzNEUyixE8JPGu0R5/HZ9tg+vBDF9hS4mXR3
z493LkkTTEKY0TGaTUB0/4NNMj8wKdxeTxQofoo4ITAv1JWgbGobbIhO7HnGdRju
1o5X6DtCmnDsb5om+e1zRfXqFbf44vFnBBliigr0l50jidjefDF8YmQoUiwlXds+
AUJLQQWkei8P3Pfhi0ux587Gq3CXw76PjT5iYigdXC7cjQQuiVg7diV1okvWkQVt
MHkB/lqvkKBTOObDLnSLfm+Hr5HN+c3ZGY1VTioDL/Ccra+x+unpb5ca09WteKor
hAwQNIX+fHB9lAt8vSPov4bHk/aZdsxEfTspgsUNsooekwU05qv42BjNYotlGUAS
G9jlFjIcKU+w6X/O0QPTk8eHAroSkN0W9fT9/au7EQL4t7L+G3WxTvtjYAy60sDk
kVCNO6KxK+dG46IEJRt56chiFu+RNCJARbKgLD/zhWriGoRNbPlcEySpRbNe6noR
vcPTeiuaB99f/8Gs5DYSueiPMQFpXXKRhm2/E+hznMBcqip08uZeIkvsE09I5ZME
jPQHkDCPnZOoclMgFaYY5ujepF66LQoVI4Hlg4e5fKSsr8DLWHvemVKESWWGenaD
gt9UkHSsyxxri9Ad4wDXe9lbQ2gzMjHdTLCshxAvSYXUKS21eM4RKjBoylFYGmDN
uaEUcghunSLLFCTAxv3myuGfcAby39Wxud0xIqAs7z585qYibh+qT2grAQeSNzah
fb10M37APkPxc9unq23bDBLBM6eRJBV3Tq/uDFZUVFx0BVlXtJGVoFzt2gW6uJoC
XUSdir8jIhqHLBo5Q2cnYzz3uHveFWAmgSnYdJRqYUj6Vk3HycJTu66QoLcG0AGo
XKEE2c6e/R1P3LD4MKn1NpLjDkrU9VB8BzGeUTyzTYfpd8WfMD9uYxxysvkSGbEe
3SH4vS4W0unvrOV1fgFxAJ8SL4dvisPTfbX0gFUAdYADD//H68nKuMQ12YORCm0e
4sJ+QIPijncFm1t5v3nX19j78MEPFismvYJT4tCSwr5fwnNWZDPpHoNTpvDNul88
MD0u0Z/weR38YgnYcNQ2BCW5FqXBgiH3JWg6tL2ylk+1NGKzMnSZbIetsQSZV4+C
2HF1Ab5Uhy/IrCGeB/V7Poz/iYB93rEFh/GHq5/sIV2uGYdbCUeN10KtYINZnfGU
TdhRl8pOezqXrUTqwbbYxjO6PPm6oRmfc+zDfQTfZOBNl2hXdRqXnHYnS4yU8CrN
q60Z0VvQo3HOzLJYbg18jYRJb8FgZ76g0uhVinAytwtBhsxzyksceGv+OGx2igPk
Ttwdfk2bHkfpDWeHMm77QaMt+nck12tgkmPXERgDLkTfB9xFB3jFH7kwshudKaHa
OmngQryz91hp2XImfbqsqq70nYnrTohCwp/nLaxpZbDB/9AFw6vKHKE63Waw9xfd
agb66j3nZIxApCrH5kpyLrCrJAnngQCghVglwKzftpCzoq9Zs88uBbOoaEHvpQC2
rIl+4gyF7mNDKFuQaBX1TGIWva1xE1MOQ1AmLa8OZJSYOnHsvmsgfugeza2QoW7w
brbHUZFa5jkUlQwANCRuezIgicKlxx4oNgsLHwfmWBI8evID/e7pfoBidxpRuUL8
aY3AHnvetK8TY8EEkG3J8RJylSK+dIQYBQ2amLB3REDl5zygyAXAPwfCC26I83Z9
jDfw/33CfHikQu6Yjq1M9/2P+Hhrnxo1MFmc20gD/bDz98Fj5rngjkPzwKWHAvDP
gQYDhUSHSGu2AaaUHKaH234D0KHmStbca49sQGWP9+MwwVkLvQerl/oSFckd4QlN
4DxK3H6C7TEjE3C8KaUXnpQKg7V8WLKei/IZOBqFIV8VL2KwouUCfdRhEqj/xOUR
G+3hQIhDn/SueeB8gyV+Rk1NIrwy1bSgCOX4q4+IPvexZ0D/OmwVx0czxFr1mCQj
3DibM7FR189cg1HEbRulDKIfgy3spXrPXj3DzMrevOFTlhJKRZ86tAganLds7R4b
UZ/gvdGCQS67+iRWuOm1IVxxaVg3XdRmuq8wk/aG9kP/RN35BJGiYlDIVVBsD53g
5IS2JKeqiYOvLCur0AGwUlZubJCMTK5Hbgy/PYPcTZFWbQFerDEuBknyjOwvgZOG
N2Li0EUIiE1zzbIPMt1yZGl2f4TtBGXqrP9zm2ODytbcFo8CwPY15hkkyaYL5OFr
bBfmxKA+iPOaeyoLebFV0LDT9JQlsZW5lh6W3xQtnQuN9mPzUHBc77l3Vgo3DvhJ
1Fr617tWkeAFDoTchQNV16Pmn0m0EbzNhP0y7+qY6nhBVLIWOC2Gol8De9FCbfZ6
Mr2Cua+XCQHqRVTahWYz5JNCQI6ZLs1mIKF4BSpWNm/oBKjHleUz3yKhMql6iLTZ
I2NzbiFFSPZtqi0h7RtCBudRlhzXpodHgPcZsLSnBw6KevbegI53d1UDCXdY2mDn
2sfpPgWtJcRfo7P4vdsH/UDDuDzLoiTNT4LTnKp1j5x1p/9VD2XlsLmQDAQadkQk
VZvC1O/wDjcvG5n4+nC/RZis/vT814k0soBdiucuzBmR8NnBXTr2IlvGtQQzHHtq
vFk2ScoxXYZKt7T6vGrYsP+5w4e8s8teIe2JQT8VHUHWV4xLxJK+NzWSxX59YLLA
QB7fqUwN4/RcotY5Z+xeRcDuBPYMoTlMDgMR4TzgSQ6kG7bvcVepcqFA8qDoiJzv
5TEiqapP4dYA7QCctk5Xwdq2AHdU61nwp0dbQ8z790LhflhcPv4V4uKfL8uV/ovf
ki6bmiTeOa132Jpg5jlPrM5dvLRxbiqmVHvPTW0diW5LfbCU73QSyM/v/uU20RRr
FiHlRpW1r4TatsCALcZIdJN3JJ6Y8KBWzdo+F52beDjT19YIM+62653wc+99PLsd
RPH/4L6OuQcn9CISve9Ers0sxex0TtM0+NLL72UR0yU6dyFE6hYrjeVBf41X5oPl
f7/VaSWq2RUNtCKNcUe3it3laXdXpb7o89B3eu4g0cuyVd0jB6oHYIjxe2Y+Ir/0
u/FIBmdq3SKiCXg2W3/sXQKsss4sVYZonxfp667vOjAYFeWd1iW1KuysFFV2BmPz
3ndIng6wSrTV4Dm9ZrrCOqPAXLaMdR5wzQfmxyI3ulAc2kiy9K5nyzUOwlx+4SRm
obyy7KV5hBiJlK21iIpm89g4ZNUyBlOzOQlFm1yhsjQxPnXA5Vkjl9pZYUz7wm6d
EX+nTm9KjxT/EvV83LGAG4vL/+nlz1ZO4gl0XS1fl7z1OoPhP8adH239sHB3RgGX
P51mamflprWAI04uXlUozlI5nIutYc64li8TFDNLTJFMnxwD/CMw7IUC0t0mDl29
rplJ3VgbtpmwNvusztPnXf2QnZmlfB61Aagk7MKM+yqe6qC6265OWC/DeLd3kfNq
7oPLX4F3iPOfI9KnosFSxLFCFhiZg3Wb72r4911pU9PS3luSqxyHzkGCjrp5wazb
6o2oAE2oTyd6wdTqDRm5J49X7cEHkCa3CqOlojeSu97htOLXrHB0dy120JRbPry5
9BPAqd5c7oOeClRIFodQ86D4ux49q8ajevgRn0QiK0BP+aHY5l5iEM9lgkZay21X
ihJEeWF+xR5MHm6DumE8gBd/iYpqvaSOgANNagj8Mho8t6uE9G7C9acr/S1/Yc0r
G/XDj2D6AN0TpCLi6g2yADqw9hvMfo6o67CPfp21wzXH/cs4bMm02Wrq84VvGujz
P8hbFWNZsjZnPBXDI2rvRfZkINxklTc7QdNV56SNbaMYO6Yb9Ji2th34Ws70ZAZp
6FJHWv2agRjk90U9d3h0ATWUAZTCPQxPbuV5DxB2YNBAnNfgrlj+n7HPRxjVxKHf
6Z68WafsAqwmFin7QW8C8wvv8iiCtElGHEf2VQ7Ey76s+qdMLQ6Vqnj2PWv3PJXA
DMTVfhSrT8ZouqLD+Q80ayssDgmG8eX2rN3R4p5LU6Vztb/gq5SHmDEKitOMSSpQ
ckUL+7iGrPbzo82H+75WAjWC4INREohDK+PbM9snyZa5pyHTPwMdrv2IIs2e1dQt
UYhHPOdL+tdhXqXWvETbp3wUQhRdLPR66S7VXp6p3sOi7uGy9CPvgTA3ez2obRdy
qBJl5y56jGXncMz99+zhkBuTfM7QxkmTYq1p1rZsfFIBS1ry+XwnBMmPUzOCVOQE
JXQzoiK5NMR5dM59uMmnQLJZM4W4XwPNkmXavvzIDkbi8033rSSsyCZ23HHt2NGY
Orey3R7x9xvZHPo0V2A46WWe29rT/5DyxVLbLZJaiyHzgjV7M7o+4hh2nNDhlOSr
+1Ry4bVfByvCSwLBaKkBqa3ruioHwaH/zKLD9v9EWmjEbjnyI8yNDdOBwoyTwiGf
boj+r385RG4mN9o/eI9ey+R1Kg0yQmOqYY/UKRcop1iQQDFVzyGMk/UYrvLi44c8
eZqshBTbfNcgvfBxwgYIj50E3h7HuDnLDhO0S3zywdbbeO9vZqSp4VnlfaRLE8eG
P2wyu69A3UyHU1n/ZCRW2fIK/L3CnipfKymOdkUY/ehTD+vaf3zEIc93R+nIeVVB
AOPysFNy5yXO+yDRnsF4SDisffeWY97IqrMX36PEnPtM5NVX5o5atpopsK2dhKcq
/gzTb4KUsqra6Oxjmfg7ftkjRfcvj6BKCRpNzig3YfVs6SGz+t29NZf3ryr7HbhV
nLMeuUzk86SAtoXhlRvqO3WWItFBTUCrhhDx5Np99sVWqSPZ5QEgAQkTF7XjW7z/
xYo5yxLlb6wyla7lyvA5LErwxyPOUOY2oXunqaTBom55vUR3/McXjQuY0Xv7Tx0+
rOtxx3j6CWqoAtJLgy+dqzQHIw7OMHS9M1KbbPHrfcqlan6LglUUoarsp6BsI7Mg
ESTfRwdAQ91MeDScCM4twbjTjOj/EOTf/yRCGXieUC0pA3aDOzvGBurFFF1f3s/D
W5w4/7Q7F+z7RzyPnIdn+jzV3zV2Yd4RjI8AL4orgBkwgGs1rUlxu2mnCGESuGZu
FP6hFXF4mpdiOpL0qtZLny6YWe2qAdWngEp+WNRLBFg5PdiZOewpBt2prSh3RJej
YK65iR5apvtF3NrXEGY9rLJVgxA3Wrwknx8FfRw+rniPs9JGJN74WYHVaNZYhuXG
v3LhAIMLpsFRB1O9KP9HX4Hq4ryKMTTzDw9NUUHyukP0VV4fwAbSStiiA7SWzoEn
lDZw6U12F2JALTrkBNloxgxeEoEFTnwRhWpdHou+SjOYJio1ISdr6bMJkBogz9Vo
Wvd0vUuA5wiTTE2VA/H4PaUPRIKNTPTWtKBFaTGARpTSsy99tul3LLpCr7NXavRY
jE+Qbq4xY8FTwsZsTcPGhpJASzG7u6/DRk1py+U2FzTA3bnKuYaw3EVm4sQKHoty
cKTFhhwBhmy7XxOl/x8CNJ+ROeDXgugQQjgHb+OQlClsowDbr5kkj6/vI5PeVJzo
gI4eO0PKyLHlhqmYtTKpkOQ+tSqoZqJQRnJ/XG/UNzKN3/H/McGzbaRQyFycgeyj
pQY54TyHtmR9hfrpt5beuTx7iWko3On5Su/XMaueQCd6VzX/6zS+/xK/uaZ+IAo/
fqlBN27JeFK6SQyZvRN7Bpxq8m5RJk+PHxRdnqdp6d9MegX2/lTRlTD+934gKMM+
Fzyr0Wh8dQzLGqvM+zRRMpqrLH9N6D3+w+bHdtNqbTcY28ZyQJJFcdKpuppvqEwC
lWK/0R+362RZqqgcdD1nSJOqTSJWxy17Xcd9f3q5YxWTomwQM9nkRJaFKAAMlOBZ
vmQBt0FjhxBkhcttTlIX0xCcHw/LyGjJjBKANFNWSwxGDplYkoc1fiAmjaMK2H3P
k7zRfzIQGoIsdoKUfl/XLDJHyLhz0bGmC0uycvt73fKuyu7p6Jip6vCZYJGqSbCl
7O/EeOMu+vygls1tA0DyVTS9FGvH30GWtcgq1WiUjtG4svmrGGjrf6yveyyd5aEj
9vc4c0UbcxfhjxxMApoPdtZZHUTmjf0zeXiyubMegkaqkzAaDzYiONjCWZPomTar
8Qz/Mb0GeTGtiDAmSRRWtzZwBqVaNhJmkRJMD32/CmIWyeBAbb1widuYvIidXe6+
b3W1HIu5TH3BLgTOtXaqyGiZ555mXxjsPZaMeM6YqC7rykYAVO1Y8Bmlt3gG2Lam
6CIjFwJGXh6YEnG0FMb4E+u+0dDjF+0KnNAgsXi19IhcRGVtnuAXZwpBnLKe4GfP
YkLwb7ETgHvhhO/zLA7hbxKKoW4bro+gUHwrFLvpfibo9XiGs+p4aaampYY34/Bo
k2lek0kuAe3KMiiSONjP6xcdX68qgzRnZ4ShV/3y01dB0iMfglrU5qLli6Q/zmE2
+oGF2yQRzQFZaDk+inIewKnQdBTJPghcO/IuZVZACGNxcC4WsA+pJvAkavcTnCeT
JdCbwitFnYz0bdM5JpViakNdKPUQLPV5GlRytC9Na45Ry6viCmPV3fjDxG8drtRQ
hDRrCq0kqZqCie2rxmzMQRjSxUadkpb4sK1BSJlxfX0z4aXTzfRnsR6sR/jBQljb
IXQtNF6AhuQ0d4w8BypD1aevhxn3OwqlIASUMNoQ8qOycihshqIN8qJS1Ela+LUA
V/FUbtl7G1d+uC0ipRovT2fGAmkVM6Jdyf2fN6D8hEXfQtJSJqQ9Ory2zv1U33BE
QfRnVV23Fj/bgcg1+mUGOX5VesKYmMk210OlXd7iyTeHhaujlQrnNzrGYm76RQAg
kvt9XevGCtePrcXw3R4ilG0ffGLtO9GzycMZ+QP4gzAMFVdgFaHxFMoKxcMONAoo
Zh6D/u7bUxv2Pacmfve5HtEZLEBDw8Eak7cg3n3ObzSeLWDoOS/YQLiV8RMe99NO
zotWyo47z14cdSo/DniXGIRS6RWMsXZbxGw1wDOORJVCgC8+Zg6v8LMm78XIIJ6R
XCYxewtnZDQHuPYwCGJh0CVk/4aelYjJgaqofBU56rGtrWMx4fpWZpoC9bcVBiCT
UrtsTM3GCEAjc3mDEVFzbA6qWkHMc2gUpZeMbkS1OCRCAU5HLVEYJupy4MZSjsvv
qFrCfB3xPyqcEQA5508KF50BvX3VWDn7rsAf00nyqmk/X+aMypkgkUa66ZFsfK0H
2XrmIutz1PM/juUj9IXY0w9skMSygcOEz9o2SAHhOQBNw4S/kldDaFxipqhylHk7
ywSOS60ip6NGTARixCsf0bmfQX1pTeE6aMlHw0WUCNJWII/iQOFg7HZRuc8ZszuC
VJT7n6EoDdTQZjBA+cUblRLoW9kdK3wd15QyW206AQl6TIkdJSrjWauWT/grnH7Q
lmNVZMVp5cBgUXXQCemth7B9MwKaAvwOnbP1q9bowKQlju4Z2dAR7E3bitMr8I/d
Z4JLKjS6O+Z/G+bzKZgbyORK+vUL7iuQZ5SWqN7YELxN8Sp40hXib5lF1ilqDu4n
9oQ8JweQYP6M5DNhJZACBJVl4rgXWLvd0h+SlcL3N+X/JGRn4civxWMVLj6rNazf
iX+x9ue7FtCtJcnzH3g4uC9Ot4S+LVYVtoYaRxXeaqWtz1mrbtJ8GIRIQBQDKcwk
k9WiT5Gb8E/93L2WZi2AnfAMOWCPHJWILQ3LQCE27yujaI+1VBLWmBVUPGPCMBUY
s3ipMhZHNSvMI4K412rXKFuWpSwWmRQPtWGoBhL0mm/XWbkSkOpnS5lfZb6Qe5JG
SYGMyhVEO8OvaFGE918sQXb3YxKWldjIoAzdUQ7QkPVZQEmt4kumgQJ4FfRRAITh
mrKzPAxxMeXRVgBjjpZx5CVNyKo9Vn6vHXb2R+s3Wns0aGFhaoj2iZGsq56q7ud4
JF6tBgkscXeuJiMvuwAqkGpFeDE8LfJG8RpOVQx0hUAuuUvtm08sJw1AVSKIFfTh
uw8jE9j7wJIn790uqNFS23CsbrlPceWDsKeRDFOXaHrCWY2rwUEWeKwJFT62lDAt
8N2s1plOtpM0G6tUyUpvf1Zn5jYfMYUwY1hb9qMSWeibnFcG4S1jQRSorP5Nbr8c
FYPKnJnx4FvvbxB/ftRzgJBn56c65shrNyCld1aW73KqrQ3QweNqMbWlXMhUujic
RaVYt7Qka6/pQuLnyF8Bf11ee84cfIt70jgQgpOThByDHpZxy23QbnYjkBKXxGC4
O3SzALpaH6X/Lln+Rf50SM1TshK6znMy4ZaW4BHTLI4gpb01RV97GBX8hDiiHblt
W2Q/ZaJRpalNdbPsIoU8YBdwuXql7eUvzKq2htGFwppEGeWLoWgZ/v1ppaXhUn0y
rukvD8ParGcLzyI109cRuBX6B2BfjGphrskoHkbJudlnzOblx04JUR8KGooYXIVM
fU5qUwiLqkft0Mcw/r4unobpmyhy6Cqi86lB7K6pkZHI00tbYnXor/4mk+xQQmqz
Gc/ug86oMw6nMZatV/xdDbNdtXlD2ySF4r8f3Higb+yEsqC55jKQIbDgnyDZqshn
w3u6/JnX/Ief20uF4YWe99qp0CK19UPkDMIGixB3OJoH/qt2+fBTfnq4PXnXfuHS
Cdc009lErw56/mRclyil0JifwIosB1NX8A9cO4b/OEXJqrlSYAox1s8NsCy37j9q
deXc1CvGhVytdhJCg7ekK4k7zD1PAHCUNOTvj4zxXARS8eFquNRLBERB/2NeNHkc
05qOgdMxc3m3nxy1VRkU30wqpyUhxjgjsct15ypODyEF9w0uYu51cbg0xbhw29/g
PhqcJ/LdTR/cGWMG7YaoUKNnaw26lKOrfHroIZST22VTNhVoQFm6V32DBeVIf4hx
q505uNSIg4uayzbSleEYlWjtGJns3XR8iBBDyozlGiIBYnT0JPYF/yUU+06KXijz
BBzYftr4ovpsnfAlTH7pjyYWfeu/LCI1dN5wAdM9YhjztvUjkv6LfDYpFzglDeYB
CWSgVbMI/p8UvgErXWyM8K1SAj6QaL07kVEwijryM900ExBJT3LQa7ha96sm+dZ3
y5d8NzVsNpTaG3d1CHJ2+5lYo3dwZrTIBuCnT1AW9Ym5EPCd1Smj0ETP8ZTMfw0+
RWGu83dJE0LtbQsxcTZXh1rEIiAugIV4/emz+JVx+4+PEuiG09npkGyLw85xyE8f
CFO2LvQguPfTt5+JJJW9NW8t0GjM3UwcK9aILIro++8coZclAREoOTv1ff3ZAXEy
/+c+7mT7/zK0+C7KkjCceHxqOqoMKQ9BRWEPGi406HImn8diKNKVbgYYe80Dhnyv
u4dcPoQzvlMxOwFkr6WYQ5zZuK1ROinYLBzUqxXwqvLUYro8JuBPROzjfz5XAuk8
+i6oQyoiVJ8uklAU6AzWRgA+PIc6zGLra5xw/DqpKduITAgAca5agpQkw64qXbiC
rtr/jyjyRadugOs0dNrPgBLnQY1eEmoY8UAjIaaOWZ7H2b254gplorOIFHw9Owy/
2rGVrB9gNwEVAVwV2YC+JoCqKKgA43xvlNIuP2nmOlf56ZRF4wUjV0sVlxvmBDO2
JSn0GJzoWl79xTzCShmcCaVc123xJhdi5tHqwZ1uqLb0UylRT/2jFmS6tEbrmXQp
QjMLc33fdZQQvavEXUY+itjSwPPLMnyuNzvw4hiEWP4IlA7GhqoUIx1Jq2TqJf0i
NTSWjew7cPU+xw3jZ20JEgqSAPzJOJZQ+dW530P3tjPrz0T7HNyXNgRPO4oloWP0
dN12f1nbfpl9mwkE7m0/s19/FSDpvHhEIzczbjmwEfNqo4S5yyLYWq3/F+YKioEl
4gKSdW4p5JPEjEOGyQnJ3WQFpXXiZy7N4JhinBgrUHjfAUCLUVBSgxm2w6/Cj5nO
53EPZ/5sBGqKibeFSzodQ4RKOA/0wkRTguK/m2bafHY32si95WLLtv8Eq8WFO0FQ
WYX3HdejpEEjpfDeicMJujpGOHIW+8EKD7+SLlJD4mNp2FinnbWB/HrvMgxfmKxj
ZYijUD8RBB4LYEFHtwwLFK+iX2ZsZvaXvlG0o6toDRdUKJ+e13vrynympoDwCElb
jT81EzXUs/377BKfGBXM2Mn+RSdGiSiHHdN1SuhM4OnphcgRX6Dc2lYrx5VNu8wG
j6QYkL5UZ1Li9Z8P4P6KxnSj6vM8mXlAmmbrQFm9j7cCyf/EtkxOYNUPbBBLIGJ7
DF+Fh5i41tkyTX04VrtZD2T6jcw7kRbCa0QIoD8afDcY9+vWKlEiHRCA1E/vpffE
GdlfnQDGxfcNcrr7dUhbpWP+7/GYMAE8aOGaffeHtE78iACQx3zM1OxPLpsZqtq5
+IVJ0Ubo9O6VP1RvMkqFS969YMUD0HU2Dwn+QNnTnLnSTeQ1DYj+zPxlvcRlktll
1YDBqiHb74xRHjRVHYPMD5Fw/mFTvEsW9i1g7nRYddC5hu04wsOp4aJIgZnMotiY
IPrc/cOOoj4dOyy2XCLO8eX9NoYQxmNuThy4IMT9cAEapbWJd8ZQpRx8r/4kJnH2
4Q5FZte+Ye49Kugog5u293rB0Jji+X7VwuJvH8rjGQ2473fqC1A3jJkuRh5ybLLn
iptNY2U1qTVwCob724YeNeyul5B7Jkq2jJGsF0ku0O/aKxp9PGCawQRH7QH02/Xv
6eCSeUklPMWxsnPmc3BJlPb9W4wtCFsAftvTcZFWiZRJ3fJ6NDsxonhsMQSBDFUV
Rff5QVkRXujoRD0Ysf2dBsFz03P1bTCxf2CcDdHj0ncYkhtLLoFxXcS19RlmmYVM
IFJ1Y+1/FPdUKhX2HKkIgOF+AIyDJyFtMCfUXK2VyhgAY4yVbMHogXHlkPRVTC76
0iBC6tBwg1cCbY5AqcL/USaZ2FI7oWk7o+KWoSLofY2ZwbhiRfcPAwHrPNcufVfV
Q7z8rrsCNg8nJUQIStS/6qHYfIwXsfCdJRrHTPnVlxx441+tiV0S5vKgHofbQ4Yi
kAe5rvId1dMXjX5LjvssxTlhjREqnsU5uSswaoNt9YBp4tcC6R9Zo9H1dC1Xo8uN
cPAiUIPNcrxDgd0hrnblNm5RG1aDOyNGnjTwifabHeqU9cxRpBorn3UVDI9AAKqF
CPN49zPZyJx2qJ1EBJH2mK7a75AZSq9O2R4b1gluZlMYy67g4SKg2J6goM0quP4L
wCvJfJNW6kyJDI07/lGpWh1TD1DMQTIIhuJaYrgKjpvYjcy35TyUDDMYxVpfimvX
llufoGOMU740n61XTD4spk3aO7o4NcomWBrEAVJKyC6dKIIJdrlkaSC/Tm7e9MNL
qOqPv0muSKlnIF0qJEYEQazD3LpzjfrChCr3lczp1eTl8v9VrG8LkVPOo7hHC+ys
0l0+9d5B/VSPL2FAWM9Q3DygHUMWAyUfrn+ea959Q3dwRWuvO3kQG//nzgChfV7A
psko+tonhAgv9iT67nSgQWUR9NSOBZJYBdymf0s5j/TGixWd/5pi4gezByCSQNlx
mWt4L768rakogUr1IsuuH2D+oChje0siA4SoP9e3tnlPUrh/80lM54+ihSxf6MLw
WLab0qjXjSbhC27FGyHtONY/12w9zJlLAboa42bfyn1AwgLMHhnl7O3b5mlDJfMd
Az6pyPJcH+kCIVQM7awfHAscZ6CkuzCzj4P4mwE+4GSSKD+PzGolcmSwLDPntwQN
n3H7kEY9mrUc8SehDb8dYydVrkyMK8UUzs2jbBCWrJib4U9s4vnyHwJOg71IkC9F
WYtgvTt8EoddxAUjDXw0rb6Hv7DWh5eYQznad5bgz+UUeUldAXbKdkTLp2K3H7aj
bjBMu08k9uN0vZo6FWAdAfibkfRMCtfnr1/0EcY1TSCPPUGytTnC99B/ZdLThcME
5BGgjm/Qp4TWULFT8xQ9EwSWhRhC/z8lLx9m4liR8LuDnMi2qtEqIBX3TwbdUdRV
vCyvo6oQ2xc6Xo95e+/nwfgkVY4wt4VW3TMlbXigXkqAbBh0mMiTUq1TDoMgnktY
JRmbSDAqfVkQFAk3863fka23tl+lbg60bAhqzexzDG0NvYs2nYaEhQZUE+FVn9z/
EBvK9eh07lMMYTir0vdLWg9ym3SGaCF1vTo9oNKtycMrwym75QkKsKH3aeUGK9hS
w4OqYnxICGi8J7Map6u7gBQ8m1ezCd/JR8mtke1GKP6c0DHT9jmHVXBzjUmKs5wo
E9i/Ia9HkkM3LEPAg7pS211Xw0BPwEcwamGhVWr6AJAQf8yqr0Kgr87aA4pLUw6i
XfUH64ZrvOlm4HhI0k50pAT6CEpWnAx6VUeRHAz/+BQ+hpsy0y0bFz9rxm2w4/7L
tnG5s43LnoGignr8DTB3imlv84OAjCt2wj+wZZvqY+iClANaBIJ/SFckk59zg94e
7MVCwoH8UTICkNVFIYi+uRY4MmPHbcc/UBCaTIu/yw899hrGUR/BZmuFvs455qCD
103LuC3iAY+/WWPVgasNYweQxHpP2bBrzHtaT8WCcN8QQrZCMU8PpbUHbFfxwJEx
imDrT82yizc7Lh5FCgLyLo2RUhmEeZcZzXJtnaa8wG56Rvxbhm6MtAlp00pyEjHj
LWSC2SsYvZR+5n+zc/80tJyKnV7YdQ+cYxkDTLtkwKUih221MbhvhxKfehlVeMHx
OjEeehce51EQGqoe+JNEg9ThaKyuyFlXlerFKL185KXR5/byCbTn7x3Zypbmcs2r
SxGhh0ZpWDk4FVREcOHN/0sUAvMQ4dvnx4et+E8LWYUmjnj0qXYFGmFWqpwxvNLv
vm4e+6yfqDZaTOA5MxmMF63wH+6d8Iq639WvdatfIDx9aAfDHpzDzVWmhImP2T+P
BYa3EHzkd9R7NyjpOF45NdEnzwIAPn71nFjvAFSk8mUUWKkwaoZFbQq35fbXK6Ng
ObdtOaSj4t6R2y2lVHgyyIGvRx/AhgRl0hysoyDqJN8D/fxJ1JSk+vs/OXIVrZk6
qLw3Ig5xHcRFhFl72VmGPgJ3bidSKCJPih+xa6qAMEnlfy+4D4wJEw77PiwGFKTZ
oVXmpa9z8vWpgaF6WG97zxfQvCYhipBfmKeMlfdwqIXNx2kuXkQEzEbwvBbidlVV
xQjQv1iZmlIPubEu4z9T6ITt/fCRiWGapFK6esumzK1H/OcqxSr8pI92t71Z7hzy
H6ijHpX3G1TVqPS6ixhbno4Hf8AeQvcKetbfM9Iq+fxmCCAMt6YkB0QyT9lMdVae
ojcuNs9sKQ8TmQ83IhWeu+XnjQgVFGKCBBh/Ey4Bqo+rY5v3Ws98beuRp69gVnB6
HEfPzTUywDKj5Q8ZMtCQmAOQ0zRfmwnsq1C7xnQziEuAefBrMl9mccZoRIM05kfX
K/7AzmMg6PD370GpeLaCc1LxyB0JaTMQIfVJbRX8M1im/kx6sCcmTm5Twy1qV3vI
ZhrRBE4P606ZMJZvDNRE3r/MoxDw8KpmwjdY+7difXreLCI/VdZNHNNYEm3Gaxdm
FONkSUJsinT9BEpz/kMUD2RVoCmBtcEdmw9QkPMj6OV0aNU2/+sDG5Mph5PuV4Lg
PJmFyMXWN4e1gqcMCFqkr34HbtzInZ7er5SrXW7xD8uxWr+i5fu5+EwKf5NCRQcQ
fg/WJ3/b2WdQRtJAcbUATjCVMSXSunt9RJBfcj5DN5Iw82BPYP4HLOW92wNnxE/t
6WtZl+7XG46H8gW3OcZj9nzGHctYMnY0RGRuAzWYHt0RL9lc9tdHYDk1oj63NR9R
NDg6ltwrPZ40jmA0GIJGtd7r/441wGF3M5mLu8IEyNDlmVDKUZ4HA4kDYa86v+EK
L9U4zdzHlnWw1irzg9R6/LTa+cVO6NmGUvwYtE3yBuAgubeI+l+44HdQAMxZosB2
0uUlH7NlWTQdwsjXXqdcMjPmChED91IdZoIYhTRVKg8iuRfjd4qaUO8w3qTdOArT
ftiFmVpkjc0cv1ftxHIDwmhvi4dTi/RXCM8NRKHG3qSuUkotLM8tXpLhc15xcJ5s
OJaUvPSXIrlLKgSd4gbtM6Cej69Ech6dZKfhIXyMX/qIykq39/Dh/D8n70DR/tHp
SzaLCM6t6HKtuT0Wr3yhdEyTyB1/uKBG33Owb7Vsxc/uD/Eng/VmZOJ9C4VR0sku
m4xNqcwT6ZXpOBTcwQTbVozk1eBNtA2yZzfEj1eODKKXWAg2WXY4ezQleO5vLU6Y
dXidZOUx8IlwjjQnARqYUYpqfWV6meCrvXtVdGqcnGtmU4MSswzIFM9/08QegfB3
jk1GALk5agjI2Z1QpurowiSTAm15JqxTsPsDU70t8Mc9SmqZJMVrWWpehuEVtAPx
qIyN1rDECkpO3u7bjg/Uitb5nj444kXVLsXmFlER/GzX+MKAemF8Ivu6tfyDYGC1
e4Ju5p2B25WC5Gim4DCQkbGA0Ipg/EixaFRBb5W959Da0DEXMssOf/YDXlGpx+lH
H4nZL9+4mkcfS9wireBlyiPbSVusZ9XO3aDaDlSOHpDOUdhLydS8WrAEbHCy0rkz
Sr7kYBHuM6hUelUFZFqePfXntEuH9wk1M6ePJ9zXkWDVDa6cwPC8XM2yyWvfmL3v
XS38OqS3FB92KnCzL9S4PItOU4FoawkV/fspuyaaFDPtn9V8x4NJoGSdO7PgIFqj
tQJOO9zrt0DNBMDEtKD2oTR3MWCOclcIn2ZdV8WR+0wPrl9RlKJofyZ+vYtcwiyu
VvrpumH+e5ZgJQmYwG4GRWi+xw8gYSHTTp2Ph5HW0parbHJCJnn+jQBmd0omvmHJ
qH/qKtBxCtQ4lGbIlRZQgSEsSOP3bbdmulCL71dV993SRE8y0rnBMuyse3pwXrO2
zCPi/p5s8oJY6VhFnJ5wdpik7+yy7LY6Uo38gCcLDyLLq5usVZHtkUyhDhgf2DjS
3RNHCeJkCPG2BbIU5FqNlwyrXir0NMN/e3GAwY4w4EOC6V/fgOuiHJGy/iIaYg2q
Z1oWkD/DcMvumNhB2ZD/Z3BOI94e6Pq2FF/OEMc3/afnoWlOL5aiXdIZfYGiM0KB
oiOn0AzqovsO1QmpKFs7t2z9Ot6zImYCcEoXt8rxkrwTXuh6Nmok3FTO63Ywl3u5
Di3Iqzs3Iuhsji4N1JsILuMYnBAhqXkDMDH7M3m8Ve7JAyrHn/U/QsY9eAk9IPD7
z78C5r2Aye1zy/D57XltBMDhbemlDkvbWd2uB4d6qukAoJ4+Oocr+/BDf1d+S6pa
8yDxIlQgC/ufzKQooSatiI1teVuiJ4Q/9jAHbKMPrEnnV6VEPbipv5CihdajNWNI
I0wBJnKYiDZ+YejZgcpokVPmzRBcgk9LQZtUiPQBWbExQncpVsbm5yelabkdgqFk
I7Onn1q71es+wDtkYZPlFOeAFXMQ6QoyaDV7vrSJwYSNinTclVEnzsSpf3FXhBEk
PaOBpMTUkto3jxkgUXySn4CSOjzcyskDKyeI+qbd9uaoRe3P1Z+3gzI/FJaT4g4G
LnizUJ8PlAUIzJquBGQbDPR5E6l4PGSuX+FDudobwsO5VGbZZavcKHrzDqdn6bhv
CNWaOw9nhx91MCmDyjFsWQr3Bws5zC2AbfjSc0N/pg2Da2IyvnUCaJl5kngqvp8g
Vg9PD9CFkAt7MSdR1aXdvykEjkjMod8i8NT5EaETbRt4BPNnvTU9IlVXWuPVLJ5Y
eRnUMKgL9mYdMjYUl6mkhoVgTpSxM6v7qN+YgRkYnDc55Q2Jx9bzS2s57uuduOpM
kSy0QNr0foFYuYk1FO8Nlf+t7P1CXQH0Z1DPlGyz3Lzdisum9jBoxc7l9mDmFJBM
e8Roe5xYTs/IMx00j0ZH9BVq8rLZdNmSjfHslMGZuRGObbrrWzsu5+eNEh9Azygm
4kUy5z1UdV/8rn5rF39lqErK0W6wUEnHPI/ljohs/sq9CfSd9DYoBBsw74ctr3bA
4nq3sDbiHJBKhBzU1vHw9dDJ+5nRJ3kOgWp/xbRbUk2VVfDQo/ltIktUiHg1GESZ
HUWNiy7tPydoG7f7ewRW642bSKEL5SvXftr4axO/seW9R72VGqdfYbJqPPH9TOqH
pNqf8FaRCb46ut6RFx23brsIYpsachFOiNW+DyFPtNZZxX3QMl+uL9uewjUTitCz
Rghy8zjTlo6F+bCEE8+Zw5827VomZZg7WQTpZIWsJHYXbAvz5thZ7n7WV6ZVFyPL
xWMvdeYOOmf1J2yV5/AcC6XBdtGezNgodFajRicZqYym3RRRPVD+hvM9KHkN9vKi
iL4ANSF/sDWcGj1OO8AXZABl+w6Vqfxk2hUXQm8F6xakhqD6lCpJ3L3j54IEfVOQ
vwIBa1PDbreZkl93dQGbgIRymMNXOaCIY9aBcQyMd//IkaI//4RfBHUdUs0R7pBb
CvyEGJdI52hjWEYmIXQAgWOMO6wfYlycunl14tcOAFNl9DYnbM6kWyQjutzj8PRg
l2y7lY+BptwlAcnH0AVYdWYGU+u0zC73AmyuJ/HP2XKzUPuzhv++xpaUoOPerdhB
W9iFYmQe310eO8WoyBUnqST8VDwnoYEjrk9XAhd2P0Msni4bVEinmg6V6hGTGwHP
gJUSM70yZq1TncJe+8nBmGSOkgABJOkCbLk1CQXLLPXlHSQjbMwhG82fffTx4hkq
uGKI88JkkX0iDaX0Gh3u5C+RQknnTrQkaZ+5NN8PBwQGYSXIs6RApHojwUrvkh1F
CFXp7GspEdY7Ot6ajQZD2nu3JQD84UJIAC+zYsmvWwyBaDkSSmOKsTp7BIqhBLka
YYHwxD8GF7cTjlceiBO5YVdxB5mdF4UYL0pRQlYe1DMLkChhJeGSUmnj4hz/xATI
rQW0w2YC2Nlop4Ob4yqDcTvbHLXpwm5bym+V75OA0EgF9s3IFmnVl7PKvpUxKVUc
vQ7gYf3CKiO2tSlgTxVAE0gA0GUY5hqdAqUHBitodNt+V5hGGP5sUMqZTzsiOF3M
hq4FXVx35fkaIY4VfAVsD/92mtIoZBaoevTAPlcd1BBUyT6RePmMLbavmRjaOOZn
e5WAoYValZhdFfqyIBqXMqvdDGgSiDSQ7dFk4VttAoI+//xrgWq+8GF/1kuNzDui
0LxHCwehhDW0/myJHWSxpI4N+KOXBJd8k0xLVZLafXykgizS8LYTOczRxSFNiABP
iIVhEiJM9Lx+ewPYDetJJyPXqNq8cgi0c7nXU/+C8/hBfkr8scV+wvlNYS35nY20
O/+EPckMn4o7XQ3RPB6ZPIImmW/auaNu3RiZScPZXXD3HcjqTB7rFLwIc0mDoU2X
RdallS4f8nMSw9eHKLt+/SA5eoiHf7gDNxrk6OCOFJR8LTXnUaAlMaK/O1ByQL1b
eOsshA2MRt+5oxXxq8y+SHgmBdwb9KQvErATDgNSaArIZdY0CqSnbFrmeX2pyDYY
MPfWpthh15Ps6+bZjM352lwzHewQB2ZYMRtUh5gGigaA/WziONedv+/An65gYvEX
RIIMbb+AhkPS0e3ktmAuTUSSuntKi+owj3iVC4Msde1mkQ58OQkEjgz47ouZvZCx
n4q5vSt8yq44KA5Dt9jH5rc9pA4+2qpFq6iGvc5L6EUfO0SblgRec0mq4o1yV4Xl
gZCGb2ad0/YPy4m7ETl/5CFEW+Q//WA6cbwk7I3NmKz7fou0YSaQWzvtMyP3smWW
q1E9XHZ3uYNC2WdrNTlQiXiluiltkBpsCbM0lztfacknlLp7/YZvCsdbEAt1LrhN
IQfvzonH35595SByWJ9H/f5FdgFDXBpJnsGh41eAhfEdWg5UAHze/E3SMbFMEaNw
O89f9jB0dDbVeOIeGg1aaKyW4KzEJqrlyCV5jfydGcbaLKHOHT29ozyX8OSE/R7O
Sc/4NywFVEUr+RZlN8iL0+hYZZRhNjSsiMGcUO0slwu5/VyzU3X6tvOw+CVXHd1l
fZ9PKx+Nf0On8xFOzl24eaS3r4DbQSTRPOYuCeELsEoOZkAJkeDuGSNSMFTRjv7D
MhLzTzDfTea7enYNooUBH2Gu4mHjGtlWcdFL2zMpOc1Odo9muvljB/Xi6u9dnstJ
TigyBqwCSCnqxLAVBPztCYLZfBetvcQF0VNempauJ+UGzfQ2V+Nff71MsKE8AUPq
UwFhviY3wd10bKfmmrfXTYUirq2eJdqId7eiUTin472ZoYLZ5kpqZoqU7hwuD6Hd
qSoC+0KK9csoGwjmWeyVammGyhtS2F/4/dI8YuXM4uais90GecY6YQXD5oHWmRcq
eussgXnNYDNP7amtPZTIKXwIcPUXelD0is1eS1Zw6OTg0hJhngE/vod3sIIKywzw
8vR4f82ezaYkvx/SxrXLF7a2HKmIr5vsYPbO2W08OH/x6Q8t8qVuqRW73qvjJWTz
i6YhfoSBp9KH+dO3pxWOlSPcIyJ/Cfd2nKF02cwAGrxx5Z3IPRpS1k4IaJDAik7h
3Yoe9WvHhimCOtQW7rJtonyxNvAy4YoiwvNWv+9L4d61edzmP3Exg/l71wADL/g1
R8UpUTAl6gZUBl4DRG3Npwv5G0/qF13105w1YsWS6o8pwugmUFMIkh5P87EipVS+
NvaISrRbbcwdJAzyd1XvM0kv885R3SQqntQO2XSA1SWRaJ8AJd6Sv1bKpDJy+xcj
+awQ1fuEa2VpP+8p51HHJ+BXgVPbFpU6ItRnjtPlN0lhlub4vPxJxS7fgZei13yO
V7YiiGWnBZy5Mgxc6fK81TN6/Fl/y/AgzTf5MjVfCm0W7H7Ad40rcHeWmWkAP0nN
uC8G1offMAnvBrEIjTY2kyCiVz+9eWIrCqPCRY7nGUM020C3cQdPfbQ9NLsCPbrn
mAwnHbcL/x7q7NXxOqx2MZrbm/f1Y9evpOBix+ssLq851cZjt4GNu2fDLBKmQuc8
rYCtsPOThg55Z5h310tX0YdHOV+4pYDk2n2IzlTTLrnjQYvV4rLNWGDhkG6g+UhV
ItnQt5jYzexf2ee4K/RQd7eGpHXWhm5cYLeXuJj93XUAbxegP1D2RcBUtUD8lSVq
/En1dJbwhjdx2dYqe9ekv407we9ldqNLjF//jGAfsSYkmu25UcIhK8/gbFaFEC4d
rfc08kggS7o4KpohT9LA2Cx+v90D1z+KLOKg+uQQs1BRKcd2k/yx6VEveYRYDx7V
woZCGwW3OxqyNwkYVmLbmN4aeBZ7e/4FGVXoGSUWVPBjZGAstI7gX6NRr1RIaQob
`pragma protect end_protected
