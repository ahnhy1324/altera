// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
rsJWBkdScHYfucENyH5KOFCdqYXPfe1umdPoF7NfyQwEyeKqMT4Hwo2TB1aIbtAjODXspGOD1woO
mwykLGz/9tCYXlCw5bz4lZXndEYWBu9+qLPeBunE0g1kZ4REDjePgcj6cDIBp+I23vc3nvwKfaGb
krHDL8FWr89wdTL582xX8vuSiZaoS7fZ0pyUjDGDuf0lT2eFDrrQzv0qlPV9gHSTd799wDOUE7SY
l/LxTOvUiPrj5uSgahqIcGXmRo6xW1SzAKe1ezfr3BhjUra9GPlyF5gzsWLfFhvkVLOEhZ+TgHBz
Kvf+RYu9Orv7Tg6rz9axYIOfBaqrcG82jx/BDg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
YnlmhnE9RvPFRlyQWAfpM8inlXAbUOIJ0gB+aUhYLaoZHjpcSCJZg4cBp9QyvkFekp7vuQEkXXfb
UCqKZbuIzZ5p278317apZ7Kq5JSg7u6lbkUAnekAcyO61vNJ0pWG5wtZaEuQ7jsFdaq62YmHcZS+
jhaJZejJabaRcKeitISDJjoISAhpLiBKb7GlP2+P/d1QQ4UhhOcmtxFwKZ0IV7rHlXUIupiFW5nP
ZdxLggp//sCCQ+3jmMoIMEopk00zY9YcJ9+w6epsupQNy99Zas6duwCXuA2DlJr4WPqa3FbrPVM5
H5i3VzwrT38KFIBM9CH2uJ4h1NjVIP/T4dznMWm485K0d2+S2dKEv4myqkTpGrpAorUjyUN/YdH6
bUmScvzjLwBVBP6BQc5kzhr0JRz7YO1mhZZfuylqUxtPr4lpFQY0zRfn3a96i7A3QEME3aNqvNKD
tMRuh28upulv3C66y1F20soidUdQI+0FlfCbnsOHMdErm5PYBQ7gbprGTEroaeW/H5RidHjbzrDz
Kj/KueZ7ICb78cwP608TGO5jYUrufASoxPoBaxhMqSm8cSYsOIjJg0753lg62+XJicXZz4zl5mGS
BGc5uoBRr3N/vEaH888n4gMH2n5fbwmev7Tq2mDceBTM1KuJM+z/qjwCRTZ7HP6hidbp6fGwUVEj
x0HG0DX0F6KqwZXP7RrKKHBuntBhN6jDDYHh0yDBHGV5WYboENfYgu0tU8bllsLrPYHFtbguL2UJ
DAoxLy7hBiaALTGCaTyI1DFwQyECMQ6VuOFpnGVUSrk5ju4Md+oic8MJKWmW/p9JhEh1jlmAk6Xi
rAmdpOBUm8Q5NSK9F/l0DlMkdX56P3RrF/NmEzTMmubCUMAiFHiY9ykGiDw4fhLAEXgXNvWZCzUs
KoPv1KuiPLlP6dmePPBjRfLhf29W+9NF5NpfuAOuPlCRFBk7e20AXmyaQDHYMYeR/y4tGs2M0kjq
Is2/z7I9Ri4ppBxT0tb0b4BIcavC5Y5MUArO3lbiXmMM541uhMilVcIcvS+/4RCSzW2vSRMwa6V+
rn7UxYKhKTBK+YbiZwOwFhFI9sGV0aJgT8DeqQ2V7ZuphKnwvoAP0PfQEGs338z9gwdhRJvIPryH
Nic8U6fe/oQA2fUGKi07tqm2LYCJ9jKcwBgegOBVYKqKkyh3ndSbn2fRxTTwKM+yyJNWlyCSlRmL
CdmqVxpglHj4N9pjlaGVmBq+cDCH3u2GgqHjDps99aO44V2VtD37eaH+wFf9FELBAlOTOKhMUx+S
CWZj163VpYerlq8XjZzqJMeK9YEn5cf89OGt5MejXiajGbJRoBdQdHeOQd1RhE6lzvq0mmTaMvL4
SRoisQhbnlXaC1RCfswiWP7qqog0okTG5V2WYgz5qxuvlifsn7auhZqRedp6cG7tyyBUewBW+0k3
vxngvFbhbNSF2+4leBUN1vaTSLaqyuN1lywUg229n8h5Pl1cozIGrdh7Ojm5T6OqdfcKjzOUsIu+
Yeistn/VAAFj+eoZz5Hf22JOadlpTUzfLtMKswkgWv3BXVdPNHyzqtALs2i6WkmbR8qQSsjXDkGc
pmpb84j0r88VKvGWvlboG7UdNjnaBkDSYhRQCPLyxE7bah3XVaHQyMfHBxfRXGS9wuZxjA1P7Ir9
G51iJX2+Dmhb9nmvEbzRvwhgR9MEdW27o9l/5bSs6gvNpOpEthMm1VsNpx7f5fv778t+hA+Rn9Qp
EcQa2INGeyOTXSB32u1HL2+CEZZEDZ0Z0euwAU8bS+v3puYkn23hYkZPLmxhbKULbFpyJOBAvARu
oOrK3+UG9gQE7/vizpzQyiyERycEEPHGnI5f9ug/RZ3bvtGyPeMhissvaqEo5BlCC0xxFEiId+/1
mLOliJ4ZWctAY+6ZL8wDqkKKVXu3xJMVrwyJ+XRqLWgs2DYpLj4Tnz+waJVJyISMYzn0WQ6Try/H
9vN/vqWquf1Jxu0vP2C/Maz19THtEmg8i/hqL4GAJSeF4yATykIjOds3quVwq7o6k9AokzPMNcSr
VClDK7MgIIHpg4qjfRjh8FuS4MWPNxVszsfAyDSiQqX32z4b4uKnbwlGOcP8tkf7pc/PHAD/hlEz
vN3wlGEhmqkeW26D6/tw93gtn/0aU4Jcax9ivuVWHa2YlbFo0xN9MNLTcbxXWkXh0IiilgYIuiZt
MS2Envzu6PlTdv8yQUjRPFagIEb+u4942zrdtWlOmmnYIhzmX5AboBv9vAf4tjuPG07YDqnSSqH4
nrvLyXlJrbEhbp3/ySkgWZ9Ak0rgoc2amjszJm1nfhnKXmnRfSE702svGQEl+Fo6CCH9Pf1+ooTP
lWUWGfv7/QVHug6xlPCUszr4bmoiXXYbD7Rxs0AJT7GEctdNcaNQFWacETNa94XSfSuv/J7maZmV
3Uvw1sFSvKwAkr2s6361Bw9Mx/8sQz+hyVgxirEe7xmPKC/ew1s/Zl+WJbCA2OKXMUvKntSyAU2n
oL0UPQjDoUMgDJU9sQLYm/ebSrzmbrz1cps/TM9IB52xzzBPIIX/xodwW6l9EzEykC8jPDG9tLpB
5YIh22cPf9yCU46jMcZFJhFkqOukI3iXoY2xFBfgImRM7JM/EdosE1P/BlPe16bBI5RGJ9ZAoVvm
V4oS1U6EsCd9k/qMW8XSr46UsjoxG+rIuhujGyc750jMRNSjuUUHbJwI0Bq4L05IGOgHRpSwRsOI
TUzovkIflP4hOeuaWOF2IaNyySDRFPYRi5uqpadG54/Kjq9nsvFwbmml11aewe0GBdmd/ty0iW8o
ZGm6ijey7wuA0ae3hwrAUcbA02xQ9eJHPSSQNjTxcdDA5lXdetdUcL2Otxd5dftOcFgB2ntbIlbL
VlxftGlImOxCoOKqpchs/RcNV5oOLbK6/tiWbePYkK3xsXEo+/AQQTqjW4aFVh0kacudK4k20oOo
kfZavknkKmErCSK/L9RCqpY4OvskLUOprcqDLcwCgkPxJVcW3j6xtKQA4rLO4fTohggZNJPYo458
dTDgcuk0IjGAq1zEviQdfEioI7gGEjEaZdTPa2HOXNpZAghz/FNKRhF31MM5rClt52ral/+iLNM8
JX3doI/fh36QSSXnA3Sb4ZtWORe5Z7G7nfxNV8syjMnJd9h+rkVh/RZFrQPVMwrYJwjPVm8yZH0u
nthXxjKB4LNXj5lFYT3T7Kdi2QDNfLDaxadmFZj/6lyDLZx7DcWkqMOxiZdeWjpEuUh2efdMrTxR
NjskivyOpwgXC3/AkyB1gk+FowHlQjVOcHNZWpSLsX5sb5x/YvAoupgWJf7Qq8dT2+99jn0eHjMF
XiDVspB2Z3yODiUMcf1xkt1l9t4Hd9/vTR+95+k3Grhznb3t/e7dyHiATx+i4BnqqDPtLUVE8EcL
+86tpveVHPQ4e9DtoPCEvOJ9CAIQ7Y04fQzjUMVS2YeK886oYAxgdTqDRiMo/DTrN9Jc0WymDrZ0
GrII5wccYLJ68m7drdK17eHQljoqNA823sOiPOdvnS1lc2WOEQMG5uat24bkXfCEaAMuINcSeEPj
AYYRIayVlB3zjGx4ujrkdRxZb6/5bFxCoKPsmCeayxrwYmuhtiPlyQNYBNWp/hxIuUmO9/jPQZVI
7Sm6RFPbYMmR4c1nsYefOXHjbgLv731Lzmqk5QHwSMq1wVJdEvV+oKWLUx7/SPXOm7UEF+0a6pN7
xmTeI877zPvI6JfhW6Ht6U/pPjG5WSF4910hE0uQaI1FVqd9wN/HuxDQxgehQ9l9lnGIMKxSd0UK
IqaocpdZ2ZNkudMwnOh6nEX/mr6ArBCSI7SkP1B1KJ5dT762LzOWsk0+CJhA9/+TSmIaDcc1Y88h
JsQsZQe0jzJNWBAGISQXuG0T/wpHMxPncuXq3xMhfoML6m/9mfg3ByH3k/JlrAIVFZkJKLnsRRXT
ZnrkJDywUZFfB6BA4zKEg60/TyEziXeHmzQxt0p78AKgqElP514LlnwxygH6WVo0IJFqBJHCyjW6
HH6fvW966wqCS3BixCA7ACC22bC/XbhRsdR1oSVAjn46fr2AfFg+sL3Jx93OfNAfSoklTx+1NNAG
sHkSkqiwX/MBXA1y5yCfwGwaJU4I+VlPnLmwnlutiNwLBP/u2oCGMbKNiTHoJt9U6VXWLxDRFmEg
ksxtK7SpyHH9ZKbL5VdCN5IgPNFY0GaTIa9/W6AdBInN4WRjgs7LTs1AYn6pB6mxueSwRSB87Q7D
c1Q93sDeFeGcO/rfTAEyuTQMJ4bIV5mV/9Khrb02BMJnSpbe6xGdtQ+aOVaZHlagA29VEKuSJD+F
Bo0CaxnXdS50pJ87iWIBpn5I7dn9nP3RoerW0lOOHan4nhizel1Elo2kC4RnLtKEn2VMBUTRtlVL
gtDsAb83EXdEueP+MmesJPP1xmZ02mMPegOyFUkaplSFbO522mAVY99EghIBKAUVIyyq+Q7T3lgB
6x5OS2f64Ku/Z8oEs2PpJIwoRkU1wvH7DOlsHna94HbDMrhbxdw2v2I2QdeLidNnv2PXzmztGqEV
Sggq9corRSYo3kJb73Sy7mhQLYtR7pT4HM4LMxJQXs2w9TPNeVxlXnuzR7mlAkWz1C2QOIVkFNYd
PgMkmQRgeaYehpD/oS3UefWixlh6dtc9xfYCmocpYkmUMZUlkONq/5aBQzKJRNbjiF4sr+wv7k4e
EUYc9kLedtVAzIUCH65dubjdW+x3tjiR65VA5s5ibmaYK7pu4UCJ5ma+Esicg1xmeXZdDz2ZNW0l
VMQYJJbKve+1Y54SiMR623/6in49IP6h1NdxXr+A6MkP/6dk/HgdpTbovs2n+DdZu6yNm/OWLpoz
ZIQJbTHAHw0uryAtXUlEIjyE3owuIPO/9qiHynGosQBnInl4f70YiMR9N0VonqfDlCsCLmFnQPLL
2uSy0I1JMONIhtUfrU3ZCy63wxt0G1FIqQcmIvPZ1j9/w6Zskuys7xCdlKKklpO3H2ZaAkw266Sj
xvl7q7CzckBPJQHc/dsI/bCEIhbbbb+l+dxLbCWlyOx1z0OWL4+5/ei9ys3q2+YHiAxWjm+7U/0p
Zpui7pSzaZyuqHxF4immJx5A7viK0MgPQgy5gJRF7jvATIhsilC+WvZMs1MmiZ9IT7LzYYFqGAt+
v4dajxzxwaWouIRWydITxO+8YJvxqQQKGP52Z07bi3OWxgEJeRgaXG+iqQ9z22ISNvcrrQKkSXii
DlQITINmRUp7rbnkDM4xFSli8uwjJYkuns1JgSHnnFexbOJhxIOWHGpH8pSG2TPXrDoibRl8vvMm
IC3KnYaapjNw46Jb8Foh6gJ6/bnfCzIxrrmv77Ow1CuJ3mCiBPCHbNvITRSXBZlXU1YD0zoSEDug
bthe+T0Y6hJ865gB7UlUEY8emla4d17vxW7uxbO2OAZctcebXlfQoPELjjrhXi683GDJ6Vx+V0l+
HnecgHGD8B3bwiZQMO+FJqlh96vmgNgst4ZWrPSe/8puaJrZzfNeH4bC/4sMAMXlTktPKA8DMiS3
vIG4Oxhp47v41RV7zl62Bo+3hqCr4q7h8poBFkiUaQkF+Zn0tOrgqvpHKomidyCWiXXiR96+4g+v
muX6nrzl8mha48caLoOMzBAjD9R/09kDl7W+Fv4kvYe6WLxkSdw2O/hGKwYb4C2NoVvISexwC+ow
/53UdJQqluGVFXFmGX3xJP4Ta68pl0rkuQ89veDIEPOde6HBvZgU0juH+XbSTE7wstJ7oVBmZUy9
TWox8tuYjdPKChJDZlmBt6HYNMfyldD7c9GoQRTgzxHQStQ4npxTxF6NofvA5wtviN0Te6qu0Zmo
donh1VycoqQa1oXUOT5E2QPA7IKswp/q7YluGQg3E2AemLWH834RJfJq4Dtn/OcskGkp5YhCsPu9
52ud290jdaYqnj/l89HJfpxMMyhSCEgGY/kFLtKxnMdZEVHF5VxrfNiYRwKhaDvcopBuYS+nkvJ5
kNYqfFFSCXzL8ba/zYerrvXFUYWkK2sjC38+rxLKyDtDa4m+HHCvMtFQTBMMiMFsI/I/3dRd3vQ4
jKsKv378sq36/PZO0uCU9X6sIuKEfZil+AoHUCHVR3cLh0FdPP2Xhng55RvbMb2m0/ixvyu/kCMT
hKLxrLa7zCCSakz4NTW3o0OnVfrtpyjyv7hu0PjzWQ52wh4pWIt/eRmQS6QnXyjXd8zLQSZ4g8or
obqrN0+VJA9HM7CXxSRnotkB4U520UC+jAjINhMZ4+W9w4DwV9YPZncOOquvYXEnFgZqV3VnOkn9
X3lgzzilpKt4Z/Pr9rQrx4itXh7IKecIs3ViQFkxQhmnHNi/MsnQaY+ACcwa/rhLl4VY6T/lWfU9
pyX489tHXeO7vWoexLaPMmY6j+x3cWfZp+AaLHZ2PW0ihofOhmuzC4/x7qrmetfHvSaD1bqT4Vt+
MHPoLWnryEjJMdwQydIhf+AFxBN6pLpug8LbTn6hn1HSXho6fpXtXjAboeba7TL1bPIV8GfdndV+
Pq72GwXWX7QkgXY2Y8zl0YN6nEQcwJ0rfsYUjtMmtMPUZ0oO1jVXcaP1VCs921idXhIe21Q9uCIz
gtxLAiINLc6y5zBvPqilLjcfcBz2fdOXumn8p/Da65qta70dBk+CQERukvqjYMxEQxt0UHWW6LVe
uY4pn89HX9lWte5L2dHZZ+pFrJujcTRZfSNyiRbMwNkRY8Jqox92oIUVbj1emDe4M4OecfWYBtVX
v4Ki6co3h6/0pDQ/WPsp6RDT1A0TD7spvyC96TWuNDBfUFL7HKe04XPxQtZJROIlPSiH8HaCz0TA
YInT7icX1kT80W/6IIft8hqPYW7fGdgzOwOXekaIflypf4rkEN6sHPcPybWapySOJs8cgMWw26dc
kdWO3XHA1sZTpvk2vlLGKiruZmMe3NMxR8MWQ8dML4T0hOGL6KPrNCI0qQhhGa+OrLgexwSxrfCw
WSGzgHwvliLxjoiIhlSqMGDC4qnMtNUyG2dNjFIsjwaEsrExx9dGvPI07tv72Bk0G5muW/hnrRpW
WpnfZCa0ygYABnN1oGCtPyyrJw5rvJqh7ly2st7b7cq3rbeUlE8c/iT9ga1gSzYQa+lIJpMMYdFJ
KgWg/ccxbecreb9R28qCdhzTT2lPY/Fs4odmk//uC2XRPBho1Gr4rsFiuihRO0yuxHSppSjvZXwr
o4NroOwVK7Rj3++UbsFmAynPz8TLw6zxzYy0XHQhb43ineiEZ2h1ZqFwGaIAzaSfm0x7+bAo1lPc
RtjsucX8H+Yi5FmqKUKutayOz9FuoYLzeVJyKzrhJKMUertOYQwR9E5je8TldheBXPxbaOfY9NSO
hR284oAt1YnLtkuAbB6Us/Iy+RrvF7pidSgvUWTpFtw71LxlUuZgIPPNUBH4gRgSmKGrqpypmh+R
8nXq7xOY96Jq9obj/FWA0AqjpwiFvuyubAjbYoLYRqjl2T5tQwa12i9k8ojS8X7MWKcBQ6GCr3Cj
UG7Fw+SI69L22AKaeOXJdvzra5p9XcFjaJ4uvmWqYrXFo0KHM9+T/qDjm//c+v6QzZsDcm/ll5GL
JG1SwyKPrqvXjHXYC4DQnmcwJzzjEmofwDy7HW2th7qQ5rXxrk5yG/AXorjab+WU97ftfu/Khusj
Hx6smGmCdFF/Wz36L+wK4+aSa09N71N0f+pQuZBauGgQ055QDZqMcBTH2JH0h0Y4m1Antmw39U3t
cuNHVFDiondSbrNOqcmWyVEgi0kUmua4PoGieVN1rjx0fB7Si6OaOAlniQwkZGVYQxw9RLNaw5GD
zwYO72E4UkcbA0oQVCH+5/anOxIcuQcessMgztKGqqfnR9B8zmRqAfRbdmRGYZybnW6GjX0aAIR8
iWtk9EHXOVsAjdoMFL6i7zejJE5ENPtIN2A4RYtGDax1h69MwKhZ+QvAdj5XjYOZJ9g2Rv62ihn5
qL9RTZR3V8//4R6rTrW2qqqcrZxHI/neqSOApSlHgrnfKNmmUtnmRroZclHHfkSkPk1CwgJ9I6Dc
9p3AMKle0ZHiSqk0cE8064ap7MIY8+NpTi23p3fOqJRydc48yTmFIN3e17hKlq7aG6Qw/Ijn0HEu
121LNxdNk+56vXhC/fmgQ9ZADKR1DaH6qGtoYPyn1lSBy2TFbXS5f4PwnDBfcMuMmO89fHeZ88k9
5n5fkQLYy2Shl1NELuRmhikrt68jpO1K716F0JtRiyhcclueo8XflLp3ehWH+071HfAR1dUpoimO
6s9J9hHrUh/ulGqPKf31shhjn3B7mH/r+SloyAk704jZ7z4v8QbSp/ZAGk4iEBbWV0bMZNdGFeDF
tSReAMlN/Kejqq3BFf/Qv9xNIy/0duPk9KVStuecYAfG7EJnMUTmoYxvQm1cQ35i+Z8xjaE8U96x
GmK6AQgHEr4frl6Oa88ZsReXuNhSyKSSz7MtjI0oFHVnYxcoySLdjyL1gUydKFcAB0cattrMEytT
dmKtgvqEJRQkHcLQ1aacrQnB60huTScsLx0VxJd8MpE9RwTUCMAB6oXOjfOCWuGNN7FpJiEwj7HQ
oNCTM36lY4C2lStcfdxc0iG7U1P1/GGCJem6Xe986IM805wd+tRtNx2TAOGS0bjAigDIjcc+jTGD
ZP2BmMF/w4NbGURXiaq6bhw9QEqFjWt28zvguNNm5EzROsrD8jK0aGeEORLNKt9zT5prNoN29zLd
r0I/gMP9nGDeqp+hrPmmQLteLBfsmw9UNy1AGk1oGIL1QJ6Jkqldy+D328UGLUzMVoQuaH74AOo2
EJyUYvMXvHUd4bS5rdSoMf3S9FzxRVBI/Vaat9JI6a5ANN5dM4QKiEsSb1rpZI70GP0nXUp7GtRb
pW37Sj0DCtqq7WbFwJglxEwObRSnbl+x3jUb0DdsU0v3+Sd2okE/ynJodnL7oxpKfvbs0RGdgt7d
HrvqFNLSw7RuxXTZaTHmHxbKH0bNHal6zIJZshEAIvPG7jNUdSR6pnfotTiVBKyV4nEv4Yy3Xvuq
aAb5g+0yxgR50RSmxx5czHBEVWDZxr5MZwsv1e1UEj8Dk5JMqDGNZSiHjYVYkww2BA7o424y6hWq
xastRV3zE/xDtufcBfh3NnxYADvk7fgD3Zn4c2LDM1bRSUCax5BUbu52XTFoyT4o0p5Q0Lb8x2GI
0Mu9ggqczEvN9Jiqf/+YtrwxY1nNVTSswWkip+flM+70VPakn6LCSX/dpmk1+Y9p84xasMyJ7znh
CCF/XvbWbYJkQ3W3Q/+TBq+jAJIoEMqdZKa5EZbR17497EUVpancHpPSBwBpcIQSC46P8+tD6pyK
63OtiwE6Me5u9AiP25FtJxAa+m5hjeeaEzjPHiOwQ9el3zhaAk7bB9W8doW1NjmBAPVYwoRU5dqQ
DBbXKTvAj5Yih9ZT1rz3ccqzoUHERJH9K+vVi3OxJoW/TP1R3ioa/kNfHVrM+3IDm2gQCQ4vXhdr
OSCn94Hd+qbnzQEnzHNCs5TYd2qNsZQ8RY6ucCtStNyo1JFrEoGbeWthaVHk76qyu9061u7MfSwL
r8jN2VkWbtrx8Ne/ibZjH59KCXMmtrM6XbKwzyOP1CgYzmO/gjhGrSeCRkJ+Z7C/jceuQt+Qv6+o
9zez/DvOzpQltOGVN9DY47TQ4W6q4FnLbzE1dsMCcBxUMbraEhtY2S4ZoVg6KbqWPz+Mlv6CJoHA
Ih+eKLOwTeYS3kPKVgPRgnNL/eopD9ZYqXevsaNHS4vg/X5NkEPSb+jj4YmQaPHlTI7fbjzEIiLO
rveZPSsZcSn+zBWXP8R+Vylu/hM5Ye2epNTjKpuhjyWdvo3G1YNnxf8W9xanZ1xh2HNhIA414KWP
Rb/hBSq9oP6iMTb4U50j5XxO5W4JrFlJBVrqclC+wR/NT/7Up44VoIOQPdLEYPEpHbp7/vYRQjcp
tKgp8/XtVEceDqz5YMh112bG0M/XjZSSVWEzhHcjW1Lfd+ESH1DUczr6BLCaLHCcK8RbzGRugMMQ
MQyNDsQ0J9jQhpbKtPawdstn8tFLsRQl++dh2KQkmNOC77/rq2lFCou25+xEUdbSWEM62BZWxvq7
wL9KSLrVhiSATcsfFI/DEEFVR3IGQmLMG6th8rwN8wxbVgEecnWKNHB8ESToFPwEKDDblEs/Iv91
qvy3p2NSb/PXJK3C4J1ONKKgEk4meY9Ht2tFDIOMv0BrY26pTnkgGxtw2tS7PrPqvfjrlMhYy9xj
hInEV3mhXXHxbEp9NwPuHyvUczBk+p11yd/1Z58d9xYp8Pzd7mY403je7uRMl6OZ29n8pj6n6Hab
YQiOPmQtMe9ef2hJTy80NBj9ELSNKXIoTGhIf0u/qWX+OmbMrBZ/N3sCpsj1S/COIa4H09Q2KWW0
R5Yfj67W7iPqSIoZgYXhv4GXKnJb6FU2iBTEj+Pb4+VdU14lRk4mZigJMTTTmcwewnJw/wq9NZj4
K7uKD+WEf4kKcnICL72V6qiD6k8R/0Xrk8K5jFWqlbie9awKP36Zk0hg1CTDsrIshXTbD/nOfyT8
n5//aKgM3nZ0+bxIPzXTAvL11Fuv6UTxrhdyAA7qtwQu0GwH/5czFG+kmDSHba3T/Dd27Niw1CYb
/Ql9TjNuPWTVDjvvJJmn2gwNsCgP/rZAJn+6XrGsQfZeMOHCpqKSg+8YOws4smIVx7FI4ZM4IsNI
VyTMD0yIgYeY+b0AzCtMABO69fkUr68RSCmmNcwTxx60uNP2BsGfUf/DVMqMe7lelBFJl4RUNm7D
tOxkKwVFy5piV+kgWz/HE8KFcKpy4ND7ArlCgChWmwn/SFFOQRjfKJ3VLLEmZ6e46TykRxG4rVSg
FMco28nl0h+Cc+yQf7f1iQ0W9BXiYD5IL6cJFakCJucxpFoXeFcTaOWXLTyeQn2G5WrWHjXBSjyS
jxF+RwPt1nTbZ4Qg7h0jUafKDIkeSKK9o+b6WXSmVxTP9J1/K53n8bHMfTI352WpxkkehLftCPY5
jrarjnW5PecIZZjSVw0JtixDhxDeRzhuZAkEKT8yR1ryVUlZFpqXOxsg25ZBy9m89ngQrA9vyJyx
C2ajqKH++u5Bh90FyeckjFNIkVH2F3Klo5Oq8dXdAYCA9X4x/fNAurMC4INaBhly/MPmm7xE0pnv
YMRGD9JY7pdXmF0czpjdGDxF9w98DxE9idADGw1sV4BzLt3kNA9vmklrDqNwiHoaMoHooYXXGrvP
+op8m8cC09gk4pudYmRu3nEkDlF+y38GnU3/9TNqRRChoossISGj9VCTo9/cC3vXJo/OllKU8C/S
QUT+63sLesHwrtfMtVTpQEQ8cBmrDp+njA9w/3cvpj8vRh5fA2VzVvMQNhCKqU/fGBI3iy9G0qZn
RuGzTqbwox5TR33Q6ir//Q4pSWmd08aUHoM6keM1c1g86Woydp56bhL3iV2CSa8KwIBz9g1iR2wV
GjxUcsFV0ym1rWSUhg0loKhLgdUOMLk1h6bTtDQIb/oRqs4dbKeav0KWHRL8o4mLAh9i3+4UCPZZ
m7DbIsaDoJoxFQoqPQDGyEsKXv2omwIsLzBSuBImXRwFl/JzxqiBP+mD9H4RUFAsfcUUB6hTE1Ue
BGUq1xEx7s/o6ruNEOHZRHU5sO/ot8KcsCuD7PQunqBPtPs6dm9GO8W0hT7XohAzZDF2vxwnJ0T4
WR5Y/SG3c7I4AGF+SYIRSbZ1MUVYJ0i8Cd0awvPIqpRgxoPIAzmNvulCxoO4pOMOfZIaaTvt/KF6
TsBaVQMNWAuPIl2C6fTDXJpIf4nmHGS9UP9qyo05+toKOhWvnFLftDWkjUvT9ng9sdGF6e+VNKAy
9tLHB8BVGTvj3JZMygcBjEjIoF0ih7gsWYL1NeWAOmYHs/gDaOCuTvLZWb0j6Bx8mXV2XNB94NTU
FVPnw7x7Y/bPkDXmQ2u5IM87pVfBC4sgQmv90FLC4qojDakJz4YzE7Tys5lTe/jT4RyQsOAkRe9r
yOQETfBZLnLMo4FT6TPW1McKCAAOnd7ktx9nsQ+vgA476tMsmugpK/oGw1PSr/Inx8CO5B/ITG3i
HiW8iReJNvQXJGPBWW1S2rz0VagctNM/LwHmoDFfvDKFwRVqyVvbYzPo+hQuAVR7/Tfl/hg2/uyH
6BU4IgSK/tIvTfQx313mbDLQKC4J6X7YcsjysMh3nedx8smIcn11G/rQQTPfILHdqCyqTqjDaJyP
KAXH26eWmwfIP5SAr3G7KM75e3Dd38pffhVe892QI+1oIWFZstIAxV6l4vR9rr/xThrvGYWC66CF
QZ4GSnaBkZAUYy+9+LIAHlrmAJoVnQMSsF/WSvPWrMarHa616Jj9U0gT+6tod9GhBGAFgnEe97ED
fm+1fbjkDd/bvhhQHpzrXQ/QBrF5NO3bE3JhBT0e28rUqb75kBUOGj9GztJSYCnQQlZLiknGnX7j
Ag7NMOuqrIceFZV7Xv9cQMftLYJIaoG2d0QzikzUum5T1+iiP6w/vITQc4EPj9SAqg3aUFUUIbTu
tRXOr8B/CPjEowVaG+GY62nvzUT42bW8wZ+OsxrNCuuTkKV6U769U7ennpdKUXWW/CHgLABXo3dS
S+NS0idEL1vF8kgxTRY9Mu2tNgBlCqcEISSLNK3Z7mWEnrIP7fp3LI+eZ3mZbFWSuRtlrwfsPoSA
SBEPUMwgubdWrENlocn4X6KwIvM8FAbwNJkokvirYoDPoOCWHYO5XwZ3VMwvjZ6dbHqXZJIw+ltj
QwuhLvFJzxS9SMD/mOxc/3PiYyZsOMcmuDE6zaQrr8NgV9HdvkoGoDk6D3QE3W7ICalzl6kpnSIJ
4N0XhFaKCd5F+cVjw6Vo5JTr5Um/7pVLWlpKsycrmKjB1AcDIqlMefjFeKjltBQG3v12kCm9avGA
j+8L6ikv5STi3852IhnGGFcVAJNOqN9GlU0Ri/2vxM0r2DyvmScah5mFyne0J4V8cQCmytjH95A4
BsZjG+C7NizAu44K717ownQG/aTRxz6+uv5W9iApm3O2mkwAm37NvSWnzgPy2lgKwZAVzcjqc7g2
APXi4u5V4T2dSYADJtKpA2KiRAEuhFmTRgP9eq16tBFZIVx/uIC79IGPZBErvF8sYErDvsPWnT2C
ojlmTF320lE+z7HnCux/zVigFuRHTftZWB+KdskS4kKwrLHAi2LIMj3FpPi3AQA8as1Bpph3Y4/9
+KPK3p/JUogMKbQrI01fMCyV1GKF23GsT1r8Le22jUXOdN3S70nSZmn8xjUdwLihY7jh55C4GSNs
ikhB6Uobkgnvifdg5aIENVHF5s7vvd3w3nmJX8t8yCqxYOoCp4z3SmczNJfZd5JgfEBlT2oAhN9u
6hW4v2o2/fOAlmHbRZMTL4ncpar997doMc481UoAvM72GVi80Ifvh01Q04brzZRD2gskbj4gpeeC
cWBTvurNfK05z2LIvULcf8P9+lXyCMpy3KBKM5r42tN3+brfNlPQRjCdZOIKXx9pmEQcMvV7xyJx
M2BCOOJd41AoBpCKWK1jNEnJR/Hyeuh+9Xta7IBPHb8SoW+7Wi5sRykXp09vZ82tP9NqeeER+VhZ
4joKQjtPvcBbk6KkHS25WOMKokP55HhWysEFgqj0KEwWkzkxIkLTVrP563q/4lFrkp4ude4OMB4f
9dE4IAd5Q8Ifmo8TKFtvx4XinInPnZin0xA8QVoAe47HoXiuyuXuzrGsDKTrEI3oFI1I9D3u9oEf
d212VhP8Fuf6lWUUGvu1XwSVpmr1em9E8Sa+QOXZ55xf0nVuu8bxhf5NkhyK8LBf7QZ6BKQiAQbL
5FyP07FxlUpODZ4OjrtABrABYbwesf3N+cnmVFFzbMsv6I8EgAKXyLBalpJ0gLWsTiVVou4KydIS
PXkKmIHYRVFUVmp3xcljF5AVeWup+e4ZyMFjO6O0/qlOl4QnBINhKtPZh1KJz7eQrCVMUVff1Hzl
uJji9akzPk2N8fBVviCauhEdsrKeyx95LY77B2ijiT78dMFo1+VfYfKfs0MNEQ6T1UhHQUXjG32Y
/kJXNPe0NITax3QP8LZ3jsDggS9RcRcFEk5obyAFc2KsDMs6F+0JJQoadADbnbarL3f/rqaCjK9Z
ygXMH/MCDqkyPZ5dHykHhOEJyKlaPWArHGq2vAIyHqvy60fpGU2q7Iti1Hdh1LFSc2Be4cMkKFoF
Sa5wpzCQ6Xi6GU4Ev2p8r8g86N9K0BqSjqUTl9uozvXhOtUEBMWpQ28hHtQjcE28fZPicQ9CSQQw
qusZNt315MH6tzyLsQslsJBxCvt6Bg8PLpZEVWr9/40YHgYbCoIItxL/JyjEnZBf7N48WAz+Eh+o
scKRNq9XwabHObYpTxRK7qXHD+WsBBW6PP9Hf77sps5V//kiUAu59SMZPH3i2s3rJdnS6dB0t7Ka
bs1pNMPxUpESrWsbkgqxot2exmqizhdiptYCtJdeRQPconJArgxnyA0VRqIFowhh0ykgADt+hiRZ
qs3jXp7jKG8HVePCxkJ+82exDx86+8fqUZnYUMyq6cMPnlGtoOVeqDDQeWQRtY+5hLXkGQxFJDU1
UqYUPBO/oN9mh8sO+vslpmNDwx2ohj9XZP3sBFlOZpQGEGttskda+oHWJgk7SC9qUmkkOHMT2tcV
AOkz0E2SsjIWN1eKGYcghyMm4WN1FifAalXMwa3cG/wP8/lmEDmU+y086kAVgKgDXsmmilHK1i8t
QkNSgzrQM87CmO/oXVUDEgWAT5DH0XyUa3EWNOS6u2vl/pH1MaMdzG/MTgfdPGi1m4vxpuP/xJij
ORIaD21e70YmkqRdYzl05I/QWiVAQ4Kn47V3bPgaOikzVvg03Vqa5YFjLhOzTWxAFfaB2YeXKjxB
nZaHB4Nwu7vLFUBLco7YaktfEVkvEvBIHEiRGdua4JJUTrF3LtXU0KvJG+ASH8fGc5p3Z8BrsmQZ
upqphmGyaJZMpvIGJnV7HBCZ1Y7m35KLTLXfVUkZm+UL8Bsw8tbHUJJxN02AX/hTJ72kw1o7JIZU
Zvyp2fK5sgAOUgvrjgNVs8Q27tfd7NtUCNe6I7Pkh5/szfHUi62WSzlJ20zyhnQx6uh6YnQf0DEa
KV0R+Df2PlbeLxFNJouGW8LgvSOTSuHDOY4/asffn9mAL2MYUqoOYuO0fOEoKrkFSaIvtGwU/+ju
rrWqwwSPsv4bCwvNvX4tDwyoHfcm2s+vkFpjyL/BCwUHVj3MSvCIG5TcqqY9Pd3O7H6GTov7XDPj
bq1kxU/FhdSRKpB6wS9/OTH8bQopRJM0bDDSFxkMudh0NefTHOBX74xyN2c9Rw8APNTAhIBETS4X
QnR+szXOddkBDRKgwo3F2RrgnkJPuXzk/rNqE6bVdaT77Z5JzAWlqxUSX9H6421FOKDdmSMl/Md9
Xsl33va7ONkvKmKmKPGzwJQryVFp4GMZV24Sjbr8aYnOG3BntmBqa3HjurywfvOFzuPrcfXQdgnT
ZdFnbHykVw9cCws9Wy3eA6ilFTG0bwqfhU1/PTUKg85n1zTEMckSJPpsgyp14OKjEoDcuLSHjJ+e
PhhgZTXRLihwJl9cn86Y6DjyaUyxm/JsNh1TaEhzgiF0Fwmz8TcpSsastTS70GkpUTbAvtuRsT28
zbQQNdR0Cq1CQgSAA28pm4cuw0wwNBMvXEcqr/vhcQgVKFDNGd910Mvcan45I7f87//5ghzUeIjh
F5I/jaQjxC+Am7oxRe2+y/Sh7Sn2p5Zu2auofSdIBJqj4GdCEt6LCOTL2GnlEGH5rlSxSQ3HGNjs
uMIjp/ezFRq2pQjE+9CBaVtSrIcwm4hNR5K2pgwNDGplS8UxAS3UIhe9dvBWf4q1ZXJXMMukFUeE
dRPuBXPJAhlVoC21Z+kNLign2c7R4JKBRSJRdEzvYC0S+H+ws2kI0rcxZLhw7FRTfLEa/Py8qFiN
DTNEMUyql2zZ+l+srSXcvp8vMOjR8kuLgyo7G0MNAa07gGuYcid3yxUNCRfaF7fwd3uEQBugUATA
jglGEYuMbHmhkc6L5/Ufps7VdPu+ezGQet0/YnC+T24k04iltUlzjiQVTTEf+OHK9STzc28s1GI+
c9+a1kifNwniPoVZYlfoqQZAwWhvJaMO/RyL6eLy5K5iCPtvZSHk50w3YS3osbMM7MpW9zz5MSm1
9OpGIvLYPVPqlYxIeBcUVSNgCxD9cW+1+a7YhwgshhPdR/pf4YhpnsqI07xI5gB3qH7q7AJ3R0sG
WsQ5lgwacLttBEQRN0JtyQmIB9cGYBm5JECaYRq2M15hPI0HRqRPqgvMKEhx7YoiHHN4wcyPcGDG
mstaA3WeraobOxhE6yF6kwnAvRiA14rakugse8TJh37yF8LwSPyiF0UykdR7KxvAr1JTOl3TNLAK
P/zGGr7THI65QJ06zgP7vAjq9TbNBZ9OUyKeexzWbz6iahgrPCKIKqqnVoDnTYZ2NVIXQmdGCbYj
TF7pcN34zXUF60gDfz/bEjjRS/miETnLtOsCm7KW+FnILsYsIyVERBjTifJ2Lv3x3Y3Uwonp01tQ
ISbbnOjI+8D+nGplJ1VBRa5Y0sb21Rjx2YOpOYpmEt0uAKf44KhVEyL/NHzG3uUGN6iZmB6qpEAw
IViX2zMLKJuuDLdcNSXg6HDtJl/i9VclnBDLh4qOfRtThpuoy+zEh6SBGUN6bbJsaJYvbrqAN+ZX
Rqm06h6G6sl09Gqnat3pmtl847XxUYv2M63KpWwyjOMN+ITZv4Anv0qXl50AlgjXx12DgxeSSgdS
/nBqcGDb9/NlvRMI9WLZxkwcXyP+qyrFJYUQSy3kdSdq8h7HUdK5YlEHYrJ7rW8zvtrRjcnn0Zaa
ridcOV4YoW17VyNOP05FCI0T74iUtTCc7k4DoNnn5ef2Hi+AYqLPRoT0JaarUWtt7t7jDBvmnw1B
mRbjiNHk6FZXjqOmdg88e+8aobc75rViKQefRzZpJ4rvX2bVmVWQ22N2PfLXho1NjObZGwOzvm6t
1jbWHnivgqtKLHGg3SZotZJe09fgIPFlzhrvdaSZ+AkSwoWXbRoAddi+kjuwtT69nWbV+wEKS6oL
Q750JlsN+NVElcNhqtfQeLFY+DZ5lZSpT82HrgqAdyg3SAtBVJnkLHQlTEVxoIKvPqspgwq86HOd
/rAYuWe0acXENPZmewmoEV6eX0r1bu08OidIPsHSiSo8l8zop2qTJnirfZmQhd0gYMCxP4+6SivK
7kdlviz7nBewY3rU1GALo60J20Umi43rZ77Wu+5RijbUqz3u9xSBp14AHAP3qzEK+olvBAAA4zpg
T6uDxagCHSTLiV3l/0i0i32D54AXQooUVSP46YuIkPvoePtP9cwCii90QHJ+EjxBsKaS8TBw3h51
v0AnGUDsCvDUHDxA0NJBtODgs422v22RHnqwjO6NC/PHVo2c0+Jviu2+TBqV5Anaq3EZ9d6WkQTF
PAby9vSf5Cw03HXQobMmsktkcll66XXukZ2Aw7LMdekcgaaf1OyypLREfxg4PhL3C1b8BQTWT+gh
jUlbW0alJcPhmvl0cf6cmdWYk4xmOpmrLY3vPtwBWuHLcwCg/T4gJdJLyCdKoRR8ZNcW6ezHK/Kz
UN1m4rg2rEfq05owwjfOw/+VwoFBGvHuxA8wQTQbwOFGHiSxqCO3R70qhKjVTUOKFipl1NgkGKH7
dmwrceFxdLZicxiv4msXZoKrwscKTFkYHdKk8frVGbTe2sPg+aaCZtbj6inmx4lN1jjIe84SRPHZ
89xqJqUf9zfAXT5vgbb5kFmRnUPyVKe/nJX2iPFmtjpF7aQJUrcPJDeCOUWPS2bKawe1iMRjg/Jd
0xu9phnlCTp2Msmu8jmYgzDpIL9jMFSe2G5DqZZ2DQHGFLJ2OC+PWwtsNASgcVycYkGLKGbpFRL3
1PxvlF4k54AxcV7hi2o18EqYJ9skAdVHzxOtmwGSsEvmxsRmRc0iRpEgNktJU1QHMsc08zLNuEdS
pNEQNMiYicSunLTO8csYp0JqqpZGldlm95lFUq/wvF4AzPVU0/qn4Ex2QxXRlATDEtU7RS1Rk+H5
9Ijrj5lIex95WjqUhIdnQRTxPcOw0rupQ4ydpx+wMWOANyk0tI8NpxtYcBQe0ML/JTasqkVEKIhi
H5rU0r+t1+L0UywjjW0qYSM/N8RQtEqmrpTxZAzffgnEHK7mslVlAH9eewSTMWXiFCRyrnUhrGhi
DBhytYC1W1KrE4wgbdgkcmI+kzuzv3PsEDOV2tX/2u8+RzmYqgUaaI4h3UonGZJFcstai/7DP7/o
MXjt1JPocn+TyiFRhDGLRwLyqPLjr3Nw1TcusC/ncE83uNCs1LufGR8VogXxCueI5XHIfBv96sZ9
0wk6GYuAvh4rK0xd6fW+bWpvTGa8V5EFlhLkOwujlsm+wmwSFTo/GPS5dKgqgZfDKUYm0zIYkLAc
68G9nbraVH45ECWxg3HxJq+sg6vajL29a8ipKms4m1Mp3ybn4PrlfErbyHPLyEuAlrXMjSOJimbx
pC7JXw6IDiXanMyTqgY2qQK2JLCVW/65fVgDOZenHYJb8JzVh3EpP5AUzs0GD7z7ukX5yXqRSGfC
lpLBIrlVHcdwppl85tSUoo++sgLHrs5fdTjIlXDk7k3+5n/LK6O7p4TBHSol29znMrpZCDoHHnEJ
ybMJXQMLAjdFZmfUSkYuPRfLRG2w2DGfww2i1EaCfRmMVWHxHN+i+kNNHkUZNSvMcK3ZeltsE5Vz
rEaPr+h1ETdreZun2UiqixxPX+Z42DWuWyR2DdtL6rgytkD7yx+0mBpzCh0IWKeHLp2ZVkN4+uOe
+f9yYItIIFFGLLhubcOgzBwH9ci+5KhGBjNzgr7/L3N4ysQqCSgH7vKDPBmDdOZ4wxYG3ZyTPPvE
epyPgkHjxw8zvNyWo549qVZz6GhC2JUGZf5GjcQJqJ3SyZACOu+tT+b5W60A0gT37e6EERZUD8+S
MxV848G/vTY/ObNeirsPk5vx0eMMAN+hRXF2vofYIgdpqqheZ8+NJD7icmAlIPZTJFh42JSZeSdh
YUzx7i82jlDvjOxB/6Gmd8stnpty0ASAkV5cumjVapz+2DU18GdfroHoKb3w5eu2QzbTN8m2J53R
s51pDhE7g5rPzNMSji+CNGVmT9ek24lCCqadPuALfAduW0CflWGkukpAak1xtodl0qTS2Sd0J3HC
saB9fB7QIiizomq/UgHNAw/Vm71RjGSkf2wG2nqnrtgzECQ6bF80ggNhYZTAdUbKvwhdo35giQCX
rR9Wt64UytkJofPUheBZtV/l65VFhHZosdprYOzHamOEAi2hz99v3qRcw90wkE+buSElP8ya6sba
g9/kKPOnJT8C4cAIkZncwfsQ40g38t52YV+3K+vHdJhLOhrOwRv4lRo1mG0B7qztl9GH+AuCMN7+
y6MfzKFsqP2TkxZ208TjqxcZ+w0PqIMMKaYqbbx+1Nnu02IzhWZvQP9MntgmMPKRcKGXC63RxD4A
H4gA7xFQeK+BSUeKBihWevHIXxkRAVZ5HrHCwKizdqbQv5DVFREWqcKydtyEVYVz2TqbjhJl56DU
i2P1OjAVrb+7LjzdpgXHTJAkIsuEETcB+a2Mq1zBq6Hc6tl0WubX7H9LGVIf0ou9Le5gz7L/1zqp
0DeDs4B4QGkDAjTsTScDsX1Uoz9g9yTDpKv0QHnoDQlPnGH9p8lcxEEn4ITs2iU8U0PjctxxH0Ok
tQyLhFtWJoYa94/kF8OEfRTorGACS1KhlnFHGmWGZeyAxdzlezjDvIvpB4H0XDryfBpyfAYFFnJp
5jJvCRXcSQdMjeWUW3+VJB6j5xM5B6US+mLwsUsOmrx/PX0Mt3qHN/JZ/7wnbWflPgtSwuUCu1Yz
pdPNKn+3KuLlqdKeLA23oqWm18WK8U6sTJLUt08U4mMhwSKMPGSLUX2PArDuXEl4IFA3CYCAktv9
aD4CHl0FCBFcFv9+ig2VeNDUaPJIRPPciQYwoA06x1K6RfXjM81jn5odxKYvivxI91vjK+jethND
wp3rhuw2WybLm1iIGxnXQGAEYQwcgXoWQ8GMWjXvLEp3Bn45A15QVUo5T6rmXXD625UoDab9hw1W
3pRoK4B9KsJNAzl+5MmJes56jLgSZ0scieu3jQat6KBz/Ksr7Tkjfs4Npxj1hv682WXvlOWH5bqW
mQcW+iRJifc+NvnAxyGi4z/uu5yBYHMSfm+3cw1bCwgbrRS42JqOHzbdtZc+F5ZfGu/tS1z/A471
iLKpeEICJM7YVa39cxRjstNhE0xY0+siH/UNOK6Ft1/cvK9ZQXOa57LWrFpu5haEFUAHwdpIXgpO
jKtHP44ssTyYXSsGu5eoWBvKNVXPgVgP5B/QiLlkwk3viWUvxdRwLt4zL1EXAyeCRmnwCPnnIidv
tqo7CrLsw+NCavoroWyN3hfzzgO+mk+kW4VJEgat8W0ZJX64T5EBH0QleCrFIM/C6ncEqSq5EPmC
D7Kj1+ZBTOvJrxDQ96Wweqr1+HDmSMuYSDbH+lnKDvVogL3dQ8KAJ9NFV3DMjxIBHBUyggpZaGZs
nNeY771exqGdfLNzw/MvyDUjKGL18ZzJiXN+PKOQQ0ACDzl+fJ5Kg8vYV8q+V6LEveSXwocuyp4b
04Zn9ONIdHrGsc/Hwe5PiK59JT3rO5TphDZ70wqlM4zXJ2Tv8Ee491mJmtbtB43ed38Uon20FQPA
xfwt7bDOcaju08jsUGpHRqgAyp4dm5XvIZNXjYoyBcxBeHXOoTEZYzUF4AFTRay38wSissiDyA1o
3ey7K7ZYq6CIE5ujoeA1RMp8N3m/6DDjQDkUq3fuAdjRflWPPB7ui+OnIBPqrSec16grm5GSJVsj
tne9ipqA2veZVhXOncmVYYKGHlH58U1mTDIG2GrGPz+sTRErm+prrQGniriWPqVMdTz6/KyZBvvB
9R35hI+gpIRqxSlwwke+1XaXR5tYvOePnfdIX1iQWaIMqRyS3U6q8Fg37QK9iMAwhER/PoDs1wh7
j3/sBkXTClS7BQHwtPczI0s+E4oXfkIo7M6ZJI7k5/XxK0oUhwObyq+V92LWHKpUrSBH/LDeqjIm
y+pVygk0o7NFhKGOaDF9mi3Tubvulnd7K07HgUwXlhZ3C08YuFmLAHNyMxlHT0+A/wa8DenjzLF3
KLPGKjWJ+z4uinhq8D1HySMDQRHiVjCXdiGtHyuTbm4wq0d6W5ZfDHFOG8PARZ5LcFFPQlVQpemR
vVlFYN/tKXrfDlSYlE21h4iHKIp+1USCh75tAjxd5q47/0WFJZwuXKIRd411AuD9NuJR8nLAOpv3
wzAbQheK2LyDtV38wF5dZH8qjyypbK/CoL50y+xOewKHkXngrjaTEEX7W0g6D147uE+IBf0mewQn
AQHxi8BtOfRvZQ7zWxFQb8f9HA/qOchfuKBN6IUMe7+TMh3100h8Kxzax9IlRuCOUk8A+Y/IgYdA
N8RBwsOLd4ux0pR3XRm7qHahVKA4gN0cj53S40Uas46YR7trpZq8XefIMnzmuP5BennGWLADp8PV
3/9d6X+yGymnl8woR3ohf6cIjcrTwoJ8P/cLo9T/vtqaqyelu5C297vRhvGgJzRVV95FcjEZQ13k
sKaLCpqGgLm4cuoUIcqMj0fFkksYSe0dPNgUTvmW1ZgZKGvLj3aWVfz8GDCWy42n6AkGhfGB7os0
dVNT5GsXTlWj8qn/I2in4AMAw3a/faoSsQD9sH/jnaG15dw9r1vDqjHc/M5mQUF4/nqTeKwLcyxi
hvG2pnOvCPEesK3kGPBJaBbt+iaHvvZ7EdwwbujpcfG0vc3pxJXpMjVPBQlHuR2cYqQJrUN4DLhL
/z41ibfbWbDpn9NjWJwj5QFlkiURJJcFV3VtjBXSVoSlPD8RReStCaWPQTl0tqTDuyBBQvVAmryf
NPXHofvGEf97WO92Jp/8a6JF/THJtHfoGR+/ukQwd7lBumorLdLxbg9/mXn7IENRgVJFYc0iNYy/
lZ5OUGuDFsMxYzD3SqdndQyDyJpdt8UyWXRWmD7Ggn0T6Cf7shQT7ZFQLC1H7/PEEB6mQD8vNojs
TkaBLkT8j+pd/SOPn5wiHvRKB6I4gjzT3WSxRdRYdPrfVJlZL4VFSAJ0L1Lh0PGXOmIxXiCShQ5M
4Ros3rSbAifo9lDrdz1M1DLohCK6vI8GnM3Bhl9Z8vTE9Rbyg0KwcLg0FN0bJGMsBIfOwHwHP4NP
sO3rwUw4UX5jDWBTQatGKx76MKXzVPqXfaqG1AXv7+dUIPCsFrP1YG+eUL99+iZ8aPEeXaPDFplP
lXs0h6zYnuMunkBfOu8quCRXRuLsRSi35Uh+hYo3inK2Dtcj6HcJS9qH7GDw6j4LArJDMZHxvyy6
dFFvdLHaNyDXsRuQREXbAKG1vPK27igfT0FIUx5osMFsiKVlQWwzz//3vuOZtWCf87zuCVfjfFcL
/N5fJMkUTSg8lufL6NqY/7d5iaEx4PD+KwtJv0BWS8Ct8RJfmoNmkF84sXE5TzUsIpv6MHvsNJsQ
CJz8K/FBjjYD4fHOogcGH39dSM4BDrjARcSHvWpwaQ+6VYXEFeNiGN18a7hRddetdzvku/yblfbe
HsXgO0xSOrbjhbn3xgd9Pd61DONM+ibiOJQfMSPUpPYa1qiMDGQ+jwJvMZBJodMuvLf6w/w8lYsj
fvGLYMrNpp8GB3I9kt3tPzXDL8WkbEFkdU+Pfx1hoz0jO9pLxReUVRY512nha204IBxvgcSj81oP
0FVwT7RZ5BBZ/qLoDnhKUiGGDm9DAv0YkRSdT2QsZVTTZSEIydqVxuIRio9YTF2YC6Qd12Zzpgx8
I0KeVV7DUftItCdcc4MWIRPw2D1g/W9ORtoad0MIenYT/D+UVK//g53GZb+R6NHyT1Qs+SrW1jHF
MMole9eJVe9THAcv17d+fQRCT+pCmG0V1daNQaTLIOBSxVyvKeFcPvwg11BqNZttjI4XuuyDVF3i
/c5XIpQ8q2ofCdb8WIJYsAslVY1rvGBFmx8AW7JP29SgkUlFL0nqNx34Bz4cHcUSEFfN0Qw6ojG2
LlQAUXy5KEFWmqJn8j59UokuOFOQcPY1FIB8v5NxvKfJPcyMdhjYtW0dP2Jyk1NNuh9hRKpOzxuJ
mWZDptsEMaJwLtgBr//AMyH32lhDxeBTd0T8cueC7hD0tgb+ew4MLMtoPY/06GAqveMZJ8/kYdKN
bs04IuMfAjiTmCE71O0DNz7uxsYUqzv2Ixofe4+RhI44RLYb2fES2nliCFKS4CAPtKO6Q/T0Ou42
qPsy0E0XCrLTdf3VulYvecXTnDm67IO/dqdEJTwykxSfAOkndRJZbhKcifHrTRg0dez/dBfSr/r1
VM4JfSTTcuWPycDR/xSYIGVDFQEUb7BpQG19BwRaFAlxc95dLQ9EqPNSWVDXjk80Tk2J+P03xtKN
lW/t3bk10uFbScW2V9+fkA5UnUYJdsIyKsGc/ZcWLZwRO2Ic656rlqkX351SGKzYkSeWkWKOPF9N
VVxL2rm62VRPlpaO3hfxTsDASKfIR8kwQPu4HKdnlza9VEBbpF7Qtxinrw/PW1MpyndJ320a4ZV6
6dSVoWih+LM+caR74hzVmiCNEIRRq1iFwxqUJfiwvQY9/R2W0187z+erRG8GHwrN2I+XPlpCVqDr
p4G1uy0751OdKWQbpLQEbHbS7w9OBxr+UF/rOazPTrDjX0LQnbYc5MaD0qu5bhPhNzE/34OvIqYj
MEHvcN4Oo/cwILun7oaYKwpUkUbySTYYErHVpR3+k2HMSG+i4bJLaMNTS4orBpf1Qr0TVtwkiqTY
4pOWd86OR1kr3xIpm68nz6EH3dYqr85FRwy7GUqfyj/2ApHdNkimULmaGnugqMLolS/VUFkYcHpb
v9amNE9LnTkzKgdOGv9pzCSf3AqucOwle+atQFspVjhal8cuuZ5f7ou7dJm6SQiZpyFNGPbnMpIr
Q3BqCo1aXAABV6u6FASJJhKPytAGKI5Zwi4ki7ZALEmFwbwN1vXyXYR2lS+uxlAWatLmXg1T8hm5
uYS2Zthkli9Wd0GAS0RYhACVphbj4EFA0WCU2EGFzCFnOTk3+3GBiWw/UfpVvQIdCP2d38BNXzAp
XB4cFYUo4Sr+9OGcF3ZTsM0fLdH2zEOunjrjBbZcddoCTYbd9yu77TANolEB7e2+fZkDmc1BXfbz
EvelU/K40XJfzoSnIF+4sb18HXjUPFdqkv4FQ9AF8GEBbjiWSWfKm2sdXrgDqzSWHRcpklUU2frS
Jk7wUsxrFM/ivKVLt8qOVQCE2sZTXT1XS/GFkCnxJusMhZQmmXbLDR4EFTdVsEyen8vSISAyJr/L
ra7xujMiJF6CM5jQGsJ0q17Cv+VINTAUdeGsSgBynjA5POLOZaTD7+PkuV4wwNnxrA8ok6jII2MY
lgThl0j6UMyLUy0EMrVvsrdvJSKOjLJmuQYHG2CVJSHajeM4AJqIKIrk7W5bhRYmuZHNdMiA104v
gy2HKviSR/pHvBoj6H765VJXLQ7cwlSw1Wwhio0nknmuLVDRGQ1g6eLfknwSbpKuzednN1AGbjGl
q2DKTiInKVjq+0yS+jx0CwMIp9McRI0bgfevLYnT6o2GKQPFn0ixgS6MW+e+1v1WsG1WOqpzVg0G
hD1dKjcvr1GuuKApPtOCHYU7KmUE/83IqNQwwJeW1VsH4c9/OVuUg3wYWnP4h70HOgeizdTFkowG
/Nh1DIatq0rVlDoPGwHFUS7HFtNVKlmtA/tHuUw/CrAHlgn1LCQBH7H5M9NDf9Xawds6VnG96X5P
kkU9/P0sq4AZt70IkQ2HyMSCO2G2lQc0qfdfudqQ6G2pOJBOn5eYV+5KKk6386k0qsUfPbq282iA
zwgJBAGnw+RqRhvkaXo/QgB7ZrtjuQ76j8/AdPfOEsr0v7qmzRYXD/B25G/PtfM/Huuunttkb80O
c0dytpDDw/9MfMQP5Z879ysrTai4VLO80ue6BIXBVkJ4nxAMbafVkK5GQBeASos2ob4XUa/zlKTi
jBxaO740J2Bkff7N00rBNKPFgPdyd688+lFMEIDpSZHi6kgUIILRXzvl8x2qIvTfLAW+ImU1kfez
smCT/cyO9klVRCeWCEDj6zPZnVG5+xPuVqJHjA7uCtm56xR2dDIL9Re2VYgUcyS0Ja/kVEta4Otv
IMgv8bS3Q++q/suKfjnenYCQqmFmfH2WDVxMv2gMZkRg9WpS1FTyex3FhjWlL0MuFJEAFB5ZLjyz
Is1fvwWL5gonBAOd+BK9pRaAvdCprRpRbXBzNfzzYedm17usd5jU6e6+r1rUEpRGH9tRVGbFGt5z
Z9A4zK3FuzEozgjsdu9eDGNotve8yGD9zqvXbpO1z0XfZwdILzqxzKZYmkm/ErXDeZnN3OsoEola
mbIcyaM7kqgfxjKCiQP11D4P6IruB/bKRHDqmNmUuuXJE7znwuztm01h6qNot4G+OKBOlCZRqUnI
qeMv6WIi49BC4UMj5pLNYHK9oGbFr3bSEkGPKrJQ1Vnsnh/nS+qy7iaOzZf1O5thTtHoS3Niaeqz
LfxxhhBwm6rcSVeHbBlpQZtTeISgx0LHOuDTJ3+Ok0UvS0cfXZHkhETxn6Upj/Rh9I4ONcm3atwh
AiTCS3wpRFoOQKIQn2mjvLfkmlrzip1ITiG7BGTrIVnah/XYEyjPKoPn/KR24OiVhV4Kl5T3yKrs
g3i5pq+HjAU8KzLyPtXGU/ySPkPiDAD1kgzyBdRnVu7BfPzsKGtnwO8XUwzgSd13xxWQ76IE3uOr
zPklS+T/94aGnxeYs+1qu7HsoYU5Fd2HjHvCzY4QfbJYBBjdV+Rv0UCypK6KtHhYe/w0r8OWj9UY
k1r4ZxvidSvNmXPt1E6d+GIvztpUcbigPkHCGQYHZsOyApn7HIOdczd775gGVdFjB0+wNybiu+nP
STqBMd1vV+lbXrClTMVGkBBXr3Cr9BZLyfMKWByWLXrAKawRHTMr3rY8ZbpKtww+Z+fIH3ETcg71
2bCBAWUAOJelg4R2jH8O5rTClpcx1IPBe0tZpcVZWO4Zs/qFShCJuqeSOamTNwQbP/5rMYwhOeh7
fh3sYnhSB77aDBByyMS+XMA9DvLe4hfbOQ2BeXFHo3KrfHP5xKwMJQtJbr+jDMxbE81K98sGqYdA
Kv/g9bMa2b38W32keFjxsYwCh1hdEpI5KeBQCQqN2HeTmIbCnq5XGE2JTLMCKyJEF+NHrzW6MfE0
4rhYCqEYVcwFufcGafPMADphDh0hX4pcemSpsiTG6B0zIZaS27fWXhtSPmR1+VeR+AFoT9QP4V02
eSEMoMJJbM5S6wIjfspRuRBOSZEYH8nFK88YqXKmUFLsSGdGENjozkGsQw79WuyhFRWEU31oaOma
Nx+b4vcJ/mvm5F6LERUtRwgzlAxSrgg5MGwqu6pLbKfhimk7LmY/CG/kOjJ08qyPlV6DTBWN2+mN
YNXs7ll5It8JI+/uAa8rwWokgAWWdd6uk0mzzqWRBqdSOmJCI5vyM53wJuvDjGH2YTmft/0Lhx15
F2/SyrNfR5seXzIufTHDOZjdkHJ+d8sDetDtbPQaAurJI7vC2cLgfhcIZcAVNT0AfoGP5AUuSoCG
Z+zGBYj3oKuLGNSQH5yQDGsvlwxlEdB2QGKGWvsgdwTgSDGCuTdS2IpLqkqVrOoJnp6sw10u43sy
JRvwpVKCl5nV+TebvzGXPMkA7LgkEUxqsL/BYI1IxZRYj33CgurVGwQzfQKtRZg8li7QYuQ5Z8BQ
uRGqTLbWEw48QtLyTaI7tV8F1B8xl9A0l1pEeXEgFW4rJl8NsBe5ouePEUZHdXZStsMKrpa1TcI9
rmeQwjO/GFdGwQYyCGileEgxIyz0bE40jRuByYJm1BRy12UsSP72JLDsG8jFedcn24YVnu1k1EBr
M/PYTwddaFPTLOnA4LDTio/cm1Bvr3Ro+e1hqNuiXkc/NGvbDDYdULJiHDyUTLoJmKv5fQAKtpad
wP0WLKwKdMYCtgRGU9onBG8qWwsouiafIgz7dxHKIEu3nq+9UOMbM47dX8ahwmTS37L7NDvI03Qf
2goNwAwvo0W7cvAmWjs1Qjmth9GGVNTyiPO5obvxU7Nk+eCTpTE+xCHRtZHUpPqa77tdG55wqDcN
J53mdBmt7ply2qo1Ek+22kSZJroWW9yH5pEi0/8AiRAb5yGy9Go+qXoCX8j5L/41G5gdjpSFhcKU
+3CfcZdvHrwoCKYAzNghdHJRoIYupWrWb0TvXg7SVk5ptgA2pOhma0LAPCk3zTOqP3/ZZUgX6tJH
xONddbQO4IhHuCmTWnpp3iF2WG9F1dpf4UvmL+3zrXNROHA0Pxf/2BsttqU/by1SCIqKiQ0U0SgH
+chKpxzlwNWUBGNrfV40ng9HZtp6kACcwiVZ38960A3UOnja7foggRN0AHO98OZLtuY73iE5Z/G5
aG/ec5WUQdHCZiyz5vUaY2XuNEcwm6M8pCIsNMOpGXH/AKEezkVoRPeUz2eQkqLGMBiAN9GCZuiQ
Y2tJo0pnniHDxeLITzF2f0r2DEg6Oql0CtcIJqHEbk4oX+b5ZROQPw+on3QKDbc3FnOjWax7VNCB
/1v4nGctAX0yoevSQVvh4liYcJCRSD3oJEQoEPb1GvXUr15IA8Qj8MNGGSAU0zlt4p16pC6jiKWu
yXi9rw0GHotXYMVgBaFA68fPntP/glLhLMImEz5UbQ1yaHGEyA0KJoA6L+lWVvGxs1g7BAiYQY1V
t5dGx8SQFoUuW+Ec5pN3RaQRfM+UyHtdqy2QoNNCIVPRLOdCsOi94VryHBNAmdIuYavBewonLTcm
cn+F/Nr8PCIxrCIJbu0K20/Fm2M++cIW4fj+dtNAnMnoxeEGFm+jABWckH0T4V8NRYvMTSwx/mot
8k8v3L/zs4p1QNf6hiErvK8rY0PRWY+8lGlQ1Fnp3qiYNaZC78hdpz8bHClImAbh+mPjhvfFBBFc
/071akdec8VcMVq790NgT/VCWqucjc7iOQfkc9HRttOvFhViENv/rTruF46Er8JJpYbMKz+1t5cn
9Rqi4W+0FWJcBVHOIjMlD7vwhM/uWLCvaLOtDpo2ryioTzTgkj67lhAeRKOMKWHrdaQvZBVYlI93
yZ99/jGioKbrzEhe0W2bKtH/ekpiF0xYNWTmss7ITJ06hthFzzokGh/bkozFjM8NxZsAFfyWXsqg
H7gisWvu+1UUiwBbrFEBSHl+9O1E8gqB+BBE5xajyJoEHfXLPA/v00IeI78E4umSJw315br3yFBw
Kv7sM+OqUYiOus9Cf83ryUnRlJ4j+aqVqo/TZIF4MimqZkTnJtiu4wdl0jmfZ0mnR0T9jz6diOBG
iSQrO5vDwX7ElnQ4mX7cvSt/taAd3ct4JwmWlIXWKh3s6fj7fQez1r0p2kNBfFC7l81vMfJLcEYx
mNJFe6T9sMlCh8CDlW6ijjV8NfY7YC4xhZ/1ZshbqlSncF6aWbWKIapfUWznV7nRqa1DNI91OwHJ
+clDqgSNcRQk+LjTPbTGO3IClJWhQJZCM3cxqeI9UGUMIvQ8Px09671kooaC/4y/TdRzJjNUB3YU
LA3ZU1NM8qtRgk7ihR7ocRHWghuD5shtvQsW6RlAoiRU2PbNPT1pbYRALN9rtkKN/FPcvC3Osbh8
F90PbesCx0NWjZsicbl97P8mrmfmSc97cyTG7DvGa6EhDEWC97Opj+7MN14dtCPdfJUjPOWgmUkU
gv7LVdFCFk/89qXmurY05OGfb/t+mrW2J48E4rNdl4eK/xk0jHNU4uu5rKr7F8J865INWHhIUDRO
/2pTSYiNT+59O/rcKNniOPM8h6t2HIzbqeyFZrRQRPibxwSZphtGkc9rzrqKT/2hlssCRYo7zTuy
/sj17rNpJ9oq4Miy5cZYxM0WP0DZwM9pLZWoul1HmECIGMIZha3rcb+4obNWqAUoK822YtXz73Jm
e6h2pn4l9mg+L/DiZXXloYWjysrknmajKqc1mCC8Espee205lDlBrAChoh/AqhyTgJHLqowe1qmk
fKySaqqZfPloxYMYuq2Y19WAI0cJL2e7lPW2czJQwu7353UwgbD/e4/27KY6zDNLjm39bw/PmL6l
wChgzGORhHzBSnUL1i/GvKRtdXAfPda3Fy1d61FZctfVJsvEpnxTn5De1pT6i46TK+AX3gqBWzDd
CQVN/90NL4nY4uG1fN2wjf6SPutz2wiQqVB4ZkAKJ4/mOStc94TkXKtlG6BezqUyZZ6esfl+D6Gu
jTCCgVp0VjDHSimimU3kpkyRHwzPDO3SMgPoBYdlfQYtsNCS7PyHZE2znNX7cXZOTuhPy+P99pNv
EXesqR2g49Mstw5yfQ7EjcyJ+wYerIHMvZa4vzZ09nUkC06h7L8GadCXeYIcU5T1V/stlop85pPe
7LlqKE1yU+P3/0i38jhuYmTUH6VXHnLwBbvvcYey+Iqg4QKhvhaSx2jIwIiLaNJx0TRsYOQjH5p9
iLJS12GUvqcsePp74LBmXzorIX+TFcerkYwBpTmf0n9abvn+rjcZvRM9sS4ogF6hd9fuRCjKTyhk
qSqfU9hOTl06RXb+mrwROzlnlsnswQxpqUlHVyQyUWMCbJeYzq7dRLow8YocWziCwrjI16bSPxiH
NZSbiyAL7qqHrTRpERXK6XJgho4OppSTLBWMVRty2GyUKpOC0EviynEDCrpa2+0T9BvQsRt+adCy
lNPY6A6/ghtSPRO2CmRUXz13ihV/wzHVdIcc1NJsY+kpjdRTlNtTtQut8ueh3oDyTUwcQNB8gA/6
d1iGWL+vyhPYj/yhcN1GXkJ192aoRWCNAnyH8map+Qd/ejxTKnot643Rm8ZOkJtIJYh+YK9Iqc/7
HbuCWrTuFOp3czurOx4D+ws2raqpRek6q7XO+d8eGDki62OVtvDDNlbo4er4y3vt8Wnvt1KQa/Fj
6POli1a3Iz49ngQ2kchcVFaHLLFCkw5sDMoS7uKqx2IC1kskngULG+dWomXy17n+WgWUqNDFccpS
NcFpYeJif01cIPcSX9Z2yQDzSjJ5Wn9VtD8eSBnq5FeDvYMHuUkvwy3V4t9bU2JvDg2/JsMQFi6E
g47Eex4YH2ejkaU99TShl0DtCDvGDq3pG5ITwXKuvGpAN1DZIps3DzXOdYS4H1KrowaqvYUmfb4q
4D/MCkAnsjoP/MegWSWDyVo9AManvpCiX+lU8+fZEWuYWA1Ebx39ykIEoUpsDBOmwHufshvPm4fs
oiWyuP4chi99eVOJ3BEZaJRDfXSwzHbscDsfMer8yGfE/g/qrpdO0JOKPz2td+Ka3ZYtbaE5kcQG
2dYC4WusqkoLLxgz/ID9z8h50XH7PhWCXZvPaYMK6G1HC/XflJW+e3e5fFtWDQkq3UJMfYgowEiv
l257H5JY/FGwkdqWL/90WNV5dP2aBLVmSx2xj4WA7uHTZJ5GlrVmOMwhgJpxIcXDNnLG41SS448O
9bTZgcHNera2MN0F6e33h7VLY7KSMvEPKIU1T3iVBpJPEqQrz7ce38NxwhAGijlmM3HtdCOJwvx2
zw38JG4OLa/iNgnNKTqEQmD6ID+kKz1K3O3SoIKFNCGO8/7yfo8fsufVJHzZLnu96Gjru5VL7I2s
24W0FuNT0kRoJhrqKpV275/YsCFtsADMx4uPebBia/ov0YneyaecMR8kGzwU9b/rsLt1M1TNGePF
1rRRILOf02LWBAG6ls18OEO8Wpl34Sz9Ywd4YdtsPGajjP1JTxf2YattqFJf2Oc/LNgd36sRaTrx
egKEYFGgt5oLyHDpRNcRfoqB1ATuy/hN/XnLzI1V/KlgWjhAp5NF2myIwB8lOlTErOLzw6jrGiRa
jgxe2UhZqo7MpzCP8zv+zcde2Eo3eMvFdXtzEOwY/eW84/TprPV8ccoOBAC6T5qcFcuFK/oPiaTq
FrAXlNQ5gdKRqd+cUOxQ1CtEuy7TS4DYJp8nivr3v7pWYR/71xrPp4SeDJXLvV60TVR2LxPKu0x/
YINKDv4Bxwk11uGVrPWtpw+fmMcR4R7mLKiq3DZ6EnAzyWykWTdPAUfHdgt10ogmopRbiKBNrATj
Ny8E1Yj7NphZonDCgo6pyoC+dP5DhsO9tbosLKYpJEMgkT/w+bR5L7/9SnBbz8RUW34IGpzP4mxk
obkkj9P5gB05sTIE/8+3V+EzJ+RrMPwD1pXOytOhBU9DRxin/xT7UAkAYSpvDMEf2mv1n07Hk9lP
dBcy48IAMgjdHLK+pSyLhd9iRHSYXlaBu3uEs1cHjFUaGUjRkVfZ8jKiui03MMxngok4Ygf/nWIN
G3C7+xvlWB+WHAm9YIdWf+B6cunu5z0AF2av7csfGyxlUaeh9xdyfllg/0PLmn0esuTRRtC+l2Ia
1gc73T7vY2DEoDP/cwSJPqWx9fLfTidamLypRG/TA2d3rlGPqKc5w5wIqTt+/7z3w9sZY3UwakEE
VZooZgMCLscjPvkI34vor3UtYQfi7OB16dNcIKgjMhCrAD6dW/hYPq6I3EfqAKbXo5UzjFuzw9Cf
DpzDSF4+Mx6lg3FH5oubRnxh8ZAaSOgGqRkqUpjknmiEZw2IO7HOsKbn9uTStXMga+yEcBIYq6AH
dnktT16HduZ08d78ZaxOR5MBzV3OdLKT1+NcGad8Zg7+/Wzi44n0bADQ/ny7DFQ1rUyMUskZ1j6e
tENlxw7P3m2EantHmZu8977dHj5zo9LH84QPYAIhqXDmifbWrRAsiSrdnLry3po3pDghyrc48dAl
GTGbM6K4BcrPXJ/5OMnvyxd8UoTxHeijfxLySJ0+uueiHu4wE7IKxB1kiOSbO2OpILuDC2ViVk7Z
+0qaGALId7MP9apwqZ6UN0NeLCue8dv4F5OvPf4wKwd1zJgQJnILN4SEfqJCQ188ZM8g+nR9hhH1
aLKApUMdwlKFSZBUkdX8/iO9NMbzevYmI/VWA2a7EW1NtsDcUpiBYgxWib4G/1v4xvlShrK7HXiF
BQ4WR0Fp3CloTIM2VtPyZKvRWwFxaElOkyfy2xzikdOZOZqzMDrGFFaLHQ/4AldVKl8P0PNj/tsI
UV+QrWURgelOf4rZRugbHKuD0UyX9KW2S24YidrOAjwTxAjceS6qVxH+vCiprvzEsouzFrUer7GD
lY7l5SnbLTJN3Cgn24vU5HYLrqRR35d7+LbFA8rNZJJFAGi5Oe6jxJaSBIHMclNK/TDd2N2oE24/
KJ+BK2+FwlArS0mPFoPSGpnjnffdT2TZdCQBdlTPxnLj27qO3b9KgmX7h2MzRLNZ7dk/uWVvaC/F
vcwJ/EksiIL4ZDC2W8KOFup8puNMZuyjg3a2qvALpkzlQPXiBO9hJPXGLEsQGj/Y5R7vMN5kl9D1
b9FtobQG4OXGI/rDVKekHBzAexAlSYZTUIhVrudJlZeDF+rTSO2BJk/6Y+tURti5PEaePfzly/8J
1URPW8y36kauaM/x3v/kDdnqNRbbLXdAnVvhDJPGllXQar3SmABeDVHBqvi+umJ+yZugu2NWMdep
PG1dR8aW16SlV/W/E4/Sff0CxPFXJjSP5vt/zls9CBtNrGAxr3LNsdQcnE2HNxMsArSFezbmXc27
L2KCB5yCJTaIz0GKMIWFhPJOTZCjc0eVDwGYCbSvzPP49u6HjXitmHyiiXKrkP9w7L+OarlmZ8UM
4x651O+EMGzp1aj2izlyT58o3fSZSSEuak44jk1lQsAEM8HCgE9l0dEICSmsqTKsYQu2KxautzSK
0AiYTCyctHebw3UiF0IVjQxPypvq9BzsZzZYxWmNdQGml3F8ew/1KrbPE4HTby5DiT0jrx6yz+1t
mjG+U6dVLymuXGm0txZMIN4PXXnHRNelothnmjTACpddQVUvkEUkhT0wYZlDRBVLRCO2uwOIVr0U
GKwSpJiGWucPsAknJDZrvVPJs1AtbW6SbgohJE0Kn1jyK48FluHq0JGu/JbcPfvWI4d17CPQP3Ch
PPfCRca3WlcJLx0hfv9JEjwYHHpo3OItylS8FXElic4AZ25Vi8tsyRa3TUlr1tdm9CJTQTmCYQ5n
eLaaGjCqHTebYBp6+jFqgLrhqucGdBYuIdQFf4nmjSScNCvJLQAT4Q9p5U5JOcP5zFJWIZzGJV6Z
fIoT7CaDHRwXaxZP8YQRLS7s3iV2yj+lwYzKw+s80pjYtCkMI47v6x33bzyHvH8/3QRT2E+Cq5fH
3alqSSKgOfO0e71hsmSZzflWBW6NQQLYAeHTLToLMLt2NcPhg6CgdAowTh7rN/GvzhwRgy3n9g83
bmwvoARKiDpgpFepWl7K7Ln39SkEoSy6+RoCoSTrlACDmhSWq6BznP3zB4fBRsFrckJ7JBtInqAF
KFZd+itx3l40BdIbUV7X5yN2pNIttjc0kk8Vf7PVUzlaQbAHndCkappp7E/IQs1n+trzEuEu8wdD
whmZyqKYq2E52CSwuWhmZ46MpnSMfbTStssBUsEgDv0B1pPsqJSdjUPiVvVMpeYIASpRx+JNGrHB
1vXQzgDYkYtLNubXeFcTz5LJx0z9K2jUEEL2eN9ot5HJUGuX5BYWTCLLSY4x9OT7kjx4Th7MclXb
bsmcGf/NlcSu7l3+HhcTwQ6iaHX60adze1tLJYFdjVArytucNrcitp9NIrQEbC3vC3Qqz2RpaBQI
iCpPzQ4Vv6Xw8qlTNQ3q6fyJXqhc35Fi2ptUc+6r41Nyqt08cGeb9Ah5TF3PKd/eRbTwoV/KUPZn
Gokd9s9LxZ8ipGhCS5uvdMHZLO5Ecm08o0WoKg5Lhcbi4sO5AlPAUffME566GOZzn5PRv+6K03w2
tIOi/D/FsyO6LwhYIIxvWW+L5ypb/OZAb9wVtCUcN2wUr8Wl0O1Od75dezHieKTMvevQjQF+I9PS
fZ7J1xDlyxUrXCmBsGblDoqUI92gs+md+Wj8T+fXIEbqCdJJclq3LI1Yf84XquozKsj2HKMQ3LXx
EpwwwGuYShyNqAoybM449OltqdT64cXQY7HkQqxewu3jnPcDbk/R57xWQfQscUvIpOivqFXlQTYE
917rM3qm5Of2/vnD4aethUg4/ajAfIgId9eOKCgtMAaU8BSygzrofYrFHUPni0VFb1+6mOdY97iP
nweffThGg2kuAiWVppR1jDA4Zoa4SeDx4LfyWJr5QkMVwrVp0MET1ewrWoOFl6iqRq1MPIoLPR+Q
VpNaC/L3aWizkMSrvr4BI+5DXYnmrtfmu/YyXJ4gxA++jKYVDCTQMN0GGSp4roIqEd5nL8cceRVf
IMzk28b8h3DI8XWpFnAox1URgu9hKH2h9KaXFWBmodg712QwczLeQjrKk9zSNg7kbaMDpVHRTMK0
Uz3wVvSIDoeFWLtsd0f2/k7BqbBGTnlJdSPQ59HLRuvn8UETYcoq+2ZNqj6dWWEQ2KSzjijy31ka
U5DkWq1E7SAv5kDDC24nv0YwCePfMId9gn9RNWsZjRu9sZRxfusPlcKbjo2x/KbzokUwUP/iq2dF
+PGL510HBVKJur3IZqOy88x086hr6HAOLt1zSpgIXcKfVZaBpw39JyrUNo4QdeQ/13CyA5lc1BKK
rUUt6YPgK+cMk1znsAc1TKfush+9NbjY1USmXVAyHm64pUrPbX+DzH+cfmvLckrbgK8wxE69BzoR
ycnV0yR52ytq/8NDTQKSofE6Zv/Uh7Qv+AhNdLXuhOg/c0FatrvWJcqeZwyo5Z4OxvSJ/b7Eckx3
O4F6YQbYK8lHgtvL+FpzKtwM+ycDrheLvqFaZvdHIdlYjlAK19sZRJNotBr/H3TD4YL60c8ZgApZ
0PKRjS0Gh5Gg7G/5uaPKuN+l9rQK45GAclCbEsBVqfFHS8HBdyI0H8cmCq7d09UcXPSdkXL5TFZX
3BuXCu+7O2vORtHt/WChSapqGidSkfIVKoO125bq2nvGJ8mBxfgZJOoOiv3Tq1RT9KhtIkpAdJHr
MeTcVFjyFmETeM7b64LvbeuANaIhgYyTzr3QNM71ohgEXoAESji4ttRETR8y3zv7heJO0sNseL7W
HgNRvk/3a3S+b7dZb2QnrMqf2Cp+E2TvqowRHEQ9y512OVgsutfNKAD4oXcJdHLKn6qQZMnw/nuS
1cScc+89ujUg8Mqbng0GTwS7yLeBkzs2nQKU1/8i2gw4N9AATjFJGBLKtwkRb7QUyIrGECrjuEyf
1zDszy7goCe5DCcCK34M15qYY/Q+CEXwRrTDaP8WeGOxCLJdTTO+OQ5iGJL8AeC6O3M3qQGWZLjT
9xdVxKQKXVw2C7AddwvzUh4HYK82Xk5iRCqOvoIdWucqyjycgUFyaveenhReqGGolsj8tEYych2N
VfFp56Lk2fA8ElqiS9ey7F/kEoOZPC4u26D+EN/1kjzYTtcQQlkLlD9fu4gTYO8bF6yUykje1Ref
hFAx1Evs5MVQf+wZ8X3Jic1cNJ5VMFW6oeqyANvRQDYoCOR2V44fd1bNk2r3S3FLCf2lA8epT3lE
bM4Y7o/hXtnKrIVgGPPbbV7ktlXbITdqU2vV0XtcTF7/ELJIgHEXR1/M63IrBfvFwI1QmO9wX1nX
SubOYprENIAALV5PMFbLEIe3uzPeSbYAIS9hpoIJjm10H6oCvvRxm2QdywvbO/fPv8SFS0AzfpmE
9JDthNlGRcX5D/vW0huB1XfBKoybjDzXac9XLNyCfTdgzRRA6JqFbgqFxxVkedMcEFukHHZ+G2VL
giilf2wzanMK7uzyKWIqfkr5NSywRwFkmWRvbm2dvdN6Ffc6fo3VH+dFqbAFEUJxaFD/WgGJvy7o
kJdNq5DxM9JCsm6LCRUyMNHq0cMmbP09wrXY1AqQacUcMO6Tc1XO8i8ihke+VhsVaUfZ3rgZ2G4F
IMgLzsMfq2OgeAtZ3pcE3UFQgWkgHJPNgJRIg/4u5RH9iVe5dGsAE1s+DocxeHb1UciDjmNj1hr5
tOVbJ3Q3xn/Aeu3TkbUhNTxDDa5Co8pi2ZtEsSC2eVGBRJ5Ek12yOCeOLDAL99DJOFFxQl8U+rPu
FwA5zIMoj+Xm4NmUxUJZivq9UT8Y04fmyfV1FMEKL3tkShY9X0nRXPkgPei/krEKNsVfXSZvRJA0
6wXzHHc4ZXzpOObzpJrm4pXFn11QsFKD2jcfJYMz7XdZMZ2Ct41AYfzp4S2k6acCoTHpi2QMMbqV
ZprYI1r4gH8NujEItKkiZO0GU4UoOlhwp/VxyIgXrCUn+eDF4z1PtkaZfqCKZwDjaBqOKRhff4yA
QTktjgnJI/Sl+ZTuCuoihP7zP4uwxoYQ/oefAFXdzptfwigfoBERdRPBJ4sDryNM3Jg7og5IIxey
7kFtIFpnU3qsv5GVXsYEyiZ2YFHAHBehEEjhBt7GLqY3gNdrC0R8DzHh0lqdv5I9KndVFyzoB9El
quFoT92NtQtzly8cAJZrfVEKscXgw/7MJKdby/ymZ2GpLJ8tmGKaJmxQpHUT31be2BeMfmgMgPau
6eH69VMGQJdm2gVn1sYX3VS/Bx2W1sWdJPVMOXrenf/o9vO2Ch1LMAs1iGO405zGzFQIvhBLzv7m
pKsgyU4QbTfcf6fOWKNN3Y71mScP23WzvPXplJDLch3jbhvxiMoKoGXMsGPblu0tgrbDS7Y1FBUS
nJQvNZAMWwFgl/PDYe4EYwOKsxjGr1bgRvp8rEtyjQIMcejxrOGt4+fVOtjTus+Y4u6gQtIAanLN
zHG/hSMHfkRxhIrR2JuYHiCwc5cx3VStvIrARFLQnitCoFaab4QbM3OGoxqI60CfFggzNjo3VVWU
JZ6xwGtThU788FluT2+QJNwj4jVB8JoMEaxsv600MmIuav6bfHaSZRTWrD63xdm2BI2uwycZfAYh
2+4WGLtElU7ydj2bDg1VyZJ2AhgU295HkNclEC95jWA3RnqFJEaAJ4de/gYiKUWxEelZSKHbenBG
Hi6ChE2zL9GEAJNJYYZN9Oh6reXugb4mCCVMccS+XT+BPuruNL2R0jocQFuYjbFW2c01efDEfnYE
9hGMU57y7C/2EZ8MlwqvGZQpVRRG+M5LaO1PggKXiH12kaqYXsYbUdUGj9Vb3Pr/bAd4wYoUtZ8k
/trjVWo/SxjJudHtSlMdSm9aROZf8Wyi/sXRHnyUEJighEmtzzqboz3FnRFty1F8j02gIO/1L6Iy
fYcGoYEeSD2YZtyJuRRzmvWwq5ly3veWcFWQLu+ZHBINjw/A7XHeGi1PS13Dgi7LEVJ2JmYs/YEk
XVsD6ImDFmWM1sZm38e2GyFMhzbpUlNRSiv7eyJuUX/kJDzzIoZiIbnGyHnUk4fNVKi5+SP3Qrjf
SBqg91YTY5tKyrMDBCIj5BCM3tCCU5N98FKEwa5M0AzsuwQyxMcoGyL844KEjSiY+F5rVdfs/ocL
bWtXzdjYoEyTo2nsnAfQL0svva6KvWYvV7nuj5IqDAlCwjqFv6CTkOLpLvXh0q6PMtS8qaHssnB4
AIkL2XH/Mxn9O8op1l7XoIP6B0fx6umRjNKZSRXI9a6chyEctDgHzwXTmtggiIz0Uo4vGzCddVQt
6lqr3ISRhetZ2oWUWYxzKmEBohdz6SNEZ4E+/mCX/q64xsGLsaBcLpsFhzaWkAPNR9nzIhxh6pS5
QL4/IscQdaA/orCIO3FUScxPL5WCIDBR/b3z0MGPP/UbETWZDDlbZ2XfpWpFsRS/zn3mMqDlrTcl
dSseKTGsZBZ0ZghgT/QJXGdJAkCQEIDJwGb0J+Bx+thcV3KCyc9JYZRmS/gvhlbHh6S+CihFlBXN
Dun6djI8K8PYPwIqJSi/6cozcIWkckqDwbOuwue8XLypRuYcwAAX1KiTqOgZyd0u19JkFoQd1fm2
0Lg042Ny5M0wQ+jpO/PA6oq1kCFYcgqOLGdIHeqLIHlNcDwIE6UEhMpJzd+3yyy5IyCMZIRhEZJH
ak1l9BtZ3ssUmpS663nkX5b1Q7Lg8yc22lpXmCsn6JQsKBC88JQDLCVW7mLVz/Qy/EYu+ysZCaMQ
9qBFbQiNvNtKDGyqnzC3ZQsN6QAaJNRZok5J6TBWhbCrmCVh++tP5u5XidT5zevJV4YbfXRAzQv+
82v8LxVOoRd9CVVyvCNoGTx5oEcGBvQ1s82sPlUHzgrlwpykGVm3mb8jhhflUuYNIGw16jWC2KcA
32f8xPDHDZ7peL0iDyqxU34F8J7cyrEJcAL0MTXEGz4sPLkjLl62IWBwzYEcJ4xJdbsjOpswV9XD
bgRRGaLQcaLjSwSq5+7zrsa77hDCrc87c7Mv+U45AasZ/TM2R5d+qNsW+dzcBJvCjhFACDMtS97D
nf+UiNwcii5y+JYn174eIJoU51v5q5e6QvmPVzZQLXanIRSr7geiQY+4wKtQa1S/8g61JQ/bfnSO
Pv1wBFNcmvZ6gKMEC7fUslos16rFqKsdaOhjMc3M84XGmZg0FonG+qcPp0bfmgqORT4FYavf+FpT
d/03EjiEUsVfXN0RkfTVBMciujWC40Xef/Fb86t68ATTP5pK5JEmureLr5UV82eKiaLBHTskf6GF
kFFML04K0Z7gz2Ck9OzMm79DWUhbCBuX5NkEDYzhD5nhPkcNhPU9zIB+il7sG43/wynI8rTGwKq+
z/d4zp6+YPAP1AURwVCQmuE+o5cvNr7Z4O6TYLnAcUuqOPkrwt5nU3T4agthmWbwp+gjMEDToAUB
f8zhxufq/0a+h2uVfkE2Aw8qS6yDdKkb9YFsb4nOFVAAYcGTzf7mr1qrj7P2R2woXWwTh4O1TIpF
KXOKrceBNaRjQIOgqwsVeetZStsI9T1wIMzyFoy/g/vLef2viTthYAkkUQ+87Gfv19RWs74bqsRB
31bs29jkz6yNWofjhlVvrHCOMZLEP7bwe06Q4ylyf1NSDtOsLEU3ZI5NdlM9XEumL2monFnSKHEP
gBcwKSSruckEJEHq9kasM/etkBfCAwxD1lWTMZXIUmmoyxu8/RhiyJg8JzeRL+/5ET/bfdWvbn3/
ze4XKMaZtu87DmauhUd3cCUWwStLzGt2G4frtlJa6i9/t47TeFYlMAmmCVG1OtQA397BETb864K+
Mz5JzCvqDR+fnH7+R6hssZULDudgiaPG7tufDG3zLgEYar+Rp9WnFyFOKNgGY54qhib8v9weAwJd
oM6DdbUWKhl8mGNIKjpjZ1COxen5uiItbxU2SUWFeEJ5mrdSVqLtFxPoiEZoq2yBcwYLhvuuVa/L
gS5tGZKL5JrvkJHgKq+5O+RXEkJcSOcybwqXUSG2oFlTS3F9Sgltp/rAPtgsRHOIZ9wu2r+AJ8rL
+FxmEAdfL9CXhgVJ7utGBd/XTiOl8kdEAAiuNr6HiZzLtPInNw7g8W8SgjRBDgrmqYOSbtZITn35
wXmPpqtUEnBlTefsaBKcJZunUm8+QNNA3kkr8ODC+WdbV875tSwlCCWZokhwpt+OQQ92xJQdc1Dm
WV3lPvOH40G53M4QuYE+hUDcBktnzCCRtm6bUiDT3awtsjxSCxfX44bbFgCCq52wUN04cRwFykVM
kH1ffNS7sy1JgjEhpnmfYKh8whGxhG1ZdwXTLf7Lcry1ocltD1j+EUOpUECLJ7uHx9PRXNNcH+YZ
rZrU+truJfXvxqWxoFD1HsdWNYU4na4HEcAmuC2/ZzZAW/ZRADS6wex5bXqnqpG3ktNeAXzQUhz6
KxgabzDSmU740Vf8KlH5WayGmWLuLY3LJ5ILqk9JrWUUG2TLhmK9SR47SzzzME58pvcnerNB8jJ+
z4MH325cj3HA0B90c41BQXkNR7EHrEm9Txks+HcRFPkFZUJK/h/qBPgbsMjkxEa8LI6XTfLva+9L
YXLsq/I9ef2Z1jShGRBCu/nEf/EspWWeDAVuEJ2yQQJW5abjoqPqcNVyQ9JQCdsW8nxnZoG8OdHG
HJpgoIODzF9E4AdcAncfaw0Kcn8qNgV0p0up+OvcobX2JPE6wpbbpspGit847sO+GFEQUKILK3gW
9Lyo77zBGdFjIfygyOvGhMGzjxXpWffinMyW5dEWD3o8hnlJXPuDwh3/ehAd8tOris52hNO0FdLN
oZoUjFSMqfvZDYrVCu3C96A/l4vrgD2l8e6nFZT2Oe5b7Mh0AVA4IHfpsLTja8CNN0NmS2Yr6zXZ
xWVQMAv1wZiabfAAMFZV6MYTKHuf3pZxTHubxx/xpICC/DsI4y9jnO96JhZ5U0tyX9vH0SVrCLFT
MJClXrIoJ719x9QqGBvb3+3r64jl9pOP/O/mL4ebWzhVegRK7s5R8uQFlh40ddfUt4vBOXrj5Qs+
LdeB4Ann42lubZF4J3UYnXFKVTTDe06V9SlVHxK2fnQR/qoj9K41MwTCvtnwwFVrU+r319DH9tqr
IvgWHVoxxLCAyNCjueZElDL62qIkylyve1lGM3dfXr3AZv1ts2SAeMDiwEyCPKjXJ2exl/y7qYf3
EO4M2iwmPmJp2ypBeU2Cr6c0xsRY3Z92GE7/nRN8OC/SlcNbGji1o0m6RntwPaMd2JdKFW3fgwHc
QuG9JwtnpycOx9mVtijxKVPXHDX62kPb0wtEMuuwt8oUIjpTy9WNJMT0s1zgjWSq/yfX9gFQr5dK
o0JcIUNA6KuWDFZKnZUUQVzbt1ULjs8m/LgTvcZJH7Clf2fPi0HXSxyUr8hYY0ZMUKim379lAjat
wJUJa+jKypO1hVi/o1T1z6sYRjUiTZJMK2SLjtRrrHT2uHaEpcKHqgOpJYjRigCVFbdNtHrq8wpU
WgjvmwSFfZTlt+ZSUR84g/aE9qRTmxvUMXFvU0b2nEMvFhAGgI3a5QvcwhFQTwUHGT/yIRPKNjzI
TidXysR9fdJspoVTr2rmUkEVsMDu4UVXBwp7e1W5MpFhyjGp2FVFBooaMePp4g3CDCukwxH3hhMM
+bGU7kuLMBEXKV5SNTw70rl8CGE+gzH8h3tYfuyyddUR36e7YV05H3XqiOrWjTfJbUc7LEZSlYqd
OPSufIee1Il3HZCkTYSdOY/kjqx8x5eUa1FeylETv7xK2PV8toHXnmS8AVKgclWaUR4F7kJloHUJ
h9hgFQ7b2SPNuFurMI69zmjq3BHCIVR8stIRInkt1X0NQHxKGvT8N+Njz6z5QDhMyX/1tXqPzu02
NN1a5NRDRaroKUwOE+9lnufvFK4mT2l1eTLFOLIIlsIKC2SSuTiv18A+HSa/ULPGz0VnUD/DwbUu
2VJrM27hj47qWDVv1Dp7GmK+tL00O1hwo+pnzXxOPlyOs2rD9RYqrj8VWsKnInoa5FohsiYkHsjF
ElRNUzhKFng7USy7/UAoKhM8fHSI14DhbM0YxIY3mLUreI6jn21AqCQNr6KnA5Ghk8bJ81R9DbmO
V+sji6qP4nwGuCmV9CG/VtrZAZTv8V7YWLxikuFjGesIK02DQSGZRr3QdCFEho5mhvpDO0bl8AvL
4+ESi55aiJ1ilGdBrNP/LUtvb3ksbkNSueF52HoHTZtlsnNFevGZR6iTvVLSyZwLc7crRUJI3mBT
1XBqIFBmVRM8/bQ6MzBVyFFFEgeaaKuRXX5TC8SepvbGYdg/xDDvoHU2qPX6gLymYaeYv4aNRo6K
toGgr/9d2kippioS4OyO78lWj2DKALPZJro9T586ipgbGRMpda0vjITAkwmVoIN+vYfv8WvcbK+U
DSxNo/8nNYYuK+TSAwkycdL9Mrw7nTvOE5TKyP9KLHYj3UJH+Kd+J2HE9L8O7JAjsWEkq+mhymRH
yWtFz3KMs2OKuEg5WroS+hcPLLIBIykaauyBE8P0aLSAxbp3IXXtGYM6eNpYY2Hk2odjXjFxrjFY
m8Fsa8BLLnr1FpN2rCHe+3Yh/7U9oea7uk315rQNLH8hZYUhZopzD7QVQ/AtV83+tmMlDz/R/Zed
yDxIYtmfrALFSxVjGtGO9sEfuW+JMVDfT08rWlX9EaRGlTRCra73W4avfrMZbyMNyFdkrGXsdOA4
hBEyn2qgM1axBXHnb+a6GcoVg31CEBGJh6wAlbhGqNY7ASLpZT2hKncqTJ3JGC7lDH4zx+AYUQlm
TiA3wnm9P17xSGj4M75ij5OttxX5VFqvoENtWHxxg8hIrsI36fF++Y+P/XmIdKgfaJpd2GfPmAEn
JwB1/z09Hme/WQVNbixKc5dJCk5kM/0w24wH712HfRUeyZgj9hAskYU9d9dzFDTwKs9Gt9MIIKjU
/DEeOKLKgOFUyl/appqA2bs1RjYPF4wjRb8Gkw3EKbLlXZIkL8I7ehSwLqNGGE0RUB/dK9jj1v5D
mQNQvcOaAhgCKY+iHaBou4n5m/9DZqkk0O86Xe2JPw2Oxz0nRozPjSDKbf644PykfL7PIwBH7l/a
Q5OL3Vfb/QYNnUUUSmU5KZpWNpyEt1rTnQCIsZ8n4vzWZLauDO6+JqMZJVNucBEfClPJnS7q0Hnh
WZs6pMuOdTUUP+xhVu0udcbXgvZOQ3n5Q0JbkZzHuwWZ87Q0toxpRV8gWRcMOsQ3qMo6R9iQqVXE
gWwGiNcqUAIkJ5eJNS5Mykd9+s4Br2hQdNM+m916DOX0vyw+t6bvytG6JIQXFQfxwqM8YuDeghJJ
DBsreDhAl3vOOtlUXGzHUgh5Ymc3rjdYhsilHtvwaeCJlZymxDwKqa70D3WFI/lyBWEEgHQ7jI+9
wd/0mxrFGwUx4TCWM2HE+29S8Ral/BuKy/4UkavqaQIuRQW5GsIOMUGxq5NzisRcN30VUHLpO8TY
HVEcvsW/OU/PSNrbPeyJwnqPUzLHMIKeTMLHltnAglMR3s7I4+UpbBAdYv2HFQqB4VGvlFjAMCKt
ezU1hCQrXqgiSeN0lS7mLtIsyFglDMx9ptEznzEwAUFUJVWn/xiEZ4axzO5rXdPExCcF21isuUnf
4im2I2qVndAOU4uCbbgjsQsDw8XSZ+K8D9lt6YY7XvHtb25Kp/VdaBqehSJ7oiYF5/ZFzGfpfM1V
lvJL+ErwB2YmpNI6Jc7hwqxKQh+JJxKl6gYk026EjGSbYT9n6jk26hhBhN2s+cVAjiAofiSakNsr
lNoFWuRidjz4daSHImqLz8rbJf/VNlrCOfVBF6iFgN5ajXULd5SnxPTK2yW8NUC0WHzVuAs0n8r+
TLvDbgi6ACW39GxoG7ZWcgVm5XWyLZghL9GGOPhEhN99GuxVPdeNaLIKwNHGt7+bFqbyNbuztwEX
Gwnq+2S/pHXsIWnv99b5odc3rF3ZUowBRwHXn70beynrOZj/OUmA+bR1pUZS+WgXqh2wK4mdBe9t
g0adyvQ0tJLZxclGXKdWd0ZWWSZbsERzV2EzBZWWL6xQLPolX4XG4vXMzIONWmGj/s+AAHAYX6uZ
Z7fcZQiPjqryzfS3s99tDa4pxo6d5/HtDIfWVMr0ntoFBNxRd9op4j6w9utI1f1fM9EZV/20jKUX
S3ktrSMEAcIh0iKcS7W3SqQqkcQNUcrd9KF048ROFQ+JIwp7wpgiFN8ojT3X+oPHjfILIVJLNF1p
PzCTo79+LujkneKZgCIxyvGrXKMtRyQ1aHQMNy3Bj4Puc3UKFwvSKt2lJXbRpd2l/cB5sZvn6/di
CXSJ+mT/HZi7aFgkuDMG96U7o02xyPf1mWKVP9/d6rQ4EMTX4FVIrTRTZMDU251Xy0LYZmz+OG7q
BwMpEpGKZL+kO01UA8JJzpvbA27+T3NtZzc6KacDbJw0yboocfh3R8utl+30QOH/h2r7/qglsk3U
uC9MLDivNXrcKXWIQFhASI9Gsg1mTaDssFkQXntyXTm080bHkkEj4nfUFwQmaCI4BSOks3zzH0ff
GrKzkMvP0yq64YdmYs2rfcWF3wdunFEtSNcT/MXbEshuaepbyecREU0SvZmZA5pc/f0gAIRWMv+B
qO8WABKJxwvgvx0+Aql1ZPYCIcO3B2npF1qagZyN8L+GoBzv9q08wj1SmL4l4//u6mLTKsIXXjAV
o2i5JabMT7WJ3NdOZhQgTdi6UaNnd42pLPli9DNKSrZf1S9GcvmSVylEA0xQV/ybICVXp5DSYvKA
mI/jVMlGne5ngnHKxaHj6D9QjlQZ26+VrP7sy55Hv2DSWK9fp4e0I11+PEyDF5yFaHbximKt7fGT
IYL6684Z7yOTZG7JV0UK5qI/PDndIcUWJXwEYbyULnywzl/awgsdPIrr3vJE3k+vzoDEuq/ZhoYu
7UTrnP1LRv4YWNg46aSnq9GkiT7phlvRNSx74VA8e+ENkAq2Op8pG+bsJoU7AkcAJ2VA2t+DAZAP
Vm3uG23v54r2ByqemA7qyHYVMEfsdtr33BxhYfoEmT649VZ3Y3eH8lil6FbjEv9dc+z6gObZxKqj
o4JOtL8K84ATIX2NlK+7EHCf6er8N7E446myiAZn/jYt+tKmhlvngc7v2xFBxSE4LnOlmao56W0V
mbK14gzWDKLs7+dPgY7/Lvqg1RuWNsBXCy5sSqYHeYVb5KpYY6inuN7Zdwspx2ryPF/0zIcML8aL
IUyQkjtPso8AbnUTHydVKkg+WSm/qDQji2AiFKdlH1IxBPZpmLjMhySJ/GvW03Ofznbs5aZDSu5b
JOW6kY65+riDw+gxBzB7P2OTecO2oonYrZh8hb4qok9yx5c8G/ubg7J36UPrZKGFFJM0vJ3q/iGy
F4k8r62xQeBOYBa/l0GnfJofTIidK1FNkkwBmfT2YOXaRMwLWgqfYo3Zxy1yto/Xke1+izYf/A1i
9LEExjN1zYGQStDiv/AL8Qzt5VmAlqtkAaixApgOKPX69Ox4FbldBeC2z7Zk5ayTUl+JfkfYAVs8
GLIY+GpxIvgpBvRhA6z3n7SmchwUAivSudDGR9EKurZ8+owvFn9UzU8dSTZf+wd8/I8QhrJn7TNK
YaLuwvxuh7kXI4C77O/d5aAbT7kzWyZAn5pZDkFDF+d46ccYS8xxduGRDs3InCNObf0kk2F1kRl6
HPIaB4TxHQllbeIhXSc/iG0S8Hv9MksmFMhxdwVw0q0WFoCZOmZbRY5XAT0u/hByndsEsK9I/+xF
g/iU/tWklCJWPaV4rkFA3LILMyGOTIbWjuI6ZgxyYMSlOO9atXdDsCuefr/ROJA1I4rTiuJ1SAoc
l/lDzltGw9YQiSFWqx95gowzVemQfpjNOoh/7Xy2To42vwYfkN0ehhwGjqLBnJ4piAYGZtjNm+wI
6SAUXaU8Vloq/dDn5lbp3bzwnocWtVU0aBAxl3TW4IaW6yCEyaDQr40DSdF8fnrlpVIr5RhYdRcV
xpekra7ivyoooD6eyr9EOibuFhAgFlQqGudD4k9AWSPKOQRl/v3WzavwmuF2UW5f0c+3h+08HcTj
Lpvvv82zlVasw7mh4UZJt845ltqTohsBMmdwYEjL7Iu+LniZzTChH31GiUyCfcromDuQNdG5qjF4
l0qjdgFSQi+yOgDspfUGMOsIjXLEIB/5djB2wO1Z8e7yS4X4g49+G9UCTAFERTe2e9jQSM9COxG8
o19N37opq3edYacqNS7/Elid6eMepdCwQKIWR8m4+wfswobolSNVehadygHuwaJL6EDOV6K/lLjh
ALlEWzfrwrWByjdW9kkAh5wZlFTQoskrXTJuwPkfIYXB5COx6B9Oa0v70+IwBopZf0FMMab0sZ/F
6NLVjixFuCWFRV1bdxS3WMBTb40UyB7OscVhumjQBzNZQdBVqoaPTpXR+/oanr6vDmDPdFVigE/D
Ia18gmshgGcF9khYH/1xMpcvffl+OAIHF5Ec9IchjmeAPa2kFQDgLm1aUqiA/VszxwRSzzTfRqXf
MOyyqDZj3ulTEL61b0Hy7r3GqfaMF/Y3bFpvjOVMG7dKVA2vIeWfR+Eoh+fFmCBZTM/LpkZWYAs6
66hgpN6/qbKcBjjicpTwiVzCPeWyMMt5o7ak5z8w1F4FNKQTZDefUP9osNRzkqtxu0VYHrimQtDc
lrT0jcDq9OVBili8C5+Mob38K6RIRkZPF23CSK/NuQ76LfI6L7+om+SjlBS9nr2QJvwlu2rUPrvR
2SS+vPHGE4bbKtVzMu1B8lF2EcYEbBU4s4d9M6s+fN1qoWnFtavKPmLExLkI9dvRy6+R3cQ74h9N
QhteiOduMT63/u8jr6hFa5tyx9fV44uLaZrNiUeKtJLkm3U+gKlsXGfzfLMwH4LrB4GIcm57JZdR
dS9gonmznWvG08XF4uBXpfikohCPzwKvrcdG3IvwJ49c9IP9/v0hzMYEvkvYw9GGuMy9Izn/lZ2o
Y9c+4+Rue9L/Rf0VHP7yKH/HUXmTL8nxwcZ2uDUAdXZGCVNmaO/VTZ2nqVbGfs+hDn5tHqcueVDT
RSIwRWh8ARnQowRCM/EPrq23UvLkXyEvLrRBDNtUhRurTyjREKJHolHbAWq68Wk42UH2pDlH6ZgG
Ni9SyqpsSemUXSfemXRklhqaxuUiyhOQ0dpBwswx+Mit4maDV5oBYWLDLBXgij1VDUaWTOcDfO0J
tKVrncf/PXreBDvqUXm1TB/Lx0/qnCxy+NaKLAW3IQO8q37ydJEY0yMdzEi6Jk26SGhJbf2EI1UU
D15JQEApUU4sh5wbGfsk3k40unKk+z9SRG85+R819heJAU7PNQj3kvNfUvyT/+2cXAWugqgXO+ur
d3gzZN1IK5XwfM/suygh3rT1jxFcPVl4x2VNQ2FvoycewqBU4pyvvL6EmzTy5kuRiOJCm5fqG7kv
TTUqztz0PSQIizjqOnUdi0oxSJWXbQmGQsLUDPKxQ2ZNckTb33aBXv3zL3iroxxYy3eb5TtB7jhi
EWvjKg4s/0uB3++Isq9Id7s4/DnYEu+XKyh4tf+Sxn0iDm8AMWVuqSgZEleojDaNcz4SPHb8/+w0
ZtNMOn4VK5vWM+j8KznHQm/fEJgrFWtv83URwSE8zI2pzpvU2Kf4wswmuQToImGFUsn6QToz9AJe
ebaaaW7DMAtGgTS9Xaoed8mHoTwi8JmG9xu/xeKOKmOv383c3fNhiJcPkhiD5YVdITDfNgXQFHrw
rPiyoFUu40e41SBYD/RImT0hoCR8y0i+a6n8ehYvKwkE9EYqB/oh5Q/jrdhKUJ3Db07em61/RsFW
k5mpcfTvLiMI9k/QqakXABCXgAw80lgu8G0VDQaNwG8IcQEVypz+jEefN3fxZ4NtDCLI+tLlxPIA
FBt7yDaB2/XELW8H+vt4zr0RKFYvv4H+YLeTolFgXfS0unclJLp5RUehSO3oTsVK56ak5c4Z1r5Q
6LH1p+ZwannJ/5NxDGRCziwuWmba0qyMvSgrKzcOjyFr2XdVqEdE3lGTTpB+CFQeTMWBEMZUTiDB
lJGOAR4636t8i1bMho+GOwsOU4sQ78XC3G/lDSGtkd2DdKofgjHWmG3LE9MTxtjCvxymIdsoLZSW
N5o9htCwKWhNBdFbNQlG8NcHKV8qaAHfu3tqD+nP1P8JSM653HXmVha7L4ybW283pvRs0uBS+rGu
Zc5fSAAWOc7qJ+tpWLRFHdK6GjMg7dzL9wiCDL9N/1TIdvOHBuIT2C9/zDMzckORngbW32BDBC7L
8gdbbT8tD+zgM80hrmkf6vFgtOE3d84NZygKAoGLvCce/2d+OjHj30o2BxWXDKf6ZkMXy2f1Nm5a
LmG2wX1SROZN13iyl4H7yTSDyP06V3etWLd8UspTJuhSqBECPYUVYJgmJPeTjoNEH2ToCJ/dpt12
pla9qCvMxXwmj299kiUzAKFhxtiyw8O1HG2MYdXRUOit+io18SfUjjc89Aac/KI8uZUlXXlDS0kU
OQ99yrPofJrOd+sC1/kNIMwsyiS5j3I3+rWwAIxi12XMeimAo5oIZUXe9p1DkMA/VX8PZQxid4EW
VSJMbj3GUqCbqMhD0BIcqlKfaFLm9/w5SNg1wXsnOnE1O9X9w05Ox20iyMJi4MSo12gv+gfdH7rP
MiwSWSo4a2jeeorjm1Kvx4EXUcHzb5qvTKm/lA8VNkIzMPIBTBp1wrGAQz3/rrmTw+W53xhuTo+N
LiS8Oq/+P1Zgjfy4bU5DNsUN1YXlP7is9rF7pMXOuhpeMdQpsRZYh+DQBA2t2qDX9XS0dhlAhExJ
xlF2OLWrYe+t84hvanjBl2U0Y362RAVzIpXx1D+eSwGbcMmsQBeB2mOHjn4mRL+xQ3z3DB1CIVWT
/63fcbN34bdc15J7mhc3inUAN8YtT/E7tEYEy81UHbADXRv/ikfyz5NSv+mYe4LFR0aY27FhgClC
AQbo378Le8WU9ZyU73bRp2qKli+Sq51XcdDtxUp3n4B4k8qMqSBafPxk3GGIjMyFQl+H91E/O6mf
vr9ap3Vsqt/2WRX51I74uex9qyyhGwa7A5xuB1Hju7qrsTPCAehc75ywRmcpFrXSFRbJJKQvfQOf
vA932G3Ovy6/mPujV1ZUx+hrYRrW3RfgasI5jTM05pOSRL28BZJ094FBsgdqSYBzljj2CLB8H3fV
Pr3u9YAphJ3hCpEh9Br/MBWIkp0TXDARg1DCv0OTp68Nc5P9HLAeW8O96mBdN8UNV3VZT0u5mzIa
fC4z3VeC80LWHsz/adzFEBKsFLDB8p7DJFvckXYXwx90Vkb8ONrb5xnXEcKi+2LyG40OaQDAeu05
oJqfJU6dgJ9k929YElHef9t9nSn3yWZ6IbogM1BCjh0GVVi2vdKrXyGp85EpPZgRJe/bIMgGpmhk
x1Ma9Qx971nFwd5jhUCgP930PyzNW0HysgPtEWPRVf854cnCb/u5hskiENWHIb+Kfkq4On1IEhri
kYx+77YbVBdiXWEmqSyit2IPGJIOys4EnIciYsBIXLZrlJHpqHyqO5ktjx32bRy6aWEJnOnW8fSD
pMf71wpTsoRrEv6PN0+LosKj/gMHjKtGbn+wdnlGTeL5CRv6dnN3bAbIeEEYA9ilESaORiuR8ckb
Mvv3Y/G5CoMsX3vBEygrrwpC/UccduMqxIpCvvyFxogpDyNCRv1NPPMpdgMvGF/o1geVlk3XBQsN
wapYQGNz9Z14LjdqwXlUfZ3jD50EYQPNXg6i9RmY7OLTqUedTgcKtEzlrDesRl8UpMC2vMwEFEDF
NB/9YSwL+P47WYY+7d7QEtpn4w8EAeF/EdMkuDji3qfZ4U+lhnpVcO3btafIF9XyT2lZfu7Vxvlr
W12/UmNdoGCcoOSDNf4Yeiyq6o5UMEq/pGtF71U/9zeTFZhY04N3o7eE5Dw4aBLyTtRm6o7CtQLe
iLzYGfyT2AKf/YdkRIel5YRzBjKj8QtrKZDCFByS4ygs+Q/Zp6s+cYrclkIQM59MPFs+LJup3y/M
VdVUkXCBflIIuOr3kxraugVMqykShSRPVFx2hGuqqCkHCwofsjGiOvRM+mIj0/w8Eo3tmMBujmhB
S5bxP8X+WIjHi7vX5fixLhkxT6CEcoDWr9aYXRDEVBD2pJJTjRqYhvemj3TVSYkfvUCCMrp7m59m
z5MZmMdVPelDOHIqbmbT7G4eVCIRNTSOq/HLonqr9HhrtrJUoO4jggj9hshC/vIqXsMhEyZM8DKS
sYns1Bw7J2IStTuf59+WW3NKPkzWmdnqHtxklOGp9inEOnyRBU8s/tEpnT5oDRJGslrINHjhoJA+
Jfw1oOGpKp+ZhMBleRcz6OGLmDSBpDFu82ZZRhcz/x77xcjjX7M2x5Tt9aYjQB5WbyetxE4n/P7s
DHf7OtriZpzxsmTDfBHZYk1mlfy89JQQZUWve5+ZezjnzTjaUJvVG9FsDpi8yWw8VISOpgcc6b1H
zaRf1LO4cj3/pD9T3XOfGRrvHFOwGrKT4JjRqC734GnMswmH9jkY3kaHxHhb7rHeuW0ZvKvSyH2a
HydicSWWQFLk2VIPVzLRpErKcv+dHwh9R7IVZ7+flCoAGXEXKHpnvlRHyLw9xpXHsa4vSAUVjcaN
pmDp2sKD5fVoeFd8+7Hr2tzVRYPtzeDHrMe3DrfXFPD1NG4MQeB0DOgVy2NoWnl0XsKNPvRHCkNG
Eb2T5Sbv3POie7/2eRhGPOYfYDMZvX9Cw+OIrqYNG4U4BjF7uR5f0zgY/RD1qpKSIEB4+dWc4tdc
BW9PlypCzFz4P2FQiYIuNDGaL3XZE/rp3ag5e1a7T5wzYmlgH8yrQ2EswRlWGlTU7Fhc0Juyf46Y
H0Hz69dtDTud+N5fViOujDMLyinkyTQTOyTyBryAgWBqnZOfQ8ZQzZ7pMNaLDWiTLpx5nqFBNAyM
dhloUxQPP6TK1BQqqXY0rleNcpTc368XAeDge+ZMcwISlEsHC5jvj96bLm8hcP7rMZGMXh1b8Im6
fWG6D6pj0RqPZsJrC1i3jaSJ5AtY1jKWAyhELyN0gZBUwJZ4TLailJzC4iDu2Wl+ivhEMey+D39W
t00hKdrDGJ57pqrcu4MlMJpaS9z0G9upRuA3e57G1G/Ia5zZRaxZ5xo42ietIB6FoM+/h7Zj21UD
Lg7m5+32jcgc/H+aGFErQCnsYjGT8gIdKvG932sADn7zejSlf7f7cTfdFpLPz5Tj9Z5IPhOpsSAE
ZB5MeuE5ATqdID6bUwcZoD0pVmYfo7JDA/Evpl8HfkOBPLbsR1XmTrBROEutKda42IlN+SOuTNJL
oUT1VIWwcGUN+uuzgVIATBMtAs5V3naynaqfyCt3qyiuMVLjna1lvSWlPcAgiCeJx7Yo91j3PD3D
UWD+tqpuAAmLiw0sg7Xj/mAjgGFCqbf7wFE/PK4ZaP9uqomyIXh4bDXUjkgz5E//K2yLDUzR0Ipe
HEmGCqvFsEofxuIc+umKJQlb53TuWFMjWX4nejmbnNZ5U14J4r0aieINgHlze1hGNV/7+DXEx719
YWix/oeDWYedn2ekMv9nlnA6I9lCG5NXd+K47P4OyAIKFxlFRVxwoii3scpfin5jZ+5iAVEus0J5
nbh6QFpBZiAOMVMBXLsSIyBgSWhcSH/D6RBLcRg3pL5YYAyW35GTcvnT/Xvc0+c6pEIur9fv7H13
ytGqyaDKclN44Nehyj1lR2535ECzf1fO3iidWZ3s3oX00EXeNXaY0WuE3ZOdV+F601xIoiqQTKPA
6zvJL7cwFxLMUY0c/vg4zcVRkMuXm2iYme08W1Kb4fwsZfaEbXg4op4ZrAQZvWtDFVSZe6TZH5Bi
CeBF6KKNnBp1JTGcfji4GqXrvWBAXl2RuQ2FGjjzVUDxItaILdnJc8TtkgslPqPeCBoHPlLjvRQs
UZyuHZWKHg22FBHQbdY5qILcqiQ7t6KNG0+p3ltjFCbLayUJzbnwkB887uo1u9jvX4wex2zvVmMA
MJm9vVNuEf1wzBLhSvM0gu/tJJDifubF4ALEsOMfwnDC8YaCa/fAbAmA8jBj2FQ8mY2cIeUZy0TY
Ne7kDyLPPIHpMpbxXIx9UuR3wrj6s+n8+npPLRBz5uXhDLQvaKcPmyWfafAjXCm3FjY9J2xrvFb1
i1JYuD2nuZCwkSjVRnOebjHg4WfL82jIWQ1HT6T49Vvwt2CBg5n8ujk1weB4AXkho+DcDrFWevJq
mV4IvbbDSLxyqedtCLQ8ubDet1k7lAdCXMz9P671z7/XY96pnU7AMQRtsW77n1Ra6pGu0pmgsCVf
lAiTe8gh8Mteacu1ZyeH9rPtV9TA6AAxEal7x2F7/8lKWliRBYT5Y6X4bNT2+SynEvDqxmsW83mS
nyrS6Di1DaiBqyPdBQbK3KA8kZtLiXy74BgzJdulFNG2UIVmE48UGfkEOkbDACM19txszBSreing
A8n7pRawO8zGTgVy2h9lLErF2VOmykE5BAzXYz2vlAWaF3GeDvHniYSbNHP5SnnjG9ZtSAQItp7/
JqrDlgKY0ATfgbCyh9Mdgezab97nu7bE7bFxDm6VYMD7/pzyOnMIs4VXYmeC9dIW6pdBCb5obdWz
kJ8O6NMTV8uFxix6m2Typ4iY+wV+zhI2u9p+1dHrEnVQeIG3rlXhIvwFnsCvhVWu2KtrODwnQrfB
ObCJIlxlGbnPlgmjBCq/13PuWMVePRmtlAWl58tZlGcT+dkJpayGxnlbtWvtlU5NmJZ1kfsLVoJs
Kg5RnIaw4FgtjGC79D4Qkm5/mo1n7wAGizcJy+x2GIRIXO3HVVjnAE7XvBXF8vzpHAlT1M0DjJyB
xvdLkzLKjBzxozk06e51PyUZecm4m0UzQR+ya89OnW2aFfpiYhpc/9gkL87KhJauPQIexvKlt0zC
p8bn7WlN7RjXyGRllbTB+skMK42fOg0Z4PTbMxlvAgSGQuLCjsnlp3kTo2+LeH36PaD7e1cEdhTj
pcfhJjAwHWhqISQgSN/o0l6Mi+T7gtasLSqCeDSow1oUF+bpYnsy+RewIqYBUdewHxnsTgi5qxrR
6qqh+SNMNhkuS+2d5CLUFUQq2IUsLWBKruZVbfCCQEdtyCYEzIeIC7lxAdODgMucC1d2FOU+A2m0
e+loHfFx07dHqOP2oDm7KLHlXi7RXXJe0a3NTt+KJR+IVg1/MghGeJrQLmOAyB7Gc65v1vnfkZaz
0fYKinlqdOYahn971rv5RQVEPFho9Ea9WW0VvVqfrjmzHzYLOIJsh9/uTA6j3HDLt+euC9OPuEWB
HYgQf3ZtsnNtPIci9uZl6pDn/PW8QOrnv2PHMOFYI6ubpD99VKIl+iS1zY1EBgtWQYVDAk5PUbqN
lJLQeLYTk2uhSx0aS2q0KxoQ0Wup+jftwLLZf/mbcMJdEyiktluzItEiDaTp1ORlzCsEgJP3FeqR
TsnhQZcsdMs/Bjf9OTCR01XOh3a4JqEV8E8XbAkDFdMbQ6fH/8U34MA1zx7TkFpHq6Bw3u7N2pwg
e3jUD7e6Ra/Kag2VRtLUrOxFeCXSoCkSgShGsA17icH4tfAuqpcJmSGUuqoLql6dOWIBudTBl3nB
Flz0PR/H66OP8Gd4UrbrSQF/V+5fc6xR1kGCYWmc4bo4lNdh2dzOVv9nQ2umiSOOJNJVJbN9mcKa
iUkzyPtobzF10x3uAS3UIQ78XfAk1RMezLIY5NtzfKVv2StMXCMQAKUOh6GxHIzOyBfZce767JtA
CFFJ1FYKNuZjaj2K1SDQ3VHeo/z6AjQUo4BT400OFOSLRY/9fKP7dEWY0hkT1usTB+CMdMYCLPEJ
Sd1WBXs5RlUnHfu31w/niLDk47knxrK2hOutGSRy2M/ODAHA38HjAatv+Z1kGBTp2lQXrMFHuJqW
SBjkinvT32U/WrOYbOVjxlglz9jNs8rtMaEXbw24KFyvUr78Nukz69cGuSZuvzUaYDrP9Pp1Er4Z
xoR+Dpeprjm9lAHfXcXKvQCIcCUnNKk0w/1/z+9crPpUtYii2MsVxbXmE5CiD0WbQMLjVPzpNt/m
YwH7fkK3sBQgY6z4Te01FFNrY++VHmHvjXirJxuDl2WfcbZ8DSns1amu+EysoTD6bvM1Hpq8Y0PB
G4sE8k4C9xi+v8vDgxUpH/5tL0XQDPExyAIui69HxzLhBnHr2h0geKUDj4/4IGNOpEwQAkIc03fS
7RngEMmkBLUBhiNSAswPw3wsasLwpOUVmB7n8bGJDcQsT7p0tL2dAIx2jQl+l7srAFYOKeFB2msw
N/eI6A53nXXpTcspV800O8zm1gFOpsFpiT8O09AKCxL3w8sCV0gvbPgKUqDEPKhxL0KttWl6pyHB
GsC0kQBKe3kYqCM5ug7KVcPTqQUwXyeB9xQ7tqXl1cG5ASxDYMi7fgwE4mPqIKi/xLzrFNRyYroh
Y5D+TMFfTQOfs3YprWk9sp1VPQkbjCe76CB6qoiSz7ExrOXLRqAv9VtAPAD0dZiKF/Fo9V1vTOVV
LnKyMgtW2EXA9KCY8vDM4cjYfaA7jM6kL1+XL/bUpOzEu8QOlwxea8FKUNTp0ACjPAymR1pMS7IO
X+/O/bUlhzoeLsfRRo1v+m/Lvp9g29pt06TKiH2jCKw61qe/ukeTIPgKyn/+bQUv0R/+fwzw+gPa
O0NpUGuyufEDhRbXo/36+BxmZCpN2kq4POTP7tnr/zJXRmLAZI88BAjuHYuTUTaM8DjyIdv8tuyg
3DpTUFXQ+Z+m4kSnuaionxQTcQcstNN5IDE6E2XNZrPxnOmTsu+GZ8k2aWTJolblQLgLrb04J4XO
K82FwmouYie5KY6AZRuP/PAJOIiCRhjd0boODHgpxTbjt9N+7ohoA07qBQA0ahKJCeczkw0qSz4u
QkQ5uSkgpoOnVkWkFp5U4z8ejdkEnkF8UqfvHOEmevyD/T/TNzudzhHzD8sHeWvpPUImc7C9hxE+
0XU0QcoRWj4YEVpFlqmZVcbhtW64QOHCbtNhvjnuV5S8sFnrLLl928mPMyq8Es9cKy/H6sYye4s/
NPj7wuFQqYXnPvyBjlgd0P96G7HA018p7Jsk/GlVkHurUwIxhmRMLmbbgUIug0R+ifSGDWTnmi88
BJoE08+QYH0nRtt3xpHx3+tnUbxObwHcMSJ5ou141WRscCjhMc571UhnHih29JI1vLXzuUQEVFr8
F8SzUkUTOM3L9qtJ50azj5NE+65LZhdX/r0Ah66k7TMqy/yEIVcOwj9sllgJTYD0XdH22QO/Bjaj
VUMw0JOdCJ4FWtOqGZEaschmg0J0Jdg3sCgg1CrESb3/hHkJ8nOiTbumoxJ7oenJxwwxzYwFZ7Ne
jfAf+ml/O7/S5i2joXeYklq6gwhw89uxF6eACDS6wTH0blwmvj7Xa3LoXd4QJ3X8XVUGyLogIF50
KwcQSgyCnV0g3U2o/rlC3YJpkvh3sL7RkHSX1JINc7VZm42Aq1ZkkWipRcXfhsq/pB+g2TtynWtS
7l5NrGIos/2KE8mfKPknUK3SL+trNzjp0KeK1NRKuClahhFHWiUSPuuIm/xh+83gDJU/D/QrGQpb
nKIksHH08Yrkwv9w8sF+GgFYj7QduIiTS2f0VR1anIpGVEBy3C1V7xtewAwb47A4P8U/2lsiEDZ4
5DLX63MLuX0szw0sRdtFUTZ8bYXaP1M79jMw085WjCVn/t3MHPu+rfXaYJp3G6PLMAbCxrVfYj6q
/BuzAeJHwOS9jZZA8ORHqaUn31/k0g+KZaDiPrNa4hVzJAAWeldKk3jCZB2sSYIIh3WZfdgwgdhY
ligRJmuI6PXwuZEAo8kPbIhkJORPP8fkvsvZ40n7Zf/Iw9VP6TDPHq2/SrC2W211HWYqCxO8WraX
YdUBsMZwazspu20fCDjJy8a9235kOu0JXL0nvR5k43tv5rgfloLSGsf7YE8ZCXFeoHwaDWtJLUDl
xXZBuIeNkWq5xGHGVOPvhTYx4BkEgzEDlF1r3m1Xsl6Yem4gUbRo0/PqZVN5I9MhtDuhjgbEaflG
j1rGcLe80dlPQpRGXkysyBrS2zTSJBG7T7K2NVErVKL4jWRjhyQP+KwpGSYV2TwfaeWhGqwpn/oE
1elcA4s0dFeRko5faxWlsn1ktRTjgoHBQlsO8sE+PtablsUtSmvpGtnb8i+rFKtdQqiv6xim9vpK
qRTpjXUSNImPZ3szX/AmnpBWbG5J9E5Vf0w7NOx1vTzS6MKrJXOwaMxoZchCZxmfmP18aYeH/X+v
nSVw9CmSybyD3Ed1k1VIK/+tRL65zLjrswuOdEXkdp5k3wzOeaSIx5YybGbB4s9TpmyKAJY2MqZT
v2PrnZWyfhMWCrkVJLJE1qcAtsFlUUVci/zlLNVaC3j8XjGNscht1+qeRa3o4deQ06N9YHKOtMrr
TXbaLULTKBe6NJ1CBEU8teiM+/M7pyoQ3XMkDD7LANo/03XZgCOOPN0Whn3cOBOM0Es9dOltvF7+
0ccrYcNfUA2XwmsgjeAFharLDVep+4PSr9rrR2Nt/ycpWDUAt61+oUZMCHuCa+aQhCZYOSOf4S5O
MCuW2Pg3NbyCdj5eswRb9A8duBobx42gBt5jsuE9TU70gYzBgDdg+1CequxS8JOs9A5f+uzsNqHO
EQKSl6cfSHyEUdn4+jQXwti3CVNP7gQpOEPgDhfeLMreECj28yN2Mn72z4joR+QM5DQzjMMZzkFe
jSPe87WDUS1ZCsEKRd3vfQ0OX+5AgrqzIlkG+7o4pXBmkcevdIzNkbGoPtRgWI4X32c4k92NrvKv
P2VUU3yBvndku4cuRo1pqE3EI+YbI9LwOvzAxT/As34A9eBnqXZsn24XsFgvdgAT+VjdwZqdP2Oz
8JiRVZmiwOdC5qQB4kwbqS2xz6tiMb8kjK6foXp2SyMavWjFsVF1t3qNSU6qL69To9pU04Sn2eHu
JePOJucWNJTM3iF4gk+8ZPYkAX2bz2Zwf1V9+zeUfzIJU4N5gf0vHvXe4XOskgAKusEdQUM/+VlR
9PeXREa50D75NqhVW5tJpY+3jEpX112mbW6SxmshD9M2oA0LWfvpZG0dsZ9iZU+skVU6kpxV2AUG
b681LkFf1n0Z2tQSY42q/Sjflrk0UcDRDhW0RGcrYKpsErlTfGIYT2YE769YnJzEIfynLLoG5Ekt
m/XFHrUrHyCEsP6YvGJbHNuUeZF9Ocni+xsfdhMBl4F6+7uFkDcNRkooqhzZOE9Msg==
`pragma protect end_protected
