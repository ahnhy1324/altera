// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
It+f0YqHmOb3/ESUK8yILr9++KsBUpWJGKBSa/So8gvyLdSeRHN17/CNxpYrqvzJ
/UPEvaftD3E54JY/daqWaYEUNUIIWR00LCpKzY/Iv3jgo0NawBlBd/7Oyby0DmM+
lDclLBXxC9GB66Fe7crouR564ZJM1oDGWiR6vNpEneI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 61984)
Gr/znL4eeFCKFMPoNTysXeMGlVSax16OKKc7bimg+yE9KkCoGmXDQnXULxAEdopT
8kLRw4YOskv+G9ry59CNm4/qrBfU5NuVkx5rltS8+ltJNcn9ewrGLyebNgZOKTot
+mgE8JasIdThgByLu2LvnucYYddhZPZPtpKcmYWano1LaOI+2lqu9WFruH0tBLaM
OCGlDYk0HNCTrlhRPqKVseYSVZ4X1wq7w9xaQYdIibxxmua7jIFvg5ix/sh6XJbf
8H0dIGnQFeejIlmmzX1YPl4AIV8dCsLgGJ9DVFJYjsx8nr3+BRdLrLnNwzFcMHze
VT50916yIu8ewpktYKVanyYr6E2swnSWXaoyfPH+oqNp4IKGWTtZhwiD2LSYBhJB
O4YtDBuCpKGDv9pCbK8ADvYypVBmC8olACmbj3LOi2FkVHKMPuxSGCCkgqGFiKNi
j5HF2XtBTrUhbKG61BJPgjSE8RuV/w92AtAvp3l5Q+lMVM8ycxRuTG/i8LDnSxYn
LveZdpQH3LjDxEf+ifDXfPbDQ3FCC634HZbpLETTjBkO4gIDvrP64S+JVRwlGX+e
zohQBu9y8WzUKnR0dW9GWDqwRjleNsAXVk6v/LHw3sU7BM/oS8kgJrZ0KZY4Nwrm
axL7caaKE7/GjosuEcIru4bJcRZt/8EcI9q3NNPIoh6dPAF/i456dgm9grtRMrl1
LT9U5xldnGCBnLCNZlleNsq8lnumkPUCrSeeYIH/yRj6Qw30sZlB3wMUWnN6F/UW
JIr6opoGRPIxPbBwYFji0sbMlO3UY0jCdAL6TkVmZKkoOQii4fp6nC37sCI9DtCz
cneJQMAkMS+G1yqaNSdAGj9va/8kgeEit5p1yqcoo9SxS7/wdEKOsYyHfM1VqRd+
J2/NrtUlSe/R2+y7n5G9CdDvbeT4Dv6INSYrdPU2w4GdpyxaCtDfmFK4aJQmGi2c
EbsgACYcfgi+qqWh5bDCnrvFins0fpnEryhHOxTp+zzjQFlsQjR5M+S+ZDd8L5tA
B6hPutD5CYIlEndKGlOMUZypJAxm6gweAwaLOcedxDelo8Y7lOW6ch3ReHn6NT6h
j+GpAYx1DVTtj7kxF2cm8RXU6+OVeWTuwq6Pm4wB50SEpaq2jsRhTgdhpHYLTKk/
LzZTwlmVK5VcolhzG8+YKEaexDbiF/yowAio5Eq6cROuxJuPRqfpSxmJ8WhAeygr
vAocZfcTJdIg5y5X57r2tpkJqE7jkRUqDgK7IKMsWy3ssI+6CI7ASWflVdxATeBU
smf6dCQeuZBjs5ugmiUeusdVz8XoYDFCvShenMw4QVtUx7Y4Wxm0qYKLgsdm7AvK
d7/QnrBqQPdGzC771uU9Bqtg8jhHFpCeZAYc66MaS76X/k+cU30qVise7UrIfXzl
Y9mCTyeZKYfEwL3Pd4+siLJFhJaIGrDfOwnoyZsDpHKoccGryZkMjYI746CSF/en
c/LjwqMihbjLz3UV0+NULqI/lmV/c0ggRRDuOxG5V+yjUabtYIhmkgPhW7/PfYO8
IFlMIVQVFR1IINFlMEsVJo4OdOVoO0+9r0YDY8tSBm+lrDoQsBYpcMuuvP1neEmq
oIWUpz41mHY5U6X+nhRJB+wMdyI6w5chMFAj+3PTyUktEBd9yCWUQcF5lJWolCzD
zN4CrVk+dMt6JRVv/IuSytuiCbyeAhaui3QAeOGjAYj0tAjPTruxYX9dADdhwl4i
bO9++9JwJYABZej4oiYWD79RTjlJWLfqnj52kwy3Oc5yrRGv9vnIMtA+lblBCn7J
9GqQ/nXyausq/AWSYvgOdtBR7rLVMH0I21iOOV8RoOhBscmIjglNuIlbjKuVI/Vq
GW6azCMBBTUrKXdcL8CLTF+BzfgaApeFSl3CM6bApJVb9GsUWwRfQJUJq5DwJrR6
9A1pZ3ZT5tIonwAJaS7sQwGAbsyMyAsMtBtxxdx7QtFlz7pv1YFABobuqjU+ADL6
vZJevnjlBu8bXOJu+b6qRAIw2EhJKbgpxJbjUMfQ7Yqm9oHpF4ksjTZYdLpEr1nP
kdpI0dIUDLB9TxRCQ8/2QCdledTMHwDhM+5Ai90y7vMQoWYEqYL29AQl9FKsZ1gS
+XGFV97SYITHNLg192cXyIuZMMnPjxycF9FnIZnaYoO9ltVK+toMzlSMSJCEPYgl
nnY8VbOTpoTS9UBcFw5sucoMyC+mpvxVDN4mQbSleSKf8x6d8XTRFDFkNcJ4162y
KITryhQWM5swEPG+cV+c8mEciHklEJR3Sof/HdUIuzbGwSpDZkBo2hH1EtJyIfzO
osbCPZGLCXNZhVdXvBywCaNz+NmoXZBca59P02o9szkXDQLCFox6QN9FhEimsuLe
8ZWiKz4YLgr4+pnXjbsubpXdXzP1m164CbH1pri84yIecijVvYWTgnVwpHOF+kfW
WRyfTKmLVD6SNdcV6bXnbH7oi594dJu28AQqBfNY485iyVnor5QETUOB7deUOxhj
wzJRdoL/IcwORt6KuzhgQ61k5zkOq2p8iOVe0KnuR6FUj8irAPP9+uty5ysDpI5U
BpgXl8NW9xKGo9d8mjyhhmA8Hjol4czb6OiUhCQOsmEPYhic0t57yq+yrHN2Evdw
S1O6oj2xnwCZUFQhs6y+vnHk4x7f5gGC23E7DoUe1rKKfo0/DrL25m+qWm57H0Ws
CGCWLsqCw8UtEOk/S+cHdNzQB8XUCLdh8kABbbXgeqJRP53VlMzUkLzeo8/X4Mtv
sms8xDfW7KUvGx+OaSGT7wzHWP2MPjmJtZ+ptTmXCDt744uXoxCipJqFkB1gp7xp
983eLPVc2+MI6q/7hp9Rld64Kz3YOczz/rd4gWwpkMHtD3lMQ6BLKa+f55aV1Dnr
3VOdz+cahBwyVSXUHVJGUMvAVbIINz7mTTQAulvDWAXRKIK4CzagJwI2l/ceGl/6
LOIvqEidJD/Uo48xWDrGnWc+bDTWETIdZNELBOdAQ/hW5SO5uZk8geD8ksOcj1WR
SJ9rPpnd3SnfbO0HvBJPkj0PN3esztAalCtTrx37D8fZBRkeUPb31Zu9cSi3Et97
1KMofM1Stc9YAZz3QAM75VSXHw7GEa/hh/D2enT2HpWIqpr/SkruULCvMT6/tcYU
ZhDT6fSL+rvTBZsIAbx5LUxHgxiGdt7MQEBGlOPeQoc82tjP2PSKLHR8Bpk4FmKu
COqScMmIAP5F76pWmqXtM6B42R5dsiYLBX1DAlQTYhni2zpXWT1ivF5+tRoh2mIT
UfyLItH1VUK07zivr7q3YacpJHqO7ASxiqZJCx2RFj9VDshwOnKrbL88yeg+GewJ
IDGZg0XcQ6e69LVcB/C37YY/mw2WXJHD1yzYHpYLZSTmhRG2VuKi84K7iQeyarjb
IXz8oM+mIBFZhCFZRQ+UYPYskdeY1SSO9rfo+pnTpMySxanD4sOL0Eq43+VP0+Hr
XvrJrwc5mfUjdqoSPEuzUnC9N98ZPf2vYU5UHejsoa1IKcgvmYVNoPAUv6SmxAkl
Z3NkAXI12rq33Z5LdjmZohhDE2d9/um4I5eaEEKytJGtxUP67RFl8rifaic0FCV3
ER/bmcciRXIXbimroTFHYdSNMO0/BKB5YvDglvCapFWWSxghRLO1WHq8jiNn2tnz
/wfR3nIQLQYQhcNBFkkqKTjkKBUut+3Jwo0RimtlwhgkY5BeSZeJ0gC6ce6cVeyi
sMPkITqljM0/n2g9gLLBULcWal6T3m/pcM1oRSo9e7eW8e/SbEM1H+uGSllAO7fX
/M3TcHV1ooqOXaIRoW2ZobwGDNREoefwSd+Zan/+4fxvk69YtW9G381eJweSLLZ/
Z/AqZQN3+lKDh90jpKOkbvObxx8mHva4rS6oOZ3h4XtmYCwGU2OYqoE9uKH43tzT
CrdklsaMlIVU9wIFK3paJV3aH+rqdllkccDegCuznxdsKLtuvQpdj39lgxFtcLbP
5smWV1yi++7ksl/aaL1/2NhhCR9cnYOCF50dptbWZOWQahV4lyrMEQQrtGro59sg
j8m5Jg5SPr3ax5J94LVwJjw/QclFwIjKhvCaLeUgHR+lkqESON9nGjwXFejoPLG2
GZvWIlaEeIQdiMk4SHxoBk0nwg09veoJGj7Nztm1nCpBlxAce2lUVErz3PkPI+hu
m484lwmZ1BkaTLSksnH2XuzQtmgxxcWBINzBWv1L+smQNec6ko1Qow6AgknkJFf6
WcN4pzXrOTaRIrn9nyvv9KQ7Yc1DxnBoUEanM5ZBr/CToHbDqHkA1GpMzZSSzv4X
CKcUqGe5MSzngr2rDtWvWGPTxqIsbJ+CoCQ4PWeh6U0yVZgDFSLKE3diCeLvE9DT
jLVKHbU4RxRHdRu5WFsT1Y1PFPh9EN6PpBEdVlQ4iRLV3bgjTnPbttwRAUNPQ1NT
XGAzSvbnxnSxPmPuU3Te/xbKsoDbilFwtAA0X4w9GG0X7gJWEyD9yPO/MWghYx/L
gV/XyxSeJlHUKyBkLk6C7fyyaU9dZdT1/TbbozCIXm/Z1oCNzjqPl3oMrJzI5rd8
CTqiib6qA+StldukGrtvtlLHtECosEmRUFStqvjqw/rUvcNv40nvyGUuIKFvjpTM
DAuil1jAtjQKKuhxTLO+PoCNaa4hmE/5WbgNOQX3o0L7reJeD1ZVTvWs5OSlP7u+
wz/WsvT2JfjkBmLqJi3e6uM3lM7oO311vR/1aRM9MSKpA4/LwzIcDSIimeFbtnKX
4RZBPKYHP7DCSvf2uz6Y1nHSG++I0KqyULoJjQBoMoxWN91lNInb3bIa1h918JLq
wa0HSb8wgISk2SnImvOPAPvhyl57C3BWE+3H2MYCs6rPUB6MKNQm9a1i3/bhw280
JBK++1nJNwtTEan6ZfFJgeuYSEHW8vngaMoTJl7mcc8ur1Mr0ptQlWT7n5A+7dxI
YRGthQvRxglltpD9X08eOajJa18YTgBbCeEQeOkJJo8lJRRG4pw72FeLPFKs6R3Z
zL9ry6e+rhy57d+zdqXOhs2cT6+LNskgi0p92yP5BtEU39R4I3QheYiLBSQ4sMfb
Gq4Zih3wugD6Lf51v5vyH4DzJEd2C1CkAPYx4GxcNbrfSIkJpcfwgk3c4eE8fq+r
qEMhbviiG/Ve2rNJwCn/oesszenk8qiwZ2HuRb4T/24o+GG5ODzE2NiQCVW1CQTP
CpNjhyrpE0abwAIbEaW8ekH2H+chnbhOxgOhn9GQmS/6taOLyrZJ8ObVBJAbx1qw
6N6ImwUuZOIyshZ5ADOlD/m2q3m00qXflJdR5G0AAfqQ3sJF+u0LT7dxY5hTPWWU
mUf5NcE1fgxYfecjRiNzza5r/oWnMxF5HfdudMwcfdxTnN7zwkua2ZF8UPQZ9uQp
aNV9R9l0mSvnlotD2VVn/hZP/2NJXGRBsdkoSlOBLbv4gyToxcMMxd1kLXSeKKtW
88WTZfEFjEbjACu4ra2TC6V+viOwfieRaf6H45v+mcEl5ZS5ravWCoxrp3E+2xQj
WdwPTEs+L2NK4gVF17M97SE46iwcL2Ez2UmlUmFnKKFyI5j/nFH5tLcdQWcuN9xn
i9OFRr/6IvEiwn4ufubLrp6OX9/JCX5IzyPGV8fsDcjWuuRqHlCCsnXVaTTUBJ5x
sk4/iHe46LQxV7ONInb/LAcs/n5oYobWy3nX65Uz0LUdpdhaP+UI5/RlC5x/eYdG
exmqGA+QN0pvNsRAdPGsXGdLjb4adQ6VKAxoSrWkjDhaXzvQ+fnIStau1iZc6lvD
93T/5A4+y90gLZyHpRCEhsztPrgdSEXaamF2Si8jxaaJiC9TfZEqlXWKXIjdXIIg
BvAe7v2RykTXLI+Lu82NBs3LHaXCNFzZgczdD5hZvTnEyQkbiMEzsL/L3H5qC/hS
iFx/HhUSsQh7Di1FZ8SxgjGjIcgQVGCUlVHJlzsPLIMAnMnjgkgnRwrPKhSnQ94K
sSETDEucz7Rmc/IpDT93haWH+jKzHS2OBfsQCT/pZ9VwYitB+rzLP1PRj0egVFn1
Tee9bV2eElbELEsPK4dWVf9ZlV4k/9c2Bsp6YbXMjwRQu5Jef8Bo91vJT7HIx/xf
j94OB5q9HWIEn6c5ilpbZQXDEjzpPAJ5HNY9fAq/bxzH+rUKTlRRo9kJIv1ue3lh
G+TYna0vaRgLUrTLuhhEUFdR6HSLO0rL1GY3arD0JYjxkRbP72gduvQizCe1MWNN
qKRzf++ojYX7/pC6gaMQKLr+VqXOmLMGhlL0gAG7bjs2Nlo9KVcGDufl1cynZqym
CJgOwLSE6HLLJbdfoyKaBU5sKHF7Rdm9GBcrfhjd3NtvmisuVva98VnaPEAdsAN3
RQYyVd6tPVDVonHV9tNW7u3fyVnacDQsH5xbecUEre75XHF7ayKsfWvE5D1NSf7b
2CpOiebLwh/Lqa/sVh2Ak/e1tS75cM6mDktZ5wSmV4XVDJwWmN3KSkRXJexCxJz1
UgIeg8yZte45XonU5MvawK/AOBtMggfDCHwOiS6oCpaPxgOUipP3LRaCu5JhGg9Z
RUD9BWA+kMID9s4l6S7jUykwCajJD+kKG1R9iYfdBGdn7ViaALxYUeR48HoCoo8p
ScFEfLFiHPYiE/TmkeUYXl4L85Td02UsjVRVUDV7hhyacq/GMNsnRYzmIdkHBm7l
Akux+rmzUBr+CHbnSz+XTQUHDoqluofzE84HObcjr7z/4PE1oDt4QK7DRlHKCtlS
VOzfkowOaWBwsgTs8mAh/BICo1b8K3Vk0lIFg/YnVBBbsNWimfFZ24m6lqi3ryOd
pyoriW3LxQzmg4nbQrl6qhkKAX8TZAgcpuiaNhYoqEOR+FH+CeXdfnv+T6+5k1HA
1Wyr4NaE6XLrciYMZ3eZ4pfUvo8zHrXQoOgcOGZBCmvTSI9Pmc8A2JBqWSH2EShN
wr6PWZZ2H+V1hxeUr2w0zCxACzSLxzrdt8iisSCKyYeGnjNT/ooyuuUjhjRHTEr8
/n6p4oYXsHD+UMoiAeMStTpzwyIWj8h4fY6Ug3tTRCxBm0NR2uMsKbKskcyXRXR7
cWofGhBmTGaGAAQurD0dx41ZDFCdC3hIXMKDs6e9UJ+pAF0zj+zl2w8CyPrmisdN
VKAYDeQz+DmR0peWqs4yRbIJHSudq3QOis/MWkU7L+uIIrV5zOZ+wdOzKtGPGGfm
IT7MsvPYYoSbwXTtr5wm9EB/YM/V7s9s4/feqhSeiblmn1EDhl233ISsibHK27nK
WLkiHUx1qASs9PJzCPkG2yP89VrtxiA3iJgNhzJpGmnoQPKd7S2sEFQzrwKioUxp
Wiog6zpGwjIC+yW6ojzeC2R8UzwxNeTmOnXgSYa566gpRc+w4dt0GwIQAnDaq7nM
z472UoQ7lS9suradD5YXRukSRfCccxp28WB5u/y4v2iV62EvKUjGupUxDEuilCYk
xC65oKcQPw3qI6xpQfo6notwUgGqIU/AkfazDNbWekxcPkgiM/8o87xP1yZJ1/VR
uD9tLMMDe0UmDxe9y+I40QsPV+pCWtfCFslnbZXONw6iHllHkl+gJ44bmvP5yI0e
QN/2M8O8ozxabv5OsWAJC9wpdbTKTMX3leZut2ZU71XfwWfHTmHwxk26Y6boaohW
/ULX03RNzVvY/dshfvt6d19OwPQP8Sgjl5nBOS13dBO4Iq8kJ0DNR0QQFJxdWljS
zM4wwuHHI2M3CjG9A6LaBIf3k9NXVTBiHMIfwaIXKDjYy7M4gTBABrEOfRF3YaEl
90itO7LVezyt5g2tSj3ss7IUvcFN1FbyxGJu8aAEq2yr1r1jbXvYXKfdZ4VM4k4v
jdmYIlZqu/Uzwn1YyKzp6sNSJeZeXGlTjRHBigz1VZpe6VdLqpJc/WjNyK3BI+Rt
CqqQXE6WUeDoz6a3eWvA6aLG1hm8nx4y0PysB3G7GYUmshVvFJPcXxRgDtGfNRtF
K3UfR6fXhOoB4L/1w0cmoaXlX3my1B8aTm29E8FXyyI5DMrbAZ/AKB30SuiYhtPD
53VCO9Fs/4YxCWIgkzEHHyyo8DEkwHxt0Ik3D0M80f6xFG4R8qsIFghKa7QXMNfU
qrLTznfEjT85zhlCRkqcW9BODqB86ICLs4IDug6KKTtMOEN/oIuTktMJ2W3G0c8t
xLJRIS7saSfs8zn7ao1frx1ArMJ8Hm5GwCA7NnjzfGhSZ4wxCKF1Rj60O7WA2IMm
AEVTydmnB6+CDwWOMhWRq86LMMsOn6c88/aEA0guuuoF02WZSGtn/WE+z1igzuqs
yPRmD79lkjvW1F97fFR73AUiMj/8RWUxppUhPXzrLd6f/YLeKK3HLG+5AaYUxypw
HtlrQWHx7g9cg83KVrtQWI+ImS5m/qfAAjmfiSEI5gwRRswjCkoSZEsdXUuiJCHj
EkfMJPZGOq7WCbzaplYm0A93x/T2MuvGpjU0Mw/wKkb/nqG4okWAOgSuLI3Jg8Hq
zWVVd2h++NkPI9nQE9LZbv9nrmYz6AcU5vZ3UyK1RwmyzWaknvfRcZ02OWGnCYoD
iw9K0gvMk+vXoBqMUh7NmO3m09h2SS7/k2UX/5QQeyidadJtcfl6g5xUfK/PWY/0
SfiAXRKFP/oGDkMj3ZxID8E9IPP86/OaUoIozZ2eccIID/5VY36cSi2opxstNDtP
3CAJxaxI4He+uR1iKTjHYgOdQbuQ/J/Oci3cusPgtyGWcORr7IQh+tCcQYgpnv2R
fZ0O//1rsz+3LMQCkcTIZFaDYzO/aa4cOxaPS/k5vJ7I0+2mC3Z0YZzMYwU/LVNu
5whpQRIHYMqvXl1MorhUZs/rChbOg2Yrc76i2+0zIScoauYz5hP/5s+PUel1BlAB
tQ4YY/DURtC8I9euiALmiqaurqgezvXf904u36v2xuz1RG5Rinu5A/Nn3n8MTqu7
kbOgMP4j3qxkbhzpruDW8KOsMzpzLPwYQohv9OiyonbuQArG3WbY7InC9Su9c+BI
IDSPhcr7Yc19EzpZKi7swXwr0XvrbT+PgpRxIs6cZ2aCMr/U//71EtiKi2jP1/Vl
wZEnuYi3kujAslu4dxrXtMF2voehvUR4ECpD8Eclsh0E8/Di7G2w198KplZA+4+w
7gHt40efS8a0BKXit8kFLXujuCQEDA5L0yIXpbPmRg6zeeK9VHZohklZajnJr8kz
jkLpG0WkL15eMCIikhQs3PBO1bk5zZd9dGjzxR5mDh+2VkNVKRS5ObKMMqFpCd5C
rmv90KvZcMAfS2i0sjxRPghyKQp7v4EQhe3LtzPa+WoWttjyStzmAIRrjKuV+TzX
VeW8DjIx4AGqGrgifvFjk+uZkGjdKnQo0NoBfTPNycNhY6ysuhOkEkxwUECh8ZKB
jlnqSqfMi9eMZ+q3/I4ABuyYU2kG+MBrKa8VEthonui7LnmP+zJUEzsHo5iRI0Vu
RdR3X5I3s0+AIHB2BeWiUPyW51Ly9WR/870XgSVMIvmWbQcqg4LUm7rrF+/TpI9r
OgnSuALE2nibyVmuZ5WfaVRVD3xjz3YU4O6ENnMX373JKnHRGGHbqqhYYli/Y8ck
7DnCkZOvZeg5SZlvR7UxviACfb5npk5eSYD1bgGlRaD0T3SBD8LW62hNsXN03BZH
TKYT6o19sFZK10npS5yA2xrxD7y7pVzG0FmpjK9z/toPcYVBcBkM2cqGEphhrvts
BNFe1PKDoMSSj+4+KrM43QTnC+Ko94h7z0Ds2bP5hya0y2nCJeixqKdXNZFOTe1a
vIoKXJ67B8ctSHS9C/tqpHcXUjXAOfCHmMxUwHpRJVI5u1eWgp95X9PlCuBC0tR7
/bsQmSIdbWt80eXfJr1S4B2Xc7hblTuEzO9xl0e/9nAUgKua42s6qihEjGHXUuyg
XpzwK1bPc0gU5du5dQu/LftBGTc6KJti+cw9/YfEHimCXuuEas1VZ6oEMuM8fstI
OOIlAF+9v+MD1psNl8wgKCsHJ/oF+2rJ0MD9jPknV/5BYDN2bSoP1CS6AP3o+Dp/
G8SVH4EUHUR/Ki4PfYAOyBWVgYaAXBfNZJD+7hIof/NOyJ/hWl4IJr4C/EuIzDt5
sJ2EyPgfGrWaCOM+6LA/amvpYvgNS6bd79ewVkqAFIJUmoR55tTsIvI2lI8Qq4AF
XaA1GWPlPK/iVMtelaLLw6cDqm5OagmlzqYoMj9vvYRzFN7ViksI//13wlQ5XyN0
bUgSI6hWKJ/2xyyJJPznqv9q7y/UO0S6f0vDUBgMoIHJjuG4O7LR94yiHZLpys+l
+RDKBuAFOGQgNazhftacQfJOqY7PdBcqkOuoIPHnGuf+Pxu5GnkYuAuFSKFiX+bl
6OvdTrhC6frDf2bybB47ocurxtdGl8uHVD4jEc28OT78ihldTPrRzSLYpo6P1VNU
xnq5NzJ5rt4INoR88RP71p4BLb9cIIN5BpP7p2Y2hF56pg61BbgT39lFUhl8b3rL
KQq/LP5c63d6iv1hLYw+EC8WC+uh9W2ICZqcf2TJ0yy7NDUAaNIolqZZlFpRSKQ8
7RN4vR9GA4ryiFeFj+wjUJ1X4t/tCcQOI4pN2VKEWEzw/zd0Gw3x2r7GvzEMtwad
e8O+xqYnUCy0Z6vyCzwj2oUX1bJgbJMxt9lhgNdnIBD6PxFra91Vw2usPviAWK/5
W/f5sIJ/6O6GDFBOrVqSxr0Ks+Wqqe7IxqialmrhAu9TRq0zB5rOnauTngOZlFRA
YsrlADctdtppX6zHe70WLzgNdHzr4QjNLbIZ+HSI1KnqI48JtcS9CF43ifUeKjAT
OsJMKfbmPS97UjE19SzE+4TD+5VC03IkqnjuIJztphZS1M0IjlbjtY+KyWfH7lj4
X5kq2Hh4C4r0NApf8DqsUbJQ0+gfi1p5IQqEIgD0mEIw4gtoV8K6N8g742lrk0R/
7TBbF963RwUSmvJNiF7iqOKoNDbmQaqX1OztU0v40hnbwmdzRkG9ESGw3TgpIeLO
LShWh1Tu4STrF7FaoJ6OQFFVp3Qi8yHvlU4+/SwB+8Wo0ID6b1AyF164T130sjr/
/yGlXcriwSykH4UbDM36wegrCS9PLd67pJXbbwmJVsMsdz720qbqe0SE/LOjWfDM
ZkFKFhLI9+5miB/DnSBGYT79vFJsGNxdZzgt04oq3C0vZXrQxXG7ghCcvz8/V+Dy
B/ioq5EBSaowmcz3zYEq0te19r1ZWhm447wM7zQBSQEoWt5CAsBOgezhVd86Oukt
CS+TKeIBeKAsOeDxlNvc4LG4mWcR/xiVD4BX4mUXRRS6526Dsd2Q2mLwyQnihlw2
V8e7ypqlTITQ+sBAkvga/y3aA1HrLRYFLQeO2PcnXL0PDhB7HNlPP8ZIzjQXPzTD
cJUFA8PBCz8u9P+2ou/F9FKKgL6PoF1ZAa9B/gO8Q9QVgiKU2605MsfOMsKoD96w
VCJdkh7s9N+jtNzj4Vt+1qSh9BXwGJbq+b+LHUNgo9Cs/kFR2cEwnviCFnbDfQci
xyy5EXgBGt+pciUxbhxXie/Nm0GoskQINmQav0GeF1MMDYwOR62+TXe2FJFAR8gW
Tnyj6HKTWqhjLIXELyDKxAa5EPv2fC9fz/uxEyKBBI3fa57lcWS8SHRVtNOaZt63
ZWt3JqpvFHR2+JOaLnT1uGMSC6jSxRT3+BRTRMUuVZdw709RrQD8jAYiRzDxo8lW
tuS1h9AwMsmvhNpIi89Yj2f2TXcICZYoHKSeZspdtgZSUvJD5NPCJX4almXhnpjX
pSqP/KDT33vp+RGjw+4aCDmQbK4MRF0pO1QsTREiWWVVYVJJ0M01TFN67mSprro5
yqXRlwNV1guZZJQIWn2UsKhw/D8Kqv1Y+JXeAW7HHOhWzYumZifA6iYVwgHkf1iX
DsBuumZu6B15PqJzqW3RZBuq3Mv7Mq5NoUkX7wU6Yq3S8T8OsmUewurUq40Tjwnd
pUyUdLLJ6lHI3PUgltsUxttEa7+IKSqitZpQtzNHeI+vPz4vsJR7WxaXaLX9wkep
xaa63nOCDE75E74PeBzCd4R2TNsGkghmX2sFfdghIJH8j0ZI6TcY0TzT4TQsn1/H
boZQw7fj+3RTsMTUUI2zwVgvLwLtMAYi0XCX1VnB2FRzAGPauLQWYHGdNe/79vve
WvbmD+SvDgnO+6P8h1TSk0akbLhSBh+wbQKWbV+xlni9fSQjOLfF0qOA/pxrhkSp
El00NQGHX5POpLif03FiFR3X88VKBM7CFS2FNlgW1GV60a2TnbmTKnUaWpcmufQH
WRKMDUTfMGYfoC7LPCkTPa0D7lq6KEf4aApOcThhF6MTOq5QGvzoXd/aomZOrJjm
uwqVyL1Aoq5UOyoKdnaYS/zKCh4BXa6vm6+gAeaII4YTOJ2I/Ytn5cu1hNP9rarB
9LQu9vsaQ7ggOfa7Vs9qQlCPWluf4d7RlFmEkqAK2w/2yy8T0iaECysxZvPYhKdA
brXAe0MqcmTyWSFX5+xOc/Z7diXbXxMT7HiJMIpl98VGmfPNOT1X3WX9JzaurcNz
4ND/tB4S/UiMXswoon6r4OIKRhLbWXAZIDDmP7ht3hBLHu7rQrEy6CaICdcKT1wM
tQBxUjtsWSPDwMSCr4eIbyNIAHGJRy5UrzXib2EfqQSr8GOZ+cUbgoxv3KoGJcch
K4w/gio+hESbGj9OJcjAlNB5ggYPXDPk9gtc0bpUs/GpmoXXFN/bIbySbE6KMhyT
tdwE3XHyzBT8voEwExeYuZY8OhbPEikSmo7MtLJyrH+pp+zV2k2jOflMdij7ZENM
uam4++3rq2T+2SF19lvd0r+qpNYlHEKi+WqKV7AoGNm3q8cmjpEfyUG3DSP4Zbfx
hYyS1G6BZVPBQP8jSvikuv/Y0kEvSx6AGdx0fD1XsK02aCNDQ2PWeVBljN/e/wCX
PF0tyyYWhPpPh67tOarDiAFTicttFwK0lD6C3pzoXTO9fuQ5eGjpXiMaptqiXMs5
062C7469XOb6NVGa2ze6QNZc/ponX5pWJ8ZDF1/aHebnq5qL3o7hidAmwPvswjqo
fsPWQ4vJMmi0fJgMyA2pROhe7ZsfHa5yN0yX/3b3tfjSqAS1eNUTO7QjKibFDNRi
nFpmja+HOXz7oTYEyGNXEj26CUcVodDXYWJwz6svl2MbkmxgcX8SF4cL9d/BLZTM
tVNxKeYo3RhtcIfySyLQzmtpW+XvLRNq6CMHFAeubFGb8WVnJdwsJ02tJVUS7xj9
Xa7lfVHduICG6sDZVUpvLBa/AA3l5tEUHT6KvhOAhOYPQxkGupTcg+RS0s8gM29M
G82f/NkIdzsD7moLWebQ4lrHunY/BogVn2RwYpPu13cXpTjchGPlW4d+6lCpv1Ij
IV59H//YDCqSiHp6WHavhvoKUws72v53Od3Skn1RnfZvgrVQZ8LtyL7lZNO9hz32
PrjFiLAzGMamU4SSYqgk9JQzo3C0dI4zes8f31N9yv/ct9We2b2sXBANBmk5JuO1
7crybZ/eqqGZNfVGx+USbhMUMGkFyNG2Kore1S4bU4GponSC/cfyyKfQmJ5o8RGe
wrQrUj8c4Oarrc1BEUV8qxvx1T5X/+l0kXeK5LX2MbeX1QgHPRnB9I9mOuPSv6vm
VCy6xWBki/6T+Dathol3S+m+Gsm/HOZF0QpIwhFcTiX1bH1O7jIO4GzdHt4v/qJg
GE+OL416wlT3BTw3OQqzKDr0v2NF99Ew6+qWGpxtYzK59JqfQ5b43reQ/rf+2qwo
PLiBbNgwd2yJmrC2itPTVBPsZSCES0SRdBChmXzgJ1NyOKakeSqsaI7aklsp6nwY
uxv4T9mEsQkFbahiy6TRSi0dPsaotoCvQVYjF3z3eqQhhxsuLJbbGmIn9uBztUnm
N0DcWqyA5amwzu+UIfTPYh3Z/I3OC0z5VghbdsunAROZiGRbh4+2Q4Jo6Sf08XKu
gnsTyn1rAfSxghwz0H9fR6eslWGE0VP5GapQJU2qc0RdNBxQbVAcbqFB+SXAFHnE
qvnttOdWQX61w+34b7mtfEojHsi7dfOSdPu5nMju7VdvbxOb/IC7I6En20kJ/l4s
ICNMsjymu811gBci+39t83P7FDwc8jSP1U29hE6nhSSh4NxXFXwgSR7wLAj6S2N6
7wHuEnsYOGU47t+kYwE2HWPt11kVT63mJl+LjoT+Uw/Ib58AXxzJYaYOc16zVj+A
+S0F8g5bx06/DywFL25NBl3qZFwtvJkBxW4OOMc67agRHkbNjRotXfc6q/RuC20o
PKqSygvpBIH2+GLxITkhNbzrKInnhjhvASJsgnbwqj9j7N9N9Wzl2cVimtuCGiC5
s3hJHM5TCLrt6/Om7aesP2v7Yz/RPgMs+Nk2rN6mxa/TNPNS0tZttW8yAo/FDZMk
GD2J9hCNEJcuW4l3XuHI6RmIDOR8Gb27ZGkl16qxZWk/9oIigiqdJZ3SHxRelUj5
+GLnGRx3freVmEXmQm0Wbr4nsODhv/wV48f9jNWCFKnuZn4juhH+REWa8MlUNf5b
fTxv0V+zmkDJYnrGa+RLTKxLuwFrPY0KmNosxLZTqyzIgedh9f9mDmph4xb8IiRp
iUY08h+FIvpgVWQCBkIKD2YOtnqOyS2jrpNIaAE2lb+B8Tb98ntVu+L/0Z53nTkf
ooXPNvhwlDgQOVl0EHTCvr2lNY2O77vwRjiCkctAaKTnu7AxcdYkC7PnrVOYXrza
bAtaHeSpNrKssXMyILuL2K9EqGJ33FUld+2LvXBip9graVLmWUvOHl3DxbJqJntl
IH4GLx+HIMjUopccA/cS/n6n9/hu59wLLOJSiwst/Ol10XwYyKm3qe6NyyPXkEpg
4+iQgZ1GmV+aV4v0x50AXl80QebgDdUiwFrRmiMoj7I7ROEaige6mzYWBV+Wi3Ws
XjqaIj3sFJr7T/+sNd5e6eWsaDHv7UwzNLRRssdHWkQSJa96HCYAt/xRQUKHUvVG
CMUK+bcErHMoojceEqhsxQW3MaTsffmiyqdLJjAr2Q64zlF7LVbLMhbad8bt/xtb
qqm2giydujahUczdWci20yCU2EXVf0ZvHipkFLcfJ1AeoHylf32bAKOegCWccbJc
VMzGmY+pZMFQp11CwcJLUL5MVw0Xt/RJqTBpzdE01ls6g1jI7xIxRlScyTNPqz3e
B+BNLfr1s9CrOw64NhllGo9xIlX/a/Rlm0gl0bbDiDKUMY2fIvNoPe+HzVFAeOlf
h3dHKhBuOB9Azx4Amur9FZ+I6M99j/EF3pI+VxUy1OGinN/SQNNxFW2LCb+wTZ6C
gBTN9ivPhJolccFk+PTonpUuzFFGuP1NlbYFj2BmbAj+gvJqu4FkVPPnQULEt++1
B8p1meVmlBvpArVQJ/ULiZ9t5n/MhOCKsUFU2cGvL0XgQqpO4KUxJyqchjaDG8C5
zBe80dT7XD6tU0Y8mjKjB63H0lEoXSneDinKvguXN4TXFC/38e0ODIoS7snZdTnV
kRDkCJ/p3pZoseeSZR32VXImE/hRYvhBfZlqiryHTMabBRkqhuWwJUfZb9unicEJ
JuE/b1TA0TW6W5Wf8ilZVG+9g388+kPP15C7cBwKtvcnyXEJnOBwdOfBWBCOn6Ar
8gf58G4uOlLVHrxLq1RcrPOgkCa2hCExBWlLW2gD64QI7uKAdMR/apvmDYYBBV+1
NaO0CFa9pGqwJO1N6oGzMYNHkFz4ASsnpq5qMwa41Rv7jkTkXwc6/71hyRvrZkkU
waveBaIdPj72kDj6n8HOHMWNJ0hd3xDw7suYCy/krU98paiIT/RM+rFQy0qhB4w5
V6GFaFINJ0ikTH3R+DOoaTmjKt3CkRhos5tDD8nvDspQGCvqjLzbLgg654RZYm/X
wDeHiERvfPygpPqNWtpceYy44XdofPykF66PyQmvZmXDr+GDnsnKV+Rb/M4nG+z6
1sh7c+6chgwp1qWTfd+YYblQy0A+ZHVR1Y4IL+BlmzGQ5cwavNcPuRluv2R6tZ53
a5dlHa6ivo7MHyTMtlmyA+vy5MRhmcWGKLVcDKAwp+y6nSNirHUdqVZzBDvrrr4/
5RvD5G3XPJmCqp47UIQYzCH+MqmVYjE4oEQpkT1pxPi6CHKlBwrK/ZspJWjllCGp
Gz/3wfYI1JyAde5tR23oBoSquSXr6N/zR1RE0rL1MTfzBDqyZzLQT5u5FedH8rk+
gKQG3T0Pcv2r/RAUo47/2hUQbBGjR6rAZ5IaSI5ODK2XRp9EYSS0H4SwlXWhtW/H
ztT4J+SmxIVYjeYyGR/mnxedUEE8cLC3PvtRPh09fNwFROeAYNEoDVpLzB+edcVY
FOQA1eEgGVX03ThI5/j3COtMlrpxARyhdt06xGorQyeP38uNCi1csW/EMor9DjxX
xDOKdBcPK6b+knNblCOQDt3UQG4EzSGu+ybCqy5gH1qty9SafwZrdrANnixd+dEF
tPMU02QGIy9t+48VGeRUj8rgbj19IWH4kYU3QqfoWLh81+LdSceBhWdS1yQvhurw
EUH34S7kAA86s1C1HNL7tCtrvvNgVE/4uoY9nUo9Z8aDctcELxkTSfAX70ZcOFk+
K0x35xjSz/7h82Kc6iUBn814FNk3HUKycViLhh5md1BPbBX/agKrvsxkk6rLRsbN
Jwfhc/KewmfpAPa4s3LhzObsC8YvwvPrD3SKKYYIefxUfAZ6BxQgeK0f3ZL3wqsl
uaRXOFA+Bm+OeKo2f3BiVhn4/7/0StZz989Q2xhSa2g8bPj9gvivEHrA+uJGC6D4
m3cpIuq/ml31srs8d7+2i/ukuJYqJAQbEQxPtgN28bU3l6NQDI8rO5Oqk/Yy53ZV
jTxcG0cOxIvJMcIOlwQtx7ilWM3gH8zdoiS+KRiM0Nvr4HwlgU9TsSApu20m9a8K
ZV9hdVVkgugVtNeEIOG0giXWVfFhvRKQMZLQr9RVWQy803ElY4JNw9gvuZGzW+mw
qn1Dva1iJmSbCev3VNRfqsMgx8KVMutu3QyAKXjr8CN4vtX10rMOGyI50rUjaoLr
sgBrPrGFDgQGEieyEH4bzGGi0QF5NRvsqDygnU/sFADS4lxM/NIlXg5Ob6gRBrFW
XCaxG/wKtOcQvMOISlbXT3MGwJKmXNmywe2Z9TGFIa61N3TapA/BoRpPVXcgH537
p2DeVxCWvtgAl8yU/3/sf2scBP9DMAdJGyo7uPgKoIaDiAM55ECy6IRmdOrSh6xb
VPI818+b98vDmDjGHpr9sEvIURZA0aFsD5vkfFxVj6WeZm6u5DJOFd4sbrjA+fWc
enA5c5+pGCilnOpS0heT1u0V06ijaTaJgZ9jCvB8AI2W00IgPR9XDkSsLi/H+Xf1
NLsHBmv3y7NR2KrQR7+x9Kwj4MXjlHqfStJaGtpAH9ZYgYm3S0Aivb2Te2b+HS9d
+nu6jb+k8N+faFsAgca1M7Pj8eIuowQCDVTvwaLA/BMel7VZKzJC3qgM/yUPHRSA
cSkai1/79jMIKcphADHgaz7und9Zl7v4LsWGB2ujFlUyawNOAafeKeZ6B/k0L0Vc
Y6+I5R5N6O4hJs35Yi5Ev4n4X5RdxkcU1nZSm1Tmo+1V/wgARR7ZY94pkLgfXzsH
Yyj4ATyr7KpQ/hDgjHaVrtsTs9lEech9FWO/Rf6zTp8MwR2f2krIbjbbw7zpv24C
RakOcxKUEqX5M7RImceD1lUpKu6e7O++cvnDufWdydcJJ8jsBmQoV9G8wgwbsDIi
fJWrXdRXwzYLCoFBd9TfsVRRrzt2DBDWPZmwOTzelCdu7LIHuIXUGa3ySkV6GI2i
wCxnoGV/z2TH6Ahrs6FdBTX8Dun77TSSlvmLi9qVH31fhIbnVeSTYtGXXUTo9Hlg
I3GUU7DbWEct6tOwxfypuk7QkI29G9hvWvDFzfm6hsS4LQA3TzSW1rVi/MqeEDG4
i5YvPn0UQBh3bPV983mDE+WEGZ9yjWAGnjRIZXj4WSavIWk+BrVQeqH808Xwd3Oz
FatOqIdV5pKR66n+TJMcg65M659gnBTY+h1+T1Wy0RxYeTRHqk9A/fV17s4f1ZeK
wcUw9lkDhPcdOFhrrz8TosJzirfTvrEtqMBLxbywu6+SctlSBSmqmnLC/jmS9wPV
s+mcmvnTTR3VL2KJEF5x7OrmDE4O3TPMwRHFnQzmYAJQt/5Nf59Ct2rSs3/lBgdT
0MX9HPXnajt6FxJ7bCvHv8tXVtszbSoKpNIJ2JdPy6fZCXvSmMbNXs+8R1LE+LvN
eUqSjOfXLY4G3Q8vmEYQlbN7onEj6s+NQGLjE858ZSLBDA6NT1C8Lb04yHlx9LEp
uewH+0mKjgJd/EUH04zq90JBxR8q3801XKuKSIIzCXAlcgZk2Mn6otqc4R3Gje9l
EWKAxkxVztwbpRgXLh5nC5awGnNDwoJez/WgmTgFgxB8Q6NGjTeannr2P28F4JgJ
cU2iC/DOSzDTw1d+8JBx7OPcFwZZE7FP+krTSbcDWRgvgFYb8J5qqBOCZwR2AqE4
ZmUg/n7BdH2gM5diCV8wD9n09DeWcvVH4SbT9qGL1tBZC7sIz4ksWpWAarPj92WS
VZEr3mZMnsFPQvaSdBqQk3E4PhICF1g/lTKcLBrHs27w4TfTTcCgdyT06r3Hj1Q1
7PFMX0KrhIESp95sRP8h8Yl0Qg1t//WaJ2rkvMX+zafOJ4tqM7ToZgc6Zlat24uR
y6pwg4WLp+S+orleDuVesfvSYUDOdYX8Xx1P9deP+rKTfMoHFAIS+V2XlenHiqmc
/faKgdGZpOqM4rInmsYWo4ZknmjOtZjz+U8UZ1EdNxbU/6HvEJPxZsWkYho8wRBT
d0ICHCMrlWJwqdOhKT0cYBYdyyWHKAnP0/VA6/GoPH/fSNqNtGUG9r1KrSuXDqK7
RJhKEOoHmYIuS8jE1zR/mdB3AbruWPbt2pwMMHAH2CcFGoOYctrANOIBiz0k+gEV
15Mmyno7pW5O3wpFs3F+rSK+UddXQXGMi5M7AhkMC7XVsPH9pXOOr/JQBtfJynq+
7LksIBtZyadrrY8hcHr0L3iFdDIYJ8qWUqn+E8Un7QWUeiNYxamUvaI7xQIiFvFg
26LOUBV4s/2rpy+zpmXNnQJwUDbQHutV71yuwZzbmC0VkZeMIZ2KwU0wvmxXhXO/
LZafm2bNmBExiUTNLvqZjIR4jrQlsERqd56uEdnRZNRPsL76EIG4sjrUmVm5CE9o
IamUYzYe3PVUFLTqUNVMjf+UfbzslX1jRk6yjBbxtEb/vyd0IqqilPpvRKWuaANI
KrKpq+bOpD3cAuJA6Qk/Zcf1+rWjmehYS/l+ClNKDqmw5Rd1Efjllao7gUYu1MfO
puBK44Mulex1Z3jboeenCTcpC+fXbvkl+9V9eezOkkuSydf2GYNeY++tT/eugz3p
jc8BF3cTDaR/5kuxII1LADVcSHK4aiGRrCKoPN06tuNr+IH5FHcwNH+zgCj8rCN5
LjzVqQaCQd3dHn7ObhPneIYsw7NeAgIuqtyexWdHdn4Z3/RjPSa/KWXNVWg2e02X
aIIf9P358GWwJT2IDG6qTUeDo3qYemuMLxcTmex/yZdmESIaGaCEFdysXTyonWDP
1Isc8o/yKAjYFBCxTIC53dwuE7JnDmACOdVyCgicuroQcBuq/o9hiJIiVpRqwzqf
B8ggrM2EiL1cmauT6aMao5jeKbC6hs7F0WjtDlqmMFccj2/oDwuLC1x21NqpKZ+N
PJywzZ1drIWCsQwMKJWNYDePVRvaybOuOR/+BAAEDKg9WiSTjJLDmEddtrPpxkhq
tFqDrS34GbH2UBQBswGAyjafXape8d1N2fFliSli6dyBjOSStX8fRtfzgVbLeBGD
AXNxuWSmhL+Z4+FqRWNSPiM4AjDxGgCIA9gnGICIFYEEVfvZfBYfku7Ffi0cYA9G
oM56ZFTPTKjT1HGHcAmi77nKyGOkliQkiAOJx6RXXMJ8Bq8QuTPzb4nqIxZrzoNz
6771CzEcmAtCYQIBnJJz5ePs/fvy9F0Vn8BTgv3kvDk8Fh/BuuVD/54GOp6Z+CCE
4HU4esBhQUXi8GduhhhuzKiG2vczj9FV3pP6TcTP/4P2WeCEtT6dPi1aeDnS9vRE
K5b9Ura3jr8OpajaI01cWKc4IXjumeiQ4Ezvt64TXUuh6DL5Lp1onB3t7xRgpFTK
9mfLL2I1eMvxZhSY/H9CbphNcN63j1S9Z9K9gCFJiqEqn1qQ7taMaaLInOW2kW41
AhziW55mn8h3RW73Md4ltkEuWHEqQs3TEUOb+7CVuhmqzGQr56HmwVLAnym+Qf8g
uz4zPrO4VD6H4+J9hq/IOUY1IT1xpngzowNjor0uqHHraegZ2Su4RG/ZkpV8wzBz
CErQm776rsT2tvA1V/33U0MoH6V/vhDS03PH3E6315FPHtPKMEQB2DxOhHwT/O38
yARaHCy5HJCg0hXB/2jPksmacRDejb7XVcxvyDnZ1XA0KlxqY0LBk4XooNysm8pL
ZoY1LH40CmCJOIM4WTSkJJPAAYx+yPnu7yQKWK1fTMJestWVOYXtkxI37F58KpXM
xI2MEJanZ6/ef4i8TyKzH5fQqI3PfFtltA3Za+RwE1gRYzx6XF6NxkBdawjYMFsD
fjUZ6Fd8jSiipX0mc+OZpTRPSVhiyMNNDc3l6z6Uu/kqWClEfi4zzNKS2nGRKoyk
Jm9nQAk1ej4TXV+tnlbSOLletFhhytAVA2I2yWKniP046NEUMJ2Rp02fPUaGYcm6
Zh3aF2lq1NZMJOhR7vICWOEaG7U+E18OAQ8XuuTviYhin4xBTFLAsPD/KMP0yr4m
osBYP7MZ4758z+XKyUItf/X9w0K1Rlz6WieVwQ1okCOkhaGFC3hBgd9v4ulp9Fuo
Zj3UVG0ag42JGR5X56K4YfVrIhqGXJm1e+Gu/HPcLDPx4E3yNj0XtCCpGJV8PlrY
30PWRPqDtBDy7Zagnp1ZRLeoxtlEn+QQGPYHxgiTJBIH1gR0fdkRk3j3Pegu4v+g
CwYZprg1+FYd3Js40TcVhPS+dv40fV6CmzKcuR10Hh8CCNK/wLL/tJByPiVDedHV
67PIyT3Jwp8yl85zoI0UumH3z4416eNAVlDM/d5ptiGA0eokkutEA4cLYlrpC1g1
usJuPr0MUwHpJu3wkwdNygW/O+MRZiL6ptqVxVEVeozpo0bdi1H+bAITj/4y5iB6
XrS7ePsuDA1DuZWj3wBCWtStbdicCHpIzRdxwhn8TeVYgkctzwvoLyXRzckaSV6j
V6H4CZIJzymVavjL4uPx7cS8BoSKn742zKCLQjm499OFVnTMqDMeODwpmHbyrhY1
EFWmeCl51SItbX/Ro7d4Uz13XjafACjiuqkQI7dGU6GCKd9A8ukVWZyXyo71MeA0
4MhVtaYAKLNHERPz09d8I6r/4u386F6jAXPp+hW+f1vqHeVrZCKZ107/GLXKYLe4
e/i0x/t1QjzijVFpShlax1HOVTtFV9ZxLV9go8ZuWqJ7BBiOoNGvsvtQYkuwyysw
dny+KJmyB1tN5+Qqn0n1VMOS1UpW1WNMr7/vcudW66qvKxCiQdrHwMGc2bMab4++
LfvtIuoWatPP4GBSCmPlrWbPcJVQzSi+3aS8ebShmaEM6soykg/0jpYL1oQh2CIr
gCxSCUa8CURywEC6D34HVfNfCgOWrWyzKkl9+VILrZczNBD1SwlH/w0xoDzYPd3A
Nvp1tyC7VVUsNi5Rto1YkhD3tQ/yD3lPVtUJTgvQ/MDH2KpFnafFIo1jvF8nHu7y
/axhq7T4sYlJnz5R4uo1O+DXEd1D3Ue3YjgOBKPI6E4eP7xCQKsQZV1yW1Rseqg/
6e8Jb+SsJgw88WmyqBDwkAkh2XtMWYgSzyw7C7oAhLQknfd0qcLzSEOI7PYC1NAJ
xw7oDDhbUHLwsyBaIBpEh0qjIlg7I2TxNbhJnIwVmpMaQ3PIpMiscyv45VQgTFy8
ayQeUYx5SNIuWHed3LyhzWuRpFY3OnCWzWPijKqQSPr1UnG9JGEIzaHpRv0XVK86
LT0trH+mGdieNl+4X4HdRl/4kPoAK0eaLIW+ynhg26currk7ZrcUs9cHIoR2ZmTk
LMBET6WQNw5lkIZUkegvGL8Oi+hEOH1DCLqG0TQnXOmorOiuHukotv1LEz7ngHgH
2iBcOnRfR5FiE6ctJv50kHH9Edgdf/m2DpgUmoZldCholrHqZWmohAu+LA+/xmBV
Ae0XVYaei0BIogpP478t5mGXE4KetFcgd/J5tXkcUfGfB6I7D6BD2ZA1dFdS2Qbu
e0RfNrNnr3roVJdKG3kJbYsvP67O6CXj1Q93n4HUPIK6SkneZ2Kezclh2+e8Naq2
baeTVhIAR+ZaMK6a0xpAtaT0A2gupQ80t3JClPvclhGe/a9WI7gzX4E40bAEtsIH
YcOshR6hH/gYOQgCu4GdgZ1dYjkg+1UwKZ8lb1FYShcKvFFNUpn976dC6i8c+ZxF
MOcWFr07VYT1jFvl0eAtJkY0POyLtZ1eSNG4/qQ7ud8FWohz9y6+6PxD8YKQYwiM
oEed9v5xCTKShulSO/j3+650IJCSJuLV5eJ81s4hCdNXQ5g0Ahwjk5/Mt7e+dpPk
KTKhBTdsb/YSSg8zz0aHI6H+9pTQftuZ6EDTc0StFvdUzgZRuZR1grPDJRiBSaNF
Mt8zcvj3Vw6EHawrQ1h3ZCYdyYu5QrhAMb0HmaaXrz3d8UJjpqdma2l2q7wOJvHU
ULC71qGGkv0UmWPwq6x2+8kIp6A7rMyt9xCzi9IaOfv4iFsepjBDhs9OE01bG5PC
jmMVpFfPN+VbhE7Eg6HnmrWVtcOQy+XN7WScdOgIaX8656I+MhxV2AQ/pndJNBsW
QUtmvkIzY9mnjMs/wbhyl2Aw2V5GzsSBQTbq2R0CD70LKx8Agxv8LEl18U2N8L47
Nc1ooGFozN6qRojHwQZfAQ/eH/2Nb3EwddgN2XqX43GvmPMfXaxa/mdjq3WItGav
BIzOfnbmrYbmYQUq8cUktZlRawaWwPGqsE+em8c203A/pw0IFw8O54h/0bS7W3hC
c+kSLdJmReEk5Qs3nKzm2DT1gtDTyEp+NQ5nRD4Qfg70H3603NbV8pwT9vdmM2wS
osmeMXhB6hVadwG1D3v+/dGRmC6MBBgy5sun48gHqil1/PSkuqIu098dfKf8ve1v
yZxFrkgk34NXF4dUzd2e1cwk6MzK1egz18gUQqrNPuf05DjrL6wQMucRowhA7gYg
coRyS0zr3/sHZYdOi/YwWTw/qDIQd2v389dPDePSJos0yx7LmA6VJqMsPdd6GkWS
6oH+sI34JPKZ9GIdgPH6Tfygrk6nSrj9jtS39euQFXNG6caUuduXRAVobh0BiLJs
RzRYbhJsEm+ogmAg5pgqFVfWCEnYGA4fGGSzUB2yBaFq9yVpwBRGln0qIKpWW5uI
OPoWGw2NnPjq1Vy15gMvKBi1bUa606ACrTbf9uZ5pWEDCd42waLobnz2XIMni03s
zz/9sHVZ2XNZNIilq05d3bNwUQWiiiMlJdymI8/3xB10e30rQ1RosM3mQD1y9MOP
viXqoizOfsiU1eHXLqXgC15BMi7zA4iSEB4PK6ME8nyNeGmI14bP3TyGeO/m2mBb
gcjTaStXULajvr75Hg6zdhcPtT3KIpP4+TPKC7Pgu6Ht2HU24Zv3ED3ogqqL/6/Z
KtVZoOPp2bGaPqlpZgF2Ytm515teq4BIX69SUyDMVxnybZd28zIVsfqMS6hT0kNA
/90UW1rQTC4rdVrvZj4wwspfZ4WlgvBMJGSoUGXpbUnwbz6RxBlRla3HEyxVLZvh
IvYy1O2lqW6/ija1AK634iwQOLumkB+fnE/EFuZfXfsclqKOB+keG9L6//rW+Nf/
mRhvqElBb6xmt9E/XrtZmbCm319M1clylE5GZCXiOhNg/jkUzufX7CE/uISZ6lQS
ImUy4RnRXevQOkzf+ic4ac9eqWLzpviHX/jRt6eTYZRKJtyRISlXC5IqroWtmh5Z
s2tymt0dz7CeUsz0pM+wpECTSSJ6qqltzk5YQfbz3gRQY7/mCJ1CIuvgwVmwzQXw
qoTABVkANaVvVomHnDfY0Ui/zslAuv30AL68qJ4+qQt9ywpaq0ghd9iz8oolp3zV
5FFKIATa5n77nVw/eDCnFyUCiXa7pFo1j1b27pdiPc5XoHXLYlJgf5+f0B5Vd8Ma
bc7lbWaGIEw3i9hRDPis5S33PVmCnJJYrYZpBKNjxyZS7EA9Ay3Z/3cck84KqBg0
lcbT3rPXWFdeRDNDO9eacLZkHzdpyQ9DRcD6bu4ZE/7y2Q4AfxP48Dc9JhE2uGeV
JDH8AZ0WGczHwM5GvrxvQYSND5RKRX5H2Jz+I/Bx0bet0gmRLrseRFGzbYXcssgE
fTWKtbBKs/qZHr7bD81AYycOM+ze8+qzVgkNE2IW/Rjy67qWn0IzixPkpmHfbNMb
N1dFIg3T86M//k3kkfqUQYJKquoRf0N35xpGcquntgLTy5qtsTcYByGflj+AaDLV
tLEI3gCdpv+95NsDzGlJfRijCNhdOVr9LOoQQ1iVktvoRkeSabnJ6B7qdh8p/gnB
hwFTqwSChhYR6F9SBPsuoBbanTlkhxPSPOjSHFt4TfJynb1b0J9GaSQ7OuDYlF/V
C2LbFSs41yirT6z4sH/so0AJ3FscEUuGc/N0SHdfWHZ3Y+P+b6u0L0lgQIrJG8LK
GoF92hzzuoAVPIYa1cqtHmvRVf3ip40dlGXNJZljFaCk0tH/gySFU/GGTrIbcxaT
aLuaNVqvfNOzsyruKaOlpFlLuCAFOpjG2UmLeJHjdRu8xGqZvQ0qiWsgbNmD3uu+
hhp73M6eDyu431u58kcHdSvs4IcNKFfBUSg/+R04kp5bhI7nrKJ+ivgVgq9UiG43
vHrwsD1Kw9XJkz1We1uSE7/yWE70+6ydOS4TwiAlqQLvD4PjOSMvwrcHmQ+N6eEo
0fMIF/pdXAyM6/l4bs07KmaIk3qQNiP/gBjTk+rK8ik5ye1jhNIUxQE1+Y7pR6OJ
1AmdxEIRh34abM7Yf+86mk9zePQWC5N0m0nI3e1FlRGeziXrpRxXk7CmKvbY4cx3
dKa4q2T7iAA7s1cFDVBSh1sJdMIwEMVzX3v/0plI1rHWBnwHNHINtgS/jKtaLT1u
RnghTsPj+mTplZoE9jh31tI/SiMkKBu3zgHLpvdpuIxsQtPtNpakspZm+cdLkb79
tLfSYSP72OY3USXhczIaRRIAV97O2RBI5B511gdXToedWBUbFiNqyd3Rb2uI1Pkc
3yBuhhwfpre+sGElDR4x7fsgsi3dPtlFDKXVg4zQI7Lyul01nKhWwBVW6DwVjlb7
93WIboLmdbpaTccCvZCeS3/RTOg/nwaIF9avrMA3ps5aL/Z2jp6YobJpcIzqDUBb
KRUAcdxirEhp6dNV1Xzy5SajeE7qG1dsfi7qUsSUERiViJaZYFScOEKLuA9eNtaW
wnH/0zCOIcrhwyEDpA6s6c2x1OhhBQFXzMI68UNbA5Ea2XNcH1HNAh1ycFidy/15
3K6/m7g5foRy68I2z28gu4+VDRpGxU8gX1HPuNNkIDMA/3dASBAt5Ffp9srmbnmA
5JbVKswQ+iZHEpmX4DB4RNQdJtcJFnxS9WygR8NJz/IjbCh57u9TCQITEno2tT2H
rLHKc3uu67fnujsnSKD0lo0cLLDpy2vYIOxLdBkfcwI5DPV1vddKpnrn//SXlYlR
vyBWm5/urKSOJcs2wYXw8zccq/59PgcV0BmZXePE/fbS+G6PQ6DbCRA6Xbo44pC9
vCi+WboacOFhHJskCn8czKHaRCi9EFmDDtJjWorB8MMDS5MNfat1vt3STLDITSRd
EYvO5+cqBbnJ4cfXDNRKnvpA9Bs3jqPHgUuKNd41yrr9Uz2sbdxrcSbIqJGgNT7O
nhaO4SEVOacdoFYcosb1WNPXvXavQmoTT4FJljF1TyojB5l9JU1SIh1QToSIRzf+
B7go9mJlRpKa4tzi8OPioik6xQmaa5NVeI+VUM4RpvfKOBy0Qj3Y95Z0yWyM1USM
3aFpc5ibXk5WRBs+8OL9u233J9QBsQHfqdXJnBjGS+wJ5guYFbPwbN7vGYdjHZ70
Y4aUW5piEQL2yF9eSNiEedkZ2WGUXli7KnBnB5wL0oe6cthdAjmpYl/8lajpYb9E
p5EoyLJ8XgJvqKtWSS1OX0DFtfoaX59eOG+kW2dPTM3as+BN3N8KYHRXCttU96P1
bD7jdclrRJ2IMWRNFARhD6Uc3MbNCii4/PEyVUS7QJjPGY8+3H4iqqhG2EdfB0hb
VMcx1BmXwXk0SxrfwMy51Yvesa+nqIo7INZ0VHtRROcE3p1wh4CVW5QziJfdnchD
wMNIoTYIxu/4gUvno2zNx2cA/ZYe7RHVj3pYo5For91T1+/xIFY5n3kC0SWjm/en
b5MIFqBueorDbOjrafUA/6H+Ni7eahEggCPwiXM7sGVqeps1obdcGGI1FRFZfp35
5dSN54QStcGW9Yt2HBaCXCoJO+qfYjOWZ67ezFxrj4chH4s1ewZo95xD9EzI/7yz
wAbcW6PJ5WftImv1LL9EaK3bU5OXAC6WeHZiSHaL9FcgoA1jrFGNMRcvCy4PIiqD
locjWhqzq+wEsse5nZvUSRWSqVd7qPxtgtqrQI1oERaRd936TRlduEXNNTHxi4gh
GEFOGnFZU8HEJgmjeMr4a4GLfxFFCmwK2hlUKUkN5/Se+VDFNCKBJ0b1V/1PR5g/
4RqaPfw/XeRvFYAwTuQpRN+A648++/dvadqfjbjcHys9/z5zDbEVD7xlcHLdMmkx
INESEV5yr7MHzUJ/8eG0RQLG8RwDWvArC2RWsdwuWAOD1WM7w+R2d2vlaK6rxMEo
jcquCDulhfMg+RCOQOkLSNybemDwPHzV4AHmaE9qNatOeVUZABFjS49fIgYF56kp
1dtnET+sKwcREBkQOk2METg1HQeklMWTHr6AFX2PiKXlrbOJETpCMSqZm9GOI1Px
WE6+35VmysLGqFiaREHseqzec9X400B2n42qvZ1VYaYnloBNuTKBcQWq8BdDeg8b
JdLOfTXA27EsW0iklewrcsbSF5QmOTynHgpIg2Aw3UiCYEUG1uaxnf+Ld1gKS3HP
QwJmZ/X72Rndb63992qCVZRF8IpQdBN5KGfs9YUEkL292OOMuz7u8hG/b8ZbuBfO
dRu9Q/gCuZU1Z90PB5v7pTrBwfrNsGP8qNWHDvvPsFkTzUv9YGR+Cn7UHniDjGoe
EZD3iBmoQYNzMl8D7XSPpeydaTFk/tzq061rlMQxrzDUHgMUpTJwsSudy4KElodc
+SKnmeAqKN8swAl5tOeDaCm0E338E23ef4pftJ/P2/7axazM0YB4LreJm8Rl34Vm
exr9pC2iK+8YtXMHBuhyzyPmaL+Eq78cnPpuOmKrqx6YsAn9RcCIG5v9asB406Aw
gRZfA2I9H7OZHzEm7/uDFVV0saTV2avQpQf+VE4yiJajRgt/71zdOqxNvexcpEN2
/fO94rEMkBK4QhUYhmFf3iK4TX4x82v9NdzNcHlLQnLl/a2PeAXj0dfKybsWK6ui
vCZ9n+Pr5l2a4be2mIh3ngEAFQtP6XoHp+qpxHOdqrduZVUqhyCUhPB2nYVnjgzR
fl+XDMk81KbCtSpS70LbH5f33wxDJMivNl1Wg9FMdSAm8U+Wc0D2C4i039pV91Ti
/lwaSGs+Jq//O0C/h2JsAJINtSSU0K+jrX6B1Ht30k0yQ2XAjUHJbzpYclgoAXXx
6HUIpiIsI4OPDPoyOwCPg/vtdpWHLtslGwHDJWzxTmfk7mabuAfs4tgLq+qhba3y
ocxWbYzm2ttda8smmxtp8X5U9BZwpDDdJfGoqKqJV7OPfoxi9QJDh08bxzb6IC99
beXvkgSDuWvyl0T8gg16x6S0MYQnLIes7yVV47I9yqc0oPen/hw8fZW4WqZ9T5hb
vFa973u/wt5G6EF7EdTXArRl/vNBeKunIDtb6+IOJEUxaSHNo65U3ozK3qAKI+81
RbrCNEh/Bqc0ibzqcZp5nxu6rKDlXvwiw8cgOBC+pOwxa5yKsCQz0fJGWJtYWb4W
0Yb/4sqwIlhFPgq6gpZzHmy09mbvW0fUUXF4WEkcgq+wxwQ3enHDrFN4sG1UD1nf
T8dSCGD42OdJKZkU2AAkcwB8Nn7tWu5CghpaET+Rf+SnqWDqYW6pieYTpKVjtkYe
wEXwTkrcoSHxfJuewolX5+KJolzE98WxS4dPf+lQws7EEwHcGg6Vt9qdG163wg9H
YN5M5IFU2nHM4DW/Hdiu5hsukqFuJKngbbCOyzYrCS5XH25vOqYNDZJGcWJjPIbl
AA6RZONHwiM0BJV1zndsvc84dJf2ChMVhb++2P6cM23A5+synEyJZ+5mFBbf1YVe
V937KsB8kz3/QQcwoc6/zKm7626bQsuI331Y7SV3iE6AFkKmjJZl4wXYjHbOJVQ0
dGkO4V87PqGLQFOBUSWhcJXpe9UP7m8syksvlXm+vyJ0C8mwbAONl3bIO2syqdQ+
wfwi0PhJ7XkSSjcX+O4FP2EDTfzbRTH6xiJBRDNHB7itE2TXchpZhi3qUkz9kqUo
aSlkzlE0n2hU71ppu94C8DQDJYBhEoQhg81x+jD/lcCotV455MRdQF15cKgjLkgg
MxiAsHq5l6UYlM9lfLPeJS5JjoF2hvIXNKcYn8QZPUzwLp8AdKel6Scm+U9/OGc8
ZSsINPj+s2Cw+7/hz77XsMpKlsv8bpnpEatkUxEHfNQ7JSYi/oGNceDI/D574Kxc
e28Hyj/wNKtxblT3odtZSTZ/iQrO4/HSdlPw7MsHdGyURSiba4bssazDU9Tm8gzs
DrJdtnbgzb46UmZNgvDVv8LDZlPVjMJa6ipTbsNrQ7bFgHqsqp+MvKTHVSqBOJId
rtIEllTIHIR69ydmvbbfXe62rNhl0vXlzmjTd9H867gwVh4bgc6oQDvosJ3svlIV
PMyRKJvWsWQfNmO+/h5n8lhE7Do0Z78aWjIIWov28DlzI/7biQcgzuEV9y+WyHJl
dUmwjo07BScBK1QoOVw3nVomkfVCVVaJsskvKlwcygPwdttXdelt4DWhOtV6CgXo
+wZiNEdd1C/MMMUQo26u3hHbkHD0/P7dx7NaplhWluVjaTY5sB625hCvtS6fox/C
L5pNJJ88W+i2BHl5v6j2U+5hBtSpoq6c5NTKoYpFO1DMHUFjBpjxnrqHL2+jO9FV
V4sEIakA2bkml/MdL95YxEmaoqhWyCzvC/hGKDAURHl1GtX0KU41ot6+Q4K0ys7k
taWPVzbXVMcIu1R7m8cSc2DT9Rl6UC+b/n00wkprjWqZLeRP2+SV4nUL41IhKOPG
oplfoZBcV1/ZEOYERY7jq8yoTqf45NvnPG9ZjbaR79RwZ3X44L6QQfcZPUwm14k4
LniSQlyE3txWn0A1TtAsALOSK5mDZiVzLyYr0XTiFKcMaQ8LxBQtlDmST8nBEK4w
1Gj1tWGWUhrQmUe7A3a6Hl50ZeuxhzDrenPqeQbvm48DMTjaB2T0p4eyZMLkdUbd
ChkuLLqqnl/QGgf0av7NKb5kofiDkT7J86+knQKbuy6Pt/pqIx5+clIZX94KpFFk
L0nD9jdnLYHOximQpjnFH0hLeTJUbBbiyp1pFJ5s/UIbrU7RRCa/ZNyhsQbL7OTz
n+Pyy7rVH6LrYUWFnlTP8z7iiS79jOD2N1ZUfyauuUHD/iNobO7ph/yfscBntQ3Q
B0hr1a13C2IlmRGVFYyc/T6EGhFrs3Dc/fNJPMyTallcbuUpZvTO8E/2AQuKsbO6
9KadydvQPfKj3CgZxGHuNGlcDyEpE17fR7HBEWoA0HJVDvP+uD7uZkUv2yOUFF1r
JSMsI9hn+IKXIb5WuXycx8EtSYFkLOipEOwqM5HClAW9O8C8G+Bo5bSUgdejYyKU
X5mCP/1H+48TAQcYV6sk6fk7fZJ/zVoqZs8kNvtEeivHuk0iF6e28gXmIz9tLI4y
1OR7FYz1mcJSl29PJ1asLUBF7LKiwUrulIqBD8//bG6RDLJfLRDZEZynHgT5YQT0
1At4AY7Z2zM4k/3IuJv2YWyYdiC6KSLQ4kK9HtW0Q6AmPQsZPME394pvEnKDKdNe
Ep5+MZs86gxXXTRHA7aLQ2z5TGNb1PETq1d2bh3qaqrEhmtwl3bZaNaiozejxClV
TTkOguvLenR+nl32yrTHkrcnkYi/xM+bMDFqmU5TM0yXfv0ZBaArEJJJ/3c6VJ9M
NR6Ldo1DS9jyqYpxZo+wL53My+kzh19xkElJdInZ1vc9wrbn9P8wCr9dLs+9Cbbj
KKLRt+J6bONsuOVJgb+G8YO5XpxFBQloRCDgPbWuy7Dq34Duy7z8IHFZXfjb6uVt
vILJgqYfE4Rw9vxZ4BYPhxjqJ4EZH4LZpja4yIA77zFM6oPMhXOpWTXKSIGGm0tb
UKUsmqBLKW1KMjOU3W0eip5eKQkffVKmK9n1Dz4K6UuyBssHMswHsFNophovg6Fo
ckBgAd6Qmke6aesQtjtV68Q0ayPzeF2foNcrIqKtKeWc8rr+9LNWc8IiFk0OYlyM
R31O6HnX+FjExEMMJ37opplR0H1+48k4UufvLdc5v9+QTertDsU7wtQ4hcq72Jx1
rd2CkHkN3ZxxY2ExAiCYEV9buDoT595xiUV8Wms/Z6SbJuHdGiffoGmFtaujxCWR
Nu/faTBzpseBLMdXmWY+xtA5cJx0kaB3duQsyXcDCw4cJ4T9RXLUAUKpLpHWkkf4
JR+vtRa7SetcpPlivk0jIsG/GEhPdr/3NKEo8K8EG5rdC+uqcaGMvpmQGzEMSLq6
Wc7FbACqNWk9ZAnlYOtg1LkJ8eg4fDX+QCQUTDA0kFImiXbX25n0rKWtrnX1Y9FU
w1NtigfgqUFT+RQlcES3mBT2XqiExoWsgElcVeKdtxx3mPDMsPZ0o3nFbAIz0oMJ
wrpU4zI3N4uzDVxJurYRbDOuPRDizGX9MlZWDyQK1h06IiLi+7b/y0Jf+01Btkh/
ZPLiWBX21pu3IoZ70LWBoGdir8KcpzGyaFySHshP6f++h0aQ+DOyJR8p1H5szJrr
//WFkSkT8kGjS7BIC9EDxsPLLJwTdFHZ0pP1kfRJvmXNJnEyPfH1ITEitjqf5MpW
cpXKsRSaSs9ZIJE1c3yL+xHTReMzy6Q0P9/WkDHgddjaOSncpMwv30sCxE+n2k/P
sK59NJwi/Bx9M/iUkbP7u/rHRpUFatecrMkCNjhEdo1bAnXB4MG7/bcYUMY6ACPA
HjrqQNpqYT6A8bwUYz7EXFWRccerb+9/BUdGe8JqhOCgewxB83j1eLk1aDhsmnsN
n1p2hEOu2VsrA81AUrWjkoST3eRK5JpEskhMk6FTtb+K91xyYe5C8x1W4nYYhsk5
W6rjgYOIfRDPKSgvBIj/Mo9ny9Nkh/kWfc4qhN16SUlQTsw+Pg01IX8BVjnLg8nR
uDkdFTUK1jjchyYy8Kq1ayx0SQHu5jzYfM4wfZ9oQ89L7CJfdznHlvy0UVD6lH4J
pih/JdxQVKpvliFLV7v/im/KtcRYUwx0YBEx8Rp8WfORxyQsBFCnvYjA7zI/h5h1
1Cr+WTsC6PnS5m0x//u2N6CvvheD8fZx2rpXTHB3/uti9CkJuKDDbv1HTY753NZs
Gg8ed8wnISMvosfvEc69D9SOougQ3jVz/b3RQFNDVPIzYpSSEtBcjXElViIMQRGo
3Xx2UgEIY1lzgJHk8IEzfoEE99PyZXp8/0DP/Cmnu+bFbPAp3DrgMMlqlKdrikW3
dXc2AcBSmpAfRrjMmz1CKCgXAy4Hm3tCijT6aBet6I4KEvUQcYQq835DKtL7exEE
U4lGPfvrRFvJmp6AMM9Ree6y5gZvEAe79cLVqO6caehsRHPx9igBqVEFgEZwCygV
Idx52zZkF70cz0gc/Qswh00YaGHC25dZyosy8+mxC6WDrJozR7NTls6PWGmkO6QC
dPOnEZxEgxBCebRhiT342QJRPlGfOUXkBS9STiSFh3qZc311lmWxpzNEvrAhSTu3
OphscQVlQx1mZ3grjjLmOPrfqGo5YGFu2hIFIKjq45KFD5QzNxrebKjIYskjALxy
ZYFprtE64K9XlxHYBBeWaPqwn8vgATlPkLCJ6VQtjkZH7HMDqE7+OreoX2M3R8QO
WavLPU2gIbQJ91nunrfeAdD5PCzJMnzmn2j4r11iXlw3Ym982GH1QeKaauoCwR3Z
gmYRRTvkMNb2qWPA7UIGh5mLaRZbQ7zlKEx/d0KSqbJhWHPouXzFfaOTOuWNNbyB
OFTZVNaFKeF9FadbfIdyaRbKhX1LUrRapIBP4Cviz8aSqF2/aUt2tgCa9dgc4xn1
bqChEC13/PgnrZwuw20MYD+w1Yfuc+ixzNIQ2hqfTKqDgPPsBg1GRI5nSX0DrT96
e4YNQjL+fWxHRreEXocE0IfauiRVvTQFc+OZq7uAVVPTO7HUgzuZjYoYJy6l1P1K
S/KwA7Rn0Vuw0VIwVkyGrnHyo6ujUjWsv1eJJ800BqjXD1GISs1PD8U0izDIsVnq
h/iPSx9EuDi0UygsKj6dGpaql+q4cUsdJl6Q9eJlKYYpPK3BlF6TQsZgxchc/C7K
z5xdvg4BDP10m2p78jq5MOmlo9AG/yMaJcAPNjw2B6ue4WAAPncDohvjL9k4hqIR
j1T4z29LTSkox941yZvXgXP7w6HZrjyhNrLmrm8RMoIGipb2kMakLeBmVzI+9ywq
KM99UM1oZzCQIstFCvsujPO92YnefmHC1tMyPs2GsSmjaCm1DM4UGqTlLhX/oKlA
T8LnAlXwMOXjOkJ4ZJl6JYR2X7S2SE8+75sswAnXT4ekrkGtaMudO//2x8xwzyLS
AB8RfP4C3IhjC6ftpRBE+7v6T2PAPFxWmkIkpP2VZSUYuTqSereguwOR7Sd+eeRR
QGQvxhjiK8hH6foELcEFsaBMH/BGFCFPpyTnS8kAn8imQP7f42Rdf3xraufXZX4i
PkdWJ2Gvk0OWfc9euq/LEi+BPopUPsfhwutr/vzTVSC4Bjmfn7Qqv0gRsBz+c6H3
vWTd5O0OeLH57IxtwehJhqH6XxnqQZEN5BdsvRFZRPegYZJNVNkCmyjnMznFf9zv
jKoFKtKwECkEuG5wkVPLsv8GbdiGGjCOMc2FipzkVfAgAGbC8o7Mb6zKU9x8pzUh
dituiYKytw9OtwlZT5gETlqIDLZoxf3/7D4NQCbZd70zMggaNwCtNf7VLJ+51u/3
cgDc0Ys1/uNIvywBD6ngzfkB7r5ENyBJmOR/42MCkrgujgTvxpOkleh52nJo3BZp
oD4Gtva5b9I1IDh7Bh1FxaTNRgex7N+25zY/ywPuyfvzPoccdQyX9MnRNqxt/RQN
5Va8e2iuNxRDdMVQC5wV7b4bVzsPqfbapv3welcYnxSUMwOtGfw1zIGjk5H4g4jh
S7WWaiA5EXoiLtmEClZyWHwforDjbaQEoFl5c2pzDZv91v7rWVQcdYxCFxvwJLm5
Dq/+qfIR75IYnPBKZeMVlp+qk9cDBoFo2Bhe5I/Njy3rXnq9Zj+2WXBCeJEZ+XXU
2uLFW7125SYdH1FxXjtr5ZYl6IhX54jT3NccRH2+SgUOkc2/0K8DFfhk71nq2VHr
z5yvTtnOXweE06dMq9Na13LDnIJgYUKVLlkY3K0CX9Gd8gped3liWUqqjTJyggSp
HS5UHQUT2JHAKPq5VN6Px626tXOqXKbCp4I+eUbHWQ8v32t/MaTYaU3ccHi3koAn
kJhXnwmws689nGHB7SsfPJnwvpvsLGu4pcD/R4JrjB7oR5rujNmJA733EDrCVdL5
say8X6YPPGWwoC1d0wJgRN42Qat1NSus2kd5pAqrkSr9JMd043d/Fa0UTQ2GBcjv
qwN1AkR+gfJ1zNLgJ8iFgfJdyzXSbO0Y4muheF90r7+E7joUYpjbP3VpKLI7qfEo
j8qgfYv83subJ0ZQVgZegSROGKxIw/V63C66HULdkwtrSwTRcQE+DXSXSYPer5rK
rgLTDzVc+jjWMuzmYwXHUP96z/tDA4h/cAsbyFlleFk9d28d1caHnOqXQd1p3wpk
Z9Oea44INkhPuHSYP/+nzpUMXp/MzQUeSDk5gEwO+Gojj8J0B0I9nI7Vr7H/up6p
TK/Nyc0KUE3xBI7pJ7a+Ad7ThOxAhk3ToYM27lakrRNA2Zv8hN1dEEBcOg14eWnH
s69cmzcEcxqA3qv3zoEZfRlF9MVDkkikodhbLTE3znVFY4N1MkpYbetSUibwlB0b
MlJZ1btlG3IqckaFR6jO4KDRQHQCrIagZlGhf/g/Aym/VofIaUE7Wg5L+e3VR3Pj
qhOyBVc1vk+a5pocHhE9kiYGbPNIFHk3QuGn+iGrN00v5/sOySJZyVNNsJzrAZsH
N60mJn4QYOVIoFQlVzu/3RZNrnIf9JLj+jmGuMlXW4q27QP87GTU5EjoEA9CQSCw
3Z0l6P6NiwboBi5yvUhjafp0PfRsfKjVgPhmqoSSdiAine/zgVN4z+MrE6mRp6Lx
UbVq90hidL27FmI0X/g7kjcLKWUg2aowACRXB9SycNLHowpo8atuiGFkJRtIS/En
+ez4RoqSedm43C+oV7MQ0sGcAK9LhqyiP1nsfVlCFNTNUP95hRBzOjiODiezjjUL
OHRemlXI+MKhMgosFqTHJSOvW4zezcO/OQJxoxSAm+FM8SEkGYAafJpOo3AHSZ83
1Y1GJOVyxPhaG3vlFriwzgSdNL7eyohGqtG9nQNd0u0pkozt8eH+PujNM194bLRN
oD8Rz17OZdiLTNihlzBIKFr1w8ulydZCpYSSAffOrRJUrYAsLP7V2/CgTvynMr8m
xZIV0NrC5hXex0e4iWu/zsev2GLsVY9pT2curKLbkpRJZAm7J4be//DCtc/1GoEH
mp5n0mfgyfWGMtW27EObl7uXpQAuGnLn41Pj8AqylT4Wvq3tqoprpls3stG0LjxO
06tGWHM469lTgw67CP74qvnHYgiHGQle2oF7Wn4PGldXCJqLWpPGrgbVygnR9Vx9
8E7nI2ZIIwFhOEk8vojXdO6LptfijjGXSCCU1SyV3zZCh9ENx1whpSREYuzyr40y
KcXStsf4PEcWffqJKoOaLRdCklesBnfY6BOVVEHIt4KcWXzyU5IoyWxBvKjj/RPZ
oD7AXoW3xfbz6k0QGqFzDKwWcMOfhOiAySfGGSh8eu6nHFP9UgUSDSAOBLKPtZAW
3gJ75Ww4An+wwTm04UOsaqquq9HPpcv1kLhJv9zf1SkfNoMn99Y1+sXS4y5MHvk2
KoN32VKE61vSc5OzIKV3UHjsvjXT+F7VCvMVaiF+Y3CHntmoCZTv4sT0gDXWhJLj
xnUcYyLmwwExUNRpW4hybmsJ4KKs/4qeqwwSZF/ENautEeS6IRLNVc14tOKzgRSm
0gpnPxvfOqEErwx/eoeTmmvYRh/1Slts51zQC3TOubL9X/lljpWsEWonf1YW9pZG
WCm4J5Gu6gCcJN+xfwBSjnKT7HeR5CWs+fYJdEuspnllnihOs+z3zfWknaTEaZbA
DO2im0b79kcIZMyZosG5JA0NKICmf0i/d9yh8rRRRqn2r8tByb8IfcvK7Dvjiblb
nE2Wj/pIKJo85TsCdSAzY6dAa9tc15DfBHjcOX1i0vPXEm8De1Yk6PfUL9Xz5XGf
F7LUHd9SkvfmG4u+sMPFTsCrgZfMk7iZUfElrIt3/SLU9sV67ZTYPFL9eiHmKHpL
jXTmaFYhgb2G0PJTa13Exb90AKZk1s5474fKTJVugjUT5JZgRVGLDr1DE7rDAKWw
OpX/Tiy4Xfq1HCLCQS/o8Hv1KMbpnBq3gMqtDQ4gi1mollt3e7GnFKa//qL+zeIT
R4whe+5ORIIdg4s9Lz6l2Rti9/jMbpWp47CYuZN4ki4BgVwwwhFOYwj1QUktZ6Rh
Lg7ep0ODEIZ0h9gTEVYsTP1/+QW+lPHqgE5RtsmMfhUaqPOxum7FwMIeVub0gGML
7pglcOYPjlVpAKdw1DFmmHTra+43CIlUdHpU1FuP7j6Hyt6D7iyoi6P6QiUpUiBf
3C4ewX+SORVtOtsXar7RLHQ+iW73tCWwQGolGB+mQ8Ie/uBZIAM9ZAqM+X8Nll86
SLcIAECnK3flmUDWpEXODkxb/IdtrvkjVOCkdWvO0Mlsr1UH3lXlzoAVRh+r0CJc
e4hKjx4CXcE7lwb6z3LqVaHmaNmfuRrx97TDUfqNjgxNqXT8nGNe5Mh9t5GQfEIl
kc/IfJSja8vO3nLs4FgYE1OWx+pbx3L6Y2PAPMiYS1ufdr4CUEofqfg+hGK3v/hR
l7bBR0iSH4wbn/187V2tJfmFcWAydhbhgHp8X8pgykRQdVyrUUo0YCgnxIXLhuVy
lQxfk85O5q+PYAxdaYKRbJwrFzBnVEbDeyuaZNtwET4PtWLV3G2GKC4uivOBGfSO
LshAXKT4qAkuFuCP0iSqB034OOmmU41adRHkMEb2W7NnITGPJur7bdluNiX/16km
niTc3nZ64BV7IZB5H5O6/Fk5yN0Uovbbz2bVWWREO3X27+CTnMlJ6djQrNDjAwYj
OcuvtrjZN22c49BIPaHuDOHyCLMKCHWVQDCV6W+lTH7XfBudukQws0nECqo2P4B9
4QdOviZw+bD4gYzhEJ3HEAtxXN/6kissq61GL7xNpPaxGs0NxXM/XhDehlVm2ixd
Ny+EU3J5PXeVKMNXt9uouSGS+FQrBxd4FUU+qjoF5HGlRCEtEvxeVuT36wM55rnU
b9m5mqAXi0yNKdyH77e48vuz7+E0JQjxrtRLOdaLYFICnDb+TuXdo6xfejhaRdZp
vIsz1SVqwg+K95+tuKGn9qg8zBwqWmlu61Ow2VPBnd1gygOC1xahMl72qDwAULtg
uphlxnX7cAZu7bWooicgeBauRna/tElTA4jCm/Kx9/A5LJ7tTIPHDOqIya/cU9ms
X9qWIEEz7/6XDz8QY9JS9MI2ujfuA3zToeYmv5fvRqzXC7tFo9C3PoOaE1lFS5Jo
VJHeQFo1AqyBGt4I11UB5A9pbtIwWFNsIZJX8eKuSseVSXorc1O57XgcRMA0rZRd
Gm7hLIaxWkeqBz2vt9DpykrdTGTfCOIikg8QGB8ECL4tuffAkNJuO43jB4QJXwRe
V98eb94pt8dTCh8Np0TO0QTTPr1mD7gDDqqaJC9jbGEshIvPUFA7gIFw0GyJ6bGP
Vt4njBOlgAccpzS5LlsVeeBpZG/OK7/GkJThvsNJbSBdmCyh6qgiL8ZxFFNHXlpP
gYWFrzb1AA9GL0l+O7Iltn8JMvOfRI8CCjNMV2QYZ1WHtc/2OHjMH9c0S7Qybtep
k682BPMphonFdxdsSqr7fZ4cKe0ziX3T+pfRENGdQ8qWjEgc+3xurNF6+cMlwN67
tn1Hg8yuv5A0fZx5RhWaPvQQqISuG2SpJI7DZZU5B4+4HuP//AJJ2qIUHdsbcsZk
VrfewZh1YLAjDb12BD9K8POd19Vz0f1VdwZ2IoxhkmuSpbMLYetseM/EagOZtj4h
QRN+eG2V+11UW52clu1DhBRtUjT4egPWjIU+qokl9KJmOoBmThdzBjwtqD33iPmP
9ajysv7jqfC94cc3flYcvXdObvxP2o5xEeoA/SVsOFUNBQqwbR8davYOhulwlwEM
XAPiFVdrVSDmA2fWcUMWg6FER/mb+I7OKU1j0fWMMtPCbvJCAIaHdr6mgj0KTEXL
F3ghGZI3GXCC2wZJ3vpjWPHeXQZe6nDFVflb6Zr0WlE3MGIJDGcryrrhd3K/eyRg
K+AVwGLLqAawtmH9qhK8PQvooNc2b1NSFNQq+GCzZdCn652Vnsl8Mrjn9xVWuqIF
cA5vZ2wGguZ13YZzaB4YCK0ns5dEByyCXdM3x40JH64sAHA1Kk2n4Iy7HvC+1t30
LsDqMBsdzXTwlMyp45Fxxm7N0QFAiLaU0PZZRG7kqH15rNA3/Z35yWhWuegV7c4M
en2543v6VY13bTOPH58xPuYEBjxKLaBb0JRgKsMLRszw6r5DIi796ph4Wh3ZagVH
niMCz/NJYwr2xjbpcPAaOKKTlXAIE3Jgsrr1cRLWPJ8EfLHtCf87k3MNY3qL7OeJ
hblXE0xL48EaZ90ufHeeR5WHwnv0IpuJt3KxS8/kB0UQlvn2it6iKT1FN4gNvIH9
izV1CxPz/kHY7et+/tMc5F8pXhJnPkhloBVwO8FQWSqmfAiE4bZXZH1ukdbkR72y
B1GzxQxys46bc6cNfBMSBkDvR8pqeNibvYiP6llVwSE4ZcisrbyVyDaQ1ym/cr8I
Xd4avfsFEILmQRjgnSyL5PAvd4n5gqa3QiApgMn537aHnjiB4iwwqjAnsiDYal5X
SffzNOOr+jnn40rIej2jqPaxEovHpxF1dBxLK6rXU7SQ/GFwJ1t0ZS3Poftnd+n6
NDbauDW6joFifL7osfxtwYtadAz8EXtTbRpmJjgE6RP/b+s7KgSkTaejqrhubG+L
Ti5n1VreptgXX9JhdC07lope9/ueGxS+bYhoqQs9v4cDp4U9O5HCGoCdek0/+oBF
edBXTpo1IVvMHCXaDKeDY5KvCEtur9wSPE5cHkkAuyetOadTkF0Iqrlm7XMCA8Pq
bzrAEayIwzxIIVW7pTLXgfeF+AZwo6pe8zWUnoc7eIav527zmbdBUAa0equAC7qI
YW8m5ZmsfW/ZOx2LmTRIwaB1wUjSfmtsPa1LSGZUPvIIGw0b3ABOWX6DAM/Mb8g6
4N72Knkr4g1saITa63UWy8WtzIj20eL7/Br+x9gHUApDDaeWQgLM8p9WBwM5KysL
BXvKxF4GC6zAIHFBqsPV6Z7ZIFJjtoWkQreBO2OldZfiBSJsK1en9k4IohdIR9AI
XygoSZ+Bo9UTmkVHXVxB1ZeXWQsT2B5K9YQAgAXLCutgSwjbJgMY7jLn4Kydwky/
OnHC3xCzwhP/SRwu4t3Nk9ms1yxmsvdPSaaHGB8dIiqhkJLEGtZ0zqjd9BqZrMEx
JbVxd7lrEe2PvE88opTycPKt7TZLQ9UleQSC47711l84ZGJIGu74dvB5reYUSE3n
v3H0HWAG7FGxp+zlnHUM4HV1AiiMsoD821YlAU68I45nCsmSIpEijsomXUUv6shG
fMx6cgD3jofvrU9HPxt1En/uoVJf3wXXLWHhWjoD4EH5hZ8m+mPHiotRZqI6AQ/D
egEsfRlad3yZDe6o1UQudgTOYD3psQsEHstUZCXnL9MMZzJ5Zm/ZR+9l8bMCOHDL
HUujXI2gLvWpA6jUxMABqcOVu81b/MCaVt2Ijdt+OdzFOUh3YmYtU6eUH2etvNVX
eofOyxmqYOOVeQ1hkRuq9GeAOdHVmqz1jnD7FELu5ukZP+dNGGJQQL5LTiKukbC8
KtyLunm5dPSpbiNZFaNTBubSfH6agxKit2ylbOkqSqKhXa6yCM4ryczre1QP2IlV
VQT7mYpDFbIh7NfLsYdsZOa8J637MS/y7zKK7DjXt8VN0hYPZHS4Y5KyxzLAGezS
5Mf+77mtf5fS7r3bJ6HDyEio7/qEc9D3XLhZ/dxdOl2RYSpNJzV/H5cGfOpZmxGA
Z/GrOs+/EPxqz/Kz4SWptxjXOAyhF/n+ksBy5Z6WIcq/uKjskf/QvbkuFJA8FeIn
jcVaCQPpYvOlntODotywaCjYlH1Lv9ZjvjZQUZGQvMh5O4U9OpW/uhwnS90VxF93
ms8kR3pQaRFnmrRL7igWqhiZ0u1B/vKysLTU9nhhGYNdfdfl/f+1ktrrgQQ9/ciG
kWAIgzyeIUGcD82uCPKIEhuFmvoUr3P7f6uEYGDx/h9Ik6K0nJL+kGEjCoNEIVw5
qzVRAUckxYjFuIFl82ApnmlOTWeiVf/P9BXz9D81uhzyw3d082u/ufhvif8YW6UP
RxQGqKC59u9jQJirJ+lfV6vkL7MW3hUKRvHCTp1t2RT5RpqRvyGkylCS7XchTcpV
mApfd3LUIRdrFWDiKQsoSY46n/vwjRbij7kWIuwXGfVi7h+QQKhCGY41lYgv0nTP
3McQ6JqeA6YmGGK1roAYyb01qvSy70uonmAQgSaDHiqbUa+/FEyHhyV1WcHyssFr
LU8nR/SjaHWTIJAGLKxiMFQsQWXpiHMay3GkhfD5ADNZ2Uan2ZINBYt7ndFXIVSj
1J3wXpO5cmZT1H6DD31iOnSBGWkU5AQqVrGDZjYTe7X8yjly0zQw3X/AU3cuirpx
UIRpZA2OHVycxtdngHXSxuZIRVQKDSCtqZAQ66c0xsREVnJnqP2o+GGixbM7KIY/
iIrrByB441dEVAJopIuis8kAf2n9B4Ki3eU7DnU6n3uRAh0e+zoEt6swY+XO2dwS
rPsT1i71vki+WFuj+EPtZEYRJhkxHib2rmDlCzY/x3aeyJSYdY0MsEoIwYOhZb2x
zecyETjyM/cdgokCaWvA2ytmhv7tpCx2yUjuheyEl6py6selI3MVGNGnjArRiou4
VtXZaM2yACClKzfZm0k7Y5UR8t0hqUXmG3KVfpmD4KEnVK+nkoFY113goM5P9hCY
IU1DkQLzC22CJZyeTeGSoXYKMGnHhMY01Pld37vXt9C3uiAjQnQXgsA3fqicWBbo
ccWGxGmr3PObL10OXlCZ1gnttQM3SRAg2J2BIHu+rTSf9iZwORpubji2PDgTl+wH
XzAcRIL5ffC/q8rSL+velmqFfRS7GGg47zhYDyC1bb4zlmFy22JFUj3/NuOo83qY
2QUHq5Mk2GJzWezFX4pFfHECopZjnOP/1vyOy2qEnatuKgNFfvztrATzcEuMETTw
VKTBSeIGD47+hlFDtV4K5/Sbro26iMBH7eiTN18KjFGSsBJ5fUY9PpX+Dr+Ib2qh
IwelD0GkZeDf1Qksk3cmQryQIEZqzm1vCsbQrSgEkmVI/pKUY4w+9eovh6ccVM82
ePPQ5NAnXWvDvZDHwcs9fSpB4WM6G+cnxPstIX+5KtND/svg4EhaD2jWb7TCj+CQ
WwZfPDuh5QSg9zA4prMjfgxe7P+2N5DwbmiKx0D3wAcrUuYSTqCMzW2lCa1FBPVz
X6n5vdb6/SWMpcdkwrAESj56F1TJQv8zZh5pPYv4+YVfJqaBVPuFk19eTAMYoQAR
i49oq3IjhFyc+KIaM0iqSf+juCNwGiUITLwR9+gi/2beh5hWy4Y0FbqZagiIkGCt
L92Tz512S/wnKskGerd22rouh++GUk0BuR4iwSG7nFWpmhY5nqn9ZigpdfZtcb07
F0I/FxwRUU8j+F0r+4JjgL17OJX4Wn5yMjD6SylhqXVlp5v3whiNmjkwRxqdwI8N
YGZRet8MoUPGfRJ3qqzODOpKOBPnvSbnhxN5O86OUoVfe8v8aTjqKW8+BCzpYjGy
UiH3qXNS2Tz61n7RrWfDR56IIg9T/qseaobCRVQLXVkFY5AyeYwLFuHWa48AVSUk
t71PnpVhtGpuEFyFIHoy0Ah1y3ZJffl7l10dOjIEMI97IocbNoeiGTc47Z6eADrJ
vvgfuRG2uIzYTrZarLRf6lAXg8nBa7B0ZXIL33ngBmNJW7JwyQs8zZXHaReZsGyp
TrqIwX68fUnMbjA7pH/4rhen8iccLRzsSyr7/DqO+1PuNzDoOno0J6KoQzrtjVtQ
odd06gnYixQcVHPX0TMFyR48parrxc4kI6ylR2wWQl+RWIWs8YONi2dPumvpalJp
NKgaKjG/8odIQzuJyr3uPEhh+M+dv3llSdDfq+9rFYsplJe2iLFlwfScXBAX30yt
munH9OpBdXLSC7wbrW4zwSBmZbjKM2g6EQHVVJ6SV8AREBoxbQVMdEw8RLmCeBM8
y2AAHANPDpGk31TH95PyHJbRUEe2jJU01gXe77elpG5Bn0RKCUs87vg5KavW74Ww
dLBd4VoUi/OUS8FLpkBuex7I/OYsm1bbYPvE17DVnFiLm1Ujk56aj62Uadb8Ajto
z9XD6JIOiMm6TwsbKcU1QnqqPDs4g59zHHqlgN8sIyxJaTR+zvkkEbcQZ68snhh4
3+xm4li6Ud+gwUSgbFsReEXL9PYBQU85h0sXBab9YfaSttpCQtR6zu2V6oEelPPt
VR4vcaniSOXyTXBGkNYgMFRr61uwJoApPHD5KeSfJLQmFSaps/3BwbEiTYPxBdpZ
eNRXzFfgNXvWchssGkznpZd+gaFGtmm3tgEnuLZuZPMFCT9dbrSKYartQR0hskfD
RZXR8X4Pt2qWlrlaPs2A7awJ9TdjRFnx7imfDuqXyUifZy9ByM/s61yzeGoj/0Or
CT0kRUPNjhwNF+l/zkk3gF8Q5StlE0OCrsW2C1XtxzwKqauNBb1SSChJkCA53RJn
35A9IDvEFAOtEZ65p2OWuSiEH4iogh9QXcE27wo59rXEoCfIctSRxdyRDnS1y/U7
CcezRaTm55QZIBkoPoW13ybNPz9e3P+MR0fiqYwOkBNwh2eiIOQbO/wHghmGCr+T
r/CauBeuixnaabeKs2iWRVEqSvA08q5bZ7tulahKFk+TV+q3jF1ZjUPUCfDDGU5a
SXw3KPTQjmlzDBMjDB2zFWW8MLDah9fTqYVLsadGUdRqS7YdtNCohQplInwQkzZX
XEQtXl551sT6jPIByT0v4689+oEz3dTMeIIcCr5xJJWXAsTqnDlnVPPxm0tIGz7s
5cJwiVAsErxcCjachNdXZA5AG7EYr2KxhxlYDebIPA4Y5eo9jyAd6X3fm3/2HvRc
UNzJzgxHECILuSwsy7taL1L8VMlYEXBan4hbVYGEqivRN6aUbiyGIpHpr4BOav8p
z4VTM6B+uESurF0fPwv672uiFAoEB7IErgtPiYhFNxBwkUIAfNiqY+q2Ia+lSCSo
dw3+UwJVZshAN2k7KghsWZ6bxsodIh1nSTQxgGtLHSDb80fFrPezTThnzjGH9wKr
L+Mq+FSK+Wjo7rc0KPz5kW1AylP/oJJUGWbCQMhUEM1G4UbO4pCowXkFuEWj5Nd4
CJUVNLvm3Vgbi186cZYAqcCAeZaUKttiIuBIcRWp4vIWPv2cv95TWKATP+jIbvUV
pqaXzlE6i+oUYKbcI9mHJZAA1yWFKLl1tt6PVXuN3qxZey8ObsVqhgg7AX0J/8o8
WOxmPIs9D5ahtovJkA6s5qZTMdffTb/j9yEppfadeWkC6nKWkKz1z9F9bHVpyvx8
LtJC+m4Dq2iwUxv6Lui5/j6Ovl8GOqYe0IoyYWAhL5vgERe/kw5oKRdM/CMuOezb
ZEvYRi+YM9INdAzg+96u6lEIcGHTDWkSVCbged7owZVEEYCbq8bGOrolqZyD84lA
LO3gd+HcUdy6pCibYGoOyzi/OCx4JO8VWhg80mmCTTCeV92LKAR9NpgNmf3Tvqns
l6Dpu4LCwdhcs45W2JzL1pxK49p7aMMq+BdqDt+WN++2NbOPu9e6b6WWk9BZlNnz
o6a1c7VOOIz/5w83/ASWmcEsAf27FmndlamVgxg8PDC4aj8GFS7a7nfEHd0vyXhz
ChFi6Y5K6y4+GM8un4VlRAg83VXFewqq8P6bBVblDzUGOlJcB4d0vR9BZVKx3grt
QwZTFi1Da7FmqWrRUeNB0hh4BOxIIm5cLGDvFYNkwyNynyaKHElRyUZUPkbf0aFy
2RKygyaZtoMpEFOvDrsvi/N+c2LIK4eGZmZbl+LgzZgxTfUmPWGhYryM4TFMqAgE
46Mm11xiTCW+zLkTD9Jczy3eOYQjWsDjTpMsPCS+89RIKplZLahPkiNGtVLcYwLG
ztsiHXOtQPADkBjauNkq932em0e6TCOD1W1KUd6kpfUGmEYOHQTplQ7nfNBINwRy
ZWiHsygqY5fSu7NoQEc0MeVnpbqInRf2x4h9ic4OyaWq8Ih1XnNWKlkg2YdhbvcC
3bs+ZmZECSR2xVUVTHCLpOePOxj447hoSCYOlGEEeIOmKvOu7+NIP/uIocL7iuzY
1zAvNbg0qyIB0LN77OlHKZVfAufHquOVltdwG0OvpP8FuF2qE3l8ppMScgoZMOHM
lLSuLvSBRNnHzGSAhBWXXUQhtumAbHaNou1k3XUIQ7xWCc+bGIkuJEpQWFxPJDFN
dDA5a1XvP2+ubC50I9qHhuC03zpY0OI0ZAv/0lFZ3OcIuq/PURhKOtxjvM60wBEg
U54K3f1psKctFEPFKOoiXDpv4FXyRSGIChEYH1UTEwTQsYri4sg3oz7Vm51u3Its
X/1F7MYi1+FDcw2GYwGsAKH+Gb+ATRN4XMnXNDYTKeeDCZ0Aum6c9PsEAuTDNKrJ
PE5ZYTNaOFHarpUZNlfmpyBMP43cy+4irsZZHXEBtbTVMsT4tyUdJbdr+iDcnqob
J9qrAkBFJSs+zLCNXiyHbWUvzOWyfLWoVVp8nJj/D8641v6iElgTkz4HGZ8dYe2S
+i/bgEhCEgDhcsYdotCGT6ntQJtZMn055Q2UsJ5eoO5puSZf1RIxN9Xc2pfQYk/y
QjKN3uMeizyYRWoeePeOOytuhL5BWE5hNfVOTQxr6zjUd4Xe7hyrREfvJ3qlqne3
+ASaYi77x0xPNRYNUhzWYxYZlFktWYKvY2ZRri74pa1GdnufbnAUEpr4AUB/CKFa
Eqdoa7tePeZGpykcooPC7sbj8rblsuisLkhBmPWzVc+3Gus7pFDKigmPT+bStSLY
17uf5OVSWTwwz3z7xzCT1jbPWq58rMNfcYthfktqMnix3PhB81M6U8jSY8MCg1mS
gVIQOzjcvOC1J6FJft9n58+3z5ofWlKavCn3DzmBoBDi+vEVYRD+zrRMyMWjw85p
Se2Vd2pOu00Epmlc3+FP2xvfaQ3LH32/vSH8m3QgFzdcIX2/edDYmQWyUQGKQY7Z
u3/Y7K0BNZU/OS+/iBAilGfdLWt+g02nypsDVrgzSZ6jqxTAHY9Q67jZU/tl1IG8
ioDorU+HWMuLzg9q1L+QmnBi6PikLoeNEjrUyHHN9swh6Cg5sp5cz2QpMmbDw5aG
3wzDVzO6DeBU0WiFGhtCTCZhnGRVFCEG/JeOwiSvnQofaA2ery2T/TtdmyybfwYS
06HglbLYdo9rT81cTaVLi7NkJLFnTcKWE488IkUtZbJOl42AW/qcp6/TeneB3mmi
F53Brm/O9r7BUmVdhhtIamL4rTCPYEGn+R3g7tJSymZRTGdWYMJ8TEFXOSqginzN
xl/G56s1DpKDHoorT1Ny5PhMpZSHQpiNKsVM35ijgmdecFKTDLp39IvuEzWvBLZ6
ZrFNLLvCSip7Dj7/1GO5ws0L0Im9yQzO5qen05cPZqcCSyhnKQdnb68G322hrlot
HPafDaA/W1Gg66B9PYCr7cWFVkAim6nJxmMjBfTFEAf0OL2GWr2MayDA7qn+lsyI
4EldEu3OnfMYbPXkVX/dkL1Y/0t7To3m3zh2Hm9DEo+KSw8LvqmOQTAXE6A0HSva
OFnQzSFQLtSshCtMK17LemXCNSrRkobWVm7U3q1LcKGwmPfkQ2e6DoffnxhJrm8z
5FSK71Z6MZmKMgEkdAuTIgsYwC3eXYEoiXX5SNNtKHSEch00A3/Ferz3yxyo6C0V
JCxr/T+3SSxJb8873yYtot9GWz3UM5YwN79YV8+fTBh990J20ActdDSLopmRTke9
rxNsDUTJjtUmNQXpJqNcXcbaxYTzvNH8Cn+Ny68ZnS/pbKb4o+RIhWCsDGaX/1fy
MzN7D9gCWryepniAsfXsVZ3PULQBFUVAag6IlojkVHy30pg0MPSSreq/qX/uhhaQ
5lCNhL1mzt/swZ0XFUdwRfHIYyCRSRjEJu3RLVr2MtDs2MyMHnrXAtqMBwbjqDOB
FgMVlc7MsoTBersUFfU0w3w/zH0O7U2IpzmwDECSnBWgwUZa7S1nckO+c6696Gmj
+KRwU+P5JCu5tF9XT7Ft7nYnJ6q2HIPl7rO77Ux4A7i1xS5Ioh7HX+uN5Tz5iLQZ
jE6rR4hY7snPSVxjPIvzQbXw/1CsOVRPHaTVqlYJt7mCodTjvLPXCFWvHtJkaWbI
veSWf0Nt3IuanEkJ67emaSakwNPTmnvU4wQGhgCJZAFSF/a66cvzuqNceXRQj8iQ
CiwFjgxjkUEPjQYL+rZHIk84QbnWIFAlr/QlVelv7frslcVurhPTmDB94d0g58ky
uPmdX2f68VOUiHirS/T6zjqDkTqyYEx/6XEfCwWBXNq9Q58Tma/W32vamI6aOts+
yt5lRdkQMOmh/urOtrzzuMkScvNIaaxRjzu+Jjxbikdc+gZsUmmdNLowv8HroxHv
2HdvKrE0W6BHR6jery83oQ9pWhu+DGmO7pO7j8G6tWp/d20sVMmsMVlvBeXIaJu0
y+ZZv4EKXsOkdXHWHq5omzbb9+2PBpl4N7HzT8KwW79toywaIBpEOfsks+YsCYfk
zWGiEuaER2h43jyObpop1SeqtgoNbc7oGHMbXpaKMx2FM6TeLDvJVVvotB3wYctm
rMxnokai9mX9cOOAYTvIm6C0/AdNMhQSj6efJVNKeb6qtGiIQDqpJkJ5cjHFedV8
e38G8v6LGB42Q1jfsyax43+Roub3tdmyCvXt0MsDcerxtrV4EY6vw0SxGhtyrLsl
6QyUxuLrd/+/YQLUisKsRGFk6j2LKkdcPtiE8XABLWgX2oQcoxlzBKWycgYtV29C
U1/lKt8hC+TR3esm+oD5rLFQbxKZhsUFbSJB/2NNSVRmPns0qFMALNehCKGObmu+
IMgcW+aJdFyz/u39egBavdhasC9fGIp/275m5qacEzi8c2GnoCa73W1kRulj8DJy
qTB8/XMohl8fH0DG/effIqS4Ghv6weEct+6/uTkIiMNFm3bCMTHo6PzrvdqEX2r+
e5PMM4Fkpk4/rLVbGsUAzQoJGVq/AEbsrpoxjAx8UGWFtPjAPT4pExSbCKXXRJhP
5i5NY6x+ZkDXE2RZ303QPr4nKXeM5IPX7MB7mhwqa5t6CiuukHobTvEEqjfJLNcJ
il5dwGBClUNqYGszAvW8q68t8Bb/1IkETHygYyQRq7eiVe2WJMdWQqQbg3kIflCQ
jbur3lh6WogHZrJQ5X/EQSvjzpVvUcoLTPhTDfyuR7KiQCqF20geI/57IJ4l7uh2
5uzZwsKCoc1nQJT2Xg0kSIGklVPGrAcCFM/Z5tId/8iYjidLIAfZtZ+DZs860ets
P9eSOiMTwKSeGl9V8NzvaSODDqS6V8gJZfy7zuoPHHukwS8eqAsM1FaCkd9mOBje
wA+JUWIPn7AomlOfjoHk8azVZ1R29TkLsGvWLTvUNZY3i8XCmIOVXGO4oucXOILK
Qn2nJX5RaQTdwlOBxKN/PfuRp8eezofooxyBCFjwF1qrZZgTXMOUD4tHbU1v9oZs
J+KDDptiuZQLPq+XtOnQujQf5OHQLhUdyzZQiNuMTE5iLAgDWpm8/TubchaBaq0D
azJvlTmUD3PX+mrem6Kx6tQbRS81YMYdPIeC8mfTa/kqd6HJ+VgO2jIVG+N+Y3Ic
gra4WPcALSMs8M31yPmmmeqhkx+Pk9VSRw2P5fzMFtbOtQItwjxwcCmNqHSaVOqh
ZIv3p06BgKM2DoyZ79PYzuDeL+I9wUI28ld+zcrk8eGC1k+FZEVzHFrkf5+uaPkq
vW1/SVUz32pm3VG6ZuFYDcd43v+SfTLr1+5xOVCIcJIWSI7RI7ccjDLXeBae0w54
VIULip8+gANvQfOrYL2z77ZPdysAga7sUkGTlnkh1LZ89S68sVCzDjVuZzzJgsPf
lG0psj7KNhgVzgRF3txLJ4GBnMDW9xdM9GnCF9yOEwXpvBrpmcYOvwIPGS908Kp+
Fce/pFeNsMaT4n2/xydsTurH6T5iUmDLXjbS0DY+uRYBytSwxsCM/zjfJ7fjwt2o
dKgj59Ad3CX3S3Ps2Jr/gD6BvLYM+jBiRql4m65ELO37Qoh3UvchrV4PtDBeQifL
oB/6bAsfosW82/FldFVWX6WoVsTbvtLSsqwlrDITp5NmIjbf3SU/MvVinJSKJxPV
ITZDP0GQNtpDSr6oF2haTeHYvvT0kf/R1rx1cIgLTrY/BsbBuHSe/HpyoxTViks6
C8dOhWLbrhjlokGDbP6y0ys0kCp2kdk1dl4G5jHaO1CYSlFA6hewrT78lIA0Yb3P
4lGvt9h0MTf62LfdegnjHYYNhXVECzFvi3cdOgD7h8+9k9HDAPQaUATUvg/fYlrJ
yOTeDRqW01KQ/jT411EDOVE+MBPFWa0iJK2FQM2mSkwI2zZKDO4+Q7ge4+uS/orI
uKgeBssvHzV3QWBUZhB8NlShbjXum2xyo/dX9BvBQNjjm3OmXF61VYd1tiAvvkKH
ifnCN8LXUTeEw3PPBmLF83tCfZkLwmP6K/apaVO6+RCjbRze5fi6+CNRpKwWQrO8
PDqoHxgKfTQApkXcxcIP0iKMFyvDNyKoAg/JXQ4Ok++Xy6jIyMGpdq/mZWA1BOsd
6yLn+U+uXyb0iDWxHcAQ58FBcprqimVL8riO5A7Am/v+Ins8f7I7UUeUJqkGnt3g
IQbbWtn5o66v/iLTcCgSXH4ZybAlMCOVjEDotdFOkXmxx/7AOSwHwcHHKQLxeW80
2sbO4dbYbc0N9YLLQk+gDGj0yaonAPV1Govi4i4zy54Cy9b1KZZTu45mdWPAZtgv
LcnXNaTmZNK/C9h7fg7gbiW+LN1gEzMd6k4PjPhUjah51+IdcJ5vDeu2wP5h2cm8
frBQY0VHs5ArBpLuSpNOy6ImFaM2zSt4xY4cUPG7sW2NRG5D0E26yA6PF64dDZR/
3g3Wd36l4ETgxw87NezK3+R3hegXzpuQLFnoCS4y2TtDDD9xm5Gw7VrGCJajCpAv
vSgDUwgDd2JKTuf0wSoAVKPSNe4/7bsNTHLOLmiQio3FvA4AmFlXOZC72KmaKDwZ
V0Kpia8dm+boQFHI73F14T7S8rjmCdtfZCqifnpODYJvQEZXlD2r7SCsRtXskK3J
CuYflcE0XCrYCFTyqH0cx77LMr53OAgGZ/+DHYmHBxu8l7qYxjiDxLIgE7aKBYz+
bwGaN+bg4s4az14yKj/HeE65wXyBair8VumMYc4oimJeDN/GaaGOlWik8fj4qF+9
mEF1l7qYy8N9ISHBpGSMxooN5IKsW3j8q5WiViusCmH3pR8krW4JXMCuuHmU56J2
oz8hYgamb9C6hdkZ8bamG72KDPwzGZk+munNfEG7OVI/1UNCRJVsqwBS1m+Cs21X
7Nw8lS2aTVuaWFSw6TATncbK2Tp+ltOwEh1/FLP8KQUVLFvxzgZZfZe4fbTIEXpu
By9ljd9ZZMVP61BX78XGZX34NQWpCpbmhHOj125z16w4qY6kHAnLA4QJJtTzr7mh
v/kdDHF2Tl27+LcfwE1OFUdcpWwt3F1PkhNUEBTh0Q3fOSe8OQhzQE3klGNq3DlV
/O5YUHSmCCrNnFuBlW4UC1DEFdqiw/2YQYv3tx2S88rOl9ENlW5HZYS2vxbzOkdh
vrgmC6rbOTzfKmOSU5DM3nXiu7nAJR+1tvNsVv8/fkcBDJetvH1gohrYbTOMTzL/
iUHi+aFjTonBfwzF1s7Y8hz5gmaSC8+LcYE5syOqTsXvCd5y1+V4IS3jZZVIf6D+
VwkBB0cssklMbPixqT22FNL8wh9bUAuZOf5+71oi876JjtytRCckZLiEIjMu9b0r
Y8FhAPHK7dj+DTixSC7AZ4D/2nXmd4ZykFhJE5aoJND7UlPOw0KPCEkMcI3RD5fG
QUMYIXTZ3KmXTufr9cfzl1Iz8SSqb57t5PjZPLj4p2rfZA3bA+spkqPwglhMMpeN
x5DxYJsRDd/WP5+FkeCQrVgV/Q5U+BhZgUYT8m07TOHz6l8NJrzJ8G4T0pDoTobp
LV26SihB1M1NHOA4iuuUggRl9OmwER+YUiQOA1Ba8A5PMFN9U9jeiCNthHOpY9Na
b+ruNp43PUSnhaju380jRUyFleEa6+G2THFp1VjTzB2SIs12wlxxNV4XlPZgdVun
EsV4QYfcJoMBhWQx9PlxTd0ltjFd3q/dU+kbbmSCofkC9lQNKRmrBE4SRB20+rTj
4+A8hL2YKPFh6+hUnAu4Mad8dAaPREz7JMRZMiA89tJyluHvDVDDd2YU8ZYYPHVs
HraPRzbI5LhIQwRzwlmByHNUVw+4ANPSmfykxRIa7YX9+ZAmUEeiWX/YDTZltmV5
uCy6p5NgUcMdX64Njs7LkMNtC/MXdxILXoYAHfwM5ETY/VvPmdsJnsSeOZR78u9O
l+2jVDyImfpuEtPDiUdRrAMPh7uV/hnpW2i+zsHjtEowaS4Ayd/c57m5hrgfwg37
84Cg3gLhrXC2VdYCFRJbz/dNQ/B6cUh8/zqSUfzszuikmg3ynq6W1xseehfZ1abN
Q7kYdmlcB2fzEAC0/VqCqxjfvzrnwcCko2mRynklJ0ZiJduatOne+U3r78rvP9IL
ymeyX9qNmokaJB5SGxuPmWU+0PBdA1wn0rqR1qnomW5pqhPEKDo4woXY8SuOjfi4
6iV7QP5CxfNJKx2zQtlqx3gYZ8NFHsudiJbsKNXJ3JceP8GE8hmsCwmdZkY+7e9t
2O8RiUY+yVsA4TYVjjN7HhAeG43ZpvhrapNOYQx9aXe9htgBfC6UQY6sfAxlyCa/
fxb/zsWDL/7Fcem6tlGZspPwKjVN9OE2KJ8SHBeRIEHZhGVsYmYy3JAyl9Dxyxvu
+vHG46FaPGgoFiEUgUduvz83i+NZvqleOQJBxDKJYleZcredMZLydf49TtNQe4aH
ygB54plsJMSOg132wKCL3lMr9HIa+WGdYBoL29gxXGV36WzvVXcjjyfUVIn52tBj
m4PGnAYsrcpRKBib+QW96KL79MmVCI85m1nL87BH0SgiF29aGvB9/W+kUs6HmuMI
Uym6dvtxkEUN2YdUUDdifFIYzINn/CPUqr6XfWWc/VyaRh/7dFyxzX/f1iCFe7U/
yQaMF6jlVD5lj+Usm0yOikte2mlGhHamMD/1KmrBjay0s9CQ5TuXLNl2Xz0oPrIk
0n05tFbHTEWC82EYynV5Rh7dCk+iNA5TzHDHAHtpFarZQSo3VjECb/MbxBMGtzWf
+Tzm54A0U05KlW/FwtIoe2JxW0j3JgQABZQtlV1uLbmSrzLuqeDadwuMColM4LNx
vzGfMYFwPXfCH/RhUXTbFCbH+CC7mO5XDtQo9eKTPvwiGru7VQ3vdYk5ENBIvb9s
3Y6xuVKk3koyb8DmIEtJvRF5pLMrF7D27H5owh17Uoc9c7SDWdaL8Cws918MpC15
u8D7C7dPD+CNHlJVxeaF2JkMoon1aPpLmWOA9kM+NPzDOap1S6kI+mvC0xCxGW7y
kGZLVKBfgSs3Y+FymH+2ulTvx4VTTwHZslIuqlkTlffZ7P5dd90IzIYdT/XRnFh5
ZU/GOacd0YroNND8PPNpNkLIrZfbF7ZMmcf0bUyiFT9B7lmFUPB+Nx8dl7TnVHt7
DA9KBdxW1jQbv7aTQrjnLbkTRF9UmM3qbPdUKFWpxbYR8lxc0wtri5efMB27hu/o
e28g7nNMn72k5nNeMAqBUKD9fn/fllcUFqPm9NnqlW+1ScyGNsmCMbV5OMuy+0jS
C1kPfED/QoLAEnA3GR4YDhbuqtDPsPX3EiB7FakQVWS7PMBTG8+ZzciVZEGLUiFG
zOg+1prjUnyZNXAQ15its749PauzVYl6zWhJjb8+66uVSiCugHN8uZxEioKPiZfn
Nmcpivfilkuqdc0f17KfYDhcZ+lK3LoHyp4Nv5i4SpvkxTxZ7TfGJ/2iDVsLuS4h
6XQRmXu6ITiY3ACwI3G3HJ4+zIO+upjhoq2Jqa/xb5K/40GLZUM6O3+tfncpHEsH
T7blftY9wP4DoiQj7Ezp0W3cfk54z9wfrhgAbKPSH9FraP6qo5SlVI8te/ANVbC5
KdOGzLWxAqC0ntePaqSDq+vHL7n2JY/6RZgyH7ajeWBfPBo8QX9rXteI3NY0toez
sn08fFl45wLS1uE+6z7NxmNFMgSSG5hlFQjY+dhYJDaPyN7/vckq7AP7dOwMRLjZ
B1GHhoTvpI+WrioTKw+nkxPLXKcB135pa+ff/Bw7XC6t3vh5kPE48zktyHqVfHKH
UXSSNTxYAFMieFRDZoZWA5aoStmljzX5QgcPpqzpzLyFCS0L1syHf9mRiJxOFrQ1
aPunm0qjkDd2GIXkRSj2/1XHlmfkuWc2xzC5bE2OmKjSOB4pdIe1/HpQWFWe2Sx2
ajMLgE2NwRTzPJ8vYeAqNiPwqPMzVlSWs1EVAa0fjDgEmadNwXSwjuw59y7Xd+E+
AwyeSpdQSG7I5tnrgRwxZTL5Ny5noPBK6gfr+7gqeGbBrW6q25P5KONeunYzBZmS
csTFpqlbVZt2NQw4RGuf1Jk54PPIZ2syaNd2o+FcLagc1ulXeU1eAtsdAEYl4Kle
p8u5sB7sETRrovRyvnsxZkHm2OcmI5eN7JTleicKWFUTZOBT44wHIa/s/nB6qR7Z
N7CyJ9EkBGHm/7V9dNeU9Fjeqkv8pnAC0DTKoNvW0gvlzAvpkuJSCPW8xqDZ591f
LPH9XBc8btFrRrBxQWU0RDSsJApHd2v6VKs1bM8El0JTwIbiMqgAkqHMMU0qfJ2c
QerbM6UmKRINzeqZoIXt6T76yZWxNNcatmf2p0tM1K0mMaCNH+TvUaENr2SWhjDU
6/xlYY6eZsYsyEQrTfy/hfN2TaQaCsBKJ33zztgfnoY0iuTQAtgsUgrIOMvYs51f
q2W8WwihB0lmm1i/k/tnI0VLoNVwfFI0X7+B3tSrQK8tx1+rx+K+6rCqPZgO7176
gs12gZPip7uA0IAzG4BsoUjJEkGSXkPcISuiZoJE1kd6o5isYsq5MFztxRbAkk1P
LsJ/EZf2Cb1tm8tfB0pA/DVAJaUTvT+GFfL5SRPynaOcq5CqyhLkPt39dVqE7k5i
w9Knh1rU21mb8ySCv3nDivQGvZ7wlTzBwv8I3BYk3crxy1MGxv94HrG4rFJg1GGs
E+Zl5HblNp7aBpkOiFMnYzHAOnUuuwGBSX9NBy0YQZtc8OK5AMX+dWfljWH1h+eQ
svtpToSdeE4bWHyBp11h96ch4AcSjVIzRiLWYZ4mMEiqVq4/Cq6SYvWDMzasZWYQ
T9t1w+vcb0ohfz4jSKRWnuVf0uF/YRtOlk0Htyy7GBWW92GqRU015wYbxE9VIP0k
wXwaSvzfUdUEk5dmlMe55WzQIddyJ7xc/HbUZX1uiB3l2wNeeC1EQwSLA+JIlfNU
/NXkuCdrGWbHBUQuvHLldXPKwxx5iMqZVFxgI0cMakUGZMDNVUxBrCo1WnCOuJ9H
Wy8rMraYC2/iWxMg6Xy4Q3rXGX69eDgyFuNc1e/o09OXoe0ameLDan796g52eetj
zwZ2hYVQpWUrTG2f7AJdpft0QQH2ljYChCYUtMUrIO+ZkBwq/YaODHSwKNGWb+9X
JpeUnRDn9G7SwYKkCavSbzy0uUHVz9DGMBWM1iTcYOmyC1V3tEUggMzptM8viRXJ
+5FibaVv62PO/QUl2oBWqsyzAEUKQ6TMN6rWHnfzxMgUD2KVB+5casYaSH1cX5ON
hH5rZQCzeZzpHBsV4RFZTGxfBUaYPSIXvmfMOPyA7YF1X7HtYNx6h0NJRcfOeC8M
svD3zs9BeVJ0AFYgnP3/Og9brFLLKCueVo2x7N4G6E7M9s2b2ZX2czs8WhCGDEbO
Xg7p3luKuHz79IxkGzduppJfY2hCHU/pfOG3Nguw1PH+CgnV6CpN9pKzJiP+R5uH
dUP/OWcecGjyJDT+6qO5XRGUBp1RISL2jw8U+8ZmQEi2MxnwEg+L6pwImtFSN1yY
mqYMcueRKS9s9oPq/Nt9NL9/gitYr26yBslkhhE9kkktQEWzeC15wlS4qSUle3OH
qpK9LGUB95qScDCMnPMGkG5mz0/UAqMMa9h6kIf8bfHT+fqLqmrUb2n/94Ze22JC
3/DiYKK28hfZtrYWWe0npM7RDJpmZM8HBXLoozI+WKfZlNiy8143Db/JACM+tn/q
47zfmsQml/7BTchbjy4ZPFqysCIz2pwkDFGn1StTt4AxXQKmdqT3hB2zhD9WTX/j
albwQPLUYQp8BUmvrz4LkDoCSptk7tofgXTiS6l4wsCG35cmVUBahipJaa0Dhgiw
BAeoo83QUjkNnUu/8KfVfKRiQzEMiX1DibcylryB/QUQhC5d6MhqkoYK34TmUvmJ
l0STTBst3kbyNpT9EaefznYDhpe4CQ1NSZCnGFEqumN0Iv0xfGZhKCoWWFGidc9x
YHWvrsuD35wtBU6bYQl/hXAMFqUUDtSmUzitiEnowg1OZCS1G8sSIXTYreTQ2WKM
LDQXwaijthxpijthdGJsgAouHHA9FXMkchMCri3RcMxVpOjGXSyFanFEFxu6R0tc
2h8avp8s/57arCuVQg17EY8HpjMD22pSQV6aJ1suzaSbP3aQ/oRYhX8kgtl09guA
re6q57/VzyimiXluQOI8r8UnBXe38jvuoxyRhPaWwkWf2a2GAvTeT2n7klbafgk7
AKnsfIzpz9+riabGRfkgtjJGvaAgAyJt8Yjuaa5BOdATfb4vH0ff4EnacraYLvaz
fEBywBULVp6C1tCXefY0d8yVP+bPBDJf6z3u8za//oniVlepbaKOEwKCG0afn4Ee
JUik0OjRRnfBNanOLtH3xTJg4voPt30nywvKeTkHmFNwMD9RojTdMT2NoBUo0pKI
IaUEkXizfDb35cS3tYQmbj2/BzGVZs1YndeeHgu5yL3EBIrE8AJsX0Ajmmb+1yqk
ljxDzHH8rwETgw3EafQ4scyYMUfTSczLMEL70dHy7dZrzAVlor5ptbzNFCLA3C12
MnF0w9yAuDV4rIPAFOyw83hflRIwBNtu3bI+rIyNOYMqfZnh87QGAbWPoZCv/IN+
PhxhOXr/SaK+CrVstj8hhQ75+uKmYZgmVCC7wRnj7qrQlSN3KouGHaXL7lfTchMr
SS9/Fw/cwW2aPzIPJkwfFw2d9dKSdCPlI30TkikIQlZb8Jm4KP+n243Cz7Fc/wAt
GqhBkb2cdv70QKlyGyWxeDn233w77p2vsGyRI0A+1aLYFUAPi7Q7K7j98liL792M
x8SaixoWW+yWg31gsx/Uep7SMERSJrceJct+KaOiJ5aHuvWHeQ2Laks2yBNstCun
qtwcpoBrLSDx7totEr0Gkb/hqYbI+6kmHQDENLypIFZttFEXQUG/HKvL9kJL4LNL
kPa/pW9v5tnWjHZKSrdMVDaELVJHNROwBPv6uDNg60ZASImX8z5VHRIZRH8XEBr5
EPjGLPYHZXwfgVydnPuvyBqTK/u186frkSurAWRL60KYDT9BBwlIg21zZbEDHHHS
NgGjjMRciTtvWrXc1QehQZ9Xh/2SjPA+wACucB7iFRaxq6T4s1/fObX3K6kLIrcx
7H6pK5Pv+inIFo2AFHeOezRaC6FTO2H9Wirg+pJWePW7v4u6a9lmH70wHCnSluvh
6wfTmbtffZIgWHgneFL821G4HnK/4f5KlvmbvK/JD7VDni6fIf8xo0HfK7nJ0GKO
HxzHIrqm2WKbvDbeBqWUrhvv2G+ODimJkvKj/hFG04OcIHea9qkKFsRD76KcvbuI
nCtN//lWYMph/k2ld4TyjBF6kGw61GZBI4yV/7/nZ+Ajesw7LA96CaSLQJ9Hozdk
XdEWaTAQqgc5tnFU77xmP00Qlqe8WbdrVQoyOhYxcNV/Cejz2ogozvX609QL673P
UIWWTMnw/2mYAUx0Jd6PYE/BEQ3wie2rhAlVCGdFq5b266dH05J9zMTx443lvMkD
kS0aIkA3R7y52iQ7YrzOfjKS6sKEgQjs37nOh3oVta9aVxsUAQIBIZmQVrcyVPww
4qjzFEX6aZB4GPFcnOh9RCLnI8Wyp8pr1Rm9RB7O0A5e72+Xb+hTbvO1yTBcoZyB
tC2OYuHgn5uQR1kWI+sFdj7dkvXt1e0lkoMw8JvNqqryegDqMDcyUI6sCP/ux38c
mMFdRs/EeLjgB1yNaCaavtlX9ORMXGHULNOsFXps3TBl6gim952C3KskeYp09ThD
2vtGRIrFrUL5MJRRAgpFXAnJXIBeTJZJwS8ki0mmUlvdtoxwnA8FYCakl+RpTkjh
l6Nu8650tStWrtYO6Wk2x+5Ys45cmUhx49TLBotepHVkacIw3+Okq3M12qGnhqQ3
b2UyoOs149TwYZooqet61ZEiBp9XE2EA1nUCyl8M5OeZCTtRttJrOTxzFrPqZbK7
X8zg7fomRnQUjlV6sCib+Dayy/vAhmbFkzR3uGpvq+/cjhNT8E26tMh2mFs9Qyh8
MuBYw/gODqt+O3q6Gs69MKMLLLwE5V6PpH16/1WGSoeCJj4Bxmd8DFjdmmhSZF9d
0ij2aL8ssCL0k3OfS+coQ1mGD9Yd2S5rf8LmND2+Yx1xLB+lMw1iRWJ2J8cLyx57
IQR5z9Pp1qmSidy5i1riS9szIt96KSZBAn5IK7jgz6XYES3oLxepuMjiaguYvQRQ
iqBE1ZY+aOoT16iuWPiMkSFCA4rEdTQ9NlUg2PTMJNIFIsod3lqX0kNi/l0zaJhG
7vSzgafGhka+1iLuvP9ORt7NWF9RiWp3G0co9PRnAZbUOdcfEsLZOdiBCcAh4JDT
7wSQ9CnaL/JBurdoWpTVg6ygsw9mrUzU3g6dglR8R9NGWWwMxLPL4lu57tZVdPye
NkA5sRSOIdva+0L2emb3rxjFzhUCcVBgni4pjzN6S72ehA+NuQZooQ2416ZCefy3
HDQaltoCVJBSpq2o55gVqs2nxyjoJZ6AmJyPktWJQtlMWQ3Rv6FIkbfDk1YTcmrS
Pezqs0JGgUfvvjb8skyBbaetRkw/jqehA+84DaLjizASmwGoNkFEkh0lhVkOAN1I
SSl27/P4MQBfd1WvcinBgSK2EV01eqmogrUvEGXO4P6X90gTzSaKeTsvBdXiifEJ
5LCEpwCYUwICpBtFv8mdpJggGK8yIq5FBGdGpgXCGiBSzkpjYk7X0SUH6/9IUlBK
VtEbm2+oNTizWUcsL04a2GuiXImNBHRT+sIuxpie+/o4mVQf7l5Tmkl2FSOVeXJS
M3ke/ZA7tvIQ3Cu388H6nIAscoioOqXrr9ahjl9CZIOFeDKjsca5XXBecVfApDvK
QukbftlwkPN4dnUbDy3FUVEOjn0Uv3peQpBhhOnoIVIkTMb56E4OhBhQhAJJXAM8
FeBhAcLDaSy766CCFJeI7IOzHbBuuYGVmqOpqq0WVahWivmu/qqIYC7XzT7XQTUm
qTTyLzY4l44tYU5soJv+7zBK4fWPKPwxRGGOq9BBFp4yY8nIeKYIBl7yIYnT+yS9
xHIFtQ1H9zGuEiXF5dwP4ZU1bijMiew/DwjB/46Jv09njOSosP5bBimZdUT0HILY
VDL8WR3Fwb+0NYRXlt6YWXoDkrpaPXQJN+b4hVdZgi7Rv/CWgw1xRyQhpX7CroYl
B/8bXvFhDFXXwc2dCBxfKvkWYUJo1Sl2unUbPSW7K3iHWnwSOiZ97ymoLO0trEor
hcShZW5ZxdtHBSjPqqbZ6r5aHOs9dF+kXGJUqlKCiY2k5mS6r8l0DBGMGU/YtV3P
hDvNh/4iix5RI5w8nB54ZujbSIxwaL0MyBLYK2539NlPJrqA3SMhxcqi0Kn7Jz+H
oFHaSrFbeGqSt53HyJ1QEg+RJrQ45sEcZhyOLOctoPT+lNUjsV+qiCOQeiGcwKcq
KUvKgdChKAN03yqkBxhinsjumjadIIQFjMZNNZxKrU9G0moOPEqa23TVyqzGRFRa
q0E7FIBuHYY+AGyl5r5Zi20dKQ3zTOGjaw6zt/QlDw9K0013zftlFomhG15ZBUzL
nOGrZpw0TWLO/3vWCQ1H1CY+FqscZqw630S20Olr84eSO88XSD+RsoQ4j+KnXovB
+iNVk6IHbiqLjXYXxJBALKESVyXOV2M7E1kMAdKHrxKo9ZGVLc16PYmRnHwnrjnx
vU+/mx2nAmVgMCzP84HbMGSSKlO92xYd1/YtDQr058ObJ7+5gGWDe6ZIF6DBEE+K
VKTHMd8mQ6RynCsNwYAmjuoj9yr0d+lIF06LDCthyi99iUV1HFBTPQzaO49GVbpY
NYbUt55ekRUBfwG9gCu/Jux6X39RUdANgxW9NESkL+CnUFv+diT96E8bPRmZ28Oc
HGqg8jOOssu8zYaqft8d2R5GGhfmc1CRyyKmCHZMsFfUnWvUHnIsEbVYNxDYN4ec
qe35W89QnPXNDYb9wQd5mxw+wpthhUcTIzpinNsomthMJm2WWhiRfBfMjp+Y77WS
+c++F4Zb7qwDxOGJy1qMtM03MtP5s7PAZcOd0RWx8mqC1vvDxa2bnJNoqpb41AOX
/20g2FGM0q0bP6OhQTlybsAS1ws8gz3bJXicWDBy4TKjSjaNAMKK/mmufIduWqNE
ou/+ztFE6p5Dw0u2K/QUWJAIRznYcog8gb31r6MtPsMsTs6IK6aNmGVCZ+F6m/Vz
S9Eut0Xh1e5fgVHM5/F0AFt0xDSj1pKyfwH3eEcMKG57u2ZdVD8qDtEeEELYqvUq
lUtEyJQOYbFBg1Wf62uQquwFZ3EPcgW72lyA+QaMawJYyc/B/3JVx39WvuDR/a5V
if8jhazMJf0oJ3OHg0l1xRhEhQ19+C2M/42irFzP1X5fn9hkw08SIjHsCISwqwVw
glfzK1Ngq9EsdEuhmbWLmD6EJ0VHAtfaKWVfWuaF5SMIWnRPD0m8i6E8W+cbPuhP
2mgUf2uxs+GegU4AX4JoLOw0O+GulPa4rPK0vnpCeNYymKfHAbm3rID7TFJl30fz
QmYPGaeMEzMoAzoiR43AH+Gs31Ztzt4nQ721y0ik6L6DGUz4MwQHXC+gNJ8rpwyH
ehoNlTMUvR7eyduhVWjDZuQg03UD/fAeQP5tsExrhZUj1kfq/Jb1DenRWgg7paB4
GM6FangNh7PdmHLo7O3OmFGDGWWQjRhO4fCLWOP17Oy81f53zfKI0oDCq/Lt+sAl
DBxyhwPGBds36sunQMGIW2B6iyrtDPA+L3T734Elgy3mSO0TZZlLLRbsurbKPsiO
LXCIeHhFYdKIVLpaKj0FdDlz81y7eROfAl26GnFh1/LDibUfyW2PINzUgcXDPtim
yMQ6tozr38JeSgcjvVVR3lSw50AAZr32mxQuTf23qbLi4D3y67y8DOXaIcoL81sp
a1TPYJcvmbu6lclwoZ+KrUglWItSgy9lWX3yBmHFQUMhNxyZbAqOmMlTkyAWNx5Z
8N7JMA1BB1laRrumRS9/YL1zkpCx90NiF/WezGkfCgegcqphn3rvSFp26V89M9sP
CLEPvfTgxRg0RmfvqdxrtuLO20fWxRVTMS3pG9pHEz1EnAUzphzyhIIY14TxLk1a
Hr3DswsvG/sADyvvmfl//tDzjp2koQpqBrPg+d3S2IzNL+KHuP5xz6d68X0TVjRt
x0H9uvEyHLVhmhnqgTSjIi/RId2U9fCqY4ydSPk6BBT0FCsMHrWNv1nLefLGBi6x
PjW+uY2itj3YVO6AIeppYG4LIKgdyYN2YoFlZUUPrOllpJxMAD11vyLh6GtW4fLi
cSHz9pjBHCh2udvSPomEcyUsI1ywm9NEzcJMjwKo3vvJW9oT65MSTVPhq1Hxr42T
23DOP07h0K62mSEKqy4khB0t5e7tNm7ukueelyTXMP2yqolXMvjgsvyLbhYj5ZD4
JDjfYnrwy58/dPdzi/wyVS01GQW3MDHojaLsSWocIrxBFKyCXc2Ho/Uke2ClN02K
wLn+OqY1JKaRkY39mgifVhf2a7rlzRd6t0fSRvutkxkH4kLgcYGejsAem4lCyggV
hofNFn563VLyJRTNiLpKfmI7RWV7XuTFNUn76AIZOdXq1RZgLjm43xfffH8Kvr4r
2t2eqySXRpR7ZHtdYLYBY1m+Q8l+0K01FIlOe7FSf3744yBhr3mzRodmr8OLCDG0
rSuUuWLwZ5p9N8rXEXXpzm9hXzFYacufd/f2tiNZvUjnrH6xbQBeOX44UguBx6FI
fRMVfb+ZRx5eVdvauvvn6+DmYYWT76H+cuU5LjvOZL/esFTSeEJJLejWwpKb5O8Z
Fwf914l4v+vJBhn5TWSjTWyqLH1Zz2KMluUrKT88pSAciwwJs4feK+WFVumAWbnx
qSVx1TA3+LRZknfRDJFmGp1KVQQWSmPH9f1+V6on0Ww3cBPmyGAl81QXqWCO2H89
ZCDH9y4oW+Mh4hf7uwJoui2FwVHiwyIX0rQ1eXzv1AHyVx/+hN5KNWMss5IE5Fye
XseSI4N6AeBkQ2R9Y8WBJTRcd1A6kf4Fw09KIlV1weRuqYWozXkk+J7InGR2MuFm
RBYJcy6xecuiGy4rXnkcmTK7JkUDdZYOh5JUXk1nI3PXyhq37k89pnOJxA9uzcZ+
lHw6qRjndR83orbJVAlem7vm1xh1bYmrRve9/1jVLBNhKYWF8czAOYVUKty39bGQ
hpbXRqjJksvdHln8/H0vDbj7NSfkyPw154VNMizRCpL8GtzucsJ/4JIpJF3P93Y7
TRuDQUFJhW9uioQQ1OrGuV7qR73+SXpLB8HAATvxiWhanHQN5rY2sDuQixnPbbm4
cJmoNgRzZAFwuXBy55AGma8ED7PA8uK8+fobJACj2wxLUgrlOvLSlPWFW+0dnVK3
6dNqUSQ1jkdaW9+ycqyXDlEVWLM091oU3ryAz5z8bLBpLO+C5DL7dkt7dvyXI77P
GEh1KE5m6zuiGc0A5g+Zt6zFFq6rU/49zVaAuqczkJEL9fYsPViSJnwk+Lb43igi
8dFcrBUpCz0ne7KPE9l7qGwLLWTsIg/r+CnXIBBpsI4UebcdgcqILICYgCXo9llA
M/Rkx4QtRdJ7OvTgBp8ksf0kQU/pIRXKn9cgKkmqrdGvsumR9lD4vLfPFej5p7NL
FSqreVSfbLcOwVOvZMUU2oYErlxOGzY1ENDThX33WFt1LEchPeCYHAqsujB/KAcq
lQzkXfNcMeIIvS+MCK4pbRHfmmfaFz8LFQVmVT/LtezM+KX9a1QqwW5tQUk5rRoP
YEbiIGhKPnZivXoO9YfjVztHDYnDVg8PSnk7jV836cKpBrZtdHDdD4NKu0ff+PM4
WnH826ZnVqeT4Vm/bp3uppGMXxZdr+9TCgds9DOUbj2U5VLxc+Y4F60pYyMzTTwU
+I/vXccZD9Npqb+4H/oeq5BuGJyhwb/uCuNw2x5fQ1V3ubm7jSLzPavlhyblytFr
/iNud6nczlzqpmiyYCy9AyWoaeVIRgDc4dv75eU5RASIxHqwtAurJT+/FDO4HcbS
iTpSZ415KRqFFSTo3PEyr02jGazdI6jf9DyHHh15VHBrtLuk0F7HE8g5qwOK7gNZ
MIjy6A2KT+eA1azDgBEmJgRtx6Czy5Re87aam7ZDgc4GNNYTzppCQqM+lnaw6aPx
Cxd/MOcjBOpdOM/GY4ymXrr/RnIcPMRU1p9rv1QF1LhsIsmh39kC9/6ocpjEFGOd
HBa5gMGZGcI9e3FXMppJHHOmd23RUZdtcRqf2iZHa/rn+1B7dtPxJPtq1TkJx9w7
wyAkKzKQXO0ybI5Q+CTRw5kYbEbuEcqp56ZSpRRGVV4EWhKFM+D4wAGqXMaXTu5T
kx9ecIRZS/HFnc1e5mrZVnn107NKhHM5HZ9CZNyPZfh4kX1S2cI63tnOUm4nyoZH
jl8ooV/CGlIBORnRu4Skm4lx0pIn1F9a/A/yasWKun4Vhu5AybwlOBWJ2q/e+sW5
pUM1P1Iu1px8KY98SDVcCpYyo7iAslr5Z8ORgj1sv6myVE5vT5jN52jPBPN+q3tZ
jlr3MWdLLOyV1sD9ELhSmZ8DWLBFMiBCsG5mX7DnPPeqHHY0k1qcwMxho/k3nXjO
NUBN9wPJJYStjIa7Z8M5NWRY6pHa4HFom8er28jKOJ1j3cZHWcuveriQ2QVkLStR
2k4XArF7d8z7/Cl+L/CYFWYzKBnU9xtiveysZ8K2/qN/AJzz6s9mtiNyDn4T8L7u
uP1VGkdoQrytLorwhzPTJ+/mCHUgPGHwd26MP6XC5uqj1K54KzgdshtK21mo4PIf
1v63eTvMOpLOOm+s7toU/OKw0qI4wfBsYivxLZ7BgLoi+Sr4JCBpgW+BldMdvY7x
aqZQgfP4V63nqdgBzc6ZrSMJo9PcjWBcheg1QhgHLrLPH8or5vY0vjq9urzYmJiU
EtbEsiopUbe0/l8VxDf7ubWHX6Nz331P15Qphf+JdSO9kg+adLDlALAgzOl57u65
Qj3GYlvVoEhmtoQCtfr0GySAyXdXTIQ3nxr34det/N6VdiFTcb5LySORDZOFmxIO
81jH8uqwDUsfMPP//h10bodAmkXpxv7KR+BFewCo8wLQkfKCQr7ixkz4H0c1E3BJ
A9JiEgYaab0vlw53ZxP6+JUREsg2Homd86R/ForlxOg/mE/octoXsqCu/Njpl4mV
Bildy10ZuYQG/0hdGt1iykYQ9U/LZ8G+VKdJyS+iH1pVrPTXb6aMUIpPrXBIAbcO
hqLa1fJEeKrreprvgvuC+qs345HqSg/ZQZJvNwX6uxOEKX30cx8BUEtAQmTUf2ie
78vcJSXgg9sentWoBw/6/HzHqVX4vTpmcf97AsZ3g9I5RG0RA+X1m/2mb+p5epSF
gcNjuklG0RJrb+6p5TaYU2ul5Jg1xk6NqScDPwkiQAK9XH6AmiQkkv52O/MllOmG
C53pA+cMiXlFzkIfIHa991XaK7FAnmQLptGZ6kPhBCH9LNSKu3+7PEZ4FBY8J5tI
UJ3NK9//X85zn2Bz1tR/xXnzAj6QQIMc1qrxsFYpjS6XZmRg2RMrqZrJcGYFqFOg
ROifR21Nsr2BvhmIeCYs+S2IIymlotZUISfR+E4U2nmuqA1VzwzId5cvoK2C4S61
W+kF+l7JtSyKZGX1PRRBp54MBY9B6XeETgESc8X68mEeiKHfMFh7hjYo/Jg9HzUo
ICWfLMVisymQ9ChOR1j99Hc4Uz/OwMpepSSHllSnF1HWbadr7z7yluQ6rhxm3EMo
MFJXU5YcnXf4A8B3r4M+HjHo3Nm54eytAnLSfwN+BxZsrvkd2aQftUsxSxD2RM3B
SZ5k1KTkBO3vDrU7WwRn4rd/FGTa/ClJSMmbSAAtsiWjSQ3x/8fwAnlSEBvLo2Nj
h+vGX16s9FBo96rKONzq2ewDUjTbnMVahLg9Ff+tGcCrcYK0FcaG0u/9oiayAMcO
StbcVxEH89IajBzmakQrUbcaOSr6rITsDJxYzjfw0OGVBKySOXsosl4/l5a0TEyI
Bbp+/nRyXln4p/04sWNaTe+Oy1n4TCsqqM5TKGZvoC7jkqnSL6545hYzzVPT2iw4
nXFHjb3HHSLSMWaBIDXu3qnbrgCTEBHOgBDe2J84OAN9m7D+jLZlVdGuMekqs00j
P3KpYI9rfV1gPIoSsXeAATx67ma8Pq3Q8gYoR3xWeFEhSkjnSPTWcAKcE9pMmsjc
nZR3z6qXSIp3Em8Ssc8TEySOZa4sb8w4Z3W5s5NWxeMG4pkCQ6J7NmJ8VZx0ixz6
EUQnbf0pazi5pUzbsgsE9fj0Y+boFCMUyzX/e2DXwTbLtR8mf9AaZ3D/DfacV6h5
fzFc4zhJMrB/wisuVzG2ldTAr5V5kXRLFTL+1J8V6cIFsZx4FYibo2bszVBWIQ38
QiEF8dgxrfb72sUM+P/ut9Pzdtap45byCPJSRbX46gP0a5W96c+zakQXTO6LqLUq
N5sOhHYo7SA2NszfSrv/rrhb+s7ozp4w6MLnCkXZ1Copj0IWcx22eVSDfU9tv6Zl
ZMW6BP1BHqkZGa6T+5Pmtq9C95JT5EeOkwwUS6uhOhCP523dJ0M6ibONi9wGv7Gl
QOC67dKET1xUq0rLAbSYSaSKbqsyUQpLqfOEsEVh3jjadIDJOqMAmMU9Smi6q0B9
ITSLIDJMoKPl8b1JvcgMr2C08Cl8OrkhTJhEQwYersIA/tVc9luCX5uR9Zw0hxJ6
HNlW5Olp5SCRRBGj91KQ3cIXzlKYElQohBb7EdDYkVjnlveaFoZhHvh3hsBEnCUK
0PYbfDEODJFcV4v85jZNTEduDU5A5kk/yHA3cFrrXtXr+ZTghKO1AkeLQclP8X8A
6/E/+9P3XWNEe92U5pPrTjAKk912U1E4kHLX4yGGXl9PTh9n52hRUIN7H1NmpPfa
XuK0Dx54y/56tN9eGxwFaH3NH/tjrKuCfromLzjiYIppB+hsBjlhsdbUgI8fW2Cw
ERakZsc2c8OtAX4h8PSkTteXB40Bg9Smw6iqSrOBKD83yE2FNwTo13XXVh19KIvR
Ml+YyXqe244fmLYq5PLY0a/wHdKAO10NSbCu9cgg5E/gey8v9PI4IwCpQnqrstny
0EdNwUZcwHXocSS25fhaI4Bu9yP5tp2TLgjlRhiXTw3pU29pQUbVukAGeVndwUqW
CFCldviVZiBmc4VWuQtHDd6KKHEDznEgaxeCIt9og3rvS1/vyTwbBwzG/uT2BX6T
3nKVduUDnQSEXOLTt/N/matjWwGOwy55meooxbpslNlOuO+cQO4XMZznBob4oof9
jIFlSWo03yts77SHST7wG4haY1B7pv/I3bJgB/Z1E0hxlY/klxBerLOo3bkPFej0
0O2wx1dus6i0R1xTZ/71esi0fMVHqg5AgQn6b8+xWJekHRLq2VrS9QtATwOj0kh8
yNV0tX5UHaepO0oVsqGbOST5Qy3eNa6gs8CfiNljodbf8MfwJDbgFkZXbFer6ytK
a6boGqEp3MPE2d2Lr8m/+lqP1YJbDbUMW13Xd88eJbodS4cwlN/97qUNL76VjbRw
RFGughqdTgaz6gKNiurVGx7f28Td7vdXfO0bskx3bPKgQ3avds8OfHQm0nZWe80W
n6EdLw3IdjJz26cGxw1lLMXd6Z/WhSbD5Dsy+VXHzXjlP+0UcPilxwIgXKn9gafM
jS1uXO+k2gvctd0b7fcARvXWs9PlGNfDcbDz4knJMQHE0mf6l9m0cN5grzemLiHi
3qliM/7/DBAeQgY84WWM7rHddlHNmZ+OrOZFiJKQ2d8wBpYlU/s3Rua5qt97YfrX
+j+N8VgGbnTomtQvixzFnc5d2jLfuwj82uJs3zdgGnMWgiorEASD0LPN/FaVXHMo
cKqsVKVW+C7NLM8eckDrdAfi8golzLHo0Uvcg4Fl+oeiG9SXsuDyE7UQDYbxe7r6
t8RmeQjeWp/ccpuvHPg859LureHgjU+G+RwvPv+JRb0eid8WB/95R9FC+YoJePU9
EJnnUkrpL0kAnpUfemP4YRBA1G3B9YbYRuOAl+VewxKDzyTxVlnzl4qJnEp5fWmt
ZFYPFeoX19NE+mJRAkcUe8/SiyIrwsO45XvCSj82QGNKj5COgC0DpGHU4Vr6uXo6
0f9AqBPbAr9jYt41z4s0qpsm2fW83qltdIKF4YHCZahgizRSsXwSmyh6iF1Nd/Lp
D4Q4aHiLm2FwN4DJ6D4lPBKOpxkTe45a4of0wpjcKOUHhR5fhx2ypUVSPVaDuiok
HtAyujxD33rA4oviHJUAmPa7OeMGrGVJMbPU6cBKzVC+42jo0J3sHASQ6Vt3LCKc
uru+zslliNGHCezpA02UmPW3AlkpqjcuTCx7khtp17ALToYElHs31Q5B3sUtVeDE
OseuBcdxC0Cq1bGydekfMi2n9SJxvMvO3WCbhEnrhrPnXG+t3gZzZZAVL1v/BxxW
NFufiWe5yUg41drEJWYCpMnVD+PqKHkTSxys59jzDZXluw7tHieYoSwakfIQYniN
o+Vrx/vsV83KUREZHoafq6z8fTLTJv6eJ7sljRFGt9bpGedpursmndGtyUBtPdTd
ZE1M9NyVcGccWNQY2+pLZ5lULa0r6q8bpkLx3HkfDTjyxtLaz3c9iAbWFyV26zkC
vNH0GR6R3eSvOTIsUvg+Xtxuvr9AoB8Txnaj/1eI/PRwsYxt/mzjihyW2GXgXtcy
vBKuwDSW8AxHwDxxfPDDQFEdzxpDyGwCUduBSDbzP/A6EQRpPAElpk0MdheAvsgC
b1j2DUdNB8ywgR1K1ltUgCq+2yhZNOFvKe0sFtLbtGy2GbFv5j9Lci8J1U/bWfOr
VhLqgOJbmUea4LVlQirzRyg2xKTwYsT8KLRh/tpbjFcbVAWOnKXfvKCuA/gMHvqD
3knbVWFxKybzlYEdyLz5uklLNwejmCtpU1t1mBG4J47l2pBiFCxWryunjGZ84ydf
u61D1mKz94eI8+Ge8uy8/k51CjRqTpNSXyPw9oTCe6wmmSbNAAKdN9mpFspv4EAY
r6c/ANWKNt10yXFxx0wXlEIz7ukUPE5gLnUJGU8BisjCm65U195frfY1gaMK0N7W
mwGNpeWfBonT8HNNxa8OnqVv6vkGzbCiTHywO1T6Cpn41afWaY7SAPyswyEaVKaF
Cy4AI1M5rT5PNOLTHkSTLOO9tsFGyl15s3c8D983BAmWGtS4uIJJ9vNOfQQlAJiM
Xs7aNBW7IfqC9Xx5xQZ9HPyUMjRghFR0iyHYnH4zQSkoBLj9QJ2hIzJTgqWxhzVv
lP57eRVLJx1JK8VC/ul0qkWtPDPorXbqAxP1jSvyToh89Zld5YrCwxsOUa8qpLJN
Invq273QDn+XdKS3FJsgazxe+Vi0AIkZreGMwnZ2YVaRpmpYdAXbGZwPqEonTYj9
Ct3oXNgCk98m9egmQhAX6Ws1OK5V/LOytUqA+DuZEnPji53OnKgv3Z5EIKxPhC0y
4KKz9F6e/9YW2aSCfF3Rt4S0FNRh+378v5z7TB49oyn2kS6eb8e39f38r2YmElXz
ui2H+UmrJuna5nFkLfKNDqW6X5aJSfkPeC3wSSD7INhu9pGekeSJQi7NNla4bBEZ
GfJBr+sd7XdpzM24tnBn4UUiFzzH4a8np/pckoIqryaFwV5QcdsC/t4l3/LxpnJB
MhauBP7+FD9Mcy62/1gtoRj69l9SfErZgwIojEIfZwFYDHb2rfMmquktuUjbghmB
IL0iVPBq1Gfc/K2Z3PzZ9ZMdp0xBvobk8vLyf14/Y2Otb78aadDZIoZXQJCV2IBg
uPskAZrY8+Tc55/B9z2WDc9b5zkr4BsVtZbsKarxS2NbT4bvNzve6J7cPHmyUWvJ
DUU6bOkkhPngJOkWzhQrTJDvV29WK3iGpVT4BtXcaXCDDI+V/edGWq9d2TEBiFbp
ZOZnWIpV+Na8OwBAXvUE0h5qK0e4kl/AxX2JY9FNW91W94U8n/pXOp9oVgkgeMuk
/ofZb3XQBWxd+7rWqER9xuhLB/ldX2XVPxMK0bFA7et6BXjJY+BYz0j0ZeTc9F93
3FtKysyMC43KxUo/IXYsTKwyYG9qCl6pr6zfFtf3kdGrYuY6e9qgAir90WvM7Ldf
UTY7c2WOytkhVX0FEG2Ij1mD0IqgOwtISLXPsLcxRbY+/XyZgvHM8j3PjbmCp9HD
BPJv73mDvWDfFrYMmnCTeStUd1S+iAh8FcCdFjELOiBgse1cbitPiJiO4jP6ByGb
c54QcI8PdczsxZyLCy/CrjbJVAwtmtr3fB/tgRqclXL1LmQUaN8iMHu8y+HSoMd7
vFV2j6WgHb+iILWtxByIzsLnShmyyEt7ucCgCni2CV7kqWyvCKgDbNq/6qyZ3tkK
MZ5DhgWEN2QhEgJ+H4NNwJG8+91Pl9RC5Q1nTfp0ZfR/HDsHI07uwelV+sHexU6j
kJf6feitvmzTXCRBnZKfQD/TZTOs7Z0IhSPmJ6cbimIzxoSaxduSqRHg7879G/D1
CiqemMcvrq7kru9kVQgINjgHewWLaZSAkW81sg7J/N5E5Oley91ILjmwtO2NUS57
4LU4ADvUdcE3eBa30MGAmEIvlHpOcMD+grBFro2d8mPtfU5nfQr+X48lJAonetYB
yb2fug9LMb7yLeTre/5DvqKURFk0MQJUdg8DSjko5XgQHm4ZbTqIiPb/55IpoP10
LdSdWu0lGxZIYIeU0p23lYV7OGs/9WUt+27mfEWMydNP8bwF1n/9YAcGdiKnrbP+
ijVpWtRCrwknCB5KWkSKlb89HW4jbmuobmODYSD4XrNXHHG4bJnh0YMDIwpfpmaw
4rcqmuyJ6RmsP3eM9icwb1CXK3anxXPN8BLUEqNHaECYxBXD1V+M7j9/kJaBgijz
F7/Fosq2g0b7DzpHYrwQrqm4EjZ2OHQIj3Z34h2aBrUSkm8KA8nnzX0PFutmX5Km
l8gBelvO7Odr0t//kbgu5eFvpiqS4BOlzAh6g3xyaI39UOh8ANYIBx+YCMQ+bNNw
mlmYH6Vug2fGQJIXMAQM6BS6veRv7cXCxy5ZyYsOwmSmC7Ij1X8nlryh3F7i7Ipw
k5RHQljUqONEE2zPZva2C6Z9pB2jcOjsztk53mOvCFyIE9O8cDuE1UbKL8cLnoOT
wIs5pMWN01nRI+rHwZy2B+HTF7ar2I6LXhuwoQ/XaishMK4iRv3EZG/dWov74RfQ
hcyXT5rVte+GUQHHYy8iLZUMId5ar4PBKI4JUrCeBS3VJXK2/1BQc6wTMdGTB6H3
NGytmPP7PMSEWYwflvPdJOjn457efc4EQHxZ7VuSHQq+Y3xzvMEd+vRrVjzGp/F+
MlFkU5i6RaKZMJCHP1GdyRL6Qpi2ou0bCQQQc+pCJtHUNmvPZjGxyfljiGgcEhn5
rlzBznArjL1xXZbbgaoke06dlbcsFPLiAttmnX6Wkc+D3AxvZks8JHnwUeHXJuoX
iIxZGthH8EolXAk4a9rRiP05OXbz9yAaaG641gjMPdQSfIMsY3xCb30GVW4s8U8W
WKsFSU7IJU9aD0l8ft+/dbtITDXvPyI2SI8bZoahDr0HWjAMYOzWCnrwfrVE+zb3
Gd5xwBEfpjzbQQbWuSPr4T8GRjlar3dlPPHSGqafX5sOIxz5hrycFYX0C9mFyGcy
zSdebWF4aw7PvKSQ+CCp27o95RQ1eO4KvQxKanfwbjEw2PEOP97xWhwfzXURbP5X
v7vRzFElF6SOK+eMnixFQeZW0Ox84B8/bH+Qyrz7t5cCyKXbQLzY9LrxCZUXr/+D
KPu+Bp1pmaoCCveu62ZNi0vGmI/47P94abiRwAn2xpnpHrql5QJAjOeGB7/jLyyz
yWHfbTS+a/LPLMYHgoKpsaMM7q0UwlEROZcmYYSR7scZ4TZclkJ9RaeRjwd+DkTU
S08cXsAej0R+H++i1It3j/f1hkXcsaS5UAv2dzKz++j2SzmLCsAVUS8V7cAp3BBA
T6Nqw99chp87W1jZ7v15BLvnY1zSf2GgzHDAO8T/9v2mmu7E1/S7v4d2hqlUnaHM
ODr6QOHhczhAA/Blx7zEThrSgb8TUpAAyG6cdNb7c9ifXE3tbSTyAoiYVrtp0Mj5
zjNrDY7t7eYeHfShzTRpKNapn0yuZgKhmwIduk+1nE+cjBJhCEBEgPTmW57eGxEk
QqL0zQWqQNCCCx7dtZow/g3zFXu8houAMamw+ZjWec24BqaFCTrXnSccpwenUfr5
bH72EACQ25L4prZYNYAQgVeHP+QLvO4Jxkic0S20b5tSWuMlzX0mhjXlPHEr1hsG
00XCBa0kZRHtPdKASV39thJvXr8yTL0CsHO1X8yiXLwTcXiJN44JeU+5rzMFrbO/
orkkkPYYZVe49ZGfwZUruZwJRbHjlyIx/esFxqTDyS2eGxuwLZX3YM8Bvo4u68hB
bYEzqoHmPe/LXbtmt03XcMS1vbjmTn9JsMtRvQ4k5McXIuYju2L7453F8swdk0IB
XK9LZDZ0pFKVpVXbTFjSvbwtnbzgpy7vWnz+BXHlR1mKKQOqhObdSEPPI+NEepEb
6Su7p13s5hB+CqfW1kBRGemMdnZ5BADLyxrhzGdd/3jGCmGrHPOUUkFfg5bEp0mn
/PjxZQP5r3X++MyUiNmg7xXSnGhKCDlhGckM9huKVyzOtcP0C39ULJGN+e1A2By6
6Wcwxa6bJpaQJ5MFsTOwRhjbICq0I5rrUSqeB0NAlDW2muWVMa/H51bkUqxLn483
9d1VUsD+QHwFZnAo2uzwcAENapE8wqlJzjnJgVXsdDrXsUMm/5+6xYLFbg8TAiTM
eTo0gfU/EIrANcmArHwXzVopjpXr+KNufS2clkAhR+1dSdCWv0aT38kfGaEGkiKm
1OQEpqITudUmh+0sNqmhpeap6FDqmmx9OajoOpzMWE3CTRdnhXOBZ6ksiTiwpwgW
fzUvy9F6RMgsy4hhumqzSZQLeXIUlVS9d+JxqGQ1GCZDV5gwjZs9YAI/+nhm4ZFs
5M6t6iIDG6KmxBQDRINUi6HTNdmzC/HKK30E4jLVH5dM+jswKmcvGRvZFXNMzLyI
aJF36N/JJU2M+mmQHJSayqnV/Vh3oUzAJ42byU+a2Oya0v/tRxnipcBc8hB1mURS
5VKLmCfvb5aR/P3SIhkLnsuz0vC4wourJYFf9+as1CCs0XCQU+oWabOC2c9j+GNd
qqq8F5dv4ffYbHwTCi2ryUojzHdItPiyQMGwI8u/i2/AgbleXw0kLunh9yJX52Je
2dJOzUiWkgx9xB+vZfdQTRGvzwhw2C0OgVnLA3MSbc8p+YYe6QEBwKjHXGs6Lrqj
ZzfcijErHhA2w/T9FKPQwtELbQjDkj2dSs8jZC1iVNkPo+e6aIUzVcoFJqyTgXEF
9ewokEq1Cx8UMkvU8AVPl3hKFy4mtpHoBk6BzwQXl4tVDf4WpghCoV0zJx9ohlAu
lArBC3Vhw6yd9p0cSS5Z91L1AWY92/TBXEuZFpgvgT82RfLD/r6Dkr2XOla1yfww
U8R3iix+M1vBzkCiwfO9JUTZu3hCAmn5pPQNfMzv/xuIEiR3+uVCidlUBzVPEfHr
orVGNz4PWdRyZMO18y4XWhyw9p0qr/LYMdHcEMbZV9gDH9+Q6LsexyyKCE6PI+vf
E+RiT/N4ZepjQQ6B9oe2ZvOxGL33LFsS1IUkToT83PwyMEl+EOUsivVMdgnfcw7U
AR4RN2WDADrYeWhZxr0Iyk1ebqKUHmMwsFMogpIr6k591Uqt0E6o1H2VddU8xMZ8
+m6hbtrH/m11Rg09+6CzKVEv1DHhwbG/RDn1iwYOK43ha24lCLM6ZL+tE+Czn+pN
1MN8rCTmn3Myh/5XJMil2EDlH6vhtDsEfaYyqAwH4eBRdwROCAoNoRpQ7p/t6pWj
Ej5LZlUlrsaVcxXCIV/OESfmMhP1NTrIXHqwGgfrqL1M3xrXUnqb/sl9itbn03Td
ueC0uY8t5PpyiObOg9P3TSvQH9FuI5A0ib1zRPE1/1J1HNIJAgu05q1hH8t+htHH
5R9Aev0oQqsjDrQhbygawuJPDfrDAaF03QQD2dzB2CnnRCfSPrl5NVuGG4UVdm39
yODl5zzxu5IUNWHNcf0ittZtL3KSGQBvREcArY32X/j2qG6Z9fHnhXptZ/1/W8bE
Ur4m6Pun+FkPFpPoSC4gbHH6PDZlbN4j3koUDpxwvx++w1lVXmntj6gQm2L2f2ZU
MFrAKVg8ZlKnuEHOdYtUx9UK8E0NrCeuY/JnRNolE5f//lnYDtevzRsuGh/itzTK
yQ5zUIMW+GVMC9pBOp7aJeINHRp0wnDanOMHQ8VRsZCge9n8RP3Xh1+plZw2n/XB
bVyH1MsESh1Rezl9GdcL12T8ObTkt/ukhhrvybQGUfzBRlfJ7Na3LVkNMs2SxPVk
T3b0bH6W4bKUI9AXCfOWTjHAeXXGkssnEo114i5AgqEfLJlxJDB8UGqG4ptQJToo
wBUfLWZ6FTtgYVeLoxpOXU7E2sn+MZQz81ZcM/vPXtm5G/jm714O6eRLDlSkb8Y9
J77Af9blEj8HLpo7ZkC5EI9/MTYcNfCOqLWaT65khCQdU61Y8KAQDOMqzqrD1ty+
bbiJKRrtmShOt6NzwqXQveNduZk6j1ZXndlfTVh620Nt9aEimRPzjsnSwoGXt3AF
GihBseMXLGXRMnpssEO7vzxCPDBPGEXKJKFL1xevjYWc+HV0qQpj0C2L9kb67EwA
58bt13fs+maGkFRdWJUBLMOK+qu2wmhkepQFzAtVn6Cs9YB8rZWna8ODhKXrD99p
q51mFXB/KHWtzPxX7ZfxccfGXFAdhAszc70kOKrBJ1rA/1Htw/B5gaNpJNx+VDkf
PR5RdkiFhZbgoYTLb9pMPHUFhTxao3p1Fxa2ZKtXm+LC0Fa5I7hlO5Gyk0cZ17B+
7itYWvCcMwcK4TzNiRYOsnrsb7Xeq15N1VUuoo7qogsKU9aSbvmCJHPRD7K9OpLm
uGMU33RSPYwL2w4Q5T7la85AkNBGtfGrECYgS/hHRXF613lCkda0nhZ0YhWB3WiW
lZekF3Ahhwqhv9BSOsUJaHmdxzntqDrxKwyZIZbiGm1eNsxbMogcH7Wsq0nH/gH6
XR5Ce7Dr3EtdFQq+J5EU/d535/cZWBdJmHfHfwaVbCo2s+TvxkxTuZ0mwLC8pYqD
Y/scYJBJRtjqy0HYwvLGRvHisOZK08x81xKQBhvb+/NDGw+QTauxsq4CWj/W+uPr
YbF17X1tqSZO4PQlzZS6DZEHkw3HqWVQPTU0IqmAT7mvpwMiSisZ9v8BppwOwd85
TTvnLM6J4DLGuOTJ3Kl9xjbBM+8nX2xwmKiHa70dJEHPcL08pdiqVqqmUYb5QOZp
ERXeDcbgkyMLVPxIJgHcVwaNPLkDe2UtO+HUNDAV8Jt+yg5OrROTLi6z/hkP3E/B
wJ6WPatAhLEgnIJ7qt+Uh8aiaCPJuo4zTOgsLSMKJBpu9kekRhDA38vDeAMNTLFd
gRNzO92xiAi9vmULvIEMNRMEiVfkGUBgnV0m2wJsTHIm/kQhGmmCdIgjU8tmMb1M
ZGgjVGEfTjKEW1C0xii1qGnuqSHk7hwZj3VSFcGCj6wFDmhCKq90G2b9GaY98FoZ
8LYlJ6+rzw1yUKJuf58WGa02lMiYArU2JCFttMNBLKEabRjowqMS+7AvzRCSKgsk
rogJjILPDKCeJ+PITYuVFE1ztxAnCfEBSkWZcLZ86x6cw/BBGw7ZegkEFt1buxDQ
Cv04/uNYCKbdsxtBA1F5MRNvzM8M331bE0XW1YbyWHrRmPTWmr6qg5IUPEoi5xgx
AiIXnSYrq24JMfCmcnZcgulagBmSrg/dMnPzVIeIya2TpFwV0NkNqeAFA47hzwlU
1g78PgXVC8QWfzHE1DsSW5Wrw7ZuglO4YY5RTY8jR3vHVE8kUuJh6Hb+2HXFb/2R
vmJ7b46IYR+ZXvErYvA5wE5I3r6YE8FlwJL9ZJO1O+rDHKg1bODfuTU2RiMfZkky
jGlH/3V+gRpzy5Cw5vXW7SxgRgIgLvAF/4FSLqbMFSgckIZj9pHiSpQrvMFAak73
aUky6S86Eb6e9UzoQQD2XlUFoP3q02jacvaB9Kb4U+94DRT+vkdRC7/Q8TQEZfzb
Hhtkz1YvMKnDjZ+2hPBC2m9mrQ7OIv9oDMpoWEiiBH0/FVX/TIt/hdOGknJpgf78
l4J2ZBmTjiVjvrL0PDeDzCJ9LWjoG5x8X3hoiQ0PHqfyGsKevNvxh2Xtt3hw4Dzl
GlgA9srppLTWNXzCdKHfv9ma5jUuRuD1JkVBOsmisT0tczvxewxVOuFRvc9Hy+z3
o3VamSGrdl5OaQ+1/EhyZtfT5IbBe+1NbeyOFk1E/mgpq/RADmN0TcEmJFl7YLdi
ruvnZ3QlzQda+/YHmVw5SlqkA2odXRVWhSm4izPFQdHAqgUM4Nud2K0XTYBSpKwB
GTE8BIGt3Gt/BMo2L+o+3T5JdDz8L6xgolC1FNEsuh6vcNag3ImPoec7V3VUqXse
nW1/V2I58+9UrmTNTPtvTILvNWP6AYwzobvjdNad6DcL4tnG2xuF/ZIkkcccofgT
Q9DZf6N6jRpv9R/pafbxhS67z3keI6WevR/DfrYPHoFCb9VRskMvFKCqrxGMYyUE
EArL5hSra+KkcxPqr9uST/okgsymiORkb2ye/e2UUso8l5ZnPE84YQlJDu/+06dY
VPAMybZL5wS80xJIVClLpHZatnBZRZDOtRodDVJCJ8n61QLNtrAGGo4CalYmjGBN
Lm4WHdciNqr91vKWXu0xl/jOgFuvAyQMdudyiBopCM2Q+TVDBOK7384YVoS42b1/
yrk7WE0Jlpk5jVzC0d+MIunt4m0TF1ithRAc7cU2E/2npVQfCiN9xTqJ33LjXKQY
MfzwFGnkwgZAUuP4+F5VS6uHKu+QqU+WlnkSB3ShSDU/aNFbI2MJjG/kRsatxRln
+yu3l+Dq/kAvu130+iPY1UmH7fBa95CPzWpQWXrLwZH0V2aeG/4ZysOGw3L5P03m
Wrz4x/eCv4xrWSKVzgCVDXo+rteTrwX0r+QG6KUdTSxW5qicYixRP79yk5+smKDY
h3yANJjxcepVzdRPwn87WdHPKT+8uw+326kA685rNAHwMW8E71Ozm1QpYbjVGOA5
5ewrnY0RzFdJS65bse38qjGPnVjK8WrVSVzUszxqKCzvEO7YPqVkVf0YPCy0UOjR
T/6FBLRnSdSy0HphzJ+qQ6yAByNOhL2dp95qucbZyukwD3SCgT3SrwNf5MFPqwhQ
wgSLAQOdqznUQz1NQOwqBqIA6v9YivBsbDhiHAeeoqGuLx7FoMe2p7n5CwIQ/9DV
wlolz0KNhb+S9iTgP5lAxXaMe3xTokHIYwTPOw7qg0hi9AgxGGwurCvF7uORmZ+O
EDnM0P3+7z4C2jFzld1RzVH81if1X741D2/4K7hulJ3S4z/G9siayiCAjTFcjCdD
TsHm3Ggjr5udDr0IZIVRpvI6mBnwWKKMje53HmNrs/maxNLJTHPgG7gfdV+sps0P
humubXnFveZAnPZQp8gIaHJPXovMQLoHvwJxLuV8TlTpK7d7ojWdetoTRvHkcFut
rLIytM3b6JpGQ1bq1bKlBKfMZjwP1/cDKLDJoWnIg8bgxAAGATxzsVamTs1/23cl
cdRjP6jxZlMbM/N2SK8TBFsNKJf4z5NI1J1yrFfbS+wpolq/KT09Oaqt+PvOEVhz
3mUIYGu1+NUlFjLb1vs9O7P+oHb+oi4JxqzNzHxyr2JXtSdJ+5KOIQt0Acu6pYRo
zbz6SHCnFgYS2frddcu7fB6uDoBIV86MBHrraHHti8UzNMshGmBX1Jj9prvNtl7T
DA9KouHXXTMtUhe93wf33oscb0GeieFJcm9DktfRZrKIkJgQogqu16IlCpTiJYP+
xFqOSLabluhvuQSim9HbK3WGP1gPHTeL9yHw9zkIe4JRlCxBn/7sNlrVQOhFUp10
LzIAWYJ7m7T4Cwz3WszutfIhZGzkxqnfgGXkd7z2i2Xeap2LKqYBFswzAzoGZA9y
yifV2aKJ5MhBxR4XHTlqvfoC2XN/q42382ITme3XISFkEm6apVoOWzSuEI0bX8uJ
RmUcD0Pd4pd2wl/4C5GG0JnLUvCVb3sNEnsdhc3nsxd8467ahwYR98jGnpB914Ax
wtUaFXraGAPcULZ1Vi3QdoPttus1MCsSTYB4a7Nw8kT6kKV/D6LYyp9aUXUr8Aed
pExp67JiYNniNQLVoPMDwk8PZT1rU8dpvpwEtfFRB6vWvd5GO5PMB8N9DCWBxkSW
l2lDB7/ddYvk4PPiNBqmTkI1Xd1F2Joul/+irWGnCNi1dGPHKZQ/A5Lzbxp8cbgo
lrMbdgr9P/T3w4oPeUcWaGULai0IFoFiaSQbHT02vzGgdVrHCtNXRNsqplfYVHIJ
Z8zOjB8Lk03lkCs79uHkxfPJ+aD434kYV6c9D61l1k7CqxcyNtj/ZaB8fp+vy3Yi
PoX1dFJlnQA92dwiPLvF+ZKlr08+18lQ9I97hhNZ9Uw6/UDnExqRAk6baR5Wwq1g
r6dvj9GP4vLGyv9oGgQgvnqLCoGhLMNMh8TOEndJiBNDRM8acOWT4AyLw34CK557
PjFNNogpXuYWDn7MQFI549sQL5gbQD0eVfzJUmYyDtjDUzIXSJwxhRcESGNGgahr
u3M81R/fQSqHXu8uz+Y8lzPjZjNXq1KW8hoyS4anoGcd3UQhBnhDHEk/HUGsu1n2
Ghmhf6iKpz3abWAKxTtppEBjhGVprqiqBnc4pPwGFwG9rdBKCJhnZlrL7CQuHlrk
Rtw67m+Zh8NVwtjQEynFL2UtOBNHkRl4aaZhCpzt7qpUtmjOYrU3RQX+diNcOGNd
L17VKm1lkYLozjkl79uF1q+yafbvKKFASLHFpzYBUj/3g6P/znxRlFBd0e/iRZe5
ApotyNYruNTWNPcXOwmno9GlFonvkXlTGjtaiQ+/MDjKucligNRMKcedO6KIuHIz
62F3o1Pflcv3rpKMAD2GBrdw5uJf+v5ac7/0jETXzcimQ9cdX/bEVA8baUC2wImf
dopdLCNxPt554uUKH/XL23wvWqtRBlXKKvN1oiu2HG7Lzr1QjySFqofCFLFnzKwb
x2a+pdRtxdP6wp7nyELusH7bzBNaYsyXyvEieS7kvyYYl2cnOw29vqmxofQcVSyk
zBUJe3vtd4u4y4KDbPX9cowoks0nvYQVWJJZbq8AEWa8VdF8WNEeTUfUmr5qgrsM
uXMt+3aCOdYZNYMa8M0wufyxwcnel3UftgRITdglzO8V0elB1nI6qucwFhFXwcff
TtP/dNlINsjBqNlywODCEcc9bVPocvxmuigSPvw56P/6mfAPfkiV9b7VZ4yGcxeU
ETc6klsuXZWQqkSVecjPMlUmJJBlsKx55BTs23VHnO/F4rASbToLh0fBen29MY3q
7q2rl7CzK6ctgz9AsXdeJUwKMShJKTcrB9I6FwHG/0sXb1kFEVsB1wBoZRXsxHSY
WOaL7MdyjmDGyNLK703tX1f0alo+kIx6dhWZ0hsxRhEu6NEN7IyKMIiIsTAOhM+9
kE188nJWAQGt3icFvIGztYVS6+3ppOwdBhVLr7wAHBqveFyZtmHNnUdb2IHrX6nf
2vcPhRNHBQIbiu2DuUHsK/XqDZ/KkXdTiUMiX9rg5QFo3uMoyTxZxhWZdV7eRhKL
zf8Xfjg1qWt10e26bGRlMQGKXk3zSc3aJfgZt+B/6cX8hH2RLU9rYaDphNR+oSZV
RCbpT19ibfoBgDFkklTyINKS1JL0rb9qnO7O/S4VZLNbjDQQIDJT/08TBcnSPnHf
bOjuMqkdE5gnfzCXYt8VKz5KUigExwvGO/9mrEeY00ayD3I/rL7XxoPboFzFE9V7
yVfQb3Xejxzp3F4a3r0+HK1qnJ+fS4/Iw0IY/Fpvq+/MJG5y0IjViEvk2puthcUP
AyH9E5bGejbsXhO88ADboFzWmxtOMpAYsF2DslkZ9va54kMKbUjsPndmX2HW93d5
tBQiyu7hY2vfdNkt9HmvZIla6E7yYYSIczjbYmxIWnuOEmX1S6XvIJxrQMHaF7JT
JHx5J2Wk9E8DwEJakN4Bqp/2qUfuDAUvM+l0vb9lxRGGHLFzA9/xJzJZaTmVAptl
JWzSQJiW4rcyZYEYaIIaIcJ+H9KNVTt9QMFyBbhDKX3QUSbqf2eAJ6J1CqyJpEtT
QC9aRF8obmQxW1W128SuYAJi/xYUJmtiCbCYBqGBOpfxENhXP5UxyAb1sasQS87f
EKyXCaEvAwcD4XaeQIgaDJn9pRG046AD3sL0FeGPyl72YbKfj3l3tmJMXRFRttgk
0rxYy7I6obdxlcwDnPw8cqS1X/rem1fW6yxt+BWFQaqG+uOfWrTmmDiAPS/1AXSO
Gqkqw0T9DxYQqZBW86M4zHZgfremLQkdQ9QZqjFUPGqA/hCbMrPoKJNZZ0A4cxwt
iX44bXPjrpkv0CiERneUOQPGbRcS9+uLW55LaSAvTDmMWpqvFTPRdMr4oO8T+5SO
CNlIJZKkwREPn/Cms5hQ8t9/3MsEPoqQHhINSDzaUgPnouXRojVEInFbBbKNyhUN
gVbCGtJx5rCiJSdUTC6cA7puvGgvk1Kt6hfkuK0KM8sfuvx6GVtW5jcvjSrR3K1G
J81PNlXpYizO4Ae96Pn9GmuzVo2Xal+bqgLhqSJTe7Ggg/9fiKY72l11pOlYzzNh
EDOdmpUpEcDAQ82wK4+VraK5IDnyoL5+gt9qTgq/6NDL2ksTlbC8WbG3esmimbJC
TYtubgOb23LWb8Mp+BmVLJMC4HKvqnOtRVZ7bys/LV8MSU7qmyqY3CKtq/lZNWnm
jStecAo7YC3MWGcXn3RPUjilgJdigacENd9zyy2ieU0CAFLckBdE7yjIRPmcnQSw
vvGRLcrXpo1Xcc3rD46fyu/Bhy/x+neOyfMUHc2xfvilJYYz/qFLZCJo9HQ/raC7
CNmT/rSJ8ioqrECY52Ecf7SacbryWNNEBg562T/PWY49ZwwC/mmFPiuD5cjUxun9
pArQWUlKloZamtS6vaN4Co4Nb4sS1b1Czl6Fc7dim6tSO1xlS8aS0AkK/SBWcSe6
OcCWP1IPlDuObPEWy+E99WQK0390cgKWO2YXNb2/lOmYc0Zw3ua9TsEMJEQyPfXj
djjFsDqpoi2orycW6IX3/iK126ZXT1tP4oYLkJ/H2SFiqmQsQCWiBC91Vm6gBQAI
1sjTvS7iNnwjKFATst/3iqrZgu+tJ5WYZXHsOSTNAmncdd+CPejJWTw93ZwF12Tx
zE8QSbeeYOuCupOgXLRszf9F+XcE/WdjeU/t/cisUTVzQ1xhmlLiYImuxwj286BW
svincYHftVWMdimoUZtnD6QFOCG84+CYTEdZ2fn2oOtWyxrNB/jdAND/Her6xewe
kpvj3hEDSBrKDMKvZJKTsXRtQxnVlP0gcoGf5VyGSh9/0I4woyYAtnp+oxPcNzW2
zzHGDm1QD4SucmwYFfxPR/9vlucrew6PS0A5TigzVHyccMXJ22uJX3NB+HZI1yl0
v64/UOw0P3Rg3B3PYQG+hIgufpHnuG9vwbNNR0P6ZflZgEOP+MtXto98ReNXYnd7
yikDnvT427z2xQ3n8AFarwVc6ToihmRnKHfQHKeS8U+b3IHsAYxdjaAJ+Pc3zASQ
tkScJsbpsDCrU3dp92Ntoo/hxfc/34vYeI2NtRrSKv5qzJyGtnpOxMVhm0twPyfa
AEQT+L+vhw8xPCuudp5yfw7FMcWvI/CVbNPYLQi1afeO9Burwn3aM3pbvUzOdTrx
UCmM/UjpGtNHYXY5kNsrS+LVI2dhWn5chzXdCDsAXiIakkh3G2Rw1E0CCDcarzis
f0S+jr1PHaTFcJEdAkpijeMgklmmKz5+gFmigTnXrexOloc8yYHRLixQIeu15GY6
8rHr7RjGVVr28MIjVWn+j0LofrKJbWU0EfpEoVUGXvSgzMvmUXkY78rQHpBDNhpy
VHdYce7yAi8oSv71DmKerPZfRTBVD+YhnI7clGj7cSQwREndwBYKr2hk53q0IndD
ojtru4Tqooh65P+1kRGKz9wymPToxOfPLINKT6/LAc7oabhDSVqpMDLykoUnnpPc
FdFfL5WylUnOtTZ+EsH6fU/VJaWF65jXxQeOTwNHKNSyIfxmJ4pU9kpNQoKXMUJr
Zl8gnV0ejueOWqBCD91qURAC1TVjMK6O57kFypeDTPPJVLGFFilaPI0LCXnJ6K1P
WIjb5obZRrx3neAKk1LJ6e0nyNWQp9rXlspffkQVsK6xuEwgUogFOUqNuWDf8+b5
1auLv7RpqkbFW9pouILZAID9OaGT28AOtbzzwbc47JY1xj+1AxYWOixVFTbzMcp8
g559cDwZWR8pLnOhx7DMvZHT0KF1D6OHXEOaGcvgHZN6CGHPWEa8tn/JcxPXE88X
W7S5H3BZ4foDVbsoDMD5J2UoIpHnjICb7L1b1IAVkivU5ylx490fWua8ABl5hsTr
2bKjlZdE1pAU43rwmwZIknkA5HfkM9EJEAbt5zrKDeApZ4UjGkmqgJH9HLvHon0H
oJSW3Txl7ZXsN29+VJUlmMNH+YWq4AaZ+dZQV/k2dFy+zNZ+fjWOxIW4JSbFDSvf
4GVseLYjZbl4WSVLpS7k9iUWjGKF3wTkKaUL0Sk3TS7TKqwTRF5Cr+uHdD7X0bP+
ziqaa0ySjbRCdWz4ogtnRRAcRzla/nVHHSpdOFAZwCnLXrz4QcZcSw7BKbCZ9dPG
s4+jysjdD45A1wkOF71TuFNPVJYz4aNfiqntvpoWl/B7JNj7U9EJOqm6kkmG/Ulm
bRbElcd9sDdUn2sRR01kC3j2gP6oHH44Fj4XOVPHmYbgVK2IhmLDGsYq719biOf9
4fdz8H0QBKobKZ6ss9j3yzmwS7A3BIcmIkTVWgRixebLcVp8JThnPupuFjJd5cPo
HycswR35kFZecVo52hu/qFPmOdSvHA3R2VCJ+nIx/Wi/567Tb4nJZkmGRIiSNk/S
XTYqthINrO3+dNXMPg15KbnhZUOBVPgVzgUeYGkEOQeIzyXxU8C/cH+69lurzujK
WuGVb/4KpmAXYg5VWwMBTKxWo+wJmd84BTG2SjFFy+cUWg7yFFST6rviOHatWeBd
quX7jSxpyOgoF/yqb2wmYyvKi81BwvblWnmfAMvDCFT6VOEUl9Twk3hciel+Lru3
YKxwdCLssg68plHBUouWi67w0Pd9oBYJTAwI7Z8XXGdi2qG69tefVgGI8yK1tydP
NZNvPhR9HRbdvmj8rDEy2iBVH8/F2Ix9vUWlX/RLr+j02gH7uesIySdYE+UbbhrM
HnHssoDTuTCWmaM277v38FfuL6W9oi0yiaJ8Lz9J+C4BgA60QT+MI41P2iO7DRZQ
eAF0rFsLUoFLsWPKUIgH8UYBEmn+/uc+P4JMm7cbOIbW2t7USlbwKYp4x0GD5Sjc
C4F4sarJAdq/O92gQwoCSS9ToHC1/0UUTNTMpyC9Mp9PaoglsRTENYKdyp+CwkBy
TfPjuUoepHEjq/OavirIdgpdPfxvV1F3G6T/U+wQsV5+0oMecN7UY2FqUwKw27fx
s+Mb4lgESgataYutG8sKymtKdge9TaEuTDvkscuebmxnUHBa2LLfdjsjOG9zjLl2
8A/ylX6sLopc3kEIkCc9VfwsXLk1F40kDc86Hog41889bl8TF5Qbb7TrIry1SDIR
bMFl1MiwpdmFRTwgBB5wc6XtxeEicUjdoe+CcK/BlyQyiD6EC3eO6+w1YPL5ulL/
DUux6Ehe42oTH2WchRDI2oticJlrNMCy8VpSDwR108YmbtEEcNkK9eSloNhdfKx1
D2IErnhkRClvnj0DIccuA73BeGNLcJPKybsgWbmKvNJSYLCqRqe09OptvWFI1aJO
STM3kSsRkMx1/snJjcrsYObzOKw+i39MdKBeigC11hAyfhsTnzeUzsiSFWT+EhY7
dAMSTo49A1P+idP+Kc2ujcBhM4056DmgOQHXLMXWAR67if4mrzgRyaAaiA0olqrr
3iiTMs4KRka7mMbc0OX+sQY9Bp5ERWd4F88Rvwb/jDsLgRZPbVrNNfu+8vjY3zdN
N/65I4vo4FixigqSVVc/aIq/zalOaelY4gjg89VAI2AUh9ugi+0fdjEeZWCPSCsc
BusJjpSqpwecdI1VNhCaYtCOGsvYFTlQbiQOU5+JSJxRTU6z5few8hSzobknHWI4
ivaUvS8Tu+9FyCl1ulAcwbEC5e+CCOtQylkLX5mh+SJdFppOXnBmaJJ/6faz6ZLo
wKkuK+7bOSbD5TMtPuFsfDkO6gngOa3A020yVUT7F9UrwTC2YVUJNEFhmifcEglH
ovMLYmt5frb8iyOqaAbiYvoIVlmpNsZDf76Vn5Cz5JPmc9A4RxDw69hFZyoaTOOG
+lqpZamzd6nVkIWx0yLwqtR1Sirrf+5IvKa2RAkaP6/kCSCFj12+7YgQFSmaYpiN
155/5C87AWVH8NQRUaaj+MDBq5KrJXOzF/JEaYlkYmgYHD7cT1w5ppuDEtl1xP4p
6MRpraThDOd9bG0LqssiwefYLedZUm2Uzsd5b0RkXoxkhuN+xtrueY9lFOSsPM0Z
1kxtAPbvdQNY6qplBcYR5vKJFhCvrhB7RSRTn+IKlZpxK/9/KjcfCQRmSbnGe29x
nYAJ6LT9ekvSmqMGOo2L1WtENOsGLT9Wb95piiw1SIKde7WBvz16KisLySb7eM6m
jMTO8mdwmdUSq4iabCSgbv0Uz6hy4kaFqdohTVzqOGuFf47TgNjTAkfoqYm9wpuh
yBvItpYnnQkWREZPlntDpuLRnlAd10Y8hbe4hOEENwRr4nrUgXFcLLAeWeV0bMhc
prL1hUQlquNCOujOtES2+VjldgVAJ0Z//wwKPXyTF0sKgX0aln7e3KExfz+36Fau
6BXvUu6f4rEYPZecC3B4YZXg0Luw4a0ERq/lECn0mAfUpkRVUeE3i2ew4Vs5ZtB8
A04TnH83C84uWQjIwYP7HXX2qTcJ0XPOhQkum5Np/3pkVYeiITSVv+lg8s2OfkEY
hAIuKacx6ve4nRpiutDCCvOEJw7XCuQE0hIWYpwUCOqRTjhAI0uIiXzIMAWUQUbk
Zs9aIoak4LWJ+2hAaxscNxaAeHTUoZCjqU3neehJbrr0TQ2RWyVyoN1bIqtHmbmY
CeQYGe7QV1WXhZdfBFAAO/scPQKdGgTkZPKB7iPh7Q0UWQxFCcUbElb27IMT4iQc
mxZrEQfAjt4yvEwO656hbaA/BQO2/QBQdS0TOPGe2G44QizxvusM/8DZMVmlT8mi
LCgkIkdj5H4rUIS/7IvaA2uUpDfa6wFrC1PYWB95CL/9p32Fox8iQeDGEAbK51Vd
FRSH8wjy9ZtK6yFfBYfTPQ==
`pragma protect end_protected
