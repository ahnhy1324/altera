library verilog;
use verilog.vl_types.all;
entity divide_vlg_vec_tst is
end divide_vlg_vec_tst;
