// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
NeupblhOb2KLkOqxAhgndqxEhSNLOwtnV+J3z3XYO+COk/ZlyKp5DeVwW8ekxFvB3q1r/0iq36gu
j9SgJKDFFLncUWWrFcH8ThlsMoZlks/xqjMpWWEDv4mxF68OhQSkptG3LU/fnSVgLod+UgYy+4du
jzUemexCTcJ5u9TmWcBNBuvk2LP3XjASNTHww3HsM9EyZxLa+itHo9yBKjD7Wr4wMm8JK6v3J+tI
V4ERhVMMihFcAdnFn2RIT289e/UBZQ995zFs/9SzvzndMT13pZ9oJGGe8nIra3S5GEHK57YKOgv5
dWhJehyedsgh06ACtK/GgJG+YUJmfLD6D9O2PQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
b2o7rJBdkP+6MSVk5k4MSGEj4L5Xs6Fuh/oMtASTfFHpledMEc9UJh1ogacd9dynvd/ZUq0jsWC3
bcHmPUh1JD9ykWMB+4Ila4cRONOYw/rFnVf1iRPJObvQpZJ7bYz5oIMCkfN8doR2YD6Mg3yU+bTQ
fkg/QBXgZKUCxfKimp0SlwLG6gwddO1HYq7OPy2j5os2E6OCVmJITAS7FBPFOw7HgEcDRN9P1qtD
868B+4l4+HfP7zJSPLQRlW4RGoLASe0hi1OJ696Q6nzRH/c+2k5iSGeu4GeKr08G1+3m5a7lgMiK
hr+/V2XMjhhWrznKLKWa3u4SYAwXaFG92ILS7aIROjvtu478gfIh0gLGMvsHO9oi3ZSvpExECRoe
yLHJsvmsxol8LyxH7pxFQK2NJS5vOjnr5wKHFZUytyFPno+LUbr2A86mxgtUvg2bMsJ1OumN9CCU
vrgXGFqpT8IFAk6HGTd6e82O5Bghi+DpMoHzyCHQapcEI+J40/U5SyUDsSJZPSRY1/llIMXB/Mwy
yHOlFcHwwOJJYRhLN6jbnxtD1hg0+viuRX148ynmpD8UvRchcYVxGqAKpr1y+OIsktmHaXPpJ3HJ
74I8a9J3PURSkmhRR4rN9/0iecD6wGOwZCsCJfIY/km+0bZRwVyb0L6ZECWmYZJTU7IPGuh+F9S/
3dWnebcxStIh4KXI38NNaXp5qcUfVUQWE99QzFkeSxz+Jp65omBsbaIRVk6BP898rNhy9e2PO2Lk
x4MAEx5BcCuUJxRjTgi80FPk++6xd7zfmC9hPzYXpmcF7j/UNfMDCr5AYS/NuBToPX3VEiCj9rKX
xix2VrH/qgH2uvy3MCZuU+tXmEVxJRaqnoX+6Gl2p/9QR4EGIdEOl6ks1uw0882WD87W0/qSp0Nj
mDqZfzCH0tcqPuwNKuOtLR37spypFglGlH+ToAFG4bhbYgLn8Vi2Bg+fiLxVR//2vwpKaqCu1YgG
KU4WAL02BNtZMFAA8RECH9tYIhl32u9gRWN7+lTke/2sfZjPCretQjd+k+3u/f5pzED6sn825x7N
Ehqe4p2VrHmjVKSXamZRipNnT0YYrANVSxHglg7CsTZSuKdlQWfxva/H9Exlv88JtJqv8aXOgszo
wW4ULY6CgUw6GADPDH4xodRM15joHyGAvxfTmnNoGo6dGTsXygOqrPJGfZMhEfHVRq3qr1gssbDI
nQTNx3rSuKpO7McIPdej6OU2Nsk+rYdbpTGrTlo/xNP0zsbUtjPUIfXy2UEo9OkcXxCF7M/lt9Ic
JDQn0pq2eBilBoTF0hM5qr+EaVQl+jMk2el5LWQnMiWq2JpJ0IVQJamZEQKZozTuUayOIDM4jigY
UT2Hu6hVbaKSkFjTLqzonft7Hqk1VwMLPQlfKKfNJuW7HqrfJKnndkVjACGBiFbeYDk7k1m7c6AP
guKgtUPV3SpygtC0Zzv5SxPRPFJBEEiQbMws790+71fQT0bUMnWCThKx8yiRu3IAl2DGnKTlXoVr
iAxl12y1LEyiZOYOm/I361T203DVD+KmdTL402wMfXlzkHWOYm6p8PPO6CPvi4fQ0w2BUl6KXoh2
c8f47o/unuXNO6/+4+hLkd00WkETWPNt2biUZQxFvs2GhwH+nNClfFmQq1W/KLsbx79JLXjwCf8t
ZqvOIrQgo79Kpx4ibZqovRVCT/Th+ew0d/k6QM9U3awQXYT6Ab4P7wIbIgmRJTa/aYgXQAUKCSmc
4kez3gtGLfFT6ofpcGv8iP1u9VuospqFZCtUijZYEpWX5Mu8DuiHUWpZGW8D8kQmjYnPvO/cZqfo
o8JPDQbmMqaZ8SfFebKA/2tbuOUYICabFO7rRLtG974Ck31VD98SQ6m7yXfvcbhjorANt7PRotJO
Yt3UTTJdZU/9C3gQy3jHEG49XagH0iehcdwEs8ruwyzQuhhn+oDmgBt6dQtOC5O5YdP5RMlMsTHk
lBPbn+Wc18B5lYF5w27B52154Gik6gj5WYQlGePuYZsOlzoayx5ceH7AyqNlnnvB7hk6x4WT4lVC
J41oti1TpW6jK/piKhbpC2J9HZVPfvChxYGTfI0Z7JQJQaMTHIPSx/egUsVKB9NR9y0UVor5ScMb
+XaVGTuwUxfpg4e5QbVrZGjJSdByj7fb6AMH9Z0Y78sFPXQIwux4yfCeX9f9/tEpXmvOkUKTIjHA
CbG/TsHiFjwhQRGbFFgd6BzEFoGzifr8R55XRvGs8qaI+RIyLMmCNSvGvsVQM17tinwYiZ+ULJsZ
XxnhbWmYzLELAdjvr7MRtC3eF8ziueyqMVHUN3xptyJD3udFhD5lMYB/OIrArLlffDmjVMLYHqGS
bBEvnQKnkmYMryH4GTMku8kJOwPne/9U5mFj2eH4EFoHxzeRtnjojgnuo7jaykq3EoDkDxLOwR/V
WxXt+Y1K2W7cgtCljdR1BwmuTrcj6MAdkafxYPR4rEUkxHETF2GUFqg6qZVnKnTugKWZdelWKtEm
7tXo/gz/+EF8KXrLKZtYVNXONC4WHDDz/LQ0oczrnLDG0p6767iR/OrpYL461EUSWLOwd2pXwHZN
kBNlM9BkUGE+p+DgF8IOzkPQXD5W+uEgntWjGy63ePA0CbSHaC10OYibRrtOV9rdtomdOh6OjgrP
gd9P1bP1JsxdcGczTULtk4FUcVUNLalAwtWYYp2iDZjVZejB6DVTdz2CTvEMNB37j2zYKWObS8OP
bQmOwCz37KDYsiEM/2hrF8i0XawUtFcJuJ379XMdyUofEwrZNB/cB04owvnGZC9Q9eXTklxEq9+K
THpRZV7tdso//wN8n376Zq9PQe4ywwPMtvbog53dsT4FU3jW+6EqKPG3v5kv3nOCTEctd5gbdLkM
pQzPEAW95iLV+iqqlSGevf4UtXkF1HnP9eRV+CM0LgmSaNEpNbjS/fbqA+HEf9F3DdxH+lJYHVC5
aqO4v0E09DogEUbPd4We+HFgVsdJ5cMod730UhNQnBcpbrlYjM+vdIjd3x7CMzcVaWpLLQgSAboc
LMBIcXun9g46dMqATbdrRhGu0VHx7xHqq+wAHX71VDwEmVkWhsD3NOq1kQQrhe2vLrsVC2m7dWwQ
LSi0DN21FEDM3F3DV99Yppu7DSkeq69V7L3o2bocKBJzJAALaAmPLXKFV01cn5TJxgtNBZhbaOqD
PIUdJlREhFRJTFNbQnd1C/wPgLK0ddEl42bMsS2klnjH5wh5SDobUIyPB9G+FqWHKUodMlPtPNcb
fwbL8uKkT5qyF+WtW1rXuhxHHve8ko3lcwr/OF2epKqL4CZr9Cp8jRs8/fGAbOIysmKQ9BSuBL99
zJ86vyW2kjNqOyoVBmqyZJfdjLYCewxynXOiSfHNJzqgL7b/mB23DT9ZAUz2Mns1Pcrvb5TVenkR
287w/SqhAFfKpHgcDXaoee3B9vWvpm+cnhA+q4EH+5O+FZmbppsEJCOSdpoVonFmlYShrcfbBDwZ
UDeL+QCkMLqjcUjOQYDVAKDTEgAZ+tcZkuknB0BB5egr7u4bEvySw6rjhqeEk40h11ccFjOH8Msq
nO7HYgJNgZhFjPo06FTxiYQuH0BP0MRFgq6bNFbhhXdVjZmOfzWAcW+BQ7QaSbXYKSmYpyQrRrYb
eh2lvdzSflUuDhiKCMapJfFee1R/BY4Mp6xaccuwzASpRP+dor5f+fPs0Jt4c604LN9BeS8wQ70M
SIMPMZJkFB5W77B0DXx+ZrSXrzeMjOXsb3Nu507QdLmuie2L0VTmZniFxunlhrEZSkprAY4vkZP1
rYtWgPWb4M0LNhvUOfnkCDwbWPfPG9Ip5QxdgYELR+gUzPCVkFtgMkVfcXNQ6dSVcZ2nq8Xm6gdL
DJSeWUBUhMFvZPSkyZTGzeHfHFmcnOlfLwyw91clJ5V+dKI/j4z9W1GAac4DrDlsYF0SCl49eJsn
KRjK5q9MCGgA77R0UCNAf+Njeultznwh+WSYGJ109/7toc/EsWS6hS7V/C0p6CW12EsudoRUs8e6
fI9f45Mt6ieMGV3ZdzMuooHOXwrBEUhlGKkYuebJQZdwbsIjMqQlUgnwxOukAfL3xeCwX0Wjj5et
hlzXwXFEKZzR6PjzSeUa6S7iObk/VOYV9cMh18zE0jUDGgXBH71iplHkT3bPzSInbj1qUzeDOfvq
n99hm5xJqlSiks7CyB/KKs5AEDuAEsidSx8QRG/T3yHULiUCvkH6eMYBmvQ2+EGPgvxv6xc7mmPO
9tSl7yIVPrFrEfbb6M9VaEFNSdeMZd8pZiMGIpQCoYCddIZS9X8tk1wQywKPfbEXM4wvdX5BrE8w
hP6zyZzOCyar99ogOF5GUg6qUv2QRQMeGSgF1fcpxB0jM82wUvS0lMsfym8Gj+o8afbeFD9YaR8L
1PXVVO8wDZfdlSGWCourCWz6IwMfX1APMgyXrmJydyBEasXEdrolmtzUuFv3/CE95XKYjp8E+OrY
oca7vL0dyPUWdg30sceU4BwCIeFATJU0nIofkc41dqh8whGP20/E+GsK0N4b2EUFm9TgQ6Xo6kGH
TPvzan/qlsDPeEXQUYeAADri7fqqwaDL+OqDsuVQfqIAFuwwwHlYsNZsaWh/yI1SEAQWDcdxyQ82
C6vLYG4b43XZ35V34zDdCjqm0HIEPpUFdDfzfac2T/ypAfyfu2rGm2OoO3UfWv+ikJXNE05mHkYD
f9bIPCzoc0y+qPxqJoQJZC7Zh/HZCmp8kXee2y00ukmcIb+np1mUEfRbinMwtOMtrljXX+cWIZuA
CbjzwZiS8Q1g2XY4OoXEIUWt8HgeGlXpwHbqlOmGGI2zMn9i+H53TABQ1FL/JzwQy3I6C8xOJvYA
urg1cG7am1qrD8iZuXfsdPol60HRgic9jsHhe6NNDyLWkokx4ccHFpfrenRms7gpJHwEiD/wDQ0O
o4Ub0Rup5obKfY/p13fdymP6aexOsL2Be3kl5iZoTSHES8BqbxjdHu1GINu8Zpyuj6lpmIecpPy8
nFEB4Jpakk+IhIAPnspLPYQS8STOyoV25YyFXM++ndQWtueULWOBUTe9aiuQaEvlhRuM5tms9a4Y
bmX9AnvNBtK7+D5xA30+weUQ4+OPxbXclkcUMEkG/3Rfabvs8vjVx+BTAUxhhscyeIzreqzjH+tp
XWkpB6tt1pftD1AWX4UG+iDy86juQEttKmDK35yYeqJP37XhWQT/6bUtKX7/Q9gEIq7RBaYG6jMC
xXeYbYEifcu+OaxUs0twj3qysnnBUET2q4KS8rJEf341xyyAmuGeUp5x/z3zwayXVKxuJcQ25gQz
uyDGEnKe7VWFEGceY5SG5GcbTTKvyfLcc96xeKvMJn54/ZRairL0bYGKewNmzi4M3groAPZCvYYv
h9/JNqQBFv1M/Hg404InwhsjTibGelhBf1iltDFHnXvUUE+OMsKrqKTM4258wW2VX7X7tKmRyVM6
BVBCjVkNVT6A/OWz91On229NM17YGDlPSHQ2AzKUkWEpflWKRwbAaPjraCi4MVq6AkoWv3J0OuTR
3mYGaNlRqngYvX60EY09n8eJmw+QM/q0g1Kgna8SUBp+MaIyIhAuEBEaXXTi5o7bbp9IY46l92hl
PCGvxrh5L+H/c9Ual//c3iyWSJgb5S1emUH1p/0wewrp1ETuuFVJ9O6thK94h8hgpGCi4jzc5gIo
aXwEY4d/+OnFLdJcxcQWO41h1dSka2g4p6gtdV6tpusnZdZl+zXpXORvZsnvcsWZVQDJ6uOG+XYW
xG57ljJ4JCKE7SVgouVSBtEXDvwpls96Vm9MX8HIhMk+enoTDPE65TgqljG4Eym/1LkJ/PeGOyI3
TweSe2W0P3C4uPmYH2K2986Cy5Zm/kamDzw54G5mBHgfccdAauMjFmWTn0aRTfiC7kzONBF0dv9w
9vVicJjIjT3Athn7kOucn5QDsjO5jkbHGGFXoUQues/m2qzcGCUodGkQuiJWbw2EW9uVcuib7on1
gz68tESCBwGnLgC+E5A3Z59+kS8quM4wWCfUm39ZagDP3NxSzH4XSZZIPWgEezo/YxtYLqYOcjA2
ZXW6DYwacwJDVSd+oFdLT+avXYWjYKe5ZH59S7R0/wXmTsCnFhiTu4cgcCyEBpRTuUcLnfexhLWg
I21AEFLUjyTZAhpDlyfzpmOY8Sf66EXhV48HxDHmo22Jeakd1HNPHahllfDNJfJuOE+YztlTAPbi
/JmDEBjPzk/YJfPctUDX9Zcm9jMtrMqTf5Pilqk2AGmJND/8+hNoFVDxWZO3eKhsoSo0JJQf0Z9G
1z+cIDRaqggMjMFq2fLTwwe/aWKsPAdQHa61yMdZVw2YKasJJ4R7GJJyRdpA2hScTYjhFylFMp9o
PSRYn6I1E5JvYXwt81YuIIh9UbKKaqxDRn/DhXPZEFVwSRU7a3YvwhTxhzg/qld+eTZ79WMpFhaJ
s379MAuDK0M6roOQo3QKtIMkC7bYt1ShsjiFkFtKgNYLO+9e0JEA7UnS3kw9GQfCMdbJ0EGM9IKG
9CMepOcblgNL3qic6Ae3qrpDG6p4Gb/krRTKm5SyDyCsW2h4Nk/PxvpaXrJI46cC3pwH8G8xo7gj
65m/Yag5s9Yfaa1jDetFg78Jt2S64v9+M54n/qo60f9nXto4AYSMW87O/1fSvsU4QDbge5QgIgtc
H/bqfVfsl8ezWAiL6+5XzV+u7PwnH+r2toZSamKUO5gE3Kcaop3jhOpjpDYV67J2vTJPO36zv86l
miVS+liGTptUR/o8ueEiGVyoUU8CQxKRkGmlMOyfxBsdWMKUS/a5FcoHRKUJcLXOQRSHmKPcKCWj
XtWJ0f+4Ah9M3ep4dSmqHoP0UJhXEhEK8oCZCogzDpwR4pv1C0VS5hh3+bwTja+rhljEe4riQ5kC
AfJmpQPxxF4F8TPZ0v3mATGtYD/vfU74jS1tXDQWORtTzITsnlMQlw0xTbIn53iwRd8uCrBPhQ2M
JsNSHTPadJABDWjT5ypVQW/MsooFP+j2c6ABD12dZKwBSjnPB8rgpALr8/uSNSx5MD4SQXHBqP58
KqLGqWz9NH7ULr329vuCvUvRZU/NvD/eBaVzYTXAf+KPC4jsc0HdAWEyqTYNcEJrs810tehHl6uZ
NtlSrQKlK40WPJnn+AVFlPfbG5rPZx8c76/nZbG3zqwBvuP1sn4rH92BanL2Tys9fU/byUTa1nsa
/I/P2TGDcghQaYzvFc/hF2I1uJUbz9/Z5dxYFl4ZNZ+JA5uPGeRS6AebGrz9Ha2HGnwQ27/e2PCb
k9IQgDVACHVdC3kx5Zgx7bpOTvDol1lYUsqCKLmvdM4sLjNS1pqGv02whHcz7ts1rFR2XkckuzFh
uSC2JjQ2ZBxez5dHpalyDCoxH46/XMbh2p2MK0uUvKV65mPvTBh1DkjP5EsHJeEmayUy3ZsHjHcw
1jWzrUOtK4eFIaPVLjX7MMHX+WCRY03CmTTZ+0dJdH61S02ZvXGe7uY+thhq8Ijk9j5cQsq6wRl6
WtvBuOD0my/fmLpyjvKy2MHPjIup4a1n/j+KSFMPLk/F9wqGzd/YIVxGxPSTnBVWue7PeM+I/56W
/Tj9r+pGpKCTPS6q7oT8WPMWNaE8snFZSa/SYHha1yczOw8TDErZ6CpeF60gqqIb4mYVYrkcEotb
Y1/4wQzfQ28247QRhONK1jQAxgm0w9IEWWXqnYf0RJX+UZtHu9bjeEA7tmEvSiaeuz/upCtsxTpo
pagfUfHOHuY1IzFtN5iTfs4c0AKz1CCuIv30+4ytsdd4HQWdyJlWfD8bHe93AumfVC6a05mYEYK3
fYkoC9dDA+xo4HulyYr5XQDzD5sYciBfLcnoXRMl6kgXhNpt1Yk7oYcutP9v7fyGWx0P8NCuREGI
Z7RU6Su0xRSfvnTr9F4FR/o4RVMOL32r4L9M1P9boJuumv9hKepXCTumVVTktyajoLEEl6Wzo+yK
qREzWkf63yjj1EAT4SOYZT1U9Tsv7EW5dSoRIOUpSh8kQdKlJcVbmRNs4Rl1LUif1ZbzyW5JnMMH
xFrJcIAJG4/ceK30TUEj0CowbXumrXL40lJ5t7RTpe5VpebR4Tt6OvXtk7Zlaqci0E0y0085MyMf
AxynSI3FG7M/c2QzHJSwmquxM9Md7hqyEjh7pZvKAsMfukAJZzav6qlfLXvrRKY5Y6a2eXYIXfgT
0E6P4lbQAfqM8G15eYfaZuZIQ71l/CvxtTSLTst7MRyG1cIAT0vjVYn9dEI+ooyXn8vDt/NG2NV+
mT/tckI3ufyxn1KdxDzNavXcUQVgxuxQGs8GuG9Ryvj6mXS6f1Oe/M0ZTBaG9pfiIgiER+O/nxxD
JW/ha6Tm90jrRv4CrETaReAivmONUsfougpSOzYkGUcaoOjQvC+zAFUTayAIIe11nKGDllsCylTI
yZPVfQFzYl8NO6O59dKjZL015QeOkf3M6vZGTs8VEQhC4ClnbcHiLJGB7OEpcx5aj27X41DCVAWZ
xOVSqIY1Y2pNvhbv/PZuFmRh6ZG1ypXjxgnsTdayyJZrNE5yn4rKEfhHykbRQ/Z1slWw9CjCDY+l
OYtUCZj5CjhVhl5w6GCcyBBQSQy86GaUpZLY0cFonJfwrMr78wzHyCcMo0wTxVP06PjEnGykCaMw
nsvgzHdXLtl1DrPfn8g1pPlLBe9K5g+cM4DaIR32vRdlfVu0+oMG31NgUZEsYhJ2YUKwXsYnjEUb
rahxdF8h5MiW4UYycsFRe3wVuIQRnhqG9k9cDnd5qXOdiUdWX0xD1m0a+8MetQXZ8N37emVHc0lF
4jhFTB34J8bOaIzhhyp2HRpZUWFnRVIfYf0RDpx4bBQOebjJlTm07iE2JBSyOYFcdkSOedKbabTd
u9WXCwgyjkTtWP93QVJjDrsgdu5A65VSQ4yX8KY7GN2yG91a/7p3aVPFmnmeDUkS5njix9+0pN0f
CECsgbJ2x0LP4KWdUa1lRuy4oT6qHaNgzvfUXbt+K8sOLe9p4C/HUBO8vi87rfC06tmcGKfCjWiz
BvE6/h07dMfnvERf2i0GAAbT2Nbnx++iU4EXM/otCSRBI2shMAgm7xyArnOPbDnqiNoPKpL8RXqg
7TmbvNLZWZrIUjvSz4VKlFIfe2x6H1jRV+4fVFB9bO5h9AlyTKaw6nYSxSFmHS2mfXuYUgjwd8jD
bQsOjeIcESw6ZrXffBWzPnRbPPU63jQqNEt+rArV/DtavxxMnUlUo8/u4z9b8oqxYRvt+J93Te4p
tlZ9jDi4mI9qR45EpqX0gpvY4uHjlpRKMyFsudxnPGp/p9NFPKqIH5eAUnAD/1QQg8xj4GathxNg
x6DOsrBihwYrsx50Mm6qfVCx4QMFxAg1ZESbYc8rz9DqAxMA1RU2PlpB7B2/eaqqTjLR5YJYnIl3
WDSFF+ajZMUsPKUr2+pDVDBM0JAh1XlfNN5Kg73zwKU/jKymWM0TPaXFWrc69hD/Ctgppg6Nh3k/
/WkJ41LPOXZ+cyYNFLIg6LpuNI9VvJxbtMZRKQ5Si7R0ZdMHNLI89kJU3JH6vLUoOcECF386Ry2H
MBG8hI31GFoArqDbpyMe68FZhjoNb970O65fLrq9vL917AG5qTULq5QdVExZygUfvUS8gZAzmqPZ
BLvNVYSf+BYKcE5ZE4kyGeV+yJGLwBESnfXvFZxo8ulqMS9GRdzWhjBY9Ru9Hw4lVR6QmPBf9n/4
TcNJ548LYFddgV9h+KCLX+R4WhMBD05G8Jpk509k5TkojWfYD1UMTPrIjgDTQauQDM0mLjGVLrmI
cvxQyzQI050OxkUhYgImiNQhVLm/OOYY06WB3vEQnxELcCofgHpEx1zWc2y8hiqUUh44wcAaYNuT
COvJD5665T8O9hmejPthx8M/H/oeO/RgZhJ/ZzJykH5V+u55iR5wCk6XgVDtCUmgoyIhZvHpgL0u
0AekUzwFIyk/myU5Gw+c6wPPY67Y2jaPRCN1VEnfNRJvBocQbYB8b7PAynjjA+ODORcDL6qj6k3x
0RPHDGoCF7nQ5gHyU800OjwO5vu8woUmsPEgkonHWSlm9us41bFBfdqDzD0HYdFIIqb3AnvOx5VZ
6Ny6bwIHfAzAkxvnrFgwoU/UE4xGErY+OE7G9G4Hy59NuodV3mttXr8lD4szrxVM0MP5Xq49bUuO
RX6jPrncIE6Zjm++Ewu2cRX2DIy48JSSTqRCU3bVLbQPvmYQddww2b7paLBEoyGEXeAASVS3PCHv
+UhAK4+FyO2wvfmIrYMbfL0/WlaGVuIOAYj3pZM3Zemo0/LlGoEM/JMIJwpYzjUiJ/nuhirIqXpf
pvUGKxtFZ9kkdHBP8Zq+1CrIIJolfOPZ6JgtoajGaJgAWa9Obek2A/dkZsgI6Pan1OF2BkJEYJXj
tu61IHMGlvSIW1h6YjWnfIbxGWmoz6iZFbZFN8WLmAmuUN4QzLThTVmb063iz6tYhmSj6cvw+fib
m9lgvFTIb0nAQdt3TWm4bFx/8JPJZj/2lRx8J1mAwJj/Kj8nJ4lCsSC41RfkYQHnwbqZXU7lEuy/
TpUtwNrUJn+ajT63X014VNTUpodJu76+40raHE+GMtsc8ArBziHvWcG5IH/Ea62HmCuV9LY4l9dG
iSG6ohFK8P2696idreK2w0v9wSdzJXNPMbKEuBb2evMjlL0wzJQ4YWkADtBwOCXYCQ9rkHU54G0H
6zQNVr6ObyZ73VSQIQ0Rtsktrs5WOUtnLcntsIi0nHaS9xr8UzDEfislNdka7E7Zmn804EhWDaR1
+/b6VafxCfNzxF0dHnp56CdNn5AhLmGum9f7NFwUQpRp6WuvES5kX85OmM3S2rXS1NX0bSKaAwoA
0vFutiZSNphy1ELWs7mj0qqegmwZpkQoh7jwQAaJtoCCJFPA9RjHRuT0aj4Sb4XbmERT8g2l7ldf
osWhEPvLW4wZuG9StfmXGztkRv8Po7E06dlaZyt2kBz5UGL4gWPfFMkpHDU7iFHHo4kDG9e5yAOM
1g5zyHBXHAqdntLt82rS9Nm+TeUoxJ/1B4tMU5TVRuKsIIAOtrMcTsDuXMconHmc18JM/wDzPgjf
hnn2v+zlOjsRsn6z/UuKQm6zyCFVhNbVyWkj0NlYxkJyp+xAV5ZWTltqaYIMM4XyhnYmwLRFo6SO
+eV1w9jkLQn3BRdvRABRpGEWhwelHInIDlw3U458gIlxTH2C1eU+YMfx8DNmcBOcd2P8jc/aDB+8
+JBrFa52Gjd/Dm5PEAk+nqhQ4UNMn7dePT8uE9f9EPCQXdv3Iyg3ado7uL6fCcCqg+1euJM+MV7z
ZPiIKblUtSd/wQe7zToYno1LB0ujZld9+tR855zCJV21g5moQZfCB0BdnMyuPvFi40vbSOuZjaC4
QLGtqtCJtoBQJ67RDSMQe4uvyoRu7yVgxT+1Nqt8jscqIy4/ipqGLLAe2sZRiITwr3UNG1hTFsLO
HnpDSqtczTbQzuqMvlEeFBirTn1ssxN1s2B6Jqwh1QU9XJ0aGl80lxlFTaeIS2m89yNY7Q7Sh6np
3trQUMcZ7Zo4BeeYlJYP2sNqkoeEvAuzPULISn6cs0w0vj4IWPpA4MfRdiAGGxs7t1kOM5kuSjua
QN1X4S+6a5nHUlAKgQU8W1c2roYUCUu00zhujClG4/YS4XIF0h9oJ8dq5kwEeZz6lUXLMTvCkpv+
8whOdrxbLYk8BvWnAxZrimIgVlfRyww2q+OKRXH/0wWTzMwMgw0MfXuJhIS8C3o60mpDBeir8lX8
g9TbZlbG+4I+Oup+Ka5hFiMAYgj6ezvGvhdtlbJOkjHCMq8wR2sNaF7Lqre00hd+dWU/sBpBlfWz
Ijrfl3t2bLb3NVnS+LWGNGGkj994M6GHaWSZJhcQNJGsWpXdjGt/6+ruARZ0udKqndkWAdHjQWof
K6NgCITL6yqQdgXdWwVTlbzwsbN4miVg7JNhW1Sn9P4UN4qm8e+0ciE5fvQk4/Riuzhhp47mxm/h
ZZDOcJ4/arGgDzJpLG9zhqzoltlyKbpEBIQ9VVB41kbXp8KDfZ9xPgWU9Hni0bE5O5mvJzaEGgdg
XgzR2LDWJyVN7qxJYeZvzQ04d3wjiLpYCVBEU2EtLMU5idi5I16YKacXzNqShVQYYr1KYng+kZ9L
LB6K6IImEb81znKCcax/mGhVpypEgiyTeOfAJ40X8fBJ9+JiSh5vuK914jrz+Qmb9oXulxofbcWo
cQ8KacU41VC3t2MfmTPENORhrkWLBPt5gZNKbNHxRKT+ENOQ+WkaYejyX3XbIJAfgBS7VkHJoWmM
qcZvpzCS3uxQih2SCXeMt6MwHmk0/lH7ljmeBVJnnNA8G8LcV4655mTdsOWTtQd9Ev/Aa33dgcfY
nhk6iMx52RQ6sCTgNWPehRa60ay7d1sCSyTacKCxQyPgTb6t17hCe9/eogP+7i+KSENC1kauCHik
5Qdoc5VdR6TR1XnBnoUd+t2zxZPOY4yHOjBm2fjfgvUtG18DYJMMaCl2EjEJ9u5/4WMqU6+Y0Crk
5r48GZC8po1rZry9fs0kxvwl/BNob9Nf39555K0rLz9KDizvMSF4n3LhTulsZOz2jqS8a7mgtY0B
dtQ5JuGBk+k5Ft/HqZF7xRwxdlUXr/dDQhgYolPsw7gqlim5TzxlkttvqMI1eYhaeDzg8sYlhF/k
G8h3ATAw6rqlQExY7BwQFLSakyJNDdXo078954HhHs9q1lS9n+uetB3Z6gUIc0J2/ZWEFpAuoPze
7utqpZi9Dmk5jBY0Ae4LZicJGyqMcC8Fr9/qinIzHVgJ2qxR3bD9crPxGVsqV/at6BI7re6d/5ln
HQP7LftydEvEyq5hW1ocO7BZdWVg/FXnWDyB/5MJ1a0BIN27aT9aBiOZsK9M8+ghNMr3Yw6wKG/k
03kM/UCXSPrvxEIrvyPOSekRh6r+ycXT91R2pkjtKzCEnHgRTWsyVyz2NvNscxZtD0WffK/eR8/E
hoG58hqPh4s4y5A2OzEOJJ61QNVpcN76m2yHGY26tpk4xLnHDw73JnLdQoppqTh6Ml81ysnQAa5X
5PM2a4G3FLfxPFD9ehJVn+hHfj/GKG5Jum4Q+C9ni97TN59N+Yr4mTUN7b5RYUM1+74Slch4Hvr2
XxKencDzy/SffD3g/63NFNfkbhetS0pof+TxrZDwQRCgMnvWFv/S1cZfHpsN8eeHnOMf4ejoyJiu
+mVVldXa0svvspP/MeE03n44Pr4PJre4cAB/Urh/t8204s63mNEfdPpiuAQxkL7otUq5BG1e1KeN
y+vr2xGhaTLcHy+/tb+d3oDhiFIEUl5J6oAd3ItsFOtCKXBB7E5xdIruF2vpOMn7/9G8uy8oZFEa
H0Yt1h30b2GGIBET+vokwn+nvabVDL1LZWlk4oop8jjhZUYC90dSZPKAJOVf6tlB2zwS8eyW73pi
Is4N+428WMiFkMX+jFl3kTd9IWyeMX0Q6znZPjSYEfIISifwP10i77xvaI/cKM8dUeSsCxerqXLH
/ncWM/B81ncj9K1ZWTQKB9wWQuTbhgerc/C5mAu5OfKe4Rcc2ABzfbAAnn4yZ92T6krpARTN0Y08
4GT8BOoXRyf1APBBsXzJwjdt2OPMdZ3WnBkeJigJ0+bs6cpp/JacGZX6KzDcMinpEJHuG1MBIpXb
fFY2XiSVEwUwYgKivf4J3q6eC293ffOcFUscR0aFuk85u5rTXm8sJVcaQSMV8t5WLGOp+u3FK1y7
TpKjBzstEXLvhR0iTqcj5+wLLXsqT1QjAeW+lEy+TwOdjZ9DOa+YZKTAZguDdG1qJ/jYWCB38353
69x2eSftlgLywoyYf+K+CKP0a9p4S+ydmlOMD65BgkpgCIrqjIhdgr2b82PFhw1SZUONEcdycCOi
8v24UlJo6qso4N6Xmutu8qlVqJQPRc4Ssfsc4svPUlI/+HGkrg3fKz0AsWDEuOOjMOKmxaLEatx9
x+AA+vE2QQZMH7yQgwmX4Cxasg3nCfqdJYoFEASaxz6rduaMhLqJ51u1ZRYouGZ0UcZbn9v9G6Vc
aokFoURN4eKkp/HSdYNECPEBidPwx5sySOqRjwXcMqb1XhmsgUuLqfCoczA87vgimxtx0UvrJ0oi
FUwRJZ4gvKo2KCkcNavi4iUxphyMA2ZGjRmZdKeg9Or0yq1nWgsGZ7Bw6mVZIohOzwl1q5/CGS4X
dP+nC0xxGhMgKobegaN5zqW7HN8TSbAzLxsuD7pYdHsOL2kpagzHdWBpfLDpD3cO704sCRENCz7N
3Mx8w7BKsUFmX+VvrIS/4GjbmRTXea3cUpwV9hnPpXEkmB9nLWYWRn/7AlGlUTbtOX249a8fNoog
phv5BNHsTDjvgo0qlDg5+OqMF26f1v3b3V8xbYVrz5Wcg/bqkIbu1mljClgQkIskFmNtH0UL+0k4
ayOIDgjb2ecayixISQnMjr1BjBeKu7JijEaMdWjVdjPZyk3Pe/eKwukDpBaXmQux1QYn8ZoXmnmS
Vk+2beJ18RHFOWUih7f2KI8vrlR74+IDtQrn+Q+edfFaWYFqDWzGYct8+lu64cOxDeHtyYLjoayc
udXFvyAjHxjocqgJhrHZKqr5hTLfV7jUglnJ1ffCJ5BdLHGsuj8Ey/IxYDK+BEuS8cTtNoWArQN2
Dprfqp4GBruOyapqZL+Dt+7/Sypg049eyOc8nTIopX94P8oT21RXF0coa+eIaXQSIA81NrFELhUA
pdpvtwwxoXq7zAEur/4Xi1K7czu5RLnPOsG+pDHHVwoh2hVaSp9BbKPQ1Rg9Pn4yQcbuDfW8cnqh
6LSX8bxYLBCBFh/UaXo7XLbbx4PfFEx1asX9xw9+uITrCcWLhG9QH1z2B7jweMfk0MvkYBlu5puQ
PT5ejXjYXAHlI8bIR8QeyCJuqFN4NyESS3hEFgoRf02iYvM7wV69gQqZqGndkcQzILWMPF+bihCU
f7qMI7EYCH1hB+670TQ/9yCWQKfdsCrPzOuujkLdMCnkjnV/QQQUcqvaLybUWF6huqJgEFgDIWBH
E3A21L1oDateSWwG41T4XremUc9+FBjrg4aWioayXmMFfpCat3ZycDFqKi4+r2kA3DDw3eLGmV7w
ZLNrwIm+VVcZFYC0NSucsLhDZfoMr/UYLNZuFCHS9j9jkYcUtHfpQtNHf1reoCCmfaD09NPPXJZp
LrJPqQc69WXjrGvzHfws8ae19x7weG1Z1txwZlycVg75fII+MF2HRPCInAVXtd2i4KiacYmJd9YV
qrfzHsTgLU8CSKeTtV3dRyTIFZpJG7kXfs9NW49rQgAxlGj16Im2WtJ2CbFCZi9JWanXKnA5EY+p
tDxHxgxZRixR5jdE6MxfDhfnNfhqnC3JkgTutGQzUDq+AMBSBFupGheCjUr0gi0PNgN/l5YLrR7j
npWCfVSZWuSeq1tF1FtjqmensoFrxiAv5zWaF5oNtzDT9S2VLQ0YX9zK/ZHkADCt9++QlcmgBCY4
yWR4ALW0EPN9HC3cnMy936kABjN+Fk9/tcBCYT9snuu6RyHKNzgViQ0qPF/eu9sNlnOk8fPd+Mvq
fe4QReKS/LzEAZh5I5Qshgf/XPTQ5wcE8wTvJrpOuPoS4sn6NNAZH2lGoOEtZYVcgg5LO0tk3xhR
m+NSF2/gehGZPtL+DgUARb6E76KvZ+jqLZcoQTL6afS5TAg0Yhj+8OoV7Oz08dJN0nzU3Qu252dw
XrzzP3z53GZH/2MwcG6RSv8fmHZEEmyM9N+GuSa3eeLRJi7e3PWxwixOov7PYIwyoDdVSDix9XSN
Z1q2Ro++QwQZwplXd5NicBNUkA485SQzxxm4IWBTpzFYVlh8lu5PJiXOVAQHrPfxttoQdxH59fWq
wG0Py0IEqaKfU6G8+6ucLjPMXfy+73k3gv72vZjUyqsMuE5Q6AaKHw+ATCUcquFe7yUBjg6SA276
B8kOMVG/tWuKvpr9utDn5YEFy7T5zwJNGV/qm0IYQkj0fTFMWlf0vzYfGE8l9Pln/j1ZeMn65gPT
/pdtK+P8weCSWRHE2Let9lRHlHmgGP0lEhpzvZM1sBnpyTScfbLJuN1HwcWrVRRvVqn0NQpHO1N8
sedJwox6eQ13ZX9VV52XgsydtQfI46T7lTExlU+P1hOsHh6xrLcJdrYmEKqhG+208C+cUzxFQjfa
wJ6HcyU5HoJ4WHXOI0+onlWRi4oaBoGsEaX5oHbMK9A6n7yvDNR+mYPuNBO1ILplnggTHIxXpGOE
ux3XMYCLmFHUORCivJlX80fVH1N/XebISLamMXxDR45eRT9Xr62BembrrB+eQHKF0GTzcwbRgsxd
IxE1NKz1t2l1ifIrGfMutZgYASJJxoodLPr7meRajcMLhHjg3x4muxns/Uv5hZ/KYuEzGmdZT8vT
c0nbxMTyyR2MGLcSFCZodfCPVupFZRrEfcmz7g2uD4goy3PEfVCimLJJaDnAz2Hva9ujeZuaI1lb
lEORWbFcyvsoW/akUIlx3TvYO6wP813FqjJBuM+RXnQvN0UiHirS5jjkD0SondxSfj0Xu+O4uJEx
2diSdorlpyjdXtQ2Qg4Mvsa+F2r+3293dFpllvNDYoMCyv6uooe1OH+7fF14a9CsTsF/fTFWiGoN
Bv7NM+xhVRKGglLUkzHoTO27EUAqMMGOPkOasv5pBvBw86mXH6ktW6t2gFZr59U78U4uVEOC+U07
70mpxtBukrj3UdOH60Dz51L8oOXyx8DYz+WhVOtzHTsuxHvWWd+dWM4infjpa5sfsEFsZbm10cQd
FMyq6YazhzhzWDye1TGwvZngKIeZVNkfCBchljtqgexomkpJltl+UGb1sGqZsc84D7dFaDnZ+xCg
NsmgTcCEKQypGBA0la0SgVRQ/1M4LHm4I1m6Iq/nzWNvy2znXUCOFNlBdNJp5OrVRagGo7CgQbAs
gPP/tgVnI9vGPCh7rY6K1CAO33phF5fDjDFgkuvnd6WcpI5Se7aDuai0JzOLTS6y/KMpGTCEs3Ao
SL4Jk/MiIpVCj22XpzGe3Ni92v4NNFgx2oxXf/ahlQj2g3S7UtK9wtIJdGQQa1fxWBD3CJFYh0nd
WOU+1yddO/VUvMHnk+SdTBJd0rPS7EfMVzIUo7a33r31c3M1jOBMeSFTP2OHy/TDu7XO6e2cWiI0
V43L2zU41UPpQ7wSI99C+7DDsVnNT/swn3UrnBDfSW07cENUjE9N43XjuX33KiY3rDZOrq1GjU09
fDvkJuFt1PLWEUbDoE45qIFxJ30uYT4U3VY8yloAk5nrKj3S3M/Ea+PAccR6oc7Tk53R99rXC5JA
LKqzQ3LuO5UpeILnlUU2vgKdpQzM2C9rvH5SHQs55Sn/5dCPFjqAcfcHhfTgQRD4b0xYNg7xwmzS
7oB+bKKT6C36BfUnrppTYfCgqatjcF/g7+yEf4S/Ng2aZE3Tjbik087L7qnt1NyfX9fMb/+5cNYD
Ggb5/ApJ80g70M5pGLjVY62LK7/Ua9hCtDUmdm4SZsVERTjFdM2BqQbDT0IE09X6uv6iipGdjVR8
bkZUHu+mkTlM3iEKSeRd8qDkj/RW4cRSrqRzVCUNXfu93Kl3Harml1GQenl8xtTlhrJ7KbxLUVkq
p+uTH/KzAsOYx/Rc7Mxi7VJygrhmIzww6fbabZsbgAgUeYgEWMzJlJ3H8nwftuM5gkKEMYcEIfm2
K+mmEgOHfig547zJhTDgpMJHGkiUlyU5xGsG4lTR/dha2bSptmuAUg//Egnd5poF9meOy/bzF+iu
pEHzTZIracjRTT6ZBazb7jPyQxFaCzDRQvNMwUmu/jZyib7OZ8303DEq/WYTmFjh0QwBPAFRB03Z
lSFUJBoSd6MsGWcwNc3qUskqbZE9yvGEC2XDJJ1Cc76d3SuU5Ccb1sSKBl2jsSzR5u7J/Ul9SoDW
LAX28CbLhmp5eFK1+CFoJM7GU4f6UyqBTzkJhP7vXi6uTEN5szfWrTw6QRrEzOjqdlPJkKOis1VX
0bQa+0lyxYeBzaxmCK2Sgv8KCE6ZyhkyWBl1v50emzWD6Ky7/UfScmBiapNvFQ0say4Y9qQuhYhK
1wAwPjeBY3lACHWOOXBspR62EOc9+PSwDvjcJt6zklJBEbeaRc4OsvhI9IoMpgWLql2rInOejoFD
OUlgYkt9hqO+Nw6DSwEGHeK7JzqcCLHoKW3r+TMFaKpg2Kf5OeuTQDJc6zlQY6aHQCbrpPmszEQx
LJbV/kc2EdMT9F8mXqH4Xw4tK1KNNRCx2dwxxkWgSrbu3P323V7RdX/CIL7YbTGDV5La7kwKDTXo
+y7Ks2pKD+kAdCWQtUn8u0sDFzf2i0qIba4lBwv4lGEeA30WTGv4WaEI9ZRCAJJn1Q6z1SNbvipX
5dp0bfyIMFkq46p47IFBnd1twigsywfv47LJjNX7mYbgxmm5nB8wp0NiaqX6KiVdyMebLUhs+TqH
Ag+FED0cha66EQ70hkfqRYs4Rn3cYXJcdhkIAXyIPYZMla5rPwyZISsDUOJZBDBK9L2sd3NPo1CE
b8zi+VGeIl/MFCV/V9vkfP77V+4KLqRoZnC445YXF6ob8wqgjFuW8pDUo8hdPD4LYLhVNdeyeQ/I
IGjP95yoCphUU1pPZScEnhOP1emTSIXfE+sfYWDe3DNYDppCCwXNqeXQZlvYKjdfNOdvYPSttDTM
IEvjleMBG6aStyAyO3q/0BrZ2MRDYKt3Sk1lOnSYBgqE9xeUcvEfSiQXYrEhioEf90MeS4LhPH+i
jI3dVm6jHgZdqz8KPAKuseonePIAtwwsNOolvwODpLMhj0ftX680rheyuxmLPx7rE5sQ9cmKesVY
Rx989vK/ZiepT+tYJfri94FH7xgUsmHFCxfS8XQ1Lvq+9MkDN6wbrNS18qtW6g8NORM2u6vi27JD
T0SPIO8KIM1kAtnmfwc9Oo0ztkcEEo5BApXq0jQFP8YNGGStuAW4iA0Fns823mZK8VYdS76naDSh
PnD/2OiRZXv91XHCH+t5IZpPBrwA+2Yy0HGxgnDgt3UHfFfuZrw0FxouyJVNXXx4u5it8NeUEY6i
zdjxFqiMfhj1yBx1lcTQzW02GfOKbo+JhjY6iOjG2LFQd/8iAfPuok8MzPerJZEMgpV8M1tV60Yq
e2YFuWO2BpTNTKlaywtkjx8zNpgyFz9CnDfNb6s8vXqDUFNVJYthFnAUT6k+vkeeQFs02sIkrodD
Em9zVZL+qFLwh7Egk61awl7Rz+nuCVpab3dyzSZK3K4ZUGORQ8biiAlVq820rxywQKSlKHduxBZd
zf7itMV7RcLNzNX5tiFcjww3xX4mlRGxxDgUdY7XNtxvh+Mu/+aRXcVxJgeXte8ebd1f1gq0l5+h
BfWDRI9THp6IFoBTwlcpUUhsz0yZJkUA6CWg80UaQAtKSA1/O84Yob4kS9miKaKcINlWMOphsxBX
R+b+50N5eNBnNOlPvzi3fED0aY+uEW0iF4vWU22trl3QM0sUcqBlaxhNn8cXIGo2EBa8ZZqtL7Id
JnXIdpV2t3WkjBpl/rubjQ3MJMLo/iltMyZ75SWInqqjzdYUkXkVOF34i8nJmAZsv0El4DW309yB
HfmwM0hHbq7p8et1AiOvasJGbwclKFmruN8uB5Lm4xrAPKVpCLBqqhrDo+2Bn7UZwmA00pDEHsPZ
ZwOmCmAvC246QuB+1QOlVMZmaIUENVf9TR0NXG35Je5Z2B38fJ7ewi1ZPAgy4JmpYG8pXrt7ve1E
Yzxd87pFmmXeXMurVTx6cfIRUM9o4/L2NV369gJNu89t+6oV6RGPF6FkN2XqVKno3+v4/53RyX2D
/SPZ0ZiLuW223DwW3FhCTioPcGGX4vlrnA7FWdS85+kc7Ibdyd0AGdPAUOGhzLgawzXv9Wi3AQJZ
U/sHJfvEuSuF9MFf1uWmM+ibpA0L8C11yggJO6kP1GkgoM/W+p+wFxHMZccFBYN880o7Ecmpqyym
Wb72Pqdv5bNaurMAucmTKo6lj40Z+vtYXP2CQ/3lRv59oqPDT3eoF+pgEhmYZL4nfO5AfV3Uhzro
QIsEQGXpWVSYlJTx1DfGk3X23pr2INwGNLJPslsH8iNmVmzPKtDl8KEmahUQYWuRUUmAVTTbND/J
iWFSTFA6mOWkc0oEvqa7U7Bjh84ocMXrzcmwiN5U9EWhjtLwG0vZwCjyZIHjuMDoa/4UO7z82b1I
wHX4PCApJ0Cu42/EXSjj6b7eOHNES/+w6klkLHoKeLlileQyG5i1T7yvRNId26t3Vz/WEIXUEkPz
asAX7A3sR745p5BQXOoL61ebiQH0zg8MsuGH/7D0F2hlHdXCZHOR4SIR79YYh1KnFpu2pc+2V7YT
30y8Yk7MGrWaiQXXeb07JEJXVzeG4AmqLkXc3nBfD0Q5UxFy+JFjuhU7wy1+ocJAWTeIIpOWwBrM
JHNl6hVtStM10P7nFtlGE4pzNK9Tkn/7WEY9IwQA9AtN+JJ+ld4cv/05uGzlTejdjEcZaJp1ufcO
ETmd30Flq7Eo5y3rjoFV8tmP3UlkFFv+a1LkvWdoL10iwgB2QyN2NI3ffuADoqN2NRpi0WHQPKDp
zGNM04Zwk1bBhooIuOrTkSv+mQi/VAm9mLJeuPjQRTbx7v71/uoP8VWK4+CC24Srui39xP2lfBxw
M4V5Y/F/BCWnCo888rVBpP64GMht0GjwsFbpc53aGCgeeCPmwkHlGjNF2AGegM9A8orWx8O7MUWl
wTtQKeAbnPICYwm+xSCsjCYYmF12u27yIlcG4sqLy/jGen2HHfQCrlHkR6nLsBJACCHUyQZcEuWP
8UKJuUOWCfofSjfY50G+GlBQH4Fm/jZNItQhumMUCUqZxhh5GDtqARY6iqSh5rn+paVHGJtORHOt
9eUzOLJOSU/S2XuMgkD3Q2IQJusvwNsib8K5OG6XRvvywxbOvET5O32K8v1PJH63IOixF/brjcfN
xFhuNmyAtj2zW47B9tOg+oRUrqElPtE3HvzxY3ecwJs8w2s1N/WaPFLaiIhsu8CX68GueLiGkPs1
5lijDsGGSu/pCtjC/NSEeqlVoSoY7Lan/bToqWua9K74n6P/yeM7SAeQ0pheDvgu5qHjLrfOZI6F
5x+Co7Wze00iqLSED1IYPEiHIssNxjvYP5JBWDCwWIU34Q8vCCoeBjoASy4ktmDS14bK+9Ju6c+5
vhEw82g3b13aZzpvV65+m5BnG2mhhFmGOIlq6j0I5GceXfN7yib290gD+gPBN8l6+aENCQDfQyu8
sdOLPe7PvGF7jX9ASzjtFXxPP6oPI4yjDIB3iZBCpxHGRuG7Mf5QIYKcrXJaTTrIPZqzwYGv0E/i
2RQ/odWdGJIDQ/L58uX2lfOkM3dh9q7MU/2ZNzHscfsx3mBrTRhki97SgPz23ZRItX3wa1ZuG4wT
9mupBY1kFXkraqW0enhKnrNZ5MTnujMlEHzSPjm7Xbfl/z3fGgKXj3D7S/HPU260Y33Jfib2jqrE
qoN4psNyiFL1VnLVPlSvFVwb2ocdxl3fLHvKqXkDb2dZGhRXq9yrGbfVZjYWz4DhXbItXvOBPPNl
nMMHUvfTUYJiCE0xB6SCnzR9bmgX3FPKr/evHeBchxEVmrg7pK2x+RmRCszOIZrCpG4h+hYcQ7jH
S+zhUCQDkyhkecFXoSo3WuiqIEkUo/+sEBZ8Y3Jp1oVC71PWJ6/njHhyGkxtlaBmgwbhtL1YLDtP
ukS9P15BOWQujLH+oNaNiE05Gsj9wZmen9DGPjgxFl80hCXb295eWvJWaHiFNinVZQJS8RUNpqWM
sTgjraUwQIvkT6mrcyMi1U+uKtTAot3yd8cpoFYa2bAkGSz+PQomcVvDbUHHmoPg3mdO0y5wMUd0
qF7jrIltL4PEooUw38seF6Bb3XhPupMTKlgzMd77UPrUxzhZf/vAQ8B7c5TnB11v+Q67u+Rq4XX6
F0B1iEafUKHIX2yvsi8GeKnlOV8cBalDktz1BD7TXZGlQMlq7CN6YTeJGZRD+Kdnakpdn8jEhAfr
rszQUXPiQm3oVykvGDw2kHO7qOr+wr4c27nOWCicMT2KKjr9W8GHIjrwgpX9ZRowZG4f2Onl3lYh
x0pX72CCwZDe1yC8WxaJ0Np5dg8Mhkty/7g4ZZkpYh0HNf0X7tHj1jZfi7ZkBliq0nz11x0uzzpe
reN7KQ0/R0dtsrsn6j3H+nXsTok80bBTSsV6D0dg76n3Ojf/F2KARhxwjsG+74oDTHBell8LW9rj
6TCIRW7SFV0SJifUK+0Tq3jVeSaQ7TuYF7uGZACyR/5gbNfKfFOKiCnbuNMCoCEg4aPgQ/UzlrX3
ZcsTp6W3SeYfP2aH78oDywTTQHOlDA5YSG4mxHvxqzW6Ze0p8gOBAgxS5KUETi8sSynrvEUGvE+L
63/E83hS2kgzKZmdQTjNIP/RRBsVaNID+cf+NfTApGtob20W3H226MiWdfcSGELZ/JjnA5MTlYpp
dkObNBesg66FAHpeJzeLV9SZbTu0xo++RgQdw9IGagaNRGr++IEQKVytWz7yOW1gX5rcyRoZNTXG
zVSykMgGhUZ5Imtm6sUnhYq+M/qlueOIbWfw12gbKJZC/pIZjkPLe4dX3YPJPg+C0VAhIMhk8A5j
n+jRKfXKM6QzXMhnAv2MzUIEwf0fQB/4pwRJ+cZPOlmzSTSJW8x5YIFctQLOSppL/2kz1PhzrSmm
WdyVyLqV/w4nSfeFB9QpqJ/+YewuXMbqMkDtXJegSkjSSRglJpSOQ0DFCbX1ghSz0eEg6IaKI4Ze
dT69Vw1jfEWQjwCOG3zBegSKwuGw2t4gLm8+gdijhRTT3IBqdF7iReJYRCt2QS73O1qlz+jjLPLf
Po9S1WVS8TAaVKEsw8cQO0RVGWUydUbTAeE5xBmE1rjx78F75u5YDnjbhMlAhAiIwJaFgxGVS7DJ
aETW1BQexN8YJFFm6wklo2F2PYUWkw4V9FAS/tw3KoDe0+y198gi/RmWr4Vl/sWiZWmMrnUeyfXC
p3VXXGr8A4D9WKmPsc8MnfbryHv0l1xCi7FiuLmS3tVYi57f/Gz5Jv8NCFt3vO9FyVwdWVT3jjtx
24Or1VSaNzM5af1eJQAIguPEutWibGjkSEHrde2G1aJ5llz8JDOfDGsFuDzo57DjWYptOIQfS1fn
GbF+bQ6H2BtNUi1MrDurESgCrB2FVj/LaN6k2uY2Iz5lwNd+2TNlfvIfzpG61k+MqSxQOOK1UPUu
jXgKPedLiZzPCpSQxz0/3ZOXOIxfyAbgPfbMYEsjCTzlQnbm66tVhLQGm4ZiyT2mX9HAgvBUZbfi
4RLv5W84EODytxM4Mdvsl3A6bS1pO14RrYUpxke6xFyKfv/Kgy7GKE0sXIRSeuSXZ79SqelZJYPy
bHeOknTyC1Qk1niKJfJJc4PKLFDDrFHciVOG7ZUjNZ2exEdgLCgrEA11kwl5t0v92ccIbymEcWTc
RierHroh4KGaMIKdUTDeeOeveu/7gcYPkayqR4nyQeeWFcKp79kVsLFi79L6nE43aQcyQAPlxBee
2GAMK3R8uVeQPi4LmPHIj0hoVaTRNGVsKcKwdfftioWOqIM1qf0Qv03cN9qoL4OWtsOoM7KsvtDp
TtpngB/76fX29e/ucD18cTkVnqN4azhr5QUGxQZJYYIZt42edgzOwjE6tjDTjCPOVYTEE9Li535+
DGEwHHvNVIlxOCwi/WASRTK1gHfXOsUCfSAbHv94h2mBWzA4xQaqXEXcrEIvN0M30ugKBpRe81yt
S7dZnjL4OmhQKEy3SfZxtADfaPcO3CF7SYbeYamyLLuML0YyUYsgI2TP3uqTLiXlR0L9a5RRYCXh
c6iSKdjUywBC2KyUBxXAylBbxNrSU+YUQ2BybahXasxZd2J0gXEEcLjOwdjIUwFywNCoYYQYSRNC
onfbHTib+46d0yVjomVUvxtU7AO+y2mmVh22a1Bgb7c9GCJhDIGg+gYP0fcrl21FIR3ru9l5JOL6
rRiqdc6PFk1vCxDPA6kMxKylyefprWQc1ZadQMttmtsFPlEuiF1Ms5fAGnjvu2U7iStzSQ4M/8oN
qX1Jmu5OXtA+IffHd7Dj1j2+m423UMgZ/g89RM3YzFavs/c+7BFRLxtS/Y3oowcIXBtYbHsxSr+l
0fwwjJfnslu3zZu49N38SN6d537KLbFGtmpf6/XCzACthYro1J7DMdBWkKD0af/FWTQZHodZXeWt
Y+X/AB+ktUikop6h5Bm2l4wrS8GU822GvwQKgXjQabgD1/zhHLntiTof9pF1FbS5G8rFMwU9+o4h
kYIdyAB+ROId2pXXFVT4qCaLadrbUU8Q4PVfi8sVb+zhkHyOBdZDVtgBlppZELbq0uAen9cOPvhn
VcZ6T5xlCPOqW66YCIDKe9fnTbq0CCQBxwgNiFvjBLdL71iQEk9rBmgjhY6ZieivBHzjaXiDELm+
XtAMaU5jMxh0mpZMoStwplmFYqkTxf48xEFwiBnCZyuxaYFjlKC1G/DLZjYXCpl/gGrVsz2CPDcN
a2yfYY1mOeO+TUVKJ9tK+g5UYqe2Awc3EC0B1mmd5ioNY7eu6OoFGMW9cLUjRZiKh8gnBkm2pXe8
VoVECvef05kB/SV9YNGYYmwx1CMNL13McLxWG269H0xxNBRxPZ+VJne28WFj6aMeNyMtSlhqNHPX
XqITqiHSJeYZdQurEMwiI007acxglqYzs0fjCzmAQ0L07AwrEv+Y2nDeOKUjDCrq/d9mR8FBX6Ig
oqkArfG6whZ8dIcHfCO117vDMuPUmFwCwv376moDzOmgb1+JpbVFWezGJYv88SBiAn1BoHgB44dG
3BXcezfxYekaMUfrNlr5LKls0yChvjpq5CaI5V2gfodbpipOeKkSdfI+73xNxagm7+42Mbd4muOI
5yikr9oqXzvz5HXWOzj3tE3G4oY6fxEvzcPaChbM+cjCpRDokyvhNZy1cdyx6OOs3vh5I0PTKxap
9Wsa1JXbEAOhBE+q6tbNszlRCiHcC4x87ihn2IEFB43KCKNk8PSkCpcarkL53nSmJ/b/tcLLJS+X
Wl+XLPg7XHNbIikRRzvR99KdZpwWUfFSPugWfM00QbqRzsraLtzBMSfW/jnFdCr8sejOL5AEfHIy
YWCcuuMRG/tejuH4ZurHgnEs5Ye3cHD14BCX5axsLo3Bzu/qhMSQEKM4oZCtitLqRfoP4UZHxDDM
G9VKyE/4dGpkgopu6mW4s6wkMt+gDJ3laTamkRtflBKV88qkLr099j4EanoSgiiXUhMBTaqKiTcD
P0xSuleAcwze1h5/tBIIA1X/rCIPWWKpBqYNbpNEZrafitlqrBUtQjQ9klB8Pt8QH2iiqcsrRCE2
znTez0nkN9MTXg5NTpwvKPNE3E1aJeoqYEPgeCZRlDyE9akoSBWNoA8fZsnI1p6QwxVsUI+bclFL
m3gXxaDZPObXMxU7qnuTdQ2Y4VbCs1D/o4N2CgoccqQ0Gp3u2hkKXAEAudR6CPmWTGhkkWTbOQhY
iAgzGCL1CO7jn/Y2RECmpA6XHVG40phzBUwE789/Cihn3kGCpV7m7HtKOvGBxovUiz9mhSZPgpJw
mmyHG3AcGsheOSS9MNeAOxUwqOzb90dgKHNKUW5LzoMQ1exShTQ6Ut6k5EtMKa12uhV1KlWUHKDH
VsoVtjR8kHDgtgwj2KCXXPo/F5cBmwl+ZmE2FByzBwa6pVX8OSv7yMDUr0yo2k0RzOSs8p8Bq4Em
b7GALbUII1HFXBrIs2wA4CZpFcOdhiG7jJz6I6lFDFM6LfjgmdbwTbf2pej4WcWNlfPM/2AzoTD0
K7KKNVuS6ZMy+yl6Mk8vvAiJh3tB4CZiCg1ryMrccAkT/l9EV1ionae/yFjLVNw+estyXvQTLM7M
saHy6yEK6I5+huwYm7XgfxUEFDQv7PV8HoBrLHtIVpuNF97CFfF+FzmnnEcZCTEflMiBB8K6SujE
sIWXXe5GSLjBFKG5S/k7q95Q/FtAjCB21iqJ/MGivlCJMWXSvjjul//YEeFfNaqPkBjWY0eW6t3O
2K9HDX3xl762GVWpXC1FpFxlIsc4ZbuoC1PEJEZ8Sd6sKbMUb2btZojR1ONfTC40/ZHLgvOhaHj6
RYV0Yn5FcZv9aB/sIrv0Atn66Ry54jH5UMw0TwEAEbGEeYvUl5g5M6ZEY4ruOucaZiwnv+lcOXdN
UNz89u6dJESaa7gHKqF2ChtCNMe/FuKclHXZ8HNTm/4OeycLx+tlMqtQ8jihY4FlhVa/7L+cBUwE
1UI3WMh+i7sYp74GtmYENUF2vLjw5SUw6NYQLlcNb03pQgsa+/gbh2BZwrj0G2lGxUEqeV+BGXEk
SkxBpLEWMpcEm8ZJ/5wHp4H+zUVZU2NyKIhD1+gJZ0hk6uZisCywdvwuAaBXKDPhOLh4HCdXHLf/
QWAnSuLfgs2ptMeYiguf8b1hbGBVodKZE3vgfxZpEF+P2ooBO/El/CKhfDFWN1J8x2YHQ/YH9Oaf
JesqswPyE5tIDx/RkPmIDgEFX/yrGzrUtv3NGOW67Lem74aiJSBVl9vUpcU6hM25KfWRMgjieaWV
jHwy6XHnqPQhIh3bF8n/XxE3wOYutWzONsLDRNtkgD39SdTopaez8vPOVoRs59UAAtgYE+tBFSqE
GXlqVisT7gR80mL8VqXHeM32HQ9w9+sjAqHhxNxj2le5gCd0VY2h0xDtxRnozF80hT3qyo3u6GTT
i+Z5leb9EhQ6FG+JLHV7JYmIqfmGBFPc4bLySPdEuBcbBXLM7tZVe0c9Nm6JYD0fDbZoQv7Dz6u7
BRtV+78JMcKLnBU048DNqAO81olEY+qardqgmjPOhFO3KyyAFThQRPH06q8IjPSmUeC33NuPeZf7
TSuhANppK3psFV27TP1nGtpO6S1K2q0OTOCWNHkt3+zcrSf20p88BALlLf7cfAJJBXPB+mDyjDs3
cDolrmAw0l8wa09/pT/5uUOTESgxtmH4fvHKUkxORxDoKpKNxp+caa/QMQu5iAeWfrfPHSsK6HqP
RkKwnjPhc2618/Dn+K7rzxZFlxR8SI4Xl9FLdTD5xv9HJcvUTQv35NODzYv0G4dWnOHz7PeLyWpU
pGWi+rnH2Xc0fttnaitDImKmYrHaQIg0N+6FdZQiq5KSX5IzvzW8NAnOwCQ9T3IUycSJh5EAIASE
JISBkEp+rl/ewVsuFGR0Mx1zuDcNSFPAMJgkaXPILfoueWfulTGlZu05XnYWvXtQ33apuLmLT7Ir
JxYeVLeqZ3MpTs9mDsgDgKfZB1oZeFclcRbQGWb11lOBfO9BxU/8gYFtwpo+rtXJ4zC8rRlXsn4i
aXKkPs53vmUK7cgmt8aG/+SHVS4v9R7iAA63/IOmHLKe9mQSau8MD1HOdnjwO05e0Tr7n3TwdbY2
40MO9yl0J+59EM8K+8MLgXItenLP+TFs5fruzPBP6XG+BBSnbeyRwcDICjD+vWhcKPVCfSQCXr2d
9nbbwlpa26mLQ6YLDhq0wurxwRoQhKihESBFgUGREr+I3gD9g0LNCAmiuPiAdT7VaS2Us1NjUY44
xOJLfuer/1CX6v07F/uegcvHtlvU+3+dUXIIdRFn0IK9oiNmlNK5FJyH5MFYQf1LwE0w/WnujI/P
LRbGR+FDldPxGtmat1cJDlN4Zw5sItOY0yt7FEFmXhWwWb0xFBjOlKbMdEqU+4awCwh1RtAzoLPH
ySnBseA0r8LumUgfJhG4ld0zHISmESOUkfOKvEzVVVSZ6hXpmMqYl9q/9iOkMdiiKKvJym4/hWfZ
LntKcRPYBSpvrG407+ZqWN2gXzF4uRw5a673zAOUgTN3OEyp/9/mOc5xzRjSd/GpPSG5W4BBLf8B
1IvWWdPTpSQDH41J001d92ufUV5QrVVZLN4ZYg7cZTOMMBr3Q3w6DZ4b17pHYSqvr7+LnMPw9jO3
uoOqpgoTnUDdf9uUIDq3dJU+mnVIbbV2hl7mVO2+L++9pD3+f0bsYPrWC3AbgEhvWgQ7dY2ZR7R6
9uga+85lebkpHN2rv4BF/7lqexMxUDV3AFZEHl7e5NasDb1QmxOmPHG3Kx5hSlbLaGvTGUVzThmy
C5PVHJ/QhiwQD6dG7wXMrvyPNerwSkzM4Cefle4876P5ae+xBcm0xHinfRMhBIT2JZF+ieEw3dXg
HZdUb28H0vIFsO0CMEfmgjkrtPS9w/uRxX0Wv60S00MOjGAohSrMPnFP9yeG8LZzXtJJcFeV4eJK
Cn0/L9ySLgyJ6ymjr1ZKx5uQ4SegAj866aHKvBCHqF6jQ9Gh0C5pdCoAB7LJvh9eeNA8vO4rx2N+
j7BZSVFmI+kSo4kYZZ49ziw73XUMvDYptdRwreZIPj6QxYoH2nVFWRgdkluTvhOWLoxdtt81n0WD
7wjkJuaLr9KwarMUSLVwNh5ZJnf2d3VB+E/LONAbJDAMPbXWPe1MfLvJT3a1qMYiyJihNlAnC9mz
bRxidLHvs5ErMXFOpTFs/oGetllARU/6BvI70aemqKS2CeSSsZaMETAaFI4XJ7VNY1hyV2sqjjNo
9YmNkgZNUSM6w1GsDD7RMjLWmK2XeE5jJTFMReWY6f4bHB1DpmKJTOmquKOJHh3F4qbxmIFYQomr
EQNqIO21lDue+o1Hhw5GZb+G+Su9IR8ZixwNWYgvWwXj/F3HrME0/WIN6+yl+Hz4CWfBnG6eufaj
gHVk4nxcDSqokC9zcqNsDwkMBJzRtWWfnMvlU0p34sKp4n7CKbIJlmC8hkMt2uOtY2Ry6bEHlIEC
UA6dKcXLJuA7peJeztQV1c8XV5KDE4QB9vZ7uGkI0TVZ21AEOybwnMqSPw/J0SskIUK0D8Ag9nWl
wkz6gF9AWYppKr1K1grryvdl4+M5vJBfMJ9Sldyw58HbEC3CdzNmpGyVVIO5j9Dp3/FQHYzoSlXO
MMXIbgoE+YlfMZQHakeopVZ7oJdsLa2Qd5Bkju0lcNTKlUVGf+Y7oInIZ5QE8Z238A0vrjiApEdy
jIlSDM0vnC/sp012kBMAXIrFEylVCGx5GLK+3Rv67vJV3ShzxvL7+d9ZpWiGyddyyEQTNKPjcdV8
H+HIFFqgfGpAvgyl3hg7siECL3y9zquGaKXvxDbLFxWP4gbSISTDkHxvsOKl4gBpGUyycVSJN7Ya
+NJb+MvHRmjCImt93CEmsDfdWORqBNT2d6FHWS1L3boGShap/11vT89EO00KMp5ggkqB0u2kgoUb
gpNn2MF+Ldc+jEPw4mzKPi76bJF1jwoIhGBzOQU1PxvFy7EnRvreQ9KVvsrTW2L6bH7cbFFT/hAv
ekTb6NvqOGi3jr+5lYaFzAmViINZo86Wqr+/BzzeobVJP8sCxHhGwbWoR8iFqqosVWZJuntTFMQt
HGJt8aOJn1E8CK67qepZrv0aRNvglHdmcCUCm/tpdXCdTDG5mXUwgcY8/skoJhLYRFIvVNX6P7xi
9mNY13vV+jX/c2Hmx3CILaQtSLApNAD0jDRdLZ3F4Wbile26vI6ehxYNx7kJweMG3V6hVV7cWiJ1
RZSxy6kQMge+3+pEHe66yTjxDGUCnO7NrP5zSRb//K+OXcJxkhtjE19nR/epUCDu48HqB5MsSrig
F8ZgY864UDKbB8zABwWgx5f8/ybuNmdbaJpsTRNp7S4JmLdVzdgeCt4JjSmHBdEt9cI1376ljQU3
Rsi8Pz4XgVUOcWpKgH/18p/+VPXYK5u6oSsXtg1GCZXJEQ0siY0ANaKmxtvnrgj2d8rKB86TsOZW
g+Ol2NXCPaloqoNkmbXOAX1MHnh20ptkso6ch2UcY/5hOLBF3yUQoE1EThn1zQXHF8FSMIe66DTN
1/+doCUasD97G1t8OkTKqo7cOtQFhMVj5+FRjrUrp4I/cGyXopL2pyicBpG+KIk9gsWqrBmDkzvx
Jjo/ZHa/6dfZB30u6G0RaP6sjkCCajYxUhkeljAbeWI0qBFr4pHz+XJazfUkCuEcWxllhQef1flu
VTlIvPlSGDHjcEZo2S8bKzFe/0sEz+DqNv5msDBG2W6tPXFu71V21ZOsiMczMdje8u5irHMGiFp/
ZL3lVxZJ4IaFF1BdRFc6x1OBnbMtO+r3WsC+1U+deNGbVhdPAIChC0yM0T9SqoVVxdDZHHDDCWoQ
7u5gWw+201qfbJ7tjTxdLm3VMHUfO78lSssUJesdsfKrf6L5EIffPHsWbkETsltzDogADMTX4wXL
y9vwE62HWvGOj4j0imwWvuh6a3mQZuR5bjoRGl+4cvzG6ETmv2Q8A4gfqi8iJ/PHX2SradZR5ozd
3GloJzWndT6IbsCnV7bfpCiB3DP+C4HjiaTefu12Bq1vrmjmkPs+2sCL/mIdRgTE0D5Y53f+exM1
a5f9VT6waUU/SRXIBI1IdKTqjDPWWLI3kODHPkD3jr+VazY1ST8ELf+OXaE3Icj1eB/V2MkBIwAL
qkUero8UTLd+Mr6lrGzNed1nqSvSV1/qPTO4r7VdrJ6dGLp/UFiQZREzrfY6LDczkuOjzAirNha1
zl9e3bZyXAuJY13j7nKMKunYBOyI+xFfKAGMim2j8sHGUkQBdniQCKEKISIsKJTUNwCjFtpDlIb2
VVUzQxlX37tYZ0M3/r66YlGx7isa0mq2MCCus92f2LVHcvm/cZsWti9GtP2GrFC/iVi4n2KnLVp4
HhcYn+/72Bp/diRGoQbydzj2wxY7y9k4HuJo3F6tr7FvLiAUCTnfsuqiXNL+GNkgzioO7rDwQRhr
JRk9ovIqeauNoD9DzmDyGeNIqAyOFXS6V7NrbLP8HU9Rbn/jeVN5YRIqZUVwrOAWWU2ARoqUwno2
/fBI/pNwObSRrssZOQSn7dMwJWykc+ETxmbxYKrSzwlDzrhksK/V9Sxsnappn9lGiTGnahV1NFCJ
hcLDbdH3J8zlUQOSBQRBEkbRrZhpzGYzBysbq+/5gfDpyVKKYBCGXlXiOPDWQvrT/fC81Elbo0dP
Cz+FjF5TZwm2PPJHfug5XQF/t/jkSsvm5yFo6Vw3ybmwnPDJ0PX2USGdd4J/hCdh3+C0jv8AcHlm
LJzZ0OCZ6Uk+TtUvv+ReKQ534nGUr1WFkWMMk7T1MVDH+Up/OZXQj/t2WdV6XEL3JoAFprmTKM2J
A3x/foPleKNzMAyS4Kfz54UAz9o5+2rPvsY7KWqi0x3W1Q3dKu6cZxraG3HbKun01SZKJu45gwRr
Nj9igVi+xFMF0JZaJuJpOHkxW9EcB/mD3Ykpj5FxLaOnkrRK33OoFO/SnRqiJf+Waasv2p26IwCX
5xDiXekNJGtM1f8jeso4UmyVbolhGAEjhXu358yDhndyBf1bR3wpV4RbTsDLOJZriVKtz4m+QKGw
pO5ARoZ4iWYkhoU7G9bJg3UlWBG+jQZ+Qgbky9ogYBicaExXDoMyDjg0ZBpTtZI100FFppZttK9F
2rYm9c+91MhZIVWS3Y6Z7Y0VQZTu/LwBSUR10GTa912JV+m05Q4eSstL91KFQwBDnOXGOekj9B/D
CKFi9UWJbINPxY9BKmpqcR3qDhiSw4OBWDPsPuUgHqZO+Rdtx7z8ZHxhIjE///y8JiMdAkaluYTW
QkACaEG7NbCuJZdmKR2pYvc+SIT0KdRHiL3qYuFbUaBktqCWvMF7FgP4liFuQzwtj5K4mPgnZVy8
98KL7jQKsQtJy0PP1jw/WaiglStAfYD56oJbQ5hkaUK0+303V83qdvKmaZKyMIbGa/0I5Bt0EFtQ
D2387WDe7fJEAomv4jEiI9aIvmfEg2ltsv0F3F5wCWuvj6KFS1fQsiphBiUZbxB4kKaVY8Js2wjH
iXtFG/L9AgMVXotAokjaPHuYTKfZUuAqtmpXclianAerzbmRzxebDSgeSr7IfvdysE26Q/UiAO77
FcmBFj4GVvYrZ5h/WeOL3DDIdNSfIRoHt9lHZgCBHMDVjbij24USW8OkeqDAFgbhNXXCnYlCVoX9
s4oqCg7mwLpsuNMPwpGbr+Y1toogOqu6wu19xCkUSSLlBQajIE2GMEvwmolyxHX659bj8yqHPdAb
ShSKwN9tHiwgIcO6erIuflsHg0tpfpn+OcMNKxHJZc8yMRJn89O77lw653CcHNC/9gsOd038KeEt
9G3Z53qgPhkSW3Z6O5vnjeCGzHnU4ikEWX/+zW2eGzPCdruVlEo8KE7eseezQTy8ytW0FUPOhIow
wJORljTXAHYEv0h4gsde/ean468wcaRYnsDSiFx29WwK4uOvLnA4JGdwUtrV99l3qnse1XDuVHRV
vwekjsF+qfyNtlT5Jy08F7TNGbPdYJ/UusXuhrFIfrD7UYmhPZUmnvpH9/k4iDMoEmlNJeQEKX3Q
TcZNhposXRHArfxNhoXdajjaHOkLWJLmxmW1T8VeHF7F66yOWeopuc1F3ygjNwI8qYA6ZG5liHGG
RNhz99kk+0xbIm0uODbAOy07TfubSdsRFncco4onEmo8CrSA8cXXd6ae4AKsbVnXXqXvGFDcHSTB
HD9RGPiFjEHZNKfcR6fa7emFgbjLF2tsIJmXJ7IraMNPU0x8LwxBJhYpYxY1JJT1KXsWyuMjR50K
5AXuiKv5f69uj61jqS11Y6zlzCFD5qnwdhxlEnsYqE3G3FtqfklYsGpIUZQedexEk4N4JJe84fIv
cAGzzDry/qM6bpdBVz+xvwahNxDOKALLywwR/ihsKq26KMjAtrBgt+auH/cwLvXi48u38T9cELnV
dlA4agxqP1+NZL0MlOEw0G7FzHcI7DpVAhuVmXCz3EEMl5vygJtuhndwfqu7tuiIz3hhJ+DUHy66
qXPkoTvf/M/IkjOJAXjkHtWlUaFInqqbYDmksVbaX/srv8JiTq6cMjiTQQrBmSKa1WCL9QDx+3IE
lHl+ffM/PcvxTKeBRwvIuO9ONx4GEkDUaJ9RkLK9Krz/ksoqQmaXYAvU+waRoOlXxsru+FQx20dJ
sOQpBMmbgmug+7xycCbEuEcczkFKp4DElhYvF8cIFf524Jpt5wItAYcuCc8gX6+3k9kk4DJxOIj1
EpL1TvB1DkLWhmL4KtTyEvpsjEpw2FhvkoJaMRXhVfxQEX17H3niR9n940XExotiSOOqamOO4xMU
Pe5iT6AS4KUla4hqwITPbNodSreCugYBGLwwUMq9zGlMVQuoBwZA5i1ypXBob7MYc7VQqDchpIfa
rqwVOB/vEOIqun6ujwu/9CSGXG0HlMY/sDz7vQTf9siyYPjvL4ho1gxDXnU9K+Og1RV5FmVGKhAy
kWYXo8KlrGQ0gYQvpVGztHmM5aNQyZpVaAurc2E9J1cPVnyu4tuyv5wSdIP3BJsklqwhUc+0+gko
reoFjYa/KLX9CU9o2ojvRS/DeOBdwbt+7JWJiSCGPeQ+Rn4xsWToJTF3NAAs5CmyI3V+VEnMQILm
kE/9u1tCOE5pCdKx7is2pXXPl3Y9U59VP36K0nTmapYorc99hrn9Wnot3KRB4xU3iAmQt4JFBnHu
yc4zlqOdew7DHD6DjjsRdwf5/zosUV6UfEebzjJsRv2oESDtIYIRsexlHcn4YBy4jzpkVeC67dr6
jECBdbu1CVmN/7gD2NygeiQWCvUfVIjPkaQ2SBiVbAPJE7S7YLBJLn1e9roFfOWpiaBEg8F9HVDL
guEQ+tpJhNU3lxoJC1p6UZlIPTIGPxuMYsURWHRx4Nd64+q08hbDQnGBSio2phayUKZsiUBmF6v7
kmjyuULrb7wQx+6dPjPinre4UtsGYY7THhXro1J3oRLmRr7hosCNxrHNFProfTC/vBlP3V9vqBH7
Is5sjYhvpCLK0sLyNVZvi8gLorXCESO4dUQnrncrRqd1jKKSlNI+PhlqS/aL6sXRVh1sCZkZhgTH
KrV7+Rx5Eu7Q/HsrfhNyDX4FATNKKv497wUzkca1kExVGlsYJyFHRJWswbOTX0PnMWusXnTOhnFY
jGxfCZhYzZIb1FZWHg9p3+if/95goRxyg+OXZaZXxqTH08sgUCHZokK60v+v+d5wywyGJfA0O4PN
r8GuC1E+qNZfQRbLRQaapu5PwUOd0aeo//RnEbfi4JKFlWNneBD+Fk18ySO0qYExeQRXOLqyOv70
Aeyr16D5DCLy1bFh5CEvfk/Zd2JY53DkItQyMySHY63ljNF4pmjw1X4u0Hdai7ff9DnO1IcDYwyK
TUBVxzTU5l10lDb48RgBWxPfxFYhkmCbjUX6SwkHyXBQ2icmQ1pnETZp55XnPewzFDh/DIy678rF
SXmyfKJbIrGKxiIZLiXZONCKpt8HWaMAbV2Prwdc+RmOpSlSKHjrKRQOTrTwgC3WVZsOBmblp/FJ
vR4ZsMvl9RvpoGVhze2FlfVaATzZdde3lgo52O3uiId12N384EU3Zc/z5vJ7VWSyhVTjYKlEsuTs
pySkIzr3jmoJvH/NIP3eErwYyXizhMMk31BhaRBPOq93ZoXGhwhTYLasfmh/sqSY+Pi5Al6udt1M
wkI8onMmud/eyDeTMC63qhFt5FgZd6YMJ8gEikYjGUm6/o2M7qFC2evyfe7TCdX3GdH+8wECHDqZ
FC6JsUVoLO5XsS+1LAJbamo7fEwgdoUGm9PpqCLuJKgY5hyn1jcT2PJdq2xr7KJsSuiI3TsGkye6
wkbXejINbBDCR6xtlMZXHLqXOsmlMrOWnrDdqMScYb9dCotC3Xc9ryweDPRz0Z/YF04TA0NeI2qt
KWXSDcM8cNYPswsrB2JOnKZx1Qf25TJ8mbBt2bT76eAvjd+8gRliP0jmkRsnda8n1KGvywRpTV+w
Q/AFuFb0QM8sdMtqqyIg/ApHzn0P9c7br9yproaoEodqLgjO/3nBEnUnvu0dC52qY7SOnn4i8HDY
urOVkZgn1DNg5k6C41Is7yHJ7L+ciBFqwxl4eAs95e+DA6TSdWz8hCpZ9Z5z9h5h/ZC9dJlqqT0w
CgSsL4REJwuc6KjnxzVj3glIWKOn+lxO0n6O8Uo4mOQ70MQr5yRQ9XzGnALN5FDtsFfLFQNoZyjI
+FUo+Cde46mPFdYvTiEnm18AgPaKb6ZmvCttzhhLbbK3V/Xx14Zfa4iLajv8GCv2xpSHSEle4b7d
9Fg=
`pragma protect end_protected
