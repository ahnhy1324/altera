// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:46 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jRhbzF7PcSD95EYKYw7d0gqhOYI3sHBWQvXkWHo7ZNM/ntgd+QR37DnKAxIFCzQ4
2fKKeQ2hYzY+UftuAFuXMgK+VMQ1MpHXpP7bSWgfGkyuqdYbtcqpgNY7KzwvhkOU
E69pMHiYazuDksfi8W82Ka6nCfGd9mlV5MUzsHmARNQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1680)
0davWi0squpNCfOst1haEq+A/v9Z09JxplajLgYSM3P1YgZSlw87i3CQp7JAoLyV
57kRT98rHrK778E/kV8P14kABU7geLqz/Qb1eu6SnKCeUray+w+b6v80kHDE7tgA
YxoLM0kOL9v7K31043hJ0qVwmxTtcw5MMV5jG4gZ2mqnrCsabXmD8k3rkTRfgxmc
vG0yxNXjo2GI2MO5hT4txW2CjEXq5K7+FXGuvYgmAbnJOrpKw10FWrG8hRUuUw1P
if9Q2KUKoaNmevFpJWIvB2vp2tOq+/XKTMbh8RINMartuu9Ihj4SPpmfcEyVXYJm
Wq1/cQEY3Eo6NWZHGlsp7NJEEMyZYmks7nmtd6aUyl5rHle7TzaWMcVTlWxf0x47
beeQ0nFVteTYHLsE/TQSjihHkbk3AqynxlkgXM9C8TpO2wY86go9hYXaEY3Q8Dt0
DfI2TrQ1Gfh3N84l85RR4KerfjyOLPehuonkdMEgaD6d0fGcai7YpJ8idyuv8ypH
cuQWw9z4fFwgWuMluBeo4EfHePjlK/wx+mrzGn+btMCEr7Wap596Yi+MFXOMDJwQ
hoCY5yDwzMkw6IHiBEcFlMSXB2x1yvWBSIWZTv/mRqidJ4MT3+ER+67Put78IgeK
Ets3cla4AtrjtcuvmLnbieRG0i/hvBCLyLLhrlPg1CGQrTT53dNWKA9tk5lG5JIf
ixGlxmXVhBHwGXhwXmhXZmM6ejA1IEf1w/Vbff7pEgq0exXNJAR0ykG5f77uS1Re
cZ45OyZlnELZboaVKifxVqtMPqPb5hINpjAyuOnlwRmx25KaOZLV2Q7XunU/jsc7
PHR4iUKLUS38tLszRwDZlXQ3fnSqpGHKrDquPT1BJgghXpaqIpLJUorkopGGWd/b
ENn4FolSBi9bhSTdaZ84kZzP4mGW3M/33Y9ofF/8sXXKf++QfhjrQ3iS+8t6rSkz
8rINgsD3a2NRPbwxXGaQkoPVUJPg94GgCfMfzWp9YGCJ/svArc//IPADxsET7yge
J9aXp7gdrimdPEQw+7zfZS5JOHZ9DymtXpHXO8yOOFW+bFK9NA69G1fCRzsuN+MV
JqUilN9o7X5dCFNMk0lKdT00oafeaD2yOacC+xqMZ2VX0zloaUHo+VPU/iYW+4Rd
w0K2PUcOS2yGuJgM2YhIJxex5871D17fimooA8awPj3+HMhjxpd/2Ia+BHHrRfDZ
YvOL84aOLT0npj5f4i8c+9+vr+dA8JluBZ3QBGSpeOk+JEDqFnmHE+/w8nKUcOX3
0MuK8cZh5CmGSj76f8YY5gtkOXPuAAbwaEPrj1LWEgwsj8XLE12IERG1hegfEG1e
8H/J4SHIGVW/+faEsa5g7SC9K2msAaia48Mq/GG+T6cs8kQ67JyJRtND2+lr2rZr
7a/P3N56nd2sl/Jnr7VmDC1r28BsfosBymMiOdUmtuEXIbDP7D0bZkg7HRA8tOhz
a2Q4rDASZKjUFYh9jNYd8MQxSS7WcANFYdK0ZbXSthFdRtXm7oFfgjGfIC618Ohf
iwu7G0DAiK4Li+JEeQpm407iT1CmEUpt5vsdrDYp15u4s457Xf8uIfsxo6dBS8Kr
T5NsrGk+oPPJuv6bYlxTG6fO6kTEz15Sp7OHF72XR/m1st6xhvuyHGFVZ8wj1Ctl
XLzUuEnlyKcTt+YzsGdBUxlAFerIK71SbOybUmndGAw/IUNlPyrHtolj/zMfhbDb
bguRq7wjsnC5ocCkhivPXzM8fcIMGVA5ShCn6p20j/PvmewboK3K64GgaLpKVCKE
4mTkgGeNAqTcRyVDXKnS1T93zJ7umh2T8tdZmu6CiAB4taWoFEEftJhvdEds6MWZ
QFfYJTnqQWFFpkBifM5jPHpDnnkRPuy7kDYwDApHqUZmF8Rz05phkVgP7Kr26EOW
x+fTjVuyH5pzEDXcaYLONEun4fGjaA57VjXFtMO8BKscJlbniPSotJNYU7ljs1k/
of3LYprB3We3OsXHPAI3/SDiukvuTzPZGOvsm7Ht+uDtUCfRdC4/NXHdfQJZEPkJ
ftoyTkfvhEykXY53k3783IbJ5mEj75YvKS+XkftAGh2LWQ6T8Tg9Ts+vvOukABPD
m7HVU7ItkCFpg83f9/Qe3NA1PH847DsDRFKvxqBslR+UkuPtCC/kGk2RK6Asql7B
PTp2U6volgdHROiJ2ohzxIsfUEpaAeJAmPQvghEyTfQ66oApyvta4gkXL+ZaPMkl
`pragma protect end_protected
