// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EMrOjTBzl7u4G4jcu6/bC2d+v+OstHI90Dx5KFxaWq8s/NESlB334Be2Dd/zfdAS
IbXe2WMqOUFnvTo6IIMOcAiPCqJosQFZgcTnk4pMIq+gVunRrJn4rsG5741NlHpZ
nDz+44C1ghfYUO2VEQY8bKo+4vBieK6NrKK2764gIK8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9728)
O1cDQNIdJMIBT2LzfarL4PG2k5N7663V3HsjizuehN3VNHFAcEJdMc1E9DqBHuXR
rBjujvhaLF/6DJSs6X6tveewvtHnQD+L4Og/ZzLl6ASM9TVHGaP4uTe3L01HZJgI
5joYKgQp46MYu9paXHaWq1BaHQRAOt7z2bv22JPdkazLY73l3DKorIwPRqI9Z91N
txzijFh7MTOU1mdoDLH6yema4dKYR+gq2MRDmPn4lbJ20GfeQrH80e+rwnfzNmAz
G4MiSuZ62AX1mbWDZILDYC6hkzOeYA+apPVMLXnZQdvXF6zs0bReU1AqMinQlXzi
UPph9/DEjrf5kgCPjM4V0mgogahfdr7hPL+qIFPGhY1xCmcu1aB/UMsHuLJE9pLa
023NLMW6ziF1W5dyGzCLcuTRrlBqZnbvvr1ccs/yTTBvx2KsYYUypFh2mMGK2PBL
/U1JDh5owcLsb3/7R8ZgHzfhmR5oaI480Z+5Z0R6HTL8KjVNUDAuxE3gHRwHBTBs
FnL0VyFS9pBygBRIrTUJlx+J9Gn77bW1h5uXTXle3MQWOr4gTNfR98NKLsxX6C0S
AY1HehHh9frPvzcxsTMlIJy1jVS2+2n55ChRWo7hNzhbnO3wLOzaEqW017dJRO1H
RApHn9TFfuVZopsmc7Ub9nZrpI/bghb95ClNsj3OmUjNCzcmVl8tWHX0901xteSA
y2VKZI1pqKp2mDV3/uo17R3ib6wwxHbL0yPoKeciRD/zIvikVFnQ9BirUI3ULyAT
FMfQooRQO3R+FgbkgAR1WeFMfEwi4xj2bZ6LNJ+eSKElwtn+TS1V71cFPL00o3Z4
lbQRsA/TTkLmAnjrBny6/YtxgSlehfqAGUH5/E6AOmcE6rF793WsCBph+c6Wv+D3
gorAXjmPNboiAyIkwuqUyT+qqI/Q/sjV1fiLwl6mOS8S7kfY0d2a1QQXfKeLiGIF
WGSc5B712p9O2oA0CWb8q779JL1ly3J8F3yW3ScKKR8IOHi1LYWqSC3ZEKqJzbbY
PnG9v7wP7BSgxOfqxzsunfT2I8wsFujc70TBowbOwAYBM6rBi2ABQF8sjaXQgLNo
x1DfqXcRtBIc0spo4ezVn2/eCKk1cdbXvFXPFM28pCDLdfH1qYZUY6/j2aU2amNF
ZOxIZbHHOPfSX8rhXgHNuinBiVONPUYt/5qwU+DhwN/m0MtG9G/f7OiFk9up1jhP
3sCs8Zreip16EHzj5McaKIO5vcDQK5+0E482wzYJe8NPBmr/NMFueCWBvaXZT50+
Dka4HbazFclZg7inTb5rUTVP60BVrZw81grwNVsJnTZY15EUmoBSlaeuMk4Qr+dd
ia15zxIXVpOnHLswwMjISTk7PP0w7Zp3c29fEbfnBEb5R2BCKC4U+tgwXMSs/hvN
pydGSbxHIT0SvRC6mCvvH4XVOLZBq9UVhhEKJX/0dAxO9sSGpw55US7OX7OrspYx
ka/zIjeue+Qe/05+yTWtrBbnXZ8M2f98KyGPlHnn6roVFNaA6XmI4gUGgBNpfgHg
nwLIEn1Ghel+JFOWH0sFBIkhQnU88U3MAapPQqV5zvXvYHoCRoP+1JpyEneA8X4Z
T/Vv1+B2laujPXXZkJ8B6KzaXgdpVntOZBP//J5WccXDbHhh4RU7GyVwKFwYzcsz
vUu+96MCrBa2vf6CQWQEgoOH91IPfo9VtF4J7uEJdUEZO4kwLx33vf2HqNBU97B7
ryO0tC8p+TiK1+jzi/R7WwdJvKad1vm07uht9hXOMhA6AQ/zI4tz1rRMOnLmqXUt
35fE5rJnJXyhgaNdC0DOtKno1as+DF/n2E0MvR4lVDCbuiU0xMTzrZVnMGdsN0Hv
zAaDQqOxaC3OjKNP/WY5CKEj2Lha0FRESWsL//lfaSNTeREXr0hTK/Ly68eICIQm
GSIxTMfWsRUYEJEMFFtt8ChOykCQ6H9EohojJpm/kvNr51uGVKLmNP9kcyLjhc51
GzyEziiIG5bCE7W+LBkT+ZNsepBjA3kJfykGgwKb5dSOJUTlhgi329lFmnYrYOvd
8E8mpngshSouiGaM9sBURE14XXjgdGbykoWx6uRHo2n8tlplgAUkycPO4TxYA8Gk
8B+P580faCt2nOIjG3qkhlV/dsQO4+UvCmgFYV23KNdFWxIcOVf60/LIy+hJLLoD
JvgWKO2rhbLewoh6UsWMYI17qxdTGjrw99COvozYWyS8zULesTUL/lDcpeNsv8Kj
s2SmoMFIde8/GDHfuCp+skdxBLZr9assfHIDylRB7FW2+KKmW9oGszwIJsoYUDc0
fnF2Ry1KX6Srnc4qjrU8GDbhjo0Gci2lPqGbg/7Iw+9xH5PkreI7pOwu1Wg9yolU
2CT5gy0KXRoCGUZ9/hx8w2PQg4hLZX0ouSZivYc/vabL02i/SHVBKf5phGcpGobw
HA2mbYf2lT7v2Gx2vS9WvmM9T/LOyi7TWprwxGGjXzkjGh7xM+GlRIHkxCwd3Ihd
iTbiZ74Uhub1lBIqG/dfbF4vMJNcez5cCrVCIW0OBIrNZDGDKbgxoYz7RQqtkdTU
Ifr8vhO/7C3wHPSNcvwIGxLs6s6atMrKN2eTGWRAYnfgTnO84FNakl/c2B57w72Y
8whUhFUS7KdzscSvq5JezT/KGDQRuehKlx9afz8OcqKe8G3jerJS+Qb+UNNlpEs+
7QrV56FFk6fthp8ebkYnDCxXN9hYTSxp2McfXOIPqT+aMv7GaJ66jonQr4+kIUOj
suQcF3kdqwSbNwDdDZlvoXVl7jsZMwOqeVKHCXYPrmJswRVZMD4i7EInuU+JuyqW
4w6P8K0+d163CDSyWBTFle4swDmw5qqYjLFjvRKl0rN2oUhCrT1Fu1tLCNT81ilH
BSR44bypx/b5ZfR50VAvKmPWSx4v7U/Tzp2vYwVZzqijUyv9Qm9CNb3VuNuPaRWV
QY2hT50yVgFW2HhkiUkxKK/2aQE+I2oozhvebFmuzml2gR7HKVVIpZAvFjYnG0Ks
1ifwRCsk/MnHKNkwT9FTklVbFBY+OSF4kYKFVswOA41I07E2QRkEP/bY26vUhM8h
O+HsqLHxs+XN1biKLfysERttWf3h7coXsHytkFpBnTvQO5rOBk4bVJskwTPk6F2o
As9n9k2EbBGqd4YOQ2d/3maIKWYCgw2xuUt9UxIXDpXvjH2bUE59gQ4kHxYnj29t
BQXh4ILViYjUaf3UR58ffvo3N53NQYZgAs1LoBkqG3tEVE13zd1dYYfw0bsWAAR6
auM7oZ3TQth6XrlQLlUDyN+ny8j+mgvjA5D8uVgb8rfMbsqlnyEwaHJNOazPqgpd
/qjy9PkUkTRyCDJj60WvfLnHZvBes17Jd7Zqxm1QWvUUcPnf3J5+uHdAXEuj0IVB
Dc0O4If04BqhkvQjF9TidlBqFwe5UpSgrmxmjgPt/uhQh2WTWjq8kZNcGywfDrWR
zbHudeY8B69bQduiz5xkPSLgkiIhVvv8Y+GFoicrG12NqUt1oQdpL0HRrn28obgu
kbh5K4N0AKYUXqV9Z2+/huHjQlfQ3HdNMeujOCI5C0S4rLnIz6qw6YKnuYXXes3I
AnZ/Yu/T2JyEZIeVOX3o2wqH0zdzgHYq+B27ngs+jyTfo+AVEwrXGVTyeKrpETYb
e6FVHhzAoe0f+7llOpRZzIeG2ndtG2ilHjs+VzwrkUmMxk6Himh+noOgjhZVu+64
ShV5nempd0/+phv8zhHG1EmAis7oLP+t8Thn7bJH0dTsHgN46X4VMZQDw9C9bDfQ
k/DWjxHjtwv0Eh2wNncgDklbbrMvGfVp9M9ukIvrE4BKNtOu915mO4U//89U6r0V
OBv11Sf21/BpNbTIj7S02j4PZE24TFI9CkNmvm8K1uZxxbJiNZKiNHotXAQKptja
OVK4K6ngMig2sMa/aRj9OQ7SGkr5KNQyV7uPuTC20U+MuzdQcrrgKQXUbC229Lph
fUR330BozPSrtYDoYtqzGdZqQbk9hLN1Yz+xaef8FwZCfT0ODnlSEYRzePzG9WVs
hw6X0yyTSYkFHSHOBF0aA3IyrxRp25+6ppHR3+kho2xP0DVdrtwPOEAnc3sXAuMC
reR2ALSIIn5FDDjsG1jjVXfg+Xpxy4UiYm/H5LTyVZExJgaC04OLM7Bs9MlOClBP
HCqGzHTSLJBOl6T8G/xreT9kDDxxu8pMFjeat+L1RhP2hDfzA0iyHNjPdoNJnkWF
2KJbC4yGZIuepyimfYZjgUwE7efoBhVba5HMxnQIgOuDzA4UPEcf1bumK5eUrGAC
Fo0b46x+d1z//Q6NgkAR7LHX3pkqkyYoJ/4UigFwI1sMtx5NSiB9Xo1QZ2gs+p3g
VKNVn2Ca2s4Oo4vIC9iLTg/GVVpkcxrpukAZiiCp1xIcPmZHYyVMAsLFkwTrxRCH
0KuMcpRWrAi1Fgt+KdKf9aMiezaRVFizsz+HLokbtomrmAznNeqfrg7HQwXc5V95
CD/lqYR0e4LqJ6ElaB1HJqL18eIcZ9c8bgEnM+xD6hb0miZ2CoU8eJjL8E8Sy3pJ
FpKhlEc1volU6587WjtEkXep+J3Z2g8hQZzfWk6dW3x+0JhMMNuH0qurdRiseZpX
labDXV2xnoz34Lu1K3xtf1bSNB5K2PGvNP73gw/u19z0lTWV8ouZ5R8Z45U3PX50
TkbfwQw0tGcLAxtCvv9oROwm85a9oQrDoDF3mABrvUQ7EZ/CsAFfqdi8DOUHLsSj
a8AqJ/YwI2zfASsjDZ1OTCm1Fc7p23hwCmfDn/7SIJUY9BO3vISNw7sjR8B8Pu8m
g1Wm08F9tlVoTMP2uUHxReIonOiFy98tEvs6PdkIRr2hBLxDJTLHV5F1mPPtLYZ/
ameJQ3i2WKKA24sBDahoRCFxeNfQkXKly4K8FUN9zXZIs7/TUJZn/O78uSw3K8NG
e6E08Wz19rtjtm2ZkI4RZIz2I9GqR9Fk0fotpyBeUt/dKW+ri1Pg2qUlFuKzbp9o
NswgrAOd+oJzg6Xeps49iZRwhkzhl2FZlfh6mmx/1CCiE0gFioB4Y7xxRTAHP2dn
wGtF/7eqyUn7Q0/jaFpnzTHRBGNXdUIW1gtYAZR3SGD4n0zYMHPi5x9JZG2u4Ya1
l08Kdm1H/Nnws78nRPNt7PkUWQKWgKWzBnW2a179pzNLtan7S6xUY7rIzBKxbQZJ
yEnXl0jblczZB7R4gIQdXZgmnz211R3GEz9cPOdhDb2yT/QumIY+5T1y+asWnr/m
iBuGtBnDNPThmbEq1VCondIdvppJPHib/DYYcCkCVn04nshcHkng0v12MmUqmFQA
kzwAVc4EJ55svCCS2gNFeUyn2FFhchdkmWeOanOv9ZzN1wy4lRVGaPCoI7MitHeU
YkM5es0O94w0O5VJZG0xI+8+to2C3F5FDDi+Qy/zz3rSgkf7oIzwrC7wHoeKGkuX
S/bB+8XL8xsxpHzC/1pZC04FLzOUM4O4HQXA+uoFKzTVVIsfhjTYWJ0VOKEIvKRU
AlcVTVphOxMdikcZcNwJqir2ntyoCIBDOL59dIJZMHIiK5xRe742MxGmtytQ8wPH
EPJLXiNIbDg6Pq76ZGGHLGr/w+cAj1eRVc8JQy7dPdMliNFEliC3TMzSMbQzXjHo
LxZkwQEOYBbNgFySQQeE319syDESVK1TAHOkLpMOIJ4qFT1vnxgEtuyDF9HJiisD
942YWxmePvYCeicYlG9w8swaITFCKozsP+r80WBXWJrfsI+lCHeizAux7JJMqPi6
eKimT+87lB9HHMUaKHBJ5/75+FbcnxG0qoqvjTZLgX9jq9O1Ay1hx0oJZHecQ3v0
5d8x74qsQrYIyj8UI2fgS+YXGHvxtcophXPY/J6pleLPmjyFcYJNxo2uSFXUYB8I
8aEjeS9JmwH28Q8k3sPjlO48D5sm/B5+9XQ/0azCknX5vxY1Xd47EEGdbYp+tp0Y
AafcctmbenUwtJmbHrTg98pE58BLm6toEcNo37mrDyTmn3ncowCw7FP9MdAR0Csc
GfmGsI7hhXAvs4ovBjEEnF5jo+0jE5jDYGM9obE3EgpiOLrp5+GPAZ4dyf5g5ySD
nqTyCWZCAyFdptrlldYcwX2rrGLzBB3e5iZZ4qIeYbANgHSajp/rdBVw0sznKOIN
z/EqbrvB3XGbvgMuIfnT7fWEaJsbcVofkiZTKen2gGJMDIk0Aakua8hSC+J2Q+i+
cslbqCovKkbjQEPg81TyGsFCV5Fjl3420BsYW4zkAXR6lOUPeRVMKrI6MycTfnoq
zzbp0PQyWFdEOFIalT4HKBo8b3jrVAeADooaxxkMmG6KvVilRnE0t2ou4EcCeNGt
KgV8MFeiUPDqGdcJ65lGW7pwL7UQsU19fcdvnYNvRa3FUcv9tZY5dhnMYh8rfF0Z
YftKLButiIoM0Ey3QImFFxaD1WiCF0CJPOulzSeSPGvtpN7uZqhvR2Y/O9dBGcQ/
+yY2xeeMI1L3ahhH4taVfdh8CeDvvY7Xmae8jaY6jIa1Hil/m2AyCdYfQJcqOMje
cMK+SUTn8RG5hvi2vmX9mZgnsxxKyFVhaJXBVbjRbArddadRYsjMjYPSCBC6p4YM
fI2yrNMMIyaYvI5XySEy+2tQWSiM6cbi3vMXdilgFZAN46dtdPzOvxH/5JrRot61
OndvGDdeNmRUHfbRDSecEzD2H+tWpTbRYUeF7SwaLrpGt9fmc6yN09xAZpJUcy4y
6qjrVl409am7SBtRgVV8c4jYZdtcOgOoNkD9nKMsWZsa6zMK0Kyq7Dp7r4a8YJ2d
mYE3tq3RlePwLIMg7Q/uS3NntU2FBecMNaFoguyifBxHPi5aFNkpJlMh6VxVKwkR
SFrJ3vHPPSr/tsxtpF6mbhTJ4eTwKOCuwpgRAwYQV5z4CcLLhzoNCtCsg+TqA7Xb
OXnYAJPFMEn5EUw05U+bbzYHEcOoJapZyC0LEfJeaZk46QAPXN2mB3Rw3IUk+nRZ
lXlKYbvawkdkrIi0JaXoN3t/QhHHdk113rmqq8WiIA1NA4lLsZPUQz0blh45m9Bu
1SyrIE0rtuT5M1Q2aKS9AZz7blhKXGC9JdAx23ur60vICs7zVn3qcfIQx2XuwK+F
ummH2pspUgpG8js3viw9nC8NJPbaJpzcNm6oYp2ovqhBtFkNlGJi7w0hILSPjumB
KeJvSTgH0rx3DV3FDopgJ0hVZWwO/3JCigvlJAE3OnWCa5JbFDlnvjhd4S5Rncgc
vjjKAzzkB/gAun6V2JGnvinvycDZoVCe73rfFnR2DpWEAgDFi47h3Kh+i/aFKCvI
lH6uZJIQg94TkJEqQ3nkQX+R7VXzYLmaPh6BRpOS30RujuqAJVKy0yNeMf6vViBp
Rvyw5iXxX+oaznEIOxbtbz1KNo/ImbspfN6uCeroKJb980e4Soxabqx1bnigJ9rG
3RdIKbwcxKG20smOG06amF8TTQsxM/RG8ShX2OE/KL/fBHaHC4RsIcQ0ueliMYnh
WSuVi+sg3u2W6Bx2teYQ8rTvrMdg8Fpa97C+4vFy1zmvpFlyMNm9sfmb+6TX2/zl
M8/ehWbZw3C4J7R7HO4eQYohwpnW3s7NwRkczrdTY/xSBUHtl9uRd6OFzTE6DIiR
57DMEOfbBkxNQ7uAvcgaGssCzD8HpUadEFP8e5nvv99MEYVYKxfFuS838Mj9qRz5
3bG9O4szT3GTvB5AIGTsDg1PlNgfcmVLieE9q3dwJXVcY2DGSGQyyijD7QF+v1LZ
oeN6F016TR1iXCF8JeaUbX99UM7yBZX3nD8BNmom2xx1/GNG3mL30B0/LNBS/mij
fgOvES0lvyBSBbczSw7Lzeos8kWpk/Qctstc5l6By/7Nlhw3H4gq7Xa7NCcqrq94
PtI6tzxfURlfmnkDn/6sHP2IiEXYtafmhW2kdcBQOU4a9G/c9kqA+mggABuNSvzr
bpiicD+1JzgfsBAJRuChHIaRcAfkJqXF7mukJ4iU4Q40B9HeX5BpGccOPpLn7cNo
rga83xQD7jXDiz10jwKW67xb6rWO919KWD+lxRVoWOUFzk/yZYG41wKS+ITZggCO
9l3cXtU1bu8UVKC4HE465++L51uAHKGMdJJwhR4mR9Zd0/gLiaaN04WdpaAfpnMz
Q5nC8uR/+83U2aZODmFVw8KXdRSc3NUFvpBXCzfNyhXjDKKAoOPWReAj9K5q3o7n
5V3FOrxoLY1S1qgp5rpBuPmUri+cbwJpj8JPyV1mgwxsqVOLIrsoUqnIQ/RctjxP
corFvlmKbQ2hjRY6ml4Gm/LaN2wuVPBx19kMnyNaLA5AKvkrgFMc5S6b8+U/fYng
tg1ycbfLex48NLyAx342GWYfVEtJZd8nRkd1HLQTQcWNQIS0RU8tZ5qdCfYXYmYT
YVooLkYL1PQBsJvk1DkhYjmz57Hw6HALC8aSMlYb4q77+xTgpKzJP0M6pex/htIH
twhW0XgFWOs0pJ6ce8zWaMLzz9NcQuV2x6OpQkfx9oQ2iz1iBQH04T04E5Y+XiJy
n8lwHcBrVB5sfw5Eov8zghgkGk9XBMhoaYVCtSTIklLGrGBHnn3LgraqBVR9bNiA
vwMIxMWqv2/BPSwyOkDVAzfOzAuJWmDN0uhggx5fXxFjA+WyRj/hX8umIkBkcmHq
zoR2UAKvwvwd6ThZLLh5HAOnMjxG1smT63zxaFwpxJX14yTFUYTp9uKLejpOYbHD
NFj9yXjPJpiwfax/5bMtHQO05QlaDP2pA0kpuobpeGA5nBRNp0ppK/NolE6wZJst
ZkS7Ms0CiHM+7hfs8N17SJttaw1ncXpOhiYfvx6hQbiAW7AzacKrJ3eS+8r9Rkmz
7y+SmXHf2VlBXjpoMgdCQGTHTBmbVyVeRLOEx0VVZLeoHB08Of4/AdWKF7ODldIx
t4CRBRgsUaxg4I7EGgQ39hRgsC4/m6u8jGrt3a+m6ck3rgINr8kZxHKvzN7HLTJZ
iJ5SgxX05j5NaCvOoan8MiE1XO+T+hgACw9LBVXUxuSNg4dyHtIHagy135AL8cvH
aegvor1DVqgLqUulyJNOjJI7heJvHMwPPwzgpdig1w7He2iJCLxxq//GB8SlKR6Q
P7bAt41FD1IXrs7jafRm56ovSLrK7GXbzb0hJYuIfhU0aHq2mpW6YyJcF1QaOS/J
8xVbm0Lb3LIE2aWBSbdoMpUMugLejXHNvXwcfbgC5h/txrYYGvzCYmdQ1YEIT/yk
E9DPbUvinPkr/aLhdbceAnne6LD8qbgU176DLNACq2lwIZYdBwGaHN17uZAIdgJm
0Me5W28J0y44h4tqB1mvIf4FnzH6AV5A0Nz0EBBpX60k4YJaLojdkYy1XSh8AtDS
gYmJ1IJ2deRsCSYeu1avEYnSnd8n2sfz70FQWJF3ZIA7dwk85EpM8QdyfUTeNOsZ
hUZJxgSzH82v8Pk00tI+oHnKCSeDf59++K9iX/9bKmEmnz1g3vNZU3qYl7giWw2H
RkY8xEGZyhnoaoNipfOSNpGUCePvBqJ2ZQY/F1S8XS/vCOaFYnKTxen+VhV+RbTQ
9bvHl3yyd72ld9GqRJ3i5dTz5qOwtpa25V2fSyQ56E8X+4/7d2yp6Q0GYUw/9Xd3
wo8xo8eaNlOhHGaTsAce95ou9qzjfBsq+npqoIKzgWjjfWPikWTJSbskMyWezAN7
lnrInYUp8xlwkDTdFG8FZz59Ll8dpQd4Kx/cE9k/ex8Y6+fHuyjPHpYwTfwRj6z5
fnKq19QvZh90pAXJCiaS+yOSJIux7LC1M/B5mTi8v/TEU9oeXETf1cy0tKCxS9kW
MRELot3lLUtItp1g6oEVlLMn8a30Tklc+ZxP2Fnr9/1YZh6aIFso/u/+2twmFJ96
sOHpbFtuSrLZrpwyQKR5O7M7jNKcKH6zeMD4Hg1b6JJH6mkv8COfqB62ey4/PERq
DBzs0zZoFxwN9PMya3xBmjGo8tsT5dCkrULasInYKtQang59zstOSKcWCxomeoXQ
ekoJv2JQc+70krTFBoCeiO7SOcJdfDCbYAauG8niA+fmMFMiZtUtx5AmV+CUYkzE
I73mMKk90VahGf/6OaWFLyYTcN/J6HH699ICiu9+NZShNZopreANPxmwpF3VG7Gd
K66McaqMkrbzToske0fu+XSF9Nv0L5+1oGCnKMsVBE4wq3IXJDWTs8g95VgCs5Sr
3gmgtP1bJzLhDDvXNl4/DEOzL0BS9Dgw6BxvUubQN1o3FONNCNaYoz4l99pl1P5O
48ZBjH1d70jVtVu8gdkxiBN3MT/2nbeJiXpX2xG6uhKxMJ8etQTWerh18YZVMQN1
lR2/sZLQg8Bzll5n2yoirVSjSrM7vgmasR/WmbDXBiR+pWS5qYTwcESTShVmIig0
l4YucXkgoJVxT6TZhnFk2tzcioB4zZKW6Q9+J2lUjs1QMEXPOzHpqFd7b3IL+ZAz
hkD9Oocc68dNxcnsQOyKBBdENp+yJUlPj6peVyq8ij1rW68Dsa0uy44Up3o73FCu
HnZ7QYzIuEmUyy3QOIbVHlEDt+YjVuY/gmQf+kZFUKdhNCN+3zCOa6sO+vLAKWVm
pV8zZ1/kPdpjtF04EfA2zNtxUB62bqnRXG5hf4uuCHCXFO9sfQH9S7z1Of4PGaty
DVaDdk7rsbFcCjJM7mHgYFtxX64Jh8dc+WCXmYtZrB0r4wn1WyofDQ0s8uP0ywWE
uGcBKW6k9bYf7iPCKmTN560W//BKHKm6yLVGt6gP4gK9FsuJk6CGL1vK/gE9sHub
R8INlSznGlIyJH+xJAYcQXfVTLWThJ3xGmoN6HHCYYzT5E2baJjAF1wzYrAcjqQa
FDwuMspQDXdPcPkqPR9IH0xTAtCpm9GCbA8GiUSlp0ISxMVD/oeU/EQfc2of2nGa
w5KUEmId2wxj/esG0mWZYyAT+ir9j7AcOoemhzMypWhGqT0+j0uEDqepOHhK6JBl
tPUToI3gAuTwVxF98pbH+TodO/OqvuJ9UAECdW9EX1Ct9EUzLM5cRm3lazPZIqnf
E+zRRNGC0MeY/VLp9KY5qAlLXMc2+0gbhUTepVhNBihzEWIVFIaLkDiW+nq/Snzq
wVPYivxsVnPiBoApNVC4isKdnCQzJyetFyaifcduM+FN6WZ/ipXGoZETkqd86x0l
yze/55p6PfbJc4fPeZm/SQsfxGnRJ6zJXgaAauplqgBfs2H5vLWiP4CTOj/4fvwj
qMCnsBtZEiQahcCuA5W4MtpT2sdlSbBHhweAZWQbJDrW17WxekUYuUxm9NZ8oOFg
M6Rp1nYHFKjeQ+PCF5b2vWpyjMg57qhuKLyrxCsQfuL2X2fl+rYmawtgfs3BHnnI
0XY9ErU6HrPUf8QVVY35mG2AR2Mzh4ZSdhiHj/xB0vV+p8ZgDC3kd4V5RVR/ZFyA
KvoFSvSac/an7jhN7J53mZf7hJIKfY/NGCYy/R+2kglQzynHXf6Wuh8Uh009JcyL
3a5+vMi4gd7zHjMLXjT9ThTLJoEpsnuP25lEVaDlI5I2W6fr+46kJ7rDmq5okm0m
JM9p5/lRiLNtXW+BoKqCVYbhe0CdDw9twj70Ej2phVDR2zzjhzjVbxRJQXjRMT7O
k4YlDZu8YP1zSg4/pXSvt4IGyXHyYc7RKqmln5dunfHdD50d7di7I28wzo3pmQ3R
Rmv+l8w6GLsJ8OHZWj9KmG8gh3/f8pm1xcKLuRhTClp7Ab1fgDXcIIF/n76kunUt
4H2oamswpA9MV8KoFY24qUYh8xvT0Tuo8j8y3KD8BiqS6oBYoZSh4cSkOoUjHSa+
0x5ehgsl86MVNUlu7TXhzjW74aSP8Qg97kpFd95HmYbpZ24Z5QLlvxOMXRVmVtc1
qoQSlG1jwSDxDgJidO1i/08Kazt6DvNhaniK8SPX5RwqCxjVp+eWXy7099wXyJ9t
eLihyuLS9vKMh3PyDkB7vKybfp4SvgWUfdHsRDO6QX8d6OlWQ7aVxgsQ4rkSGEJQ
gckc7niSpdsAX+uJfrePBL5/I+Ifw/ew/KT/ssL8AcllIbqNZLsdK2HF7LWUoZKF
1kt07wafjXIIHW1GMtYXXKjxDFRt0HPLU5DQPAvcz+OKUkAcf+TJQ+HbnNy7O3C6
KVIGEY2qKF8WEqTHCzZmmFMd4uwXonr7daHiCug9STJR6I9CHF3Aswm5UBBm9+81
J2LvFByYjPfhYWwQyP2rqzwjlYIRAj6zJWEgRkY2pTL+Wl7dwhQGwZHyvkAqnmzd
cWWvPvpJrhOO/RPxUewlHs/xn2IXMqhI+Hwt18nM9LkGaCnGL4fqlkku0f1x/ha9
r2GHjJPVDrdF/srXc9l6VS8Jbrn188KzLAadA8CCEQ6+ASq3YRdOksEoeoL/7llx
YY8HbitwOGip7VHUJJ8VBDrUiSOZo9nl6WLzvsd9+aGAa916yW5PL1DhnAScmGwI
djL6ifJC5FpE/E45umIHac9U2Ldcw82svxs6REhPJfA4UI93T8xaUYwXK1bs5np2
Lf44SaTHzIK7tgnvCNcgp5QrF38TkYiDERhDjI8R9QxCZTfjUicueYt/UV0FJwqg
SS3kQw0afwaBgaZ4xN4/fk+jk7MakXKbvmeYpRlm9Qyx+64XvUbIC5bCe99rtxuq
gE9EFwn84WC9GefXOZsfgZjdk8COtOT4YzNjn2+kt6+3aqsXorDsVoFzAHEq0Jid
C7yoAVA37yYrC5S1dcT07a9PgNxCBuqMuWtjWbwQqoltu8WH9ziBi9aqt3DGr42W
Lgcv7ys5a4EU1ZBtJiIMlRzGTpR5X/QABkXFaC5V4orgsMmKRhI9WPp0Jyu1TI4/
qCuYs9NtCw1lNzbRFY9E0Yv6SP3+I9ftcQ8+aUsidHe54y+aO0L/LAkLcT+6DWso
dKzdsxjTJB6bGHmFcRmr/SYy3b3SWaRBNINUG7fdec40v12Nu5m8J46WozG+b+8f
VNdkQ3b75J7cEuW/DAuVtl7cz2QOWlkdDGRXURvfhBM=
`pragma protect end_protected
