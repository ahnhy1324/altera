// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FNtDkhgqiX1VC03Pp65hJE448RCCyby4Em8ysEb7kcFizrL4QUIQ7pZ0SgvUvmEP
Lqul8KXAola6YjDmoi5KPw3pSqXWxoXxFKTwyeDukTprpJAafzvswI6Cj4A4/ONU
if2W6sIroII+PO4vcdayz3On6Ayx78T8qHMa09/JP0E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 89520)
IYHC6BVHE6Y1nVDOAXYQryuMyXOn6WQO5Z8qNXeuc5ywbGUOZcTEr7BCtqFFQsUm
f/M1zm+KOIt6pITdvht5uLk4auqpNBt2AK//NXfd/hxSZ92natBuDCy53+C61Kdn
w4Adl2RI8Cysunn7o7fQ3Ooqv6tb83gcJcAr/HkPF2c0Asae481fxl+zBzVzagN1
1LFWMdBnIq9vXs2uJfgrminC0CeL4fDaqThOPt4zaLfEXHX5/BB5I+y4+RyWgNnp
s9F+iH2a2F+KM9Fu5+1NpOr1vA1ua8tRMdX1NVs3Kwn946rvLZ0OPu0AjXt9Yp4M
s2B/O5GA7vqKZatd1EBWM/2K31aw2LXKkwsQou8UYEYJqM89tCnr0LmNUxoYN/ne
3LYNZRk/XvIbImB7cRCfXBjWVUvHdNSuBCqAT54rs9bca8fLPkkRAPL23a+Ei40m
GdrPPKbwo39RWGzYB8EeHpIwfD7z9ZbkAH66V9AinPg+RR0PDWwfoeBT41pdvary
VHJLYKnpp0AX7pO68Xqdza/sj1Xf7irQE1zOMtj5jwCLijrh5i3ecAgxWDrYxFaf
oBxFqPD5jfDU1vOExo8JGuts/mGncGDEhO7zf4odno9lSHcV9lAuTxUwykrO+dtC
K0vgb+cldUlDZwAraj6F5YN2+Ds+HpcZGmZZumLINi0qkXICTbvaR7Y5D9tFp5u7
H+9nK6pk0WDLkNCqYJQAuTEwB4wGKM7Uy41hakejJ9TjWWgEL4Q/R2ExgO1Kqxnf
b2dCDn9rb8ucbT6VIkpAvXE2YOIts11u4alRsIL+51CRy5t3CCdZ47XeUec+xGZp
OmHQRm6Pn+YJOj35quq4tRMGIfCpr3yDPxEYU6ul4ra+58cJNrMZtgdeG9I2oWnO
AHgrvcC2BBR33w9e58woer4Z4rvSDZgX9JdNGt7c26NyRDRb/NquwN09CbeWb+wJ
s2oQQYr1Xj2Xp3WHk+VoGChmLHlkxET/+I+Crgc0s6v8pabyhd7FFSAhchYMntug
XmzcqsAhBh6i9rbzIgOdL9wAA1303351tCgydJ/JUzruS2Oj4KqgNlTFvm2DgPcR
MBdKpGrIfr2u7VfK3Qm3WyutUlblplPPx+i7ahFKtpOKqwvBarxzD/cs5Mlh1tlR
Bxd78/swgoPTl8MidCOrN9wBSEsaIy0aXcgPfScFWKeK8IEp2lg8JRSM6qmgmOhJ
chMhv0WfHpLM4HxSXC1df4LoJtzoIpiZ47e5FF1jFnDzC5rg5c42Pq/hEAiSZZn7
uGJ3oM6cvcqWPDoWZ/Xw9PBlr1l534CjnVgN+CRa0R9XEaPWcVLUTzC6J+3Wn2ph
8mfDqC0MUq/6A7KU3ffu/T2dL0lwzDGl/4gHz15t6u3w3vAgBiYgFAqJISKf3yY7
YqL4fk8uKBCBMAmv53l/LOiyazGUkIsLjFKsLRVb5fN4yWzT/sCwHH38c+J5CBhI
Gc2Pjc0BwucrwYeV7IRjOLEAdTNYIfzTXAIggifh1gaCkxO3vZtSk1utqwRFvkyC
LPfvQ+FbhDY3EXAxT0hcBRWvPZd7EgeMcmrzaQWXp7h6pelbbK4MF/faG/PfKIk5
0h77h+Q3vcWLLzkYpEYzdheazMFwnJEASehjvL/EGbZUnRiMvsFcw3aYoF3dsZCv
Dc9FzMoOJrs+VYZ9xuauGSPRaij920DAooz2rLL+/VpTLuzbXjB/PgKSWaWLvzlL
+JitjE3ZF/Xgt4cBuMuLgCYpvTIugQjFs0UQh/fBNZf9V3f5El9CFrOvpJpHTcig
sEjr+S6/hFYrqWsBXLRkFOFPUo5855SXAxlZFuq444FJXOD2Rn096+81jQ+IBlsA
po3Jg9+gKTQ776FivOrpgzgRfbkdLolwass3ZT31t1giVupkv4SMrxp3bXY30tnr
GPhSZLdZjtvHOT4kjKwZjBxb0m14bQcRL6+4ZIDQ1sOQuWvAwY7oqpJERVyfPJkV
JzV/Az/AUUuV/u4DEcWlB7uqBtnfQ1EtBbE207XmoMZLR/moa/8SBCUY454z3IdY
Fa3YNh9plMawTq616iC88bG+kGwTz+4JB+m7BjfphqXQTvNYNFbOvFbvCKs9ntn7
bFG1J78ZO3pD9K+1qhtxLcmKd4mZSwCf+1pH2HxSdelrwfAOSn314P0u0yMtdJrU
FlTgHyTRnQpbscZH8p8rMKDujlBhyg3K3oWCz8fsy2UO2uG5Or2XHGpzaE31uOSD
yM9U4XLOHrJETjQ0BS7tIDCb/O8T9s1ldZl9H0Lv7T57Og86KLQVe73O+J718nCI
yMRWeLyrUqwswookou1r7nq957U9pSz+ZIDTXKq/O4Z888XZ6iGy0zRPXi/6WsH9
83TKdX4IIpQSpop4d+E+qrSqoNIg1s49GtYVTz47bXDKWYLYpgPMGUg0ccKCby/9
9XPD4WWg2QEGPlkjhxltdAZ634rNIBgzFksN4NNYJi1UMWOgKw8o1KcARTGFtjrK
oqSzWvBx/zl50nS6XJ02vvqSekDiQ+RLk07Fwarkgzty+pNX6mA0BxmZSu3ANnXN
javMSrmJtXC8XBYcj55GOpusyUW7GrhkS6tWMIs3cC+TpLXw8KwfNx0CaBAylSVz
QA4E3XzKQsGp4V805GSj0UKk+JhzmGZCSSsb+0rnxHp0Hfc0Be/Puy4AJ7dRHkMe
cwg0CignckRtLsRp8xwt8zGvani0cG7mOErIi18jpoXZxPwQXU812st6Chl4xPW4
TZWw1xkE4TZE+dG2cye2Rex/mm2CpG6YpXjtb3cD5y9FplxKk1tz5TJaj11pJO05
lYLUZIYkHTLB3cKMrhd3UZ0uRmiaIbeSWLcaqzXuGmCfS82XlwpqvfWwWUuKIM4G
lKyVuVx19c7CeBe2D+gfxQDazVuJrtOisBlNC566OObsYVtj1FTIk4/luTlMNmPz
M+EGL4RKaN2Xguw8oMPO9WU+2nlL0fAPan0jCdTXLdLw8WNjqgY4884gQHESG57E
W/o1XNiqEf5HK9WVxkgUiqjHdkJW4+t7ZtrEHUVyjbst08HZAYLa7FC5HTrdeo8H
ApYq/kNTzJnNyNAn4+BqemAnbkQcmwNkNRuPqYnVzaw8sLkfLdnGjIHxKY7UlA1R
Ko1xMu/NCZ+R7c/3r/aHLxBkaZ3hgRjiQHvXItOYuvZd4tk9MtF5XvWEhPRC3lv4
m9Xn7Luzi1PgvHLkgA+5dL10C2z+CoHsFoQGM0w/vXyiElugY0DYj/b5m5NdJ2wN
mJQ7Dzd5odXw8QK0aehIfpxApqRz2oWlSZ6dEker2G0ZNz2bGR800B10d7HAJRLF
qXvt2J0Q3/TMo/kGtpU8oeO0RPaGV0SKnztZKllY2lJ3EbvW0TxyFIykxXnQhhK/
Gx3IozHVvWD9BgeTdzs+V6cHAYCqkYaKqikC8qghqMXvGi/hBCVnNwc7CMT5RqMV
SX/7pD6u2wqreD/k0cuZRx52FtJScmHB8ixEJyK7feHxV71gAfxWbF0mRd20E2nB
dj0O7OnNmJNqNA0n+sl93DF+QWirbpsPFt7SOg0fgCeWR4UbKV9NgWdr89/oRjZT
PEEZ2DYPGd4raPvQXMVA6aoh6Vcb651QM28km54ukJE6g7dAQlm6K2eHC7lF1PZx
IxXMmVQgEKrwWNbjebUwW5RMd4wImQt4yU5ACVeTZUisGagMZVGw9j7rxOTsp0my
b7MPxJ7Jl1w6GnUMuySMmqoDGagXoQXb7nBvb/N96xB7hBy9J+2BFUaCsi7Ctjfm
DgJzZMnvo2prx/P0vv2rPZqW/ECoLiOT60XVxgZzSsWMFG5jU0CioBcYKOwJ4gD5
AN1IMIg0SQDf8/VpLEGDmzHMHognWRjScevCzHeIw0Y1jyTdHFQYqyvFMOdftpwH
ySSnZQSgKJ058zUPlmszkvM3Ltnt/XeiY+yAHB4oPAj9uYn4xsEXwDZJR3fQdLOL
yDZNERV/ONoe14PAnTgpcUnikc6EwcxngB/P+9sC/GS/NGbYhQkSg8O8ouUhfVud
P/uWEXI33vOA8Dnpq2ttxFAPF7FdyMorPQVgrRo3J6QSWjJamR2243J5bh9DCXcs
+rpPAwN+Qi10nGK4zaIDFsbJDgmhtWtNEXhTqUaoAt3xj7l7WmA7+Xcql38zP96E
sQntwyhQtbgh2Be0QP6V+mVhfxQV6EXErPDPT0XQiUDsZ/75ZfgLjZTTmaNn4U1o
HQAO8c1DSD+aP0AkcTg6TBoWgZ9OxxWPRAKiDT9prYPWmuScODKk/BCAXBVAYvw8
iuJ6kX8qW7AZnrSge5SyM9CpUhlcdU8uKioFjbWRr/O+PhJvXBUaLFr2eX6ixdCp
/+q3Kp/lvqFT2I+wB9Z7md6hLhXqw0XzQ1uJl6/vnhhil6IUXw1h+Z5bepRcrfU4
N8axE9Z7Xmae1x7hDnVhxZ2QbQzYEZsVjEFgy0acnWqr+/hWz5wn6XT6kKQtKCYE
lsoASzrnl4NsvtWkQyL1d4+OxuoOOdiDkuHHOgTPwLkbOXSZ1IIyA+wJzx/fs3Dz
OoXal4PD287zpq1vbyq1A/3jECzGEtm3bJIAOXVWt7ra6Dq7je4JsSmUPnEuqZjl
h/zLiP/bKwKWX6FNAM4EkPrkco+ZU0H4wan7XYoUaMvicHY9nTypEijj2iz35oXM
akzDkNq+gvWgq4kpWYV9N12hdSwx3kOomvaHAMzYUzRIBuFA/t35Ifm1JnpRR2kL
cDuNy1nsUoeGNVxpftFnCKmurYvS05cfPHkkEZzqhcoKDAEyAduljZTKtSz6Xr5H
uPVEFJxmEhFp1mtP7y5j7WM4Bkd8ZKAramEV8PlVyHyt+qKKO6zcpJ915hMfk2bM
R471Z++Cmko8CSjqTvk5W4pe48voHek/thhWtEVX5RxW0gEd7H55OQlwMEvMXUiE
SIioCsr4bXqtuhO7sHW2u8egQhSRZF0etOWmxwqh/enkv7RhojW52vQUd2wxFfr+
ET1YiYoYYKpr6a5L4ey8ig6NIUhJq2OdwdrMHP0MVX8DwF7lY9FYdkq898K7j+0b
hY/vJZeYXaAKfzC04Lb204z0T3FzsJacvuPSZPoGC0E2upE4jorqp1ROEbzQZJ1u
c3mhIKU2VaK65ZqdU6JDhB1g1HwJpnxxkm13u7NMPVvue1gcNUqW9BC33VQm52P2
J9+Jo8aNHqwvsHwhRBZiXOPBotWiuGfE1JnMhNWzDE3+3c6vIgh8cotF/S5QuKsR
X1oaw7DeLeun1DTo0ufI1Y8IkZi0aaP0k8J9/yQxaMcTNFxgnYoQ7Hhv1EqzAMv5
vlnO+5Q4eiqi6d/pF1sZ8NCTmJqoo16iykJHqx2QpyB7wXAOpsQYqxItjbmThgXJ
ZIzDSZghjiHbSUqM3yJ/BzDPh0o62kU3XSG62f+CLSVopbN0R+iiJJR2H92P+3pb
bpcZKu3cpFZnGW6GlY2UL5jdxkMSEpjDCVWryNsIDd85WQeJduXdUpf9I5o2SpOM
qNrV6xrk1RSQS3c0wJLRooWNnAWpLWzxBFvDQxM7NzK9u1mwCfkF0+9YfrwJPFiS
RkvZdmxHkyuyX82OOXwWQ9MBhhjaYGl2fXrS9I2p30bWTqsieqk8OBExAI/gADn9
32dS3GuDrBVAGZDTZo6SjWw5A41SQuD1nVRY7oW6N/1ukXMqzOBmxxTjKEKaQgBO
gEMLgWqen+zOLR1k0QqdGbC1fVHAEP0KaPsQEIBzksIZvMmt398/3R6sZzHx3sJr
9SBQCRwpBE2evHQnUfAsGnNKYkIaGN85EY5dxiv+SbhDUcfhkou7VkcNhM1g/nPZ
f8hmyCntvhdtp2d+q5YbGPZDA7EnRJi0yor42QZoqrIdSCK8vHsmD78B72g8ORTV
h2nlvIPOdG/vJEnRD/l83oStHqL1DbVr9GSuYHEUBbpk370/pwYJKk34JKwGkwBR
IKu1Qklp2sRNjwLMSm0KlopWC12M5/3lv/nrN1Cjcmtgmak80pOlKocJTg2nIauX
7S0lXpblq7n6WFBApgnCBHy8oLBi7E+ViQMMhnuNwCQAzIfPa7USpdeEqhs68DOO
APFWERquGu1F7cNLmPoIOGhgncvMoPDhoMss21Ks+iozI9JOSvtWaX+wrC4eFewv
QhY0uOg4Yey5v8qL3sKwOjZziAEmFYdJOsm0jiCIIGCUunGB/wEbOoSScR/cvMWn
WSY4g/bOgXY2ad/sVVi7KULS0zZG4CH6pozLoCpR8RlcfTQW4gMXTfUNyqvvVM8S
Jm5vlTJc+138APumldmAPLy8Fi3mAckEwmnDu5jVQPTDUbX0lyHIdjUzMqzyrZll
hd0xtLc64EEr101ApV4LAr+4HQi0DmusFg0RKIaodTFLY4+Th0pZxwG/DdVa/OVh
0ge0Wg3LfkW+j2jEtPskLq6bJBgOtV9zn4MaoMsYieUwgvwchDY6i0dWhXDFdElM
O4d1XXEXSAoWVrgW9B7MT7nV8ZPLG4B/ZW3x6hzR60CbZtK2ehyJN8T8iq1lxiB0
9YgFurqjN8dchHt8LgUJJuA6gUefJuMx/KAw4ZAaskHzd/hQ4JLT8cYVyFfLbMDv
XjilQ6QcjR/S60m4H4pX0F8QpAbWLt9LKM4eXKDEAc9dz/R8qiO/CS8AI9+zky3V
SK5KF2Dabqb3fZHady0MCQUjGnqrU45a9J9CN1X8F2ZYCXV538a0WfYiNjncD4h6
LfYQEEoGFW+VzmVdqx4f4YIGoPuM1IEBdp7YHNdmelXMV+/ebH+4XR5ASWyRdysE
GDHQJ7Cdhzcr61SFJ+mkinF9TFVsK2gyNzdSFyHkMz/HgSEY0lfql5Y3ZfZWmbxR
G9SFLN/ThnrJ2om/zaNq/pH9ml+ELCJ2zwn2KRgvZRsh/WvabCB44qvAZZdiWzJs
uIRQOHCBlap7Pj5iw+qj0IgtrsZV5Ym2bfKRVQC+03cuyzoMDJ/JCbsHldE71KBY
5snjNpM6Q3WrnnYDLzU3xnPVyzPfLtzVNJ/ndtRAuM99CeodtxzbQ32TRg31BxbC
hYZIwo8ziFMWKE5+GZN2//VTWBwD9bOYmLkUqq0mvoIskJELirHs+kqv2X4bXuFU
1gF8KzpLMRAb43nMaOusX1VuBImH3K15dlOFsUzH9lmwBQY/WlcGQ4efh8XrzqH7
0Yx4uST08lp28B5Wnfmp9Lno3HPuVDz0RhRFEQyfBUkW+8lVHdMUvXoBUJSM51HV
nxQkyjY6eUDbZ/3oj5Re6+6MihV+uH6uM1lXIdXGSqC8MX8onuDBf6FRaHFxRr5i
g6rPH/1dZU0yibc8spQjpYd0oIX16DhVFzg1fpcFz9o6fQEpxf+GK4dFierA2wJr
bHJ/ePc/aTeEPLx2KrWBAR+jt0vYYot2nD+BclktQO+liZVxlhKDk62GNWLZYgtc
ELwE8q48ePGylUNuakR3sb6zVyRCFSfp2WytPnI4Oibg1lknL0yV9uS9yRNTmK3l
WOHFJ8Fdx/JeliX5bEcnuD+cwct2RBv4MJhj4sY938sA4tp99lGlvEMjG9JSokeg
Qr3q7vzlBg4l6nRQH4NS5ezUi9L4X4U5RXTE+RsGTAuLJ2NCe8Kk2ahjLy9Kok5W
O3/nSKoeFgjUvB23wjWfXIuntZAl+tSGEdhFlK/iC2ijxeIoShacHr4/iPTzsho9
6W6aPwGo78CLpxVr0ZZkyJ3XntebgNB8grvr89i+AUHlzCAHkXkZxz6DtMDObTfH
mR6Ph2z32mH32Zi3sHTwJoOpXksyz5AdVd+wGUIp879yGr0n0PZjkUdUZ+qVo8rc
kMrAKEmQnLScqyv8X6D21VwcCcVZdWlCO42XcKgFAqrz+l1izAmK0n5WE2zJATKM
RbE4m4KGa86QMNa6DdfdgZ32d+fIhBs9OjV5eQ0EGk31hLxn92F19JbsyAZUQT0b
v26YbT4gCo9DedHU/hvjHIjOn9Zr+nTq4kTUleIHXj2FUmT+5kJj4UTLAL3SN9nQ
e8oy1z0DRgIW9EPm+A0q6IZfCN3oWL8ztvJ6s9xNFRXJVTBua5fTSky1qwcZkzkj
81o8HO846IPFr7NUl1TFYnZi77epULtDxr6II06g3tD7jZDMGUwNcrky46L55hB3
1CE94P5Se3tGysS74WvT1Wi/bF5yj8GXconCe7CvSJ7CpWy0r+bPiwpIfZFv0vfZ
9dZzf6IwAGhgCJiYVqMGx6woqc+PRQqzf7iRYhBcguaJ5WEEdtT1QbvVEK2UUBnQ
B6P5F7LPma6jUnpj8cGqniAVX4BvRy+wmNn317tZhc4yDFmyllv8+J82hnVCHSPp
YaOkW0sLivoy5tXXhQzrUq1hSABsEL1SFQ0Nay61OEaLEyhAsI1+JWkDrq4xo80c
l31AryH0uNx2JeNVjrV/B8qAcSFW1ixVEbYLLK1DLNqmKON147Bol7B3RrSdJCyh
/PeaFBjUIFmmDJ1gdmZfutmea1QxZlEey1bzoPvwYrRNxZ8SoTXXaJCi2iiYaj6K
YdldmHvzVqkz462DQMzbcw11MlTC1U09wKqgPJQ33ffgVm5ZSNpBXVMba4qjlqJr
IB2Yz+sXVXPSouYHttNvbXUe8sriPFMjiK+x9+bs8fbWIVZ+iWU1vRBALgzf8Ftx
P12Xl9CwItV91pq0s3qHOJNaRc21v2trwRpq+oJmuqmdakr9NquwEYzxiIp0KEsx
i5Mu17LtZLTpwgTt6eIkCaQ938l95xiS0C3hGOoP5Wf64E1vZ38P4X1E2/6kxp/m
2f1p27gi4Txi1e0E5L7WwbqFPX2tkZXM3qk5FR0jU+3d+PWebxommjnXPz/9VgMc
SRx6Owus2liNQSTHcIon4nyy/tcaPYDmHL3uXcdgil+nEmHaznBcaVoA9pbW/vm2
Q/EDslZBCavm0wIvYQ5zr3QSMw7NeVTopXKW7qsK3ZG75flTriHeyI+VG191q5hQ
Ov0n4Ee2o/v3rwkbgKNHOg4l60er/yFq/B1IOaRpkcuSdML+973Kcx/tz4Uf++3b
fWwuA4ifqZHQ77SLDtwYcw6efvE5ifnmm5BCS+b2BKfAhOGdP1FY/+XCjQ9yqsKH
ngQw546QrDw/DREiaPuncUwvKcPJUZkvhN45eiamnzrTNR2EQewYhvPoaNxJ8Qwh
AHQvONXk8EonTk/N1TtzCUnLS3uXx4iJnPXis+uPV1A2wJBVPx8m+y0goXNObtRn
PmIT5KCcgSXSZr+x2/zfhaus8OlCdSX+5BDg9RRTTkTTjywYJ336OKOH1bbhk/pI
x459K49s0PCv9zCpqsXqcbzqjywn+I0phJ4BTGoTokoYqx6Hd3Br+AGdpLHgu8QA
59GSGNKe74RVtFMQ+lb4eLKr3+ivxd3TQchJi/SBtwwjHJ2jmtmdECYgJRo2FdVt
LWCq7b9AmqlKwczXsCION6pKsozDB7qK3HByOL6xYf6VEczM256UKzSyTiXyKCQU
gPfrSuoOWvHxJqNdPO+xRH0Qo/Yr8y2J/hOaF/Gr1jFiywhEfWURyuq6I05bdH7p
PXb5GlGxid15i4gwB8yVDUBLjppMpZbJtauBYfQY3nrk5nMTPqbI3ECSrbPL6ArP
VAuC9koEGOibGXZrYm4c/BceNQF6iGgNMlnnSn6BjJRv34R0sE8DElwM2lq1h6Q1
24D1s+hqFSd1rLGKMiEL26xzphJFfxpJOvg4lsBtBmgbDmnSgSPMOPAelVLUPJC9
hlMtv2+Qp+qwDtVkAYbLMxYmQa4GNLHtBatNJhXv+WW1XjkKHLxsFpjpst0kfl44
TYF/ItBhSOsqVU7S8anOWVHU3oQnbwS1xhdj312JBHHphxKAWAdTJ72hmv2EIEgt
jI/c7aw6alB62a4UI2cjGET45Ksij44WC+1SHcZ3Encz6Erjmj7Ja6VstH4BKrrv
kWK308sdtABg7Ep6Vlj+FyYwp5duM5vpkfKy13/d5cJyisJYdH4zDQH/1gz1ysRA
40pXNcXXv21io9dNgEJtVGdylKRV1nTgNrHmPnewMO6MeZlkhUGkfafTECNDG40r
EYWrtLv38qERpbgDGzAZ1eV1KkJsknqDlfWRZWN/JP2Crwla8lJ4Eza5+Vo+Wncv
ark9uPdnLcGJEyFtT315AuEKZyw6grDa11N5aTFtzK3X/JZAZegh/waKqhkNzoBX
ZjbNsmkReWstQKFdzKCVIJQWabPfRLgfiAl4TfNz9/drVpSRCffVdS7E4CCRaCi2
K86D02zfIEOdt/X8mYYvWWJHWeZqMsMrBmj/gCz+2bXNGutqJ9ESAS1IGcv8GbXP
IVytOc/8r+vcfV/v35KFNT9p4lxonO/YvNixtnTiX44K3Ug9MoDF18emHJBtlI62
37O0bTxZpBvqNXa9gayb909202vhxnWq+jlLBmpJOUnQJ2q6IdngRlRVKEp+73Y6
mKd+tA/Y8lkMm8V3xT5/ku/Ssy7GpoYvuJdP/jG7bWzi9jJKupC557wi0YxPuzyJ
t+Fr2GPr/h08HrsrOB+38W4/TmrirId6Ch60sA+m6aO5VV4D7XtNAqMJizyRbDIg
Axb5TzQR7nd2I5N3i9Wl9BbDg1uHfazAULUZKvj3UAmSB/D1jWlbRvPfOGLmYywx
N0q8xN/HLX/K7pgAti1cSeM2j2Msm+hfA/UrnIKLzQvxwH/oWWybj/KiBGlhfydl
zlVCEXcjLbA2xsjcdXLl9EPRKokZGDZnqOf/ku7MUDjOE8UDUTr9XB1or3I15q9O
+s8lkDzCjF0IrknsyTWUMnsoirZ5qmzPAH6lnfj5RdRghD3IdGVhPHmOIzx/YX1F
lVaHObpCBMoKj7CFj/s1DnmVj3FhmkhhgY9gWzP0kdp0Vd9PV7TshTnz21DTCYn/
DM2DFTqQeEsXWbHy6wBUP4yKTMSGD3KZlk7YgigrY9DY1fAw2R8m04+YJox8NxZq
a9d9AsHP7WPGJd6OsqFni+I2/sFd63+IWUVOqFIPfoBbP3VCLpZWjyD9KIHbQuB3
tWylRVUshTkICFadkQ8fuP2eEnXtkDpzETPQVhD76E1rjsQXLmRcgrzXP85EbQ6z
mKiQ0X18t9fs7j8DB/5N6+AZpcGxmCZ2EVIoUTK5m06nos2kiLdKEB/m/kgvSihe
Ufl42Yf2Kqy/qtLjJFKlqLBibHrF0aWkajYoy0JQ9CYqLWtDU0cWRMkaEtAZAimj
KqnBYcmZvi8d9xGSg1Dyl7hZIXjm09AMK/iQAl4yL7FGPYKAlpzBTsAVIkyME79k
4o1XG0O5gImgfP/lTqLCGYZHt/KRKKyOMi9BojfPfrWs+Jlumf9dqAkhkKnpz7eA
38abEoq9pQC+bLmxq1+FOtGaxg+O8kG1o1gGvmS7Lbv8ux1X6/6d+jFqorV1O259
PiqDgxr9HWa5gGe9FyjBT3pRSAvPV3rke13hVGJ3G0rlZiM5C2H2W1sXaTVOGptR
94BDUWxYNnMD2oP3bAS1ed7a2YopozmtVPclDozRmuTB/GTHKs9BPpgdQgTzasn7
9qEYTsyH/UqmtecGw3BW9/XsSWe/igLjWao9NxvXARbHUxYrwXCuCNDDBqbX01Ry
xTl2n0bn1QflDVjmhIM9jrMoiPdbG8/OgOcqyOuXPicenGiecZ7LEJFTcdZt8p3a
GBeFY5opX0dczgiQpzX7gAK1FTW20hh0dymrVqeadony7YuknfuGdH2JAB9cFUOt
jt1OtmTNhicucCbajEODfOXXIcwqqreKOBTYNZ4krnBDx2vyDBM59Mxs0YncIHm8
bS3xGvfYPrAmaBy0xLsh6SfvORUTM9dgT5h/PCPT+aFzQ8xgqcKzbksBlTg0XwCT
J/Rq43sYjDvYKsTHuOBAyqxI/5j4e5pdknJBLBKb+o9od4PZ0WIqwyNExUN3/NcB
PvvXcEvI4I/3W9Vu8BB8t20/KJQTYJ8Ldc8o3NnA51cPZyOmkIOs86KbIdQVV9ZY
JyH416D/2OPtO5HwEd4Cg27K8Q5HLoUgsuT1+GyXS2GJY/+0xYNebLmuWiZLPmpd
TUgImjIs0cuIdJt/WyZxJ5nq8R7ip+iX3dbYh7M3F0gNHKi/x85ZKfyCYcKw5uku
cKJuta1NhG+0hjrXxtPgKFHKKbsqh4NAoqAPMRVktXuyQRUj/SmXcpgJrs2cnzqi
mBqGQC7+el/WqUSqLYOOaMJKO/JgAV6hdrQFEXSTuTGDD8UPr5NZ4/ntckqYMYRL
hOpUr4sOjN4Pr8Vm775nWgbqCg1qgZ0MBFgoVRRLACZFzUxcOc/DTJ9QMk+SaMkl
77YiVOWPk1cOWVFN/uGwR/iEG2N6IzudY1n6W05eeAa0UrwZgxGDfT4VbOyNxjs+
nsRwTfPGhTwiZZExZaYCyqPcOT5uiDBmFEQgH0qtypCHihnX9SgL7KNGQNfBE/Al
gb4EfHA0wTDLuYdw7efTY8GmQ3emkShnRY0c6jqlsbiusfwtqLG9u3BxLDy+i0kU
ZakDvgamfy9vStt8cnNiWZ6lkNoIyyiOdqIo5+RQgIn4xfDxVmvTjoJbOFH+aZ0k
Oy3mEPna73fyswBsoqBM5STidFu0m/VW4zyDKjW47hmsjF8uX/2uk2zPndLEOACo
ddEByPr45CciVrzCuCzjpWWGbgOt0Y48DB90Y9ICA8tiDEig4146WbfcGQYDg2Hw
aksGfY5jIqp0mkX9S0pAwxjkUdUUaBq3sSyaCeyJn9ZXakgwGZ61jQ1EB5j4+TzN
3Rg5WH677nvYj83TVZ5bUG96k2aYY752KLquHx2a/UHUh8Mq7SqfH4jnUOQXyh2X
wyZQpgZMou+GNGWy+rj5zV+KqQn04AoLz//mdzBEjd/a4AKN8AE9uyM3Ruj/Mjtu
n1EMsgk10U2ZadMHJmdjvxTAuqSVTtMIwOcxPkqsETURaad4Qgu/w6VTIafHHsKZ
PV0uRBqwwA5EIDR89MlsJy7RWlOAgOLFkm3m5dOQPEXVr78meiMIec48AiBnX/oT
3aBrqFLYsF0XciTK/JFkcepfyFsUaHEHt1momPBEP0Iocqz6UdI1K3hmR/1Q1bNh
ky1L7jwx1vBDHpVl3ZidnLkn//LTb5tUe6/iQIqX1LOfEtTTTSEYhL5fOg9H2l4y
R5mRBV1c1VyUHMDDkNYn2KqrBE7t8hOZmCXrsfAAu/iys99z2rlJGLLG/1c9lXC2
+PK+T8/1QbMVI5YsCjPyMgyldqfCzxKnx9Wk8rkv2jzQIKTwC6ll/ukjxMClff9k
VW5NslEBZvMuEXESHC4pIvocqJUJ2nCKIYEP2X5TA7hB3hovBfrHfq21XE7IzMZz
7YxmNr24QTgZoMDBT9X3gaybevkDD2EjmEhrM8HhzxEPoYwzGzK4Co2cAtqvgFJ0
TWtk4dKXJQvO0vDIqH32UyoKTNtzrA5qmavbIYp4gaYgDJxSpbIlPM5Veqxv4AEG
zJpePa7lBC1guyMlkBzbOMr9/g16Y5orP/nO63ajt1gTe+FTmWV6YvZ1ghBETjyr
cHP0UmXoa5BpH+CKhkuAAucvJUDe2a/+PQQVrAJ6duZHh8NBkf8qeugre5BZqdGn
aGTJOldDyhA/NlgK/xD4JTTSROAfmwBCg1iG156X7806lqZz1k7sznm0F4EWn2Hf
71irle3D+bT2nIGP0VEZwlz5Ef7j9WVa2gUCBvLo6XIUo9/ZDo4ncOjL7WS5fTNw
1O6DHVCGfioOMqIP5XNddgkrFJGmustn8fN6opRwjCo1uOu3lCyAshKJvXOPV6qD
D4Lt2+/dUrAbQlLdtb39fMeRXfDvPqeb26dfGg1LkKrLJdrVWgX7S4ugKOvHMFDa
MHzz5PMqAaW2tQBk4yHy5J1yMLFwuoNxt4YbX6936LEb4aD3leAWzdmGw/PyM56y
gEpO+4TGrBsi0+B8I3vKRTsULyWMHnvcsv6442LqosGJS4A6cMIXUKwm9FJBAqKX
l+o1c18IdAjRsKvxgyDMdrUDdBsGFXEpArKvMtOfaZmfd79eO2lmHRvqqmlvi6d+
F0oFYNpt9fJzGSkXKUmYlwlpHDHEeCA+9nXVapOfJ0rILKXyDKF+uQuPCD6sGwvI
1M0WNeEdEr9ub4Ut3+ZGPmYtZCeImNv3r5lsYP5cImTaDC8HuhAN2VSlU5PTqxcV
lNBQMSMlftOCmN73N6wZk5i9kYDZOt0U66dKuj0PehfgKr+7phTUNe8HqWZtKhUe
mYJvkIMiFrHg+CnDp9y2axLUxJf9iXAAl+xoN9ptX+Mqq7Y/HUv0SHmAblcs0iJz
LFCVgd9YArESjiJz2J3O0F+j3x4lZBpFoth+1+YOoHZHMXRURTF1zoLybOaPSK2W
AZIHB166QuYcxJ7hUeiC5tzqjFNVv0UJyR0lkAwFtWD3rWDRNE87SJof8UuGGToX
TplTsPxMcDy3DFY/0hESJNjAB1Ck2rc1j33NfFuQwy6bFPyya/VHY4mfuSrU0uT8
vHZgq1hKQTFGQjHqjH2P4ZOb2rZTWPD2ZZnRexyHfHUr2V+yRDTgxdG1ms93ptJA
Ac/LntmI2uIOPZ3WWxuIezUQKB0Sb62bitnUphMeJim6aYzuFS9/JOAJ3SXmV+Ut
4ulPLT+3b+UkyrL2L5SSK8Z7T1lQMhpT94S75ArWNOMQC5rmbaRhrJiQSIcn9eHM
wm8wMc81ovqvfjBReyMRJmj5WUCRZeWVw6WyiYsol3iPBp5yUjwgRO6K3DBLHQrB
JvCPaTMzk8g2nJcDtva17EL/xsFDra3zsRIJuj61FgJVGv8PmcKCCB+Mt04x+anu
WvqAa8+W18dzCosScHt8KR5ZWyBxVrIVeMNWWV+8HtI0XH+NzWq9hWfJIoBvzX5P
XXhoUT0XBBvbDFyYOlz7pAO1NAsxao+eF810nz6iXh3CrQI4Bo93AQVYgJg7VGyQ
vlNKKQ5vPH+qVzSrv9OwCrPIWHUwVPYODSfVBiGIYoJj1zzcOwXbiLLtN1oPJslG
NpW401RhgzPjpLHwRz88M+xtVBo0pn0GAt1kZ9gxCwYLvhRSroPnfNlB/ZBcu0PR
XlXzVNeWv8A1JR2GQr/GSAnbVd7hypGouuUsyuUIGrG0vpd5exFCX8Cjk5TPm9K9
qj0ZEyVjnS/JfxEZCaPkhIIZl618Q4xbwNQVsI6NunADOAezVsD3VC2rpJ9dUvCh
LhZtvaNoF748Hi60aiTvcmoAZgzoDe3txw6/0S+tDRi4zZwfyDrri/z39HuyoPXr
vYjyPkb4xFeJdoyrsUvELlUNaADP91XGUpjJKu6lpamPQ62Sw7GOtGyDddbN2x05
dHlkUVQmEDKBdfqVklxGblt5cHR2jPrSYTl2m5TMZWddVQH4Pu2HTr+5BSTXFywO
Yje2vtYq9ev3MY7yHo/rQa5dbh9B2KvkSSKVWoXmPCll1iMYXRusPnK7F0pNEjTb
0PC0hEKx4etwC9uHjJXckioU+UvbUxMiLLCBUxNtdz3F3qsbXh1z6jntJnCX7sr0
+Av6ylk3EJ0ke275b/eRAmOHXHthI7MaBxT0eLr9N1igYkMjYvf09iwQO44y0yjO
ZhQ6KW63zs5DeBUpkEIddg4YtvZLGSv+i/kkiaTt/qnzblp4LlDyHAwBcli2e4Uq
qJnsZF4dFyUqmOUKKxzFGho3gO++1JOflXHrCvQnPhO4icctrt4rFr8ufBGeUKm3
IAl/L3yR8J/2KVtaBSp7zHXXsoB3cQRR+GTpjf/8v7KHw2CdB1YjHmLkpEuZx8Sf
RBLPvIsZ9KKCllpbpZtmZuH/DCQXCjyXFvG18cQbEC3+X4/Vcv8wqPR8mD1iNgdg
vZt2OoHpe0gQuGxZ4VwZRHEhfVzUzeDwsW/OlhRW6S7T7V9MjkPnuoxCCyzNdJGQ
FUM4BpPB272bmsPj6R5M6P3WObbCgqGcuKSxluu5hJko44PKqkWmypvr0Bej/8Y8
gGWrvKZEyb06cZe0G7+UGLXIj1u0EWmKb0Q1s6hvEtpsAb+UhRWKz3H4TdMwL2fY
qLqHOTyHB6XzBkv2mHS4VTEh0qBcY91UuU1getASsQ6OkHOAs+ApJV2W8FxT0e/+
nccNgYWRcrOL7Ae1M9t32Dr5h1HJY2kYaXGmUtbSABgoYtymiML+T8yIZJEy3c/C
Hmqyl0xU8be4WV9O2UBssuqj8T0vHGF4fI+QbPKZK8EjclSeubLn99w6PnX+lzlW
L720D2hiN43TjBY435LK/qN2eDrN7w5UiPt3k9Rr8tPDwbs2+EHBDhgtI33Mmc+f
a6M/TdhREEKkyuKmA7f/C3IlmjOrOwbdoQOT29ho6ZW8C/tg55OQ2yuDmXMv1bWM
v+wJihdIv4BpdDN8Yg2fvciZ4ATmHmYiK0HjyTbC6EuJxih6Jva91ct5giVC34xH
NsOc78qDTjSqIiUaF/Lbqwo3WOtU1CEwlDptMx2jBzDYjhhfB3QbZv0YrgMMkzLd
usIH7mU+CtH64wvLjWRDYR549G4lTk9tiyysc44lPV/dOU6kZ29nTANzan7sLDSV
ATHVpzGi2Ls6WLT4IbNG9v4DbwErC4xlT8X9RhX/3P4DE7UjUSmbU6lVd0PE4YHY
Mj/mZuQMpXTtzwQty+Dzn4TKoKqz83m2lT/qJJGtZr86HyR3/ob5v3MhUvnbp82H
EBdkWgjQrBofNEezvUC5PQyXfD94Jr9k/wCPpXNCMdUHVouGh1vEjiYERWSV7c49
LV8C7hrhVKUBn+kS2xdPoulM0Dql9YxVxthNkeyxMRKmi6tvKauIWFebjXYXl2gQ
Ugd/I9IeZ2tyUEkNyN0BaiDOWwBPBhgWx/4U4kkpCQO5y5oYej5GICnAK1DoUVgI
BUG8L1mZJWe/4KY5yKUHZgKHZDZpJcgMuhSEITw8K7xx8z7OB7O6kNMZ/iQIDNTO
QXOdm2E8ok61MpvJzY716iHZBkJY3HKldsOx1o5uzzOIrziKc05SGeJEboG0QAL0
FBkpzLaI4T0P7c3vTFCYSHzLFlZ3+sq0sWQl4KzAmOdSWISRo1dhE8L8hb6vuCdl
8ybgTo2AW+fYtaeohcW6qj3GQ+lm64LaKVFGTPy4xGy7B9y6RvTjJ1eOEUcSpSnz
XgFFetO8H3J+gOY1Zpz2bfLJL0YUPI9kxM+eySGUa9YyoaUbUiLt+NUBpIaOQeAS
uCM3Na8ah0E6sDGGB8s2g0VWTiRDRtB/hq3Iw+4wGxPZ40JNRDfYXtO09qiAF6ug
SfL85vXr7yB9lyUJ7PbIMMsLsxY/oFkkF6fCyDLRc+QYtmUf1oRfj4ZFufOD1WR6
BZ44rCAUtVKsB7ioZze7QVdzWSY+jUFxpgvvjYcRSp2EXrD2lJmE9NSI2eTDrtkW
x+03dDkMtAh/YoQ5TmQ97VyorxCbWmJT9ByXJ+Mh4v583cYF2YlkInWvQGSE02JG
GsfdaFt9zDRbpwOPMVkAAB5tMEIBAX2oKNZGRDlbMVoOjbhyNqsTJeDuttWuEz1t
RnJ4rPgKJdA1GEbEaCzt0fJBt/pt34oH1qK6oonFAR6y+Iqn+Wlrrje32RkmLE9B
GZCKsRf56dE80zhiZSU12IPNncayAERhOFwWLtr7jJpx6ezxfC0fD6ycYy6nI/gu
piKbFQf4V//lDCqlsxZ/2xYceeBqOS/RVM8xsYZnj4wchgmtDA2Zi8XC4lbDgc0K
jf5XglZx6U+HX2+6WADV1PTItzTfAkdg4tZlPUD0x+BDTN6ZNlnee0V6u8p/Tw3O
DmmfRiPkJuCE+j9lZx0u1ZQfPE/KMNuGXRaybMvndN91z8NtbU+XPo6l8pZD8Kq6
u7usDxFMBnJpZ/0V4XSenkvYO2HoYY6TkLMYlIimRr7GoQjMElYU5L2IGGhRJn7I
ED5aGMHmN1jL4Cm+6+6b9F8UAszHDcFhcFBzge/rOGIvG2iuoHEcDoPWUisDWeoc
BhKlc3asGf367BMf/Bz57XTyCwCKPsGDXRzqmnTjU+dpIa4O86g732wMKfQKJYvH
3kKdSFmv6WtrS3cHXkG10QuoB7aYFF7JcZFiPt72+XU/8O6owj/1EhDJYVPvh2uq
OXmVKIasbdyrHTuZHIIjh9kh4py7GEQ5gvNJAb3nrMPT0QPmjTDwYxv/N9WZenZD
QvlD1oRIzpO/CzOg9ofr3N5BXggDzE0jC4eXRIe8oLPGqeL7qhSrWf5gft7pfyrp
GW2D8H5hGn9cT+PIWVBs2wBDqrxs1e1uF52TLhIPL/L+EpegbO714DxHq9Cyhvw3
+b4ShrsHGGxED4Yz8OnKUO4UdBXrwiHy4vxFDRksZKAGlFzJUVkwMWPgF9eFDG0v
iTLaIN0AOEs1EslLbwQ8Tj3FyT6y63OgXWKzoEGQrMtWoLhjWB1IRBjOknb1wK5X
dSYW8eUMMuW+r3AgIB9Y9wntOgQ5uyWeQqxE0Vygu+B+85S9cBnU2i5tfpNm83bm
MUPA9HIwqh7QMDcLMX6LfODF1GtI2nJFURNaOgWA54DOMATbPcDlJMbCYtdXnmtQ
QUvkfo4wrwxPURjok4lk0dBvV4C3FTuxbTZS6litfTrC3PSkT5mC4a5h5yQQVU+f
mPosFlaHxffLI5RlRnkk6UPaIcIelE54whOGzpIbsVLtE8+5Wcs6P6aibT2hBgOK
vyMp6wkLtL4WQJ4qRigzsIprqlWyK8k+fLTskXcppDuogsClatd9R6MhAC+LhNSL
87xNpTE/JIhX3muf6vzrl4aES/0ByX4BsM5Wk2OpZl5P8vxhAdhdUew/P02yy9HF
pt1klAVvl+plOfgmjgc2nvInEtBWFL0E0emRo7I5mBJH6f1scEqgDd5sV9PskQND
WM2ShZu2L3Kyj+RtTHN03EIBQM9BwEK+p1gv49STJ9wJBOdrj3/ZwVBUX5RPXUW9
Tg4IADMPu+leSVqS5lDCddsm/1AFVAUgpiWnfLq7FirXKyXEBpafKEmvAcZ0AN3x
0IU58+1NxoBZwios93+fNTh2tXgRqUmm8wsQ4PPRA2eWYrgxQ/k74FmFy+y3R1+q
PWWQRmRTny5FoSQo+QercHI/9zqXa12nnNZIPM88nsYYWqYlt6+/5sA1lvjA9vPC
EBIOxZDo3PenvaJVHBx25MLNHV+F1BCOdvd7ACMRYmdJUQ4XcHg5d6a5msGUKhKS
1kcrwuunbfwnJ+K8DRdH4VKbFFkcwIgGKnftetPb+e6TGL78dVkitm9af46T+EwZ
AXgwsUeDdOlZiqKcQFdCBZNTCMd5TcxEQq/xpT4RSJglRwx05jfY2SjhE3OfmUcQ
2JbJ4ySN64MtJrHGkIHhLzvPq11PuW1Wd3UEpQnrifr+QjSJVQact5LJVuQhRXyL
UY/xMLLw32ixnW6Uvbr9G8rje4FSzSIJciVDEhininhL5SJokq9tTdON8R3UZtRr
XeOy8M5UQ6DTOW/PcFtgUpGjaklnT1TPIkdxUWUdQkSVBoqGUd0AX7Lc1OvoNn9F
CXCnGGenpQoIw9hK1/g3TIyK0LVtCAHyY8dSHuzwqV2f0w1X3TiM0Hf9ScjXcrSh
LK6viBmPuLyb7RHz13oAilHHdyBI6RtOEet/JnaLBsKrX2bvzVPoFynw7cp+Dw+b
oU/nqLV31dpdcf20Xv8zsXa7xsdjS71YdlDZdoI3QKeA2QOlFSyfzP/1G9psg3LF
M4xvoMN1BNfdPgG3iTnu6DTdD+WInr/0eejSVk9vh+tewhidrDSyH0BxZWswOcdv
ffNBduCg/RFpJTd7Fqf3JjliEq9eklgbU8Wz78i1/Mo2JWJexR29bBompMadYudd
MYb9YQJwkuGm/Yf6oI9BFQhKXWt8Bqgc/+HCzJcXLhNhK8qxKEhrDN5GbkIaA06k
cGID0qLnZM0VyMANCXIgzQSPCkrD2hqfZdNl/Zxbgnp2erCmiDTrohAgO2GlgARj
mDR/a6aglXkoBl+HyYJcegnAltwMz7bFfpE7LbCFsAGg8e4rGqqk+241UeHJPRma
ISbdldKEA97Wj79GreN3gNIr+FO3etJ5rEmbP99Y3ZIDPX859oUVKwDgPgz4Uy+I
TTV82S66XXA6kbeLPn17jIlKmQEEZz+pmxM2McItw/NU3o2yoR441t6daNaoyeN3
P5tNuNpY0NLh56M2uMk4B1CXrvCsRL2UJqyxDf2aEqtIq+A0+GljJGbJX4ag27LU
3tEox77W6AhuVrBh9Je33iNgD05nmAgffesZZHmKhOeXcfUlZig1ZmvgmsTTfQFt
Lg0wEr5qAmGN9NzfVWVmidgIoD3UfySakC8cxCX8Ag7i8DCtAg/sH9o7MGqq3FYf
7mhTfqz/wny6M4lE48ggVtUtlg4cAYzRe2lAytv1bkUJNNsnF84tCqNpVNjX5rf9
pq0OXujUz1PIsqSfcVTy/9eV/q/VS2RmQcVRqfTQOYY7UPlj4Zw0hAElDhTW/C1i
l4fTSG+iVUy+6vABz6wEQ+MWXeYC3kGnQgooB+NMizA3WGSVtZ19FiK9wOc0vXwg
RND/b6mf+z6FhrZfBlWL2yUh8wui1PJeYMu4KZ7sxUNyv1vYkXPf08itLFCr6gmV
RkMVMumrnfCfr5GmH+P+wkZDbBe1PBk68QTN5/ikGCdOlNp2OyTqVc2XUmzEP1F9
YNFiO8TPrTr8EW53M7uwYI6AlzOcl9Zy9Pe1Px0Tw6TXy67zADXt1+XCbHoZyNQ2
oIwGA2K22+Gi7YZ2Fd1PV+2IQHsgXEQNlwtZSD768lNPrZgraxTUaSFEgaNrNMBw
9NRdm8VV4o+EVl87gw91GnvlN9CWc06RyP9tPWq5bkfWfIn89c95s5F3fMS4USbX
GprLLK99FyP7PTMYfEvAPHPBrRAQqeOh0mjf91QD+h9INOAm/LgBgMlkWEmNEdF2
sqR0SsSyYMoepxv1mLkxs/h/s6qLyv/xK5ZuAxqUVoO7e1WN2ExYpTQDfIIDJa8V
4FkfNNrbtxkKUhrcK3j9O+i2w3Euth5uv/FveVuNRw2EFf0gr06gn1gOf8ZoUwGh
xagnJkwEH3sBWAG+i3Nw1HC/KA1EsJSSG/kb7+YySTgh1bg5uCVhDovCg2Zqt9yy
WFRUaB5VHig8xaEC/ttbeigPtjrKbjLIaPOXNLWaxRMG1wzGu3vCrva30K1WIaaE
E5vVdafcoLOtI52cdcU7p2+fFjZoAITpsxroGmqW89ZO2QhLstkw9E4UQTG9qJrt
32/2ow9IgTKzPiUPWCMOcjDaHUiRKkAZFmGDlOTrvAUzuVOXHIRRoXx046jQlpI6
If2rY0HGyZOS4H0ToutqQ02N45jZBfv6zdzCA4ZZiA7qbwifzu3oZkBAKv27TcL1
8Aq1qwZlCp+i6FR8HqYG5VouaXaE0nxpMmjL0oVnp+PuOVtupL5/9nZoOHGMr0Je
qMk5AO2/pJst0WUlc0+/zyRR787jkmkFv07MB2QszvdxEhn91LvcqTncob0jENEV
wijRKTspxQ9RzVmUFRk9rt010i3+4esyIqHEwiPGaZrM+RwOoOr6dp1/BbyBZeQk
5B3Y06gIfvZCGJ1+32b/5vWqknogcU1iQV4uK5JSV+TLaFi8dQRUZPvX29xoct3L
4UM28N6C7WcmieMDfaNg+6473rriBtTP8fSG58XGbLH1JEJ+mcfT57ANwhDYsRpH
4ajwFVRBd0224o4+kXXg0CH7nspQU/K5UF9wcp/a/trroOmRFxqZE30MwsxQ1fnt
jOoDb0QO3eBEGD5U29lmuMZjCNmOKsofjCM0wcGjm5ozzenxKNtA+6y+F12m6Agd
crfC6oc5YBrn7bCUxtLO8CP3dZZ3QIZGBfWm9Gy4s9M6ARMO8Z4lZyKlOYHRIEuu
Fy9qxkJXOKhMP2+DUHy54FwrEFZoKH52matGohuse9IShUM83Wy1t0pQBrZjzoWh
QsrWGH58m+WNHpz75Gn2R8pf6hXkXsFIbWhTykLwuv9qSM7q7y7hk5/eV0kW+BkQ
svxPpEOFXEtn3laYO5n3I/O5FSAxub8stwt/h1XCbiVswjWTvdvBHPLF4ZhmVWHm
vfs5/HMRRVZcXtKdhoWH2ouwlq4Iy1mr9+WLKaEnjV35tSyL2pZc5KNVzPYymLCB
is8uzAfMrW5gOENgCG+iF0xy9WfwqBhoLmJrF1Kg/wSXbb2omzi9O2T18s36oWjo
AC6ko35DdEvcQya7bfjqw9qxrI1g9XZPKOCZGGEt+zFnzOSvXRNtoaa3gX5pDJjW
pmKRR2M0fHD9kOYjwE9dIn8cklolWP3YB4+9AEWhJkekBU5XqN4KGfO0g6SPH3Dw
oumxvlaivOo1VoW3jzWLTEVRnWijPov4G+lfdpQ8U0EfO4uMhexsJbhcQc7NPArU
q4NAXZjOWOqsCZrvTTHIFic4Mst5s0gkZgP5KHssFjVnBPK1czf2zL0uugmuG0xA
EB8LwE3H2Xj5aWvovA4I/IXfANbB0sCXLmAKX52SvO/qlkSNX2IDiVKXi7UQvfY0
5OVA39gi9W4hjUe4xG78wQ5nGGdm05e06k/cXfztrdpCZ6KWgETIuVoByxdMelDR
ZURCUxVsD6wXKOU1PUKXqSXi3wtpzJQ9JfpC1Rflw93bZtdw3RGIccvW9yrZqak6
DrPYCyNBUMe2jP/vBko67GInIS2JxPYHtWH/UhMjhWcle4agfBl8jvAEislGd2qG
/TuEsPkKzjIzQ1T8RhM+HinJIaQOio/ChHtKHd0O9tKuxhAQ0EA6GD2RlwrvjJzF
7xETKkSdGXRe0RKsQq13MueQ8TQFe2tF/vDozQU8bbfE2U53LDT2vgZlm9V0b1Bo
39VidmRCEMceaUbN6rjALrBxHbeTykpKjdmmNjfnvj579wp+DO7tXa/XQMXhpbC3
GrM3M0hI64CKNW8nLJZa020W80TfLbswCIWkknvo4OCCEg9Qx3/BwqJHXrGyi3Dy
9sQNGXv+FgK+9LkKpxLNEm7Si4zEMpT5iqLusdqBmclHee13iMMMpD92nPss7gEQ
m30D+NbaYoeL8rckFt3bNt6K8yt3BpsI1y8cZwVz63Y6cNODRoly6Btvq/WUCuNn
Fif0j7YIWs7us4sg3aH5X8nl2lsHBvtbOlDTvtU3b6W6pXA1SiOVstz5Ttg6NlG3
xa6TN2p7jbeKYDlLlvROj9pWgXpNIA7To0QlyoM/rNkO6JLGaK6E0rxD0ekwtHSm
qHB/CjCPycoEpvnzcTvevhHbWQPjoxL9A6hr6xrzMb3FlF9ufonFZoI7WxFmsrV+
jpp6Qv+gmslsYt3ioBKsDWlDrxtAl1X5JDJCA+tV0R61U9zWeLqegLSP+le60CsH
LlFAoQCy7MF/jXHIFVLq2gRkgei4Hdpd6IF438veA5JiQTTtxKAlDJj+h6tisf8E
PZ9KLAXIYoTyyjRbA7IwvjzTyzHex2FOXXwBXfIB8Mi2hRUl6PrKBOhGk1DF6gpw
a9n7WS7auwI7rPLtdc/RHJIdTos+BvvbZVu7DFrkdXDn2e4Rv2V4ygSLBBkfJtuA
/GtP2ypzkzNin5QVEpdk+872HQzQKIT27SSOBvXDSnmLqeMqcaU5YO1qvDb0KoWU
4CbBbLutBxxp9ht8fM9/sLwL8kMXX5h+Xt9guyikkQZa0g1XxfQECdcF8REXVI7k
EFPnbjDhkFzR5+8YrrxTYRNRWsrAysK4YdHZJCeBro73GYEt1AMMKO2qJXuwZXC9
wZkYr0Favn+GdkbnM0huZ7duK5odPtNWeGYT+Ftd/zhetrr+DscY8uuOdGSmk64f
RgEM2SXvvq/wLGdyb3t/ncpb+ZCp71EUUiDHgp5Itxu/px8z6BmqjO5ImyTkj5vk
NoUtE8SBpopmkGMR+AG5stK40CxW49h6gAwT9IIv7aKS3pJzYI05OutBcdCf6hnR
/Xwo341RW89XcBtk9Cvv+ATmbe4Ai1xryZYnH077d872KDjjKwJzbuhSqorxlTVQ
vBy9FcXscSwG18q0ETqVlTgmTSNHDZoZSB7YuNPc9983iKL5RZt2SDai3hKDxR/6
iDYHfEzX1WYADNvvNIRYAJbC6mkC4YJNCnO4rY7rkWnwy4l3FCEcwm+iikuwn/UZ
jSGWzskikAledGzSfMJkBSTxUh3M7xAk7iKl7PvaNY9wrDKu4A5Aml5l59zzF7fH
rmSScVAe7qtP7ImZMEqTpzOQjpbmR8ihZR4KWVGkcTBttsfdm3tHunTscdmtmCmK
P5rSwdpnkqlsyRoARRKkAJfR3AYtNf6rOYnYknd+XXMm02lsrhvyHgr8BSqux5So
2uqCDZGIykCucPKGg7Acd9InSeyPQxQZOburWmt+0laDt6X7gA9JkUA4Covr/DZM
mps7K7jC3OzdIQkY66u40eujdp556i73ET2dkpHURA2HeOKD8T/pe7efxepqFXeu
oI8Nf3nnxbZzPWQsQWbfAJ9Nc3QuF5c4M8Dc0tmQy9NA8kInslwb4hBY4SdyAOwC
fNwQUEnTo+AX4vMPv+aigayEUp451rl9IicB3Z2A0MFBNUyl6P1dfFFb8QItH9fe
otcQRx4RldmDEYV3E2XZDjayFHvdcM4YWblUwfboNNK8q209adDHsJTq9VI6qaum
0gwHmWTAglsjL+SiMBmIjQrY3IOGeu1jf1gXIG8furIsBXnpcK6goMKJpc1wP3Mb
a71jrjQBJsZ+UnCgcNRaRwvDlfKM/XF5r4SHU8surZfHDVhcWT9nbk/MZ+smVZRP
phbAtZFgBg0yueWGUQNylVeAKN0i+ixjK4QHIhrMltGduKQVaTN0YEzEr3ExWVNr
fti4CixgFkdAl2Bh+t9i0SZAdcfFNHyRNpCrMHAh29Kvaz0HCqK1YWnr9t9VPHoh
Y8S8J26RDaoOieIwDGpC+ivhXtfgsNan5qn6A9haP2o2rUi2G7cae4uKoWhVdcWo
Gyjqz+6qo14KkxGlkYWN/sQVGa42kyFEEtgUU6f9jXVjdOVvvoaq67eZBD43412O
XNKJz4lp7KrqD8spPEtubV1WwY2n0JfpHWoTAGa5ATa7Gi4Ot6SY5EczWWf6hnn1
xotVX1nJdhhroWg00KDPem9sKaIjPTgQDtl6Q/w3esMt/wYliBoAEVmlJxeYww5q
qaHt6t08/uYSk0pAtrkpGJU9gQbQPAzvJ6asqnysMJd7nDCAjuqtVUcxy4HehGIK
vC9+rLcLnRi/6TVXBw94zAsfRi9UOwRQpl5euHg292ZxaB7/YwBvYwJ6665kjAcP
dvxsfBPrOTG5Kj8imb1+nwGaC2SNfOKs2CbIBcSBlv8rZp16/YuuUaw7/zgK6RkZ
fSuer+E0skgvxa98mluN9WvxZ3E7lHot7lLU5G7mvsysQyS2gAmMq3Ie/vWeeleX
NFOG9LK6RL9xnInJpg8CdEEFhIF/o1uNcVfytKkSL/+5iasaIrOXX/M7T1uIUHUn
s3UjH8huwc9VIm3cSjFwMKufysGeEyR5GfXGzajkw+7thYlcR0pqHlvfCBXwzSTC
01XUmJkL6Ge9lP3uXNV8mOh2Vum1OKS4gEhou9TLjiP6F6JUoFZKmNIploG5/3AA
ksMGtjr7stpBif6Lwp0NZfcKtEd274OW1w8J1OQZVmFXtZqc4dlk0l7yBbfPVNvH
vgIEavxfhoeeXOY2Jj91wRL9JoYeRI9ImGDtNWfMUjeEHSgeoMxfsMJlhrK/UnHF
ullYJ0tgN9Ppe5OmA10cmBD6eTPaVo3lplWs580QjcPQdI22asUZp5p0pYViWqZF
RwMqgxJC4G0ISKrd/753qeqkcW/hpiPdqPQUBeVN12GvaijA72YaYlc5sU4wTLnP
PoYCVZjjvifRUQU6uI1pt+yK3SF64TOStmUVAmsKWFELFygZXV2Eh+djvHdDksCa
DBtd0XvLsxMKwB0ZTsu1eFmQQP+1TG49V98mqHZZcjhEDo94i8OU3kpN7OELyLA5
BJUwEgsTeuRGvTCprFvbRn3buyiZ6d1ZYB7ZbmhkgTHPZO420K91OYkLN9NLnRlx
S+dGVZdmQzh/pKZSEDVoiv1OGAyjLE5hpGytnB4FVbcYeU7N1LGKCDHbZMiLQqkC
jMIqilTRtr/givz9HVafPCdV76RtDsuRZPgHqCDW0+JY1nLVKM5NuwblYulLBfP1
JnXb2HXJDjnZ0nrHXwAMtVjf/7UeKJz1k/c/9+XBH8nLz/0IuQSJvnKrCYxVlHcr
5HKHacuMadAgZ3Mh8iwQtz861pKQ5LG+GYqHYPo/hzpJoOzBch89GLdFjhkCadP2
gUtK444sq11veGXjuQzH4WQBK36RQpVhdJhATcWqcM4k0bhWShyrJhDU6c05rDxS
65Uoj2HWdVtPZqrowgMCnHUnv2Oda76i2+unMWMkzZR/UxSlXQDAm/RsaPsAKFN6
p4bz/cPyglSTSMXduofH9InS9d5dXXesbOHVIP6T1OXQ9hIIT89Em3L/NtJT14W3
aCSEZniFROetJRfm5gDByUFH328C6lIWUJNYneeGEQVwx+kuLHyVbeBTYO6degAq
O425fbEyTv/D/W0jL0QdOyKjgugVOLqH7+uMWSbu/zd1cGA7j7hpA1oNLorf2Tbe
CuMTTHu/Kd0K505DidqmGh4wbOgWvuf9gpBxoho6vHQmInlYYh6KwdUotpGkAB++
wCkEKDF1ExyQ7nqpiUXeFxzohUoEfuhWpTjrseOUO39v2q+qjh9eg4Sd6iCj4unB
NHnet5vP0vijlRspGda0fzAn8EXSijD+pZLJMftQWTXfEauQohNIgTcXwSZBjz0V
zqrvDHDYuYDu3rQcYroz0p8H3+DjxgTV2AjwsyqfTYUTnfFwIM24Ff0MGwKkweS6
EHYz5mTJ68hInSYnSZftU8J2uH/EZSyCvJF9TbPXDu4D3rUOgNrghIW+xEMfBwa0
mPiu2r2L6OMYJC3w+Dah15tMPpynjFNycSOGGkbjMDmdNLNoqvKBaEpLv0duqMge
MiHSCjYhXNJ+/jpReoidoE0sk6pwEkFBi2wizRlB9tnnzBRPtDghWHqtqnQYxxks
RZU8V0uA0FwpSG9VLNpo3WPuODDwCfXOnP9vriPxw51DHPOIegZ95iOmXuwkU8wh
TXZSoOXghcQJR0vqCReZRIziibjpTujzz8rP+qbNgXa7tf6cdPXOgrHnPMihttoe
EcfX+0OWyytSDlG0d4/iNBZW81DHYZKG5OMqlzr1BxKxlFbf5kvnyA/9d3WgatJb
3PJ1DPZp7l6watjPjXQ2CoQ7vhPNNzqPAsZXps/0nRqx+T46h4aZBxiS/hEfk4iF
7Oojq7qHzV2SieqjUY3vS04NwpGu/3PKPMp5mEMg/F+IHgXHbkchUEUBppD2NEGM
BYlQeQvDX7+cQRbs9ckIH+twmyLGxcSxyyOX09OY3+Knmk3Wwub8c1/0qRD4J5yg
aT8fWjWlLKRcQMcgl8MsoCUN7+vZtZEJuvbi4KShdIEVDSeBMvDzc0dq13JHumVj
MsuHpkn5zsVhAG9zbY2dPZmeKa5tfHgVV0+d50Rq2klUwIPPIkFwLmJU37mGwPFx
nE21Vllr20KbhWDJ9bfKt30pPCHu4kVM0gwAJtHVOtUB5JJzEXeysH/QSzfh1awI
drlZoUfPDT+V9C95d2tL9Rv3Rh5m3OIjoAdLIbiGB2th1mkwY/bO1lPgI4wpPT5q
oBOIsz+GFUfEyGdzN339SokHehet5+w5UgHoJ3xGTwbW080x3atz+D//XgPok5ym
E8kQpR/+CA0XrwzwzXFx86nZQmigZwgaLc03TG8zF3CmqrbImaTeZL5X+4cNYGss
eoswbFzpcqyLYQWiUb7V9bS8Dfowk3CTHNwBrJMhyJd1OFq/0QgpcZv1BRc1zT0Y
kkdEolEmOXlJXjObE6r58Dx+u2NftTrFKwLbjfsVWVFuw/Agi1QhgRrp6ORt5SUD
5lT0PG3jGHOl0f3FJlBHSWPeVLtO8dzxhZyFir2I1uDjF+Q1g6CDiBUenQrVdqLL
QoHeRVGjha3oH4Zfcdw13l4bHUxpfCEftUXesYyC/22n68v0BWajWz2NatW3mzu2
Hw0bSTq1fXJZuf0Ra9VfGRHzDeE4g73EE9pWrTwhHKh+NpM+gcRdiCT82Y9xdSNw
6BYg5IgxSQTJLk7ud5rg+qlOJEVJeGeHMmc3sZC8raHxaH21WEnjdiawbL2SWwgW
XM98MRZ8zPTSMk8DYjviNa//9boI+TnreZ3x/Eua5Bk9fB3AsY6j/ASB7HScrKFB
9H7fSzsKXHlceEiv0sDQ4QeZg8cYDIXlhc7Ml5SsItKRmev/yIQESOloccVXcVqY
wwI+hziXxvSLCjydf35z7iK5IFBhi6yVbnlBR7CWgrwdOvu2C4QDSaHVCqizqlQi
Km+x61+6WUYULnVWB1lc+59N1qkszVlCQncLVFME01d+uvHjXNi4xXYQMhC5nndN
TKeD5D1Tw3u7YbMmVF6o5o5m15+yEGLF2hKqMenTC4qvfQ6fpPy7ojItXYpg0ysi
gFBmMdAk2Ak35Yq85TCKjdOoYqSZTwAuMRO++1t4jLr/fdtsZaR9UvSp5vOKvOmR
0QYZvxW2mlQLlXfC0RjU5I8Wy+ICUVWq1q8WhW5Bbz5i+hbyG4VYLlYV7dyqrDux
iss4ZAm4LYHguFYwTBxsxow7XzDIh0INaH95rNp7E3mqrtlFsEOWo7UPrTpAp9c/
XtMMxL6RH+py5QglIvFEJoIRJW2i27sd+zAXacir58iiWO5qShx94SGk6I4GlJdY
nTqw4x5suEqwsoX9PQHduRkWXUFaJUVoh6H7rcdG+8U2hpZ3CEm9+wAwVJipTzCC
DxUQXgWo+XA6oeNpwDqWHGePgwJjUwgWPDMBv3ucFc6nebcMV8nndhfKRcjfaMmr
NOkZFlhwcldWVoNC7L9al8OZmdQuzDBddk8seM1de81RB6HJjUMauW5fpoXNi9Nm
d9UvvnFONg7QjIThGvOn+EeLurszGHpy32Vk7phe2ErXR4PXZ4louVlqzNo8X6Ue
RcGNGQbXI/LtC7k8jBlIB7CZ2HUC9fqNXPPjNv9TZlU1bXLXSuFde4bq3xKytUFr
tAXoV+37CJclJGIUECxdrmpDtoJ6r8G7RzDAYhz0ONe60KQtIpzNCNqG47jp3pUk
tX3fCacYJNqSYgkpt2O0aHJb32MJSPF7tcQKux6gsTLTKhIqEm8vvqMDHMWPwQwV
uQd428E/X58PmV7z+AvFawOpPYfCeBsXrZE+VTWi3AoAcFixwn46M4KGnrYB9aFt
mTjEU3Ipi9zNYnHd4ekxMyOSzjnradHKmsftiMFmLLdlMCecYq+JWDX08o4YIbnn
dZiAzGbIJIxtgZrjJPdgGaz+q9X3pXl3T1qyJfIedOZDqVLlD1k4szAmjOqHlmXy
ugxOIUt8+8iqd0aiSOpnVAk5UsbP+XUCeQRQRZytslSVoRXBYpTyFxUDGkFnllYY
rW0OhWfODS62FloryZegGTeiMyMOa9oSL5jMX6NYgB0Oj0awc9Znnzn4tSP9RQX8
Xp7jiM3VedNjsWn5e68alIvj1rWZD4tLA/bybpUL9JUPLrRZP9vjLnFsGOImMR1B
rgalmQ8+Xx6v5wQaAP2bNSdRqPSeoThE19SERgKyosD7nXM+tRkZc1Im8arnhg7B
ZBwGnXmdli0Qx3nmg0vm7CQ0eyNrjRvxTHmSW7S3hNxSEH5NzozsPQyrUMbbzT3U
GnpZoPnc7+joC1TUGc3ZoQdUxXZ9rI96DOuOq30MrJ3aYujrhGv+NQ/eGQYQGiql
QNFgpJG462X1vK8CFSbNVnxroPVNPwInYm0L/JGrK9tRsu5oRoV7E6ed9bKqtcNR
SAe/Cx3rTpuoMSmMtDKw94NyabWH22DuAhMaJyjjamE8PN3poX8ID1IhtBJPSTcq
jeNO3/h2PbCfmN0WS9DoTweLr2igkrfqQkXxLcieZbkq4gXCRMosvJ6SGHu85lP/
749FbWEkx4Q+Y3TVHd9uWK9/l046Y8up28ZvZQ8t7x59o4UMwYUaJNIS/4zIE0f+
QLj1egihP9kP1doYgXHK5pdvnDpXQnlnyYCGJrp4zskdK1P+D9BAY+r+VEpk99lR
UtfE/ngjd7aJqVBDRuxst82d0sEMdWnVABAn5FDmcZqOudwCUPwmNRSFku9iCE4t
fKbU6QfS4QI+yGrWUTjPIdqt+z+WZnKIauMInjxU8qlN9eX4um+pd/dk6psUHz5u
xqxThlLjKoqcEkVupZQrmUrLy2qikdyDOY7OJ0fLU7BhQtJEV8sYv6D9yf+G/MP9
TnNv1z0wrrnfLJSzYvibKTFNcSiJj7e3y38nmFwyCZILuXqgOFUpFaw41RbBeYqj
3XaRECndRVdVRBcKPtgYL9W4OyiA3lKRtBePD0w8tuPhVjqMSYjp79xoiihgP3Ao
xnb64n5MkKgoglo/yZSZAQu8xgLCRlmjRdoL4BjNHpxZrv18n8Oe0BBG0jFvXwyz
9WZhU/VBFx63CGOOa1cL68Wy/jNpMl+tH010dqulGDgd/VCaaOLXJR3c57Bn1fpa
nVlCcQRZPrqimlN0xEv48ZTPkPTXHSCtf3baSPBAlkbEecz/OWC9EIWGkQ4vH2DJ
EElFDn2fQ2PyegPZqrIiQVT7OOJjtpks6khwvK0/5OQhB4kUpXQRXxvNi+jLf1S1
dOscI9jqMkU2APNu3vj3C5Fq14D5OUZY7gv/EKqtpHFnITQGKIVf5H6bpjKrAXnX
WKQeul5cCOAPDkfwXRImaNCUuOF+/OaBq0hE0m3gFMqPFbFUFlYyNqsHEM0wQR/E
v6oSHb7zLn+86AYl/7DP22koV9aiwRiJoSg0nc9s+GUvOBSajnB6hFAyurgwawPR
2AOhm+qP95r1KWkc+Ma/fijoDuNUKaA4GcR9JAPCmUYF0rQgOy6/W3AFDpqgUco2
9jsPokKVBqEi13uFPbksLIptzwO5sSM40b+Aj1KReNjONe1Jc6mGcggpDXUF+znm
vkm0zi4hpAr0R+Y5jp+zCg9tVevxYOgo/KIaB1M02+aP8818OenvmPC5Q3/qRPfL
eG84pNcttqihDeGYgK1hzb2JXu6uFCTp6I/UmCpu58F/IwKIcQfmMS/xFfDjFllL
9Bd1QSUiDFFoVERfAgnWH+GbUjLxya2o6E8X35TbkMB1Jy4g9nrlnBAjvVrTQG4S
EQvwCAzDa9Jtg/LgwA09QblJZ0xkPcuP+UOUT8HgAksnH68chvQiP5ABpNKy8e2C
ZzczVmDiRMhKTIDFGfsdfSoTWGt/hWlW7hJdQg3uzyfNLQKRAM/R0S1XUe6MJ9q3
9jNBk6XKrC4ogeJI3Cfen31z/wAJmVdx3lqyJ0Fb8UqEoymEGZHMHKVmSextX5dX
PuWt43WP8fXjfi3SOHwaRBxO7ttR9TyWzgg8u++BD8Q3tqFPPhRSIM1dP/Q+jDF3
lC052iDZ8U6BGGygUPgfxU1VgZtNuBxvWemjY+iDimj0rVo43TJfFLFYP4Vx7Nxc
m/ObI1q/hUEcY33oHLSUV8TRaok3e7VI+2nsVQ7rSOvLv253PszTQAcpLaWusksE
GQtKTjLlCFaS1SngC/3CS3/4legBUN6T5dMPHyHtr9vwF1xYYR7RXVnmE6LKQFME
sR05Rxo9SzhtuSnv7ic9CAJfTRH/F2MKqt8/RproNYkNlbR/VKBMZAYVNzgdwvgx
M+owF/NxCwgsst9W7csx45eoFdLqyznar2c9dQA2ex9Ik0/xN/E/vMbhSWenTd5U
zSq/5tnb1du3HgL+zBRWW0gd05GQvJRRLfIhIlDDqQhj/jIAnWmrgYlK79k8zbOQ
oxYGwEBDDTOxX0FljTa1NXVdtSPBesoEEYDcLcUG3ZMi5nTRlbLhvSnibwkGl3am
scUUQyzkSq5uQaxu6PUa8WiXvakDRd1WA+4f/n6YRyv8vCOSKPKSlqY9JcFpYvPp
2yG/NQ0r/uo1vakb1Rs7IZtZJzwc26xasnM/jxoRzX7V8IRE1tMymVv6LFvJrMFZ
Qa7ZeatVr9TpIpIPEyPkU9GpY7liNxgfMWhxdPUCUeekV4Qki1k8Pzsrkq7UW7iB
Ixb2R7LhaU1gUWDSSkWLAfmcwOy5qjmopgFPanMMpoHNmlUOuuIs5hn6vpYeZ6Ww
6GclSmlycQa9G8MudbFKqA11Q662TWurq9ibc7sG5tOgdD1ydW+KzDoOlw71B00T
4EtPYsshhEu18ATLVKy5Fw/9+R7dC4wcPNgNORt6fjymneiJAwRbDW2N3RqrxO9V
TtmSbOa4tFW58QmYFen/ZmKlpuPCyy2jDWeWL9Z5/MoBh5582LGxhfrOG+c+N629
sGilpk+UiPYYRykNXxR2NrV07XDWlreKJSVGLWOy6YIW02hA7RO8fcf1fUZUoIL/
2g4Iwf9HGBqexyyOl5lWW+Lm872ux8UnSAIv1PqmejfMDNXgK7+2UQRA1DGHY+wI
QTA4J1cwDkKEpW4ZiKDpYnpD9v8pHJe4tBvx0DOhzEwDLHpl99gBq3c3gcEq5Vi8
FWZWh0Z7sfj9ssaiH75lDLh0jkrp4xnAiw2ZJnOQOw4cO+tYrnm9jqWLFDjdUPPE
1Ksob8/rKecmbLKMMAuvrUxP+PsP4L6+oQxN4ifsS8SSWVjdgZA2U+9iwHIbl2Q7
xnfE8LnT8Trggev1t9ihVUG1vMlpl+A6hzfoPhl8TSngfwB8lyH3HaHktGTr9yEW
gQ0FZd+fkG/0wjuRqQfGu1U4NJkRF24z7pcbR+na682E2nR2Mtr39VRAQAJVlrH8
h1vB4Rrg5xu1QXWE2gH8/i1WFEfSVhN/CfWhpuMxNRX2jRjzO915p4V3bpSGg4uz
XqYLmvDtY1/w+Fz8vJ6zx9nJDP2nU3p0BsZfRIfzxvEQaBVgECmN1UJdPCWGfyeD
WJ18Y1jBz1YQZHJIj0jOaPeLaW2N6mWjk4eG3ugIST185MhLPenMQT9a54BZep5Y
TpCTN/tp/f9JSD0sIZkXiI0zvx7ggDF/38rSMZ0Ml5sxi4QZx4ahvphSw02IRJwI
xXoZGWe3E5PeoHnj5LL7s6h20+tymtrqL48Jv0OVj+2yRFTWLg01i8BaHCj1FOcL
jmU4T8GbhlIEmDyDixE+XmqlMpBONIFY9m+8na4BszHOfGXsEDcMjaUElFAVm85w
DF4RSnJzOC7VAc9azZDAoBoEHrMj+I7TQf6bKStJCX9/t3S2MKzIj9vL307loM73
606E18de/P7jc0ie3UXCORefDQzfp/EqcMq8jqNh5SeZqfp/+9lwLYMuR5cg2PRL
tzLO2mdNafSyH0DzEyvqp4ugWROq6h9LiQ+/38At9deainZ+d4yTcoLXURwHiqFO
sk0c73lNpokn+3Pvfx7wRV4vN/h8q2RTuULCnOXPwSOq9ujtf1f++omQbAQAbJwB
7XYyvh8drbGXSJbT1106jrax4k5pOj9093dWPpdA37zT4j/eQuS3FoQxjbq4B8ZV
QYRS1SAMhqMm+cmMIen+GBNZuexxiX52lRg+kUftv6XE25Ox0e6XoN0zmOqj89Yk
Ig5hu+2Pm3DvuX6Moio2MVMVSFafVEcMa1BmhcZsXL76YMcsMZze+3tSp66mhodd
N1pXO+6tD3nDShcMa0Mt5vZd8JCL7pCwNIHuR/OIXLTPDqXWc0v1aehQH03iEXCn
MmfS0Xu3kwqRhsvNxBCIeUq3HzFYugk3nFBB0Kvrpyo+jad0h6AvC9R+/AQVs3Gl
moDs8mmw4U1FlgENIKdX3qDO+Pg+Qj/AR1PJZrkAbwfSFYQiYE4WziIMux9Vz5f2
Y3o8Ftj9j6k9dvVWNeHi17qlgzdUTcvL+3Qr830be7/ucsFAOeddoyLF2ZRnnHSg
1fm9uiCkzmpS/mQVYLKW/aPWHKY9DVF9I7tF8pFpmKse36l+ajg3IywCFn5INinK
rTfUi+k7PFpaf9kb4v5vD74YE5dBYEeGGJQqS0LQ0AmkgeLj34vSEYnlXQv2/YVr
DgPyCSTPEs7VqLm1fnsvDLYbsekuZr5kxZMTak3++LJUfYS8BxwnXfWI4/0rI0fO
MduvkQcOXNy6TSoqL+kS8D7Xhj9bQSKVi2L2kg8hwow2q/zjS5GAmRqTTIhUhJC2
8C+HBCacGdaMp2DmXyhaclK9chIRU0qpMPfnyK4yhcdSUszc5FH10DAIYqDrLsrd
ZHQJ6AMD0tGFhIosVP8p+uOxWwyRfTFhNOq+4ui3s3GgNmV6SiUKkJ/w1NA/Xd4Y
xr29rL7Rt/zvrqYMV0KolGE1fpq96YUVdvi72a+TVni3xwTM2abibXxSz9hy84PM
UAXYJFaMQ2jCmBMkj6+kYGiYZQ3gOrtnHdWsu1wbypf4PD4rLlE/3MH5yzTDjOUO
RSDk5mAuWTSFrWKl5cx+Noblm2jBtiuFXv8GyaXsi94tFao92ynFeejcQtklVyoW
2qhMSXYrasDiS/rTGCxJ1Nt/a5DitSmZYcs72v/h46roCNHYLtDqSJWnh2/O116u
s7RehiXpmMttS7+fcHLJszb9CSe7SBoFP9y6qILNkRP/KKmJ6RV4uZ9yqY4xhrkl
nJCj74pE/+cttTk6fsPxNx0HyFc5KwnhZoG+v9z0WOKpQ0e1ZSGZXey9P3DTumzD
Bmm3Dysd69FyN0Ogdw8hH1y6hGeFndmyAol4SsloyeBk5//87aT0/x26QsspIoQH
zjoZkflpYKcXoQoEkf99/jDHATnVpo6sA5lWkdAreXFQyJwcSUOhFyl9K7J3R7fb
lxXeEhosxbSd6wcaA7XR3cBA2iXK9fP8yH7LaoK8KpYBJjMsOZS80Gtpke3k3CBD
LF/B0Jiin/kEXxGdnGSwis6NTDaQqKFcwcAr8G8Djesp0OcL/X2oehgpVVdC8DTw
IINVQchYXfimuFjJ+fsPcXYnCTOyxRkpcYVeP8qhbR4vSg+lQE7woo271NZwpCEU
MqgyOh6GO8gpav5Y3WmIhfJF1t5ZjskmFeadm0cRyWy3Vjn04Pn+JPp7J+ETzPch
85SBwRUSls8HmF21dI6Xnbtc92ClH2vw9shRN/ildSVr5IscBi5KlVabtWh5np9/
Km+x9ljcizwxPE2Mjrzm0P/y7OeGQwMEwGNjbGGZhzCy/mYUoPFeSB0ul4iN0aCX
hsWv/hbbb2a81XzbBNgEJAJk/pY287D+W9qGEi9d5n3SMbwBncGf3+u8Kwjr64Gk
hXK94slPlC/Xth/MN+4h9oPJUNLkOBLN5LNi88OlzK+3egfYwoDgLn9WitXhgQf+
+5+tGZcFPTC6dGG+1N0yUS3lDAPqdQlPK+wDDMGXkG2Jf/3eNF/77qKGZ5Do7zkk
9x9APKF9s2EdXkQtWEJqwyMvjj0amPCBTPBWulRinrDJSbu8+wqzNC4JLUzHPcNp
bgfjcR1Lp6R2hb0bZozkzAMThcfIr4ag4anWoHmW2QJRUh96qWbGXhFkk7L+5UAj
KhDzOg9NsHwLdbUABagkvPPX/B2fT9rMeeapCnEGcH3ZL1l6urpe21kgVI+lOp20
BDRNdXkXee/xH/6o1hCgBkkdl/FVDHylvs5z5XphmPFEky85FzjGfTDlfmoz+E4t
ft9l41oVp4LU67SrJxMgDMV36i72Mfn5KNgHtmoVdS080fMZqhhe+lXWIGtxZHho
KA+qgTdV9cRhh5qRdSMjtg8PlWPX7agDW4UpvHNVXUMW1Ao/KdUT/m2ZFfObRuGS
/P9F7wiOBxwTq8Ny0Bth5MwiKWK3RULeUgbTht6/eDG/twOE1iK11csDOZsktYqv
qsmXnpOu2kwAEK+lhZcAwHeH96KOQpB+7jiDhl0g0Wwo58nS4hn3IdE+ScZrkXme
DBA6DpWM8tJeQAgh0vj/OnWeXJucrgQmr8eDDEua+Nwugxh2HqQr48wt12WttJj7
ONxBCpyYyTsBHuAOtmo47LmmiOpO7DvcNP4OAVV7B2Ul1/MgUj3xIEdhI2upZ9b/
J79tEVkc5Z5c7yBEv4qt58H1rZ93glBo2Dznvbkc/0sXuUcJeJzQ2P/lUE3WBDfX
HepSZ7KIDwetVNfloMYoHa3E9fQoi74wHl2u946MHpikMR7PWS1QyCy3RjQKZt8r
bJUEsh2JqbmmL78sk8eSxI/ezoFaZH5Hvhvb2J0orvWFWCrg9w/tGfxHD79cEdHK
8my+fOIqWT0yS7IkYlKs6oorSGMm5xpyIOwJnBSqIf/xaiqJ7UDp0d+xbFt8UCSe
+wpkBEgw5c/UtTIHMn7WiPnpka276n1X7ZUaZpDJ6Z/EsBf5/T5yzY3wSZrhi2up
NPIevCu82RfIpLzXBAh32kvfSX/Dit0yq/eVu2j6ohQatfRhRJ2fy+kE0f0hmXr6
/xxUSxwj6KOH0LsaLU+5UDFjFL1VpVOvpp9z1MpLuFuZ8SLrKdXelxMgo/pCBDoh
odzhQQmfoZGxoJM+bsENb3smrodSK6SOTZqhtH33R2r2Bn/iCkS9Qlx1kgc9pYjZ
8j40kx2lWmKj3a0a3Hch9Hv5/AtY2rgETXQ3kKshfbZBxL5MISdmlcbBqZ1OmsgP
BllSE5diy/XylCfULJCYHMYzHMIzPfjE9S/BY52uaO1DXO33wNnLYaMhPKu8S2Mn
KGEDaiPn943wsTiQHEGpI6JK5Z2TLdAlFbmwvIPwpM2qPinesFPKUVJJhUN8KmZb
7Y/2cbG5DTKfALtZMW/9hcmYHUzjdxzQwneR+JtC35YZOBn5VLQI5ryYGAAo8onb
fH/fe8HRtmOEkhNHSAhBuc6hPDlrly4nMLb1M02Q9270DdlKGlR5wDLttq7QZ/I5
KlD+lSHWiN2ZhY8AQB5Wv9HZVH/ZuMuX95c0chhaylbmYEK0BJAN8Vq1uFNhfWQA
0SnxT0uKQbytYfM4MsoP+QYa772A7MSKNV42tcTWRVrOxBxUVx1jxWHM/+axpBXu
2Yqf/CBYGXruvGlKt11ynf6RYlasF3Xoaqe2DBSqE7QawRQ+QzkcS7ygRdC2Yn0Y
YjLeDDX7HKPOTg0rZa4uUb//WITE9cjilM5zR0bO/3ejOiElLWEgjCyn5LeDN/MD
FcPX9wIAjRQH5sd3e/gPoHjIqODbM8acKCpYdvx4dgsANNvSl+nVhz/81LtvhVXT
Eo92MDpGMiJT++FDTuXulO9ykuv5nzTZu5km2wFPeh7aJppyME/4CW4eLbrOYner
1TgG1dxtCIq6as9m8rrxuyVYJTH10gVKRgNKIxxzAa6qaBZgEOC2maH8QTM1mH6g
hPr/j2zuJAwrnQDfoKigY+MlpstTALiS/lYRaHZ/QDT7AVBybS3g1d6xdzmkoBV5
O6EcnrfuoY+r+nCI7YO46gr45zSDGYZmIjx3gDDPk6J80Q4V7qWHQv1JHOpZRmZP
u6D8ae5Xb1tnS7SphpXs7eqpfRreJenItPU7ZX+q29NsQlQdukoI4OM+MzGDPshO
lGY9bUnBVU5TBQ/QJCW6RZlBNtgOZDDJsJzP3cF4xf3EEMht2LtlGryslBpc9rIW
hl+WjBkztwg64dC+iGVidz3Sh3JpF06+e8tJGO2VsNUrn8Z/3CUWxMUz3RQyRooE
x8T9M1p8PgW/Z2HvGr+l0LqUepnbuk/LSWY1mtJ9UqMLvjZ6JhW1g9ZFgvAvkkR1
5WbOq7/VVLsgag3sLlavP1l1ZX4pb6BHs67obViRHUmEgZ1Wam3eyIn72XFvHwnJ
JfYZGfP/+VCdz/UqkQE6r96V5/Pbe4nVpp2savO/SgMV+/TBoOYs7MPQallDEues
nR8G2xeluYwriafpJwQ0tWvFVVPef0YAawvFO6z6EcjSj68lZRPewHG4c1zgCVBa
ZwyknXqMneNrE1Lbx7gvQjMeJtbvOTJ+tRQuRIueVE+hjL82351W04JXg0HM3jgj
ULtG+myUkHKdhbUwpH9q4FMlip5RSI1HK9FkAvQyBlrYYmC1m1dR60e4Jl0Qy00i
pmSF2tWsP743hachr6WYY/sRu0SN8Ef0r6RPSu8z9taoYnoIyw/606LCreLA0KNl
Zd4YHs/o1P2K/Iy546JXXJqkWz6prhQ58dkAX/HbRvS19GwID1X0e5hNsNW2mB3V
HQlbZZM9nPP7BAG5UdY7MBayFLRWnj10R2VrkDSx4i1axUjbUsuyYDjvfyiMO8T3
xiqoix7Os1BPcvRtLqHEOqPnx2oGSHZi1ZLSw46HYylxzBel85yqIOkgdQ4/mmtn
LTpG4lPFUwqnYAMWcW0vZ5qUWGBMzd+6XtUsfSmqMAHiRZqm1sjduWgTQn19SGrr
jUyE6hecBhXZJTOlVLAREtUgtpPbRS2+fBz/e29BeJ5y/8Ta6mTn+QSg157eIFYG
ubKd0y6kE9usJb9dBgHo3DR5gu5cMw54rBPZUdhEppRyGWyl0+J7a68JaM08dPTC
HqQhkVx7Vwl5aC73U/zAvsm9LCVaqw0Ecg7RM4/cU4o6JVNepsT0af6p6yrNQ/c6
rqVqXyJSJeVMuHcFtgdA9Kj3fvzVOuue99FmL2Z+EYVsuTCHT60AiMlPUgIUr+kV
L+uqwn7f6FKnXy8nRSjDqlgeiqjEIqeF0mWe5CglpMBU6u2leHKTxgBleUAd5+gY
2T6TJvH/arxsVKBzbsd/ehbTkD3qG3vgsun7xiK5Kc+quRz5opSQLkw2cs4KOYZA
cb2x013thBDdbchTs8xhbU+YEj08JDWXIyOwlQVkM8jZTZ3FR/bJW/RHOeR8GbEb
xAdPVQzf4+S3nmtEiG2ZEaXJh3gDU1yAdq86zlBVWLGM1IvUQD34AyvZE5Xp5sy/
BKn2m298Yqq2uiREbRq4SFbpB3y13HrpWr2yF33ZTTRyptsPRc4QnsToF2QsD/Y9
ClGDPyLWZaukyAZuGQWMCstrtOjqzC9Ki2SNm2J8CgTrAYMm28l6jJFf5Dfpdynw
SmNM/C6z8E2/+PWU9JjWd22saGkhWfHTzvjmMA7Dw+d3B2gvtkPP6WY6Bx7BnR3U
nvSyGRZtMkiZHU1vkS4Q0AVRH7LODoL15SW/dokrEutldJf0EFNGUnWNW1Ev8RDN
KO32PeYBGU0TrMP9uLkPa6GKV1S9GHJZIxg8f59uihXZ65sC4LUwnkG0Ry6NC1Fb
J/zpfd1e1XXdm+aOmKdxnTXLx03SExQWhoIPgrXLgdygKLwrwS4YI6nyMGJDQVbd
soRzCJ6JJ1+0G+FCrHkVIFrZdAJJApqyWZ9gSL7J1mjMBikxylJEhOjjw8nJQw3c
rh5nfqwShS+XWA+r4eH1JEBWAaf9Nxiw/xJffrjc9K/uHKSiFRhNJc4STNjMsQpv
/Ue42fUcOdAbhU1awxmp7LKZHJBDnZcsa+MCsqSGckVvcjh8y1lEQspsPinKcynI
yuE84Pr5/WoOrD2EcwuKrYCUOEAhmT+AiJ+SAO8cmiLQcQfL1LSjEewLRqzmibS2
muMKl1j/zXVNGXfWknvROhnyCaa0z/WVzDcXUh9BPYSzcXKQuYxxo3R1Rx63oteu
KFgLbqoMSkiXhLoJ8w3FzggjbfMBhxB1zCiIwB7HXXE5Yj6KYd8ME+j8SK6FwLz8
YWM9QiDnqKiGW4H/3OCZAlzvGVU2FhVwC+YizdMmDiq6jy5p1LJ7Y3wQH/WQ6x8+
hTkbsiF4SIpLR5jZqMNDfj2h0Ffx7TVjK7NUBHKGemKx1mQ13lFfQ9Zyl5fQjybg
wZhqZCNSxK+TJFgw/ZfdPbcu7tPq2vTadKkNQpgcG+i23WMK3topuV4UnDWqSc9I
1AYBw1FnN9Oc/nhbrwGkTHawE0DgTNL+9cjJqi84W76S8+pcDKZ2KakArrFzC7Kp
MXw4jUoQe8tJ2aCb5Ga+VfUIKq+XBDO3gSp2w7jM2lQLiOn+paVnoOKEL7tvWuvh
WMA202xeQZFDNG0/s2E3VT8rffQCy0vIERv1aPVGiVxS0DMSmirmXPD+lxD5wB3I
ARdNgdKR5bKVus+xIhrdgVPfbVnwUT2quufG0xUJ4z8el5b7pbr6mwUx80bu1RGO
4h6SV7sZpCTOy8DJhf3YgbrFrlh88pLbP29DkQnu+qtEWRtbF2h4i9MvwZNrzn3Z
8ObnSpMZrBo7mrPD2C3cA9AI1TdiypZfOQlrtkdKh1X43LYCM07nZDkfd6GnCvLZ
HHx1pfYhiyi+lhsmd/42zA8fqoNoHag8b7W0DHf7RXYW/LwkfGvsxSPd3JRXKTMl
SwaEtwpUgC5l/XANDn3qHMibuvYYOgJ+YnApJ7GGmhwJHJkioBCC71PMFN5LjuG2
Y4TOLknpYoTWhy81jxUeNjPUUbnRS+LWMQJsn1j7Sh/SyMc+n9ICBHxafFm0niQJ
kKHdsBLYshmiKyHPPCFFMqeu1ZkXc0Snc3x+PkFZQ3KcqMEVhQabZtkJEBqVTLFl
LhzNc7OfFqqnewxWyHnZ7e2Wue1FK6rY+EU/7sE0+3MkcF5+Mo/VzNU8G92kVy2G
xCfRoCeEXBFXb3CYbvrmJaMPoMoj/g42DolrisUzTuA7YMJWTXlCT51K5oNfd+dR
4OmLLdEvNNBLoBZPAU/SKTsoJ3U4J96JG0p05GqRPgWyY6jGdjGTQTL+f9B9CArW
kD9a1uT9fq4e8hWq9KOcORHJpXY2K/q9DbplWnoDUI8Os6RDL42HbF+RdA1FXUWr
nVFJIApHIeEn6Hq/PgC8wXHuSnr6IyXqG5QG362SPzEczZer4uBudWOpjHOyZ4MC
Qade5cCJhSWkmuIm2XkhKqMNjTuGL9HJdoWcvUaMU7BZwkGKBJDwReMEAAZg/H7n
QydbUdjlVaA37lBk37htCXWd2YkX/y056f405bsvy5ZKAy8zYTPyPlcjaACpIWRQ
7SFUaT9iwuNSP8G/LHGoDkBnpokpQ5RwOdQ4nm0dQ3jXvHrLr4LXE3+mWxRx6hH0
sq89eLMQS5RdeU88PX97euSZoxd1weVsOjM0NMDgJXAHh/2nMEu30s2hAfsSt05m
QUhiliaF63F/eHfocwhBC0KhtKHKRxVvKSt81Q6w2Q1ptMIdG5y9rDAwlgFxd9ZM
TJ6aaSwtlLAG24JT3QLHTLcqLUeqdTZ4gYlX/Zdr8NbcjAvLi7iH5XgX61KeZZ52
YYvfyzboSiDSM8M6KeaByoytZ2AJyFOqOCx3OYvJdbyOETv1sFPuoBFAjPTVO4eY
srSGyILDfHszpLoaK8yECETPAqaCyPUunLeWyRsbb1ci2WwUGeTIaKE1Dp4t2ZFN
IUxjro6dM2lKxDkVRLiGAO0vLxb2+R0nXjGcD8LYvz5p/mYUPLWaV+f2e/CJ17ij
Gp/WDOVlIO390UJVqwxnh2B/0pSOqCk4sMAqc5yxu0+OUzvbN80U7lhYNJS2XpoG
KsX4PRLCGL8i+QPySP7hqXyVASZ4uZUpOiq7Gk9kwX/2kQJrDRO0+m2S8U1npRpW
7K0uYVcJ7U9VuILX1yhdG0L8h3wb4ITU/S9CUCKiP3xEcPfJTn+YMHu8rjfq0x6Z
hgJVkcqi+vdFMLKQPZYa/crl6p8+8KPashtK/q8qTErxy86Yk5J4GtHzhQgqSVRQ
EyAKU7GLMNDOqaIP1UdcROSv+cTDObsE9LyVBo3Sc97O/YeqiTgPke/+xVNixIYS
L4lXTq1SonNvU8y7i0FmTOa/yo0egrFJ+baLBOWvwFiWnZJ5yeO3raHG9EZ+Ct4J
vf68nnDK6Z72m0JKvdwHH2fHI4Zw4WdfQ+wxvxW53TxxhupTcoPGNCWFI3E128+o
TTYu0D5hq8ndF6YADguUNWPWC0LA4otHn4rjdF19d6omzmcltmHgElvPExohTQM5
wqQUqoNg715zd9ztG0+sXFZBljjmjR3ydMkMIV4ZBjzsTUkDBadYa/JFY6FyER+/
yXvMaFeXTLoFsj8NAcYeavPQImR7SQo1p35sTi/NizQSbWWTH4o8ziReFA+Lkl2k
QlUIBICIsPCvDvcOoCZAKUSz82VWKOGmHTRtq8QFOFje4GH5vFNREFdHFGB0lf49
AlU/8WaSQT6OsdAUkgwGQsj3DV/oCeeR2xMASjbUIkaT5z72H0rwYx8itFGKLY1Q
u+GkvPdaDO5DtRqQAbzoSLI5MJQLBNacrzfgtHmmU+IKcVA4P4QN4r6ZRAIkWVNp
+IfyOr1rObmIaI9gFE9+uAKk1ULmyRVNoI41WAIzUtVehXOYw2orKp/7cYmSeRnN
5qBGytlFUIaOBUmT23NqCgw84T9t/9UyQjWy7gX03mDB1oYUEc+T6PMMjYOLIzzz
p1aJl2Jd//sgni1gyWXPpXd7wfSJVW4Kav7+TxzH6vzjULVS1/6t+4n4TCmeE4hJ
8hiZCt5rCVoDwzHozLnlgvbsUlq1e4qBz9Pj6BO/emUNe815soYMFIGOZNDJWgr8
RweGyYwTDQeEkWtE49q0cjhERelNRHAqm35Gp6lmbIDLwIuYIavQ7IVrxmJatTH4
yoio/5PMYhPKoQShhMvHEok7dE9qgzX/VYOG+ntRt+Ng7JjouSMRP1O38T4NWSeE
4uKmxyws7QiKIRzpt1FJuyyGyA9VNAehnkotTSWS1x6cQ1cKwsylkvh9EfSUiIig
r/WW7Ai/kawZ3fxERcL5JoBu+fKitvdK2tfkDiXViJ2/iRH95yRrXrx19AGl+PzP
rMR0Q0ghLnreUShmsYq7ziPri0+F9M/uqpYndiKWg63j2AC6wcSmMEOumWdar2QN
6NOad65bAJNVtnd/cors1JokB0bjuUWyyT4V6GL2VkSJIRS3a98QPRj1q7HX8s2B
T9D42kjaX0VQzhH7yrONb5OQWd3rxV2zFHb86Nkbad9A0XCBTtY14jzpjmJrqksk
2wp9DKdKU6oV0wRp1eZYQ/+R6e9eSHAxOPJai2+dx7BHz35P4Jpb+KnctyNhiyqj
u0ZjPyBrRHiqmXoXNgqI1tOkx5Ea8FOZjV6zXpDIWNtcPXeTw7nnsPJqVVdJ0ZQ4
1UFhnpO8RwwpbNECdG1T8Te4owsD1DlnjMRtOA9dvdRuqBFRbnDA9+Y9t+vdhdQs
wLFRAlfKtv+whKKmRIVBIlCjvruYr5yLlvP22f/dyJsW26Qi9RWhRsKgKrXOs0ru
SevyFOWyaJE8Te8s0cbd9q3bHFi+F7qQg9Q6u0hPZ76PQLC0Pj8oReynpzcvaiBM
C/FIJZVFYDewr9ecn4JoxE/sNok4ueAGRh5Fb030nDkBEWSQXA+SrHJ/ywoKfMMV
NC61RevkRDgV/odRvSKNGH73tjBDKHee277mV0ZT300B5SebElf7D8iepztPlMDf
ebhtc6ie2re0KkLIGx04Mr71BDLZ0LlAC2FGoj0Hpf2v057EeHbjW6epbCFtlxFF
TReicF24QflkJTtwTdXwFDCC/ssT+BqG0k2Nlsr3E00YlaWA4rmqeWtaJ/uYnPt/
N+KlsZm4d1b4nCEfwYjjFy6OoXFl/F8KsxoZ8kFFQ+3OHkUkNc+ci/c9XY2XM3nV
iWMGi/GLGFGFJF3dIo6t/Vp+4fo/ZFRlYTzZUFXKXsfONC4Y0rPStCyp64dDUNg6
zDAUpRmNEOF+88Z3tnxdn8atxcj5CMph44eeoEmzO2MjA2og0EhPxe5uOnyxsFV5
Gl+Oah043g8IIPZcMMgfwvz5GNVzWxTLEB4hSospGiTTDH81bPntLdbB/8jB3QMP
8sr1iTiXSjaUVVLxkapmBKwpakcrWV8MgQ6lFn+Dv3iYq065M8CF6gNq2dZsmKsI
KapYuulysWBCfY5eF1lOuxnxON3xf0h197oFCfB8OcPtnA+Y20Nae2Pi7FvTPzai
khWCnH2V5eD+H215XqAR+Hy5+fSySWSR+hcjRh2jKanibvcKFan8FBRMBaHmA0dh
1co+c3CF5hmrfuHjGor/jz7WyrX38rTTQy1JR+y68jM+Pz1A7sS+NXYivI4UbjEI
ccqkBNF6ePdKwNGJMe9NNUjQAdA8IW9m6HK5WcsSrTpO8FPvk//el+HjXOCAUx1l
Cyf6k6eRUuKBuSyIs2HP88SjUcttW7u4oGZhR1DBrRlnGK8mWuPx1WzDjm3+Fx0e
yLavwTs0G4uq/LlBjcBOIV7nTLxubPlvPAxBACpEHcFhWJ/Imj3qpUDoW4jozRS1
ToJVGbhf3BTeEVEqrM9rOvLhpBMKu623NXNwgOqVQZutJg7BfqLrbCdr+9mOe9dJ
opFuxsXR62FtKaMPK0iOG+DiQOkYzaUQtyxmola7oc2kBf6fY8B5lnl1B0q5OnCJ
mjqaeVCegDuDm6I6RRDpzjDdHI4YZ8zAR7+dKI8R5mSACGMe6kHaU1S1+JMSXkA4
4N5G3jWQjEuc+qAzSRbQxsztxYf7GYydvxQ+nAO1pqSP0TJY4n4Im5mRxL4tDEhI
RkioeKWdNGVGQ6mV8/MSBYJbEbU+sVR2ENnxlDuCsgjEFN0M5EO9r015LXOiHSZD
o3sxGKctxDD+U0cHE5qGxUgUUPz/l9SRp+QYaQF6X4UNZhlM0sfWdUFfuDbm5+Up
MV8+C7t9/rF+o4+wWFAs9qYjLz7LbTvkAytb6bxi1Eroq/VXDqS+2CGz8TXecJCp
8mG2zffMxJi8cOWzuavOZp9W98ZN5zGWCk0JGn0UW9UHMdIi/gUbkT2mwzqv7YVM
6yM1vjdo/QLTjCDNIkScXwzy2d0DOdYU6z9ZdrUTCORv4ZuPuiRPCpnxGWNDUqVv
Ph++z9bYZznUcvAZ+WUAtqAqZCrMBp2a5RIddXrq6yM3Rfh423ABOSAT/kxYoSmo
wTtjqtDDm00q58letAXrq0PQpzNVrrldetlDz/QvtSqsNTpo6XwmkaCBbxDaPCqP
NOQTS8Km3Ye1+gDDZnSXR0HXVWgJvPDU3TX9CuX2BLLQU4TvtbAqPo8fhJRqJlHl
st8kzeJ6rGRekfNGZ/fPgHapuR2TjWIuv6QCOnYKwuqu/D5ayC88b62nQmsGUQFY
+hg8eX3sLXh67SRqgMycZTaW04KFiyMRE2wvzh+ioLcjcmKxWG1CQf29zuD8rsQZ
jZ4v0m/5CqZGaEL5CjmlAk8ULsQRvrG/eodzkpUkhebQ0pkxvAk7SyMRdhQAXtiT
s9mp+TWTkjKIlzed4rcHu6eqkt4jgPE5rESpeMope97LLAjSSoOt2Bl1AbRwI1/4
DJ6SYhaC72PeYkNK2QLGOPCnwl1i0iyH8ZqACf70tHmSWKIDxGq2dLlp2lqiGnkc
+wPHA3rhxv5iXF2SkryZzxnjQiERm71onRgwySlfpkK417acCMieZULyWQp4pfbj
mo64QpWyWcHHbPvYX8Ib9zo/PdSyVtSGC9xx6P7EWgbRe3hEPRjhQv6JYpKOTfu3
9/o1IMOHLwUNHfoWE1pAmvGwbJapfEDUXPMZ4KnUOGd6gdpUrDhecKkhpOqt1nau
ra7dhUBtl6pQwr16Xq07peCY8ZGJNNRA7hIAd+qwtlbjk7GYYqfVGEIgas45unAO
wQKmBGu+bGzHZHS7caHmhvqrWTuu8kbgwUlE2vCV++CXI4prgAOAtcIsrQ5sOEfW
PG6Oc0L7KTtXG+yTVMvfULSzi2A9J2ljA7ld2M1uO9AnzcbJkAtVka2V69U320NH
B85OiWyy/IkY3/OTgfDgC/RmrFhxQPGgjrVOhIeIQINMYo4E8vj0TltxGcLMW+hn
BTPA2w0vrHmW9tWYTFnhZVt+J9YvNtr/4aWJwyUoBcuqMwAi/f4Fg6HfZj0YOJ41
u5FPgEzCOTf7ckDuFQbBbIJrwAVh3k+cBgy+gJznP62CkhOKrUwb7e3Pes5wrPdv
9CZ2in63SqSjBTGr/ntjTkjiKHsj0oLhzOW1iYGJi4T0KmZFjDd/NFnGCITyLyzL
HBDpcpkg3UYg+TZv1ODotdOP52a01aEf4bWiWnrzl3TzVktfS7uuJ4ZKjSPEP69K
SXpJk01rmXJf33GgoSh0stDQOTlpfPfSlDAQ/XirwESXCNGcPxWDb+2jAMDwvCY3
QTHMAOOIGk/hKRLk2Fmqw3r7xhiAVhYn4YqiYx10l07ONZNp/1CUHQ0oNfz9ctAr
wUVvGlJ2ChqnibqT8kX8rPPy+FJ3WEIMfmKanHdWBWtZ9u5EnVo2BhM27LZ/3Imf
4zb8SNs57GtGcaRu8ZHUwnasmv+QC8bN0638di49EPe5fP/OeW37qjFDWDhw05Qz
recYQDwJXp38Oe6bFGhnEh380HHeIMWb/uTcXGXYThviAbrWIEkn86/zB6AOoPUV
ZVtijapi0RZ95QkMCymnWZ/uaUg/O6qvMPvT2vF3Nho42D3e+2wkQBRGuey3sC1F
G+u2sS1ejs0yMfsowho7F6YPr/Ms5ZPU6LeAAQ5ZVP3MvfGrCOdMEc71r0AbLbJ6
AK/el8iyUyFbeS9G2S9J57g1HlYHdpjLdIcFaJCIcc2h9acQaly3yGdicSuxxyTI
/qWtVaWS+MI+PDDskn9KFjxw/70/I6fv1qGr73fZy7968uP4iA0yZ+rAtO4YBrEA
vvqMs96oDKBKRrTT/Vpof9zplg1T6/dgjposv1SdVbfZPqUnzCZXWgaNsBHoE0d5
Im7ADW89oIZ9nRxqreperepxekt9AVfULjKpdPCHiS3f0EIVSyEpQLuc4C3Uc9Fu
YJRwAJ2KHC+o1zIhxzdI0pvuW3nuwv+1R7yt8IGGK8UmbQVhdvjLjeS82tBtGgD3
cJco1/FcX4pEH53pgaD1SUEtT/ri1viZdV1Gz0XH8NdvXWlaNOrFgWg5McZeBRzE
QA5r0f9TbrWDkeF2vy6JWz4jmNc54p3u1Qd07ii0GXdUVJK4FwQzxjhSAJ9CL2f4
nUal3upC6Lq4/D7kaNkZjjqtSHXNJvsvhCr3EYynvoOSvmxDzq7a1sHX4T/8Hs2t
sn7NB6ohV5+R8uvmwqcPU1QZf/simHUAUVzquOMiJ3E7TkY1rKut7F1CCQw9OQmx
jdCafkMBan7gVXB7eSSOMv0ThuwtITvPKXqiZoONGlhgSde9MkSvPnQJ+ykTpUaQ
o+gf9KUuaIrSwxSM4zvNNykq+U9PKs35jJkMQRnILcl6IS6SEO95AQ5eWAwThxib
EMfvT+PFdT9zy6F7eypRoIHGJuKPK5QvpmRYClfYDzvylRpnSEOGHdPYo3bclFjz
0M1/oTUVfrXC5/AAy7rh8+8EQt8Qb9jnNxK35WCBNYkzCLepousZO9Qfuk6C7j7+
xswMqfOX7kLJos0+MYw3NX6kf2JBCYT+n80yMzeCIO/aFAygvhNN8u1eCgAuV9ws
WHR+meLZNXQs314ljNUxM6J0nXeqni2XsBtCDaKmszQs86Vv6HVfdWRNY50J9jGz
4Y9f86bdTTh7vmLXcDqmIkCbad6d9qd0IK03PSHhOi4lD9q230sanTT/GcIamPmx
HxXH5P/wuwIQGcMfk4MrxROTc4sUZERZu5PSVo0/1/iXzclGBW73rz/jbFrH35Zj
RlCMBk1vr5pAuilrCjaXOejhYPZutlX2FagEHDaHWRk0idSzwClHTMfA/DmH5ZJ4
JpDEI42wduQl4e9+kVvcofj2ewZbqVCee4rhi47Johs6Hp2N7MmknpHjmkquTIay
4E9SKVKtMBewwPz5s8U9hTyE94KWocRjuwOsCRfqi0hN9XBoXltqQlWYHiLX5iRq
h0Znkr2tX67MGWEH/5jzQYhEl/vHvJYoDN2QaEotIuocHQ6tMtZsmPm+I+VbdRAp
1FxiH0ywxGe4MjLPZMO11CpFiEc/vm4J2OO3w7Vg3RdNDF2gk4Ynlbk5vThv4cdo
jGRI9kUiL2wnrW/UGDLXDrS+PXE8cSgE3WvF/mO2VxJhB6CYA5L6CHMuo02LjvAE
lGy+rD6N2qGB0BnePC6Np1Wmiw7gNoXEmeWtMVRLVlxHKy1uGWNiune+KXCz45yy
JaINwyWZ/tUXhPb8AjtZ14e1bXbXXUfRzUujTsRTzPjDERF5ZGfsubDhdvkugWfr
BKqRO8LWJvVrZuThVjyeJD7MOkfOSbtiEzhK242f9FNzKSkGRR5YWbPl4FH6Q6Wa
fOGAdvSNrrJHCpkD/zUV+6hQLPm7bTnwo7kcaM/78uqS0j9Rj0qW9An4lQWFflNk
ynWIptsUD0q2Pdzpcqqk2IsstL8/0PzfaWGSb72Q99NjwFftsRUh7GLUMIqZ8chY
dvOqob0n7GBUZX3H7Bnq1bS1qG/gzC+tR82fEnrzCv1YVEcINkL1WNqmzz8inu5Q
WzbFtrvv+Qf+NhBM1H3lMbPTbJd5qLQTMglJ2P8O+km8v/qA1+aqbIzYCkYRVB9r
ToPnuxeMy8j4EKvGRHI9R3gJT81C0wYIXqZM7cweknd+jxUKDl4/ZOCLvCFu7hA5
bNeDvizWBm/7mmhTORawTPjKTzMcF2OOKw3o0IXSKVxtRF02+jTFHRCVgQje/xFv
svB9v253ERuYyoJQkNrn/pbD0ee8xlvXcijR6KNiMcpIkLM36xtyfB5//VcfDrQA
ojlt8fGo7w+7Id64O62da9fjQTsppLddmKwr9zkhlAUnDFPQcYqcBR//LJ6QOysq
mos2irvynLuJfnvasCihGETJcyYus0gTg8ceis8xD8TmPQ8EYZbp7FTWYN/V7djK
k9cJvpkNab6d0yvtFAZ0ZsOrEYbnL4di+FvLksJv0u+tY/inYqEpCId6wHPhGBSm
ScSipacztKAjEH4amRwZAz3GddN+YEkVjMBnPr3zM//5uy36JIf+C9b3zKIuCosZ
K9r6Wx64KgfqRbFbo5gh8ZN9NDCMLidh+tL+4dmvibu1zbjz9W4FeoC11pMXXtf8
zqu3Ml7m3uaEHLgtGFLOMYihNqhE1DyxcCc0ZSV57GEWyme/IEr9VxWO/LO7cRLo
6vXT/CuBMDa0fg/BpTEPv7edsPS1xCaMQgxN6Ol7Zj8fMeDMxgAfqZvgkvpxFWVX
cd89Sw+kuMCDoYonPyRUyTkyOvDa2tnhx/ICxOd/AnKORlh8ngoislKVl+PGvXT+
CviV+v67+cAF1rl7dU7++Jp3Q1ccjjRX4HFpaCwp5FgjjbVb640F+svnqHbJEWJc
OequeFPaMtgpchkNiPcCGxoUf4rHVJG/59xi8hq9KTZnRaRXnpDEkmkoEiOhM1aP
8rRfrMI6rRLClRfreUQZl+l5zPgeHra61JOcOYN0sIDvg4I9a32CU157xExOv3h7
KvImnjF9nA/fGhT3whTKRiW5ciKEOTyKkUJLNeSHG0QKvqNjsxK7ciIYaEP18gba
ajPlK5LyibMYgYo4Q8qbupnTlayT54v99WrWAIIYSfMedMwFwr2pnux0dDqQ25BE
S7GVmXpFJ4FlgmN2m89IFUUmroCpZDwop2PXSBrKn+7JJt6ZGmqOcMhx+sNzq6q2
KtXeQOUulXwVMpg2kN43KWhkyiXNIaB49ud1TNZMpb7OIRMNVDEfm2/O4vCLAoLn
9GFEuUEE+T4gMGTlvUvCLy6SzDbUdB5tQ0ia7lVkCmLnF+NnIdcEwnXxtSPioVSQ
GJPN85IoyOcwviBNnpE9NAqvl7JAkTzWnA49cmTf4AB16seBeWLzEAwT4P06CF0F
Ud9EDy/nNR6FOgbNBgQgWjZ1IVFbKDUKzQ70oSzuKbHxwgVi7YN8lPuYR5oRNeQt
l73r0yM1+6nqKC1uhxD04BTFuMmmo2Q1jWnwLAGJPw34LnMKeiRNSS2RSfNkQd0n
lowHUds/dyAKKSJt9VQRbAfqAUnPTaRHzmj4whEXIHuca+QL9whez9E1ftolBZrA
ZwJfV92iVh/mq8EWxkdg/mTyQOXOICDbQsbEsB+jrpj8BkUZT9d3p+51JMrUrDn8
gq2NZWn2F/mX1gAF+Yqcqqp5BewdkQUoYhulZrhfOuWQaYoOs0MZi3XxS9DMRDt8
e3qfdKei8bTdcTLnH6UVt3CTSzzy/qNPK3/d4lSNxCVd0ekiKuGADcn6E6lALMVN
70maugwpY2WUiOX0De+mh6J4yjKveCQJyRHDPyrwz46W5IUDxVECOEaNSyUGK86L
9xxfLMJVZP9j0gyVPn+MYBYKuhLS0ZdWdXH9tOt5lmnKIb+Bh6ExmNmNtA8yKM+P
AU9Nhzzh6SB8/P4h6P/o++QcH6iq7LWeiLHUWbIyRlIN55F5qfNG+gn9W61gCeH2
+g0JYeazK/ycLhdKkVeYZxWe73NFy55cKEFtU3q6pYvEbRY1RzY2dcmcTThMIvaa
hMxlLIFSPX9/J0b54mFMVOJsT+M9HWKR1v73fi67i7/q2r+DhqWCR8M/a6SwEfW1
NqnJeJcB6ws0NQNyq4AjwF87DO+XS+msKWsnclc0VJAIP/ICvRd9dWzuYfSi7lXw
VIpyi454PoyNeWUluprDMGvLbp1ze9kl5EM5QFhvAkABd9+lu2uwhF0hj5xsnmct
gYRRjunSnUApgt3WXrOqD4JasIwv0DlprHB5LwDEQce9+llX0vsVHeM/yx0tCGbX
YFVN54x/5Oi1J2pVVqAgazVqTqg8SAccIl0HIxHtRR6ZuG+z+UmZNX73xShP4TYZ
sn1MffO5FOlYCh8T4rRkmf+KDg2aF1CPE9fUzQav3U8/bRUZaJiPTZ2UAZ0GxY4l
8n0BPpnCBZeH76lukOoLV2zvHh/s2yK/EqyfMMuHnW4E4VUoqflK/rsfavMKW5Zn
EUKvMh+txgf7F6Gc1AJ3KDBRDHR4c/jdPbwDyg34PEtfgHeFpIT4fCh7uSoRNbVw
iSh6g7MS+mx/otXG55J3JBurrShB1GmfVWUEJkgCZ10YQ5UQ3QtcpvLTyFviyrmd
HtjbS0ixbd+doIvkb2LiYBX+EDJImiPsRY5cRig1GQnt4SeNAIf32EtMOCZ8D8n0
WxLJZ512oFxzhgiUOec/8jhgBEMQLI0TNxuTU3Po54+tdbK3EqOp5xRm14gJ40wk
MEwWkzHSWQy51AMsAp0JRX5SIqlvC11ftpO3i/+jJ7az9FuVV5rZTu4rTefJKILH
mjEGaac0iPFlkLWPpdlxfzFI+zsEZuwk3DairI9fdYOlRtNz/v3ZORRt3zXu2C5p
CPP8IWT8q8wnGCLpOeW8UJY3hTBIQ76K/IyAaKJUqZBh63/iw5b02AA47NDapwow
oU6KNnP1dm8/fyWZLzDuGicUcCrhTWtWcVNxK+698szYcn/PCd8Dqj/GOvTdAt6V
PfI8XhVU5fzvi+j1g1itAWCNq6yuG9YHabnIK03jrzqVV/zZX7WNUzy9JpB+7fkr
gI5ZL7+WdJA9hG/zsvS+6+QwpSHtSsp9wud0CnMvCbcOQgVMDQYVy8DyWuLF1be/
F3vzL/eVEN1qH/RQjC1JXZoBNL7t5DMCbvPoiFt8nBC/dfIqjee1LmP0Q9TO9Vyt
DfMM4jZJeM8PoHmiWONdzALTy4lPwNgUu/OZ9IFw5AsVXeAU/bmxEx4LbzNZ4yWO
IauGCZO0IVQIzeVzEyt8OnCAfjPjd7xk4q4VkdCrvcftuOlyF0q5/JqvaxjvlYt7
Kv6S7IKxGOTObvMm18tNn/x7YmbKgBVVCbPpR2y8i1l9j4upKL72GIX3cyfS1Ykt
NMVDp6SV+aKzW8UmOmbmcl8ppT3DU/Om7JoXrazlOr3pXtFQTT6GQ7+UI+TTYLja
Wobd0MhcBwxXQfMeNkrOhe90EaLdwXGFNHbmRpHfqVD1YOFEceUope7InUMzRwGQ
Nje3kE7HXoD5C1BMAHoZt0qF/nQ3co1gbrnzg7aVUykzLYZgCxDIUDkMVsHV44tm
/axLWAXovP7WiBhzEKOdjmUS/Mchp3JKNSYoEkdhcoBWc1kAVT4I9jnF+/Y750/7
hKTYcpwZ44voVy0Hn+xbnag09DAQOPQBECWdZU9NIsTBXaxZ37wWuopLmIhvjMLE
U5akDjW8twxm++fAvBVQ2zJx1NIs6Ty8mhJ1guoV0PIksKSM1aYllev0M/EHJqIq
RxBNAOaVZCWR2RJ1dUlfAGMdC8okzHZmW4DmiakAtzd3UYTHguAPSjGiUHD+i5Vw
uoh6Sd3GH0MQ5+VTuSTL35IlXm7i89Pz6hEoTuUplTSLRa5TTVsWYgGh5brxOZhb
3dD5VTlVlBuYPZQs9PGB+c5VSIJHVYSmbstrUXArDc7tZO3RahMB+pkicgBV3ees
i09nlbkqKBfd7Uwn+vAsgQXFnJxmA8k8VqL3jV/9x2h/G+rxQPhms2LS5c4MWDrD
Xaa3gtpwp2sG6UOtszab2IMv2SXXDH1GXJ0TQc6UQX6yUJSIFVNImrdMmemD7mA3
N0WR6sHAFljNvqlgavEAEr+1oSWkiluGpetaoLXn0Ey/E4ZJX4cWRS4LAfMDaebN
qaktTVuy+Xxd2lRQ/TK0LtPH+6CjqJ0By3PsSEEJLkoQNkzJJKXfEoOX8M1LeMF+
EOtkx3KSTxZCK+C1yO/7cG9BAeNX7UH8vfMTdPcZpRgPKOvgvph1XPhdo0VyCCgc
zl7doKgxBO4mVpNeLe5g/LlNrsw4+CbM560rbAPEr0IQmO9WZDnKktemoIwfbvn3
bWNML0coWZbxjqJ7bdAm5VB63sSQAyihDZWW+j8UmyWMIYG8foRMwWGHZVNhc7De
3GXkWVfiF8umPcxLrARjUhmZwJSEQa2VaMWf8WlesuLmbmrqXvrAAUdpDH12yILi
z5ei19BF8d/G8Rp7GHfhhARQz8W2T4hi80C/7zCCvWhfnnEJwMI1/6NRz5kkUdzs
3kTAQwwvZnRhse7sd3ylMaLY2QPaIwLekc3UiSTkeJOGrm1nT0+yZ6X4hXz6QkpK
OtbezeE1JyC5OXZ1gZQAMjO0faLUW3sJvcCF5G9Ym6L3bqMaOaStAoNsAYJhp4qk
X2mFsLlVgb6cba12fbCFDH6Ewjfql3Q8iBX9Ke3Luwf9IF261BoS1D4FXA3eKtUA
pZWoDjhl+sR1H3yoxTIHgwyzbEhoURFZl12KnguMnhgEj6T+ouzR1i6ph42y5aJi
htsbsFd9ahWkYs04GOH4pPBUVVCwhpvc51IAChoVUT2znJm0BMNlzjtbcR1Cacv2
6OTx76/rc8e+VCMW+qYx+IupMXfOsXqWw/KDF5iKJj13ViJ30vqrXG8Vj1gIRTmu
2B7xdcuxSdg157isCd742crvp5msiCcjXJLMqJcOjQvKSQi2NNLgRbH9+cazsGOc
EElWjEcbtTLVTn55nILL0qbxE/nbpxOcdafYTzGvMMYK3KU988kk5lgzKSACKjtj
kGwPvVAqT0DwU0v8G/A/H1z/lfYktk3QrFL5AFMzDGsCJ9pA2keN6nngPhhQ0uGv
w1NDjNRnSnh22JAlkZ2TGMov7kAmJHrxNzQFeaPkyBW8x5Jd3cqq8s3iC/TUhtOt
f53BFEhnlBF613bZ2R1vsT591S1Rr83Zff7JdPll5s0uvdq0flC8SELi7jHnpOiO
oVwgsEDQQBuY96AqCrGqRmzEsX+KGKiDozUi8WTAO44Etlo75nLA5gS+7I+A06vX
pJsXdXTgywXLrj+9jCxVDsIuYphAowTWZPilOlT6HJwlFg0GgrLcX/iWcPJN74Q2
QUkJMEdf2LZiHyXwqfHjwsO+uGLeFWJZuPVR0sTiIUI5ej6WfbzlesDE0LkEJnfG
RenM/76ihAEhQNm0e5X4g0jNjUauJNln7UnAkoI0M9ZJ3uC2w6+Opb6uFzQY7WIV
wEQXHRbbeREJZZHo8WG1IO0MIGOxdSIxYTuhndjEHb3w9A4hwJnN4AZj6QSuJ8bp
NNfLhHdExDiDP8Vx7XWpGpJPcs9vOAq5sEXtwhCqM/iF7ZshtwFbwE4GIsRjk5Zz
Pnh8eemVgMDBur5A0XY2B/AycYyoCTH7NSo0bY+hm82MM4TfoQSUNm8Sna9QB9MC
dLVJH//J1bTeanp74DRdLeEXA/SJYDCAptIWx2HHli6WDHZntxuhX8HRbm6ZxAoQ
R/+LOZXrQU4WuDqbF9B+USZwA37+GgToxl7/3HOGXC5VLRQVlm/fadJKZi3sOg6T
w6SEIuZ+lxHT1Phq1k+4stZwdvJiuEw05TzHGFRb6BRfyd3Gw+GgZ/U7vytbBuIq
9B9IEGy+ZZazrWg8cBXVjylypvViBslM/vElZ25wLOiXtGzBrbdp3x1E73TrrmfF
GcVLkNwThHzhIsDm5TXx79GI8oU6HWb8gFmh+/DRPqsD4qB+WUvJJyoGpkraqRGK
AkqUnxJgSz8bnZh3o+bwwlGt5gx2SQHjuaD7/ns8gRyOAHUc2sc6+ToOkqbV6bLg
W4/qdvy2k6ytKOUk+ZebiREyoWK/alLChUlqhPESXo5/I91bzU0pE7CY4Jq1fB/L
wj+BehWKnbTXzkkhAerzKBuX1vvlxUWpwY31hIgJAr+Xr+zjhFGeREDOTqqpS9ep
e0cv1i4X1b5f6KBWQ+doROI7TUXFM5Pr0CfJf4t3qgirKQt3knmqCnuFVw+eOYS3
fYFW6ispe4z7qAg1VqoP+CfqHvwYET3pxt6toqXbIx+jN2JyTDxQ1tm8OtcRSxWD
i38zjoNcVPJe7mXy0zgKdbkgylLVU5S/pB6A2RpxyAKKjMVarKLkLPgx26VrnEKM
eTraS3RM+E06BeapEADCK76V5uqMijjotyIGZj2WdBoKFV/RKBgRFbwkMKm9X7CI
siH2klx9ctvQjJgAhMXhrFaB7dXCvhr1NvgyTDsui9p1hrDi/zcjvE6wMchUds10
GDqI4iCfu41Ic5I+m0QTVUeGJoV94yAJUEkk1q8AnXgHRvfldw644i/WYNanzvHu
5XpY7IAjdeM1icLAWOGDLeRXkmQWmv5nT4y77BievGBz4oOs155UJiBwuD4TPp8F
RCdpqjSlBQe9Q2HfPOYSNQOqBGw7auWGAGZZ8SUszcVl/YTIMhGP1Wj7ftOx5v1g
Zc9jvqPyul2muABEn+aq+HjIrZv9eY2U865FkMA1lgko2y9JXkLrftop9FBOg9dH
ANCHhh3JrGqxAKAxWKMHBOnpjgFAVNnc9TInBdTI8XhP8hR+NrcJFecp7RIoVvLY
1u4DzJe7Eumy10eu6rq1KW9x0PKan36eynfTH1gVoIUmVFH+/X4K+rV+OisqGmXg
4M4OSd9FeYqOWsg9C2ePiWeLJzxpE8TtJ4VcPW7iomKX3S5M/QFsKYMo0If259sg
Z4MH1H3sR59XlHYTg0R7U/b0AkuPyOvwhxkt6GYkeGT//58xlYpxg3VWEoTVyJ0l
vQ2fFKCGqm152c+MB2PuY7ZI4UOfoVBYxcsZ2IFj2s5ItdN2AJDiLl7WVpUm8+x3
KNHIAYqOXAyd9t8kg/Xa5TX5gVERklRKlO4tCrdhHeeLuxSSyT3cbKVVLCjI0Z8k
KTJxvOJ0u4tU9+lI+TsuUqj0jvAsChMZJu7EMJgp3vRFpSoIrXmh29RvWFJkbNQB
aYZUKaWZBr25Ytanx3Li1ooUB5OF/sdLq/nTb3ItQwjBeIfu+e1dZBQXgn3j+j+n
UghnQDsg8RM/Pgj2F7FgD9x/lWdIoL1doDcMShnWpTuNKXHC+VFMjyOBiFCFVZCq
sKdxikAQP4Hh5OfUmf/6XVRJVdMAWV7ce/5w9bzneh6SsQHs54JSqE9XjJhaPTx2
RRrEXVDimlBBACvXRr3+nK57YUikBcmpU9z168vrzuHYvlusrT9funcvurmPhyYF
Sm4LANAdi6EqVVBpcSljNKc3YMbt95n+EASfVV/yEv0MpeweJ+FNMEk5wLVPfNbI
Eebl9F2nIdNDLNY3ujfuTcZDg8dq6/rCWy2KH2587BhNi5OLFhg7+G9xhxY0wYlf
A3ILKCotTArzmZjUJ7KkgXtE+D9nnKzQLCx7xPTCFo9UJPr+Iz8LhIABnul714zx
OJgJ2TsYeaEMMGjiObw8OeM4wbsyviTmxobbG5Ry6G+XtMfmHuwnnE++EpflOXn3
qJMlaRh4erRSXIqow076+7WieOhLTa+uyMov2RkWiven7Xvi52ABQNYuFYZocu0R
BpJ9ZjSPV93NBx0j5W428lCy6o03GcTNnXw2KPT73rB9dN1siPpTOSCtOrnl6sXy
R1g0s90MFTniI56hLxuBVMPgDwXPbrqIXJA5Ov1WJ8P0KU5Odi4m/8tMV17Fi8ns
WJitv2zEkXanUOULbzcTDKtrzhKgunt9H9DkQdZ5Mbz9zrxYeHKSiYfK5ioYbIXX
l90KwL08mJuI31bXV/QTruU1Mfp/r2SLDw2Kc5+qGg+CNRBFJnE2lGV+/A5PzabU
S5A/6NBlOsdMWFRfwdrYtOFOcWMVW7tepwkvowHUcj0wqsnSusO3xgZz/ShvGfrU
1HJFnLZ2YMse2xVxVtCgzU7DEUTzBFou42R9TjYEzitg/gVCAdX2vZMbnwcsfhD9
jNL209s/bBfRikduYEQmExGj1XeBkOQmYiH1h/8bFDgAVnZrtwPspZT/MHzG4rWF
UWlMwDv7YdG4VKqHzDrHtvpU3AgyaWOG5j0DMWs2FTl2NPKWoXmmpucV4LZA00eG
IvKY9c584NxAutDXZiO5z0k96fUnPnvcUiar7EEMXE6+SNnd6EgTI5ZpSkwHIqlO
NKHm9fQNgi9ILtmByA5eE0qhyyfRmIizH75dE3vRz+aYbd+P6RsqEI50msPqbG4a
o3TXKjtAYhmpgwzGW/X2juin4+40lx1CHjT1OMvLGyzPtlOQ0+GBLvjVJ/Dv64Ls
LO+mL1epx8rws6eC1HlJ7G2naAwkV6X8sUt51W2ZK4dZiPqkScIor7ShN+zNodcL
RawDC+bxrzc7HTHlliWB9yQ/SM4iqlbGEO8kVcYfRgQCgOlcU0QwscSXe3sdrJ+w
nMSXZHLNWJOOnJdtnvkHH++9hISHd9igX7xTIthjzCHycZ6ZOkgWw3jLINRSt0lM
QfL8k1Mdsywvh0wAAJ4lp+JRfGCf5nfJD5zFzS/mdiNcs92u1tjYaiF4gVfxfrzl
i1WnbLydwu+ecXzLdFTwFdzh5z5PBGd4BGyzXG0n1XxkzoJyv2I9yStOEy2jVR5g
xY3X/G9SB9CVq0IxpV/bM9NfiSh5NHEb5Cgwa/lrAHMVsG1OXTV4fvXZK/nCSkxZ
ktpzA53f0PNthoh4JPQkwzDOeDDoTjR+MO2bB/0WeRONJHZcEU2VTHEHuEi4kk4B
IJsM28zT31Am8KhpgpWVdTtb9t6z741uGp4OHsIXGIz8UcAsNjgHXtD4VUps3KwZ
M3TFbKlA48NHniV9GgU9wrty3hXyBsv9pPz7gp6Us2sjuU+808U04tGSi3EBzCyT
rf3CiwSaoYlaAaOrLZozp0TrJjlaArQmKJ/EXUZVhMBo7j12X/tdqe8su/FXGJeQ
fHsDzk3wdVTN4ClDRQZGdzaM3IkEbd0rtNtNjoah2oyIZsp5jTrmSrndbaPpy9lz
35zwBQfYtD7qrfnQnnBg1a6dXZf573PZcSif4M8NZUB/wTlutXcyUWVIGUT81xW3
l8amGqqNhqkXpvWSJVdfwyOTMaElMkLp2hd+/f+9a4DIydZlq434CLu8uTrpQ7Qd
PnivxWJkgs6Uw+MJ3d/XvWrNJRmEiX/HTFvZvUKtqmr9EvEyiw705FwET+5yd7bj
oUUghUSV2VMEEHgFtdJlwHf/RUc+ITBmHyyqv+UOwO4XjiWYgLzlX2bhNW4jvxzv
wgQwtGStsbb4iLCsWTgi5DInNhbBgEnf157KGS1uvfl9QLtgRJ+afThvDQojMpTl
WJBqiERr4qByDV5lKpPwvJpvn2KaH301aiMGXCaZ8nOiN4rPE+EGiX5qQrFh77eT
SI53C1nMSz60GCIyKswf5y+Hu+kSYTDdhhJ5YI5TBRqvVUrNpVLaG86YZW2JCmdO
UCLevnZF9HmFq4iPHqqHximTjUbnrwHIksFb+H+uCXdmwz751LM/IBj++0HBIL+8
34DOKJNGW257xR0xYzUnAa9NV7gZ8EtLd0GYwsDs8SGpbV4Q72+CeD/xGJh8L4M1
D1Qp4dXa058FOsMJ6U84JVxAEoQAJIpLRuVfMXNPPZl3mXDhUWOMm5/R3tnEcV7K
Co92yGEzrRF7EEQQbGzKUx6E4W/yNyXvMCTw82NML28YAJTv/E+5fmXak+2T8/ra
Ra4ZVSMiqN08wKCi9GfXdIJCTZZC/PJpw4Dc4WdjZRSl56oawNs7/cJjbmiUYDay
6c/sHpkAzj0jQ8sQvCelWNLDezIaPlP1CYxVvywGv6ThY1ICcGzSC0kazucxMI1l
ZLeIP8aXbV/htThG6MbQUKNdKz+o7Bo53MunY2IZPB6Z2OwUL/xgVx+Gf5iN06ci
dBjoQmr0XmLQC7/IxdtOlMv3SxXUjTNDS2vyBVX2psL94yCnZOqneYv/RWDr1ZXQ
DebZkEepAKs5PowP4unrgGw421rhURdMoY2WEUe6qbf5yh+VQAmGRfb4dBVaeXxO
RUcSjLBzmjaz06XZoHmrHiAj6yHuH+1IP0BQV+34dXxzHZheooQGQ4d65gs2VDR2
f0wJdymx24k0T02d8q4NJV02Hc+R9VNGW7dNLXjOfwdIyntWk3WY8s5Xur2ZR2Yt
QcRr42WsGqDunUHdqcqZOp6KCDaUF+K8rzxmidpcK/S4Jbsth5cq8xjqDSJRRMUv
r2sSL7bWSJjLeP0eQljOfl+/1hvg158C8sBYpAz62NFcxLkS3iYTzp3XKRv86inc
fTcKnhSIW5nIcZzegYT/7u7dqSIiyZrT0N11R8i+gL3hgxEgkJMATA7D3+pK2aZq
tTROvZ4AxZYeSvWnPDZBughDh/n5lCKdT53S4uFIlXCQN4nOiIi3AvKqaeMr3Jva
daCVXtkW/xe+bXUB9nne0KUdIt+ghcNkf9MEadFZhrMDGDH1femSmbF3x1aj8fZn
gqvXDhN/bJhTAlMdKIMXwR9PooUHh9n20/ToNjq5N2DHE0ZzzXLYBjknFmJXWq2l
SMiULLhDsnEBGtoODLmxkoDvg+0pj79bACJFMDNPX3NDVst0Wn0s4POxik5B3LGg
TLcJ6JHrD4sspzmpdK00MKV7CwQL8MtnwEhcXDMxXEQYv4loxef+rDiPF1WzB4CE
gMzVK1SDQjHLEwPLOa4w0DOmTMoFOz57V46STZvcOZrTi98aCE/VL9Bm6n79hF2k
DoWNZEPR6WeOEFv4OngjMHzAuwdd0mi3V+RgzxluO55McygaoJt7h+xpmtOvLwXX
KRzhb565ojRpHMwwUBwttodbVySkMJKk0ILCXqdartscdrfI5roZdMRvN2f8y2K1
J1QQNMf/1sahXy6tf8taBdOUIKMe1chx90vgDB1m86Bqknycu/6FEcCsWy2oxau1
DBEGbUrOMaKxjt/Hzkl4YUOh/u4VIUqoLS0jK2Be1ksn5Nxdi2NgdpZxPDLjXohl
UUjxpwWxHkoWRvmjRlMWO3Y3lvSJtzwjEfTyy0l9TTN5D+S+5GvkUmjaoTwDQcgl
pyxK+E4qyWGH947/aelwzNGEjcjrspBSFCytGgPO4qrhA0EeCJc83ttgLK/nVXaI
bx1UCvZpFITf3Gzq1/D0svN9WjuO4BXR4dFkS34R9QwnrYnNwKuVOt/BNA7YkdJR
k8o0YX7AvYILYZyDycXaHeYeHTQR96cKKabHePnNdWXU45ezfWqTvMHM+M0sOqlD
U0h8KeZgNvmbioQJmYJNN3JyXfn5wRQLbhHHvFz30EnUaK25HQqDk1q0+5p9T95i
QwZ0uf8bsB3iyYJdyejSJarZ91FRBRXCupHUfR7Yp81bcBzUiZ1egpVGwlkLjmSn
WuXXvnXA0LB9GTM8k0Jhv6Tet3DzCFAnjiCu232BhZxa0nQYtppbGozn5Jx58Pk3
mb2u7trvZHd66Kv6vCWCA0EiFsc9JCwjGZQERm8vsMjRX9S+pg5xLOKGOh/ns9B+
VskziJnbnd7+W08UF+Bn69Nz4wp11Lxfw7LZKzCIUBY+dEa/LZgXnlIL/XUoN2Vm
O/0sS2PHsEUO4hH97RgflsZ64qhGEeffBwlVJ1pynFImLjZ++o+ogsGbV2Geo0nr
KAFGRmvLemo0O0+LpGBSxGf5jTBuPsSjMdUXlOXwX/If89sWdPve46trED5Ixqed
hppJmotOxReVQ0i29f1z4baMeZHmjQdMV/EW3R7v93SvqbUfnnvAv0h+ekovpNS+
04AtF2N59jKJkue++M62zQRsGvk5npuAXs8tZ+sjwOp7UPjVv/Hvi4KSJRdU3Jj2
2uhq/0sDIyX933s29lXkCG6BBQ4i4TXB1BDQD4syEQ9HkNw7m8Ta1dplsw2vm1o0
TA200sYyyCc0TvpTXAd0HkNZVfUyPZZSdvHvqiPcyBYDZJmS9FxnXj4F3GRyz0YP
PUVzSI5IoX1NolF1qhFIW8ooYlgX9Uc+lzo7elNTRxYyc8GVuTNZ24+CF7rI2qVX
olP2n0zgla04N5RMKGhZ6vFKSH+5BBwv9ZIbNWQei0vygQGWPyMphj1c1uFpdhxt
DkZXm8EDDNN4UnQv26JN+pVxI45FiKHu8WnKsncFY84+qW76RarVbSMW9Z7+9/1X
vOA6QsSpFCduLN/BuTOzPVzau+ypRV34Slsy5NL8lYPkaF0KqBPB2fKqecsi+Xwa
4lplfgcvV5Q/xXXxtqxhZoWd5s6M0RJE2FNReNubVDIu5DS0yrqsdLy02UnOwZPA
VcFuysb5DGrGS8j2RhqU846Oc7absN+XkusRnH6XOQsCipEpaHgveI0KP23AjjaO
ykn6qHJ338EorLtNdqMT0ABFuAOXj6O96qHGJGAfR4+0Q69xJd0xpWlycMEubDHt
aY4z5OMtjow4097TJFsT1Ia6/ZXdMo8/htHYNF+g6z7B/E+oSe9S8OW44IsHgqfT
A6BDdOCgINTHufxAaJeqn2P9q1XKi4oRvsBFxAzflsccCFTU7qvdj198izw2Shu+
ktyoK0QtrD930kYuaBtdGzd2Q1ga+1dS8Fbjha9lSdd7qZGSU5mn7uoDizfUH+LS
6RbJ05exPeQbB5NSunQFE/JNBwzb+xLhCamyQBISqBfIFB4UlLwZJSTl0XxlXRJJ
O/OgiUsh4+ourcmAg3knCM8GJVSdsO1V3deqluw+zF6IUfBsxVDWrv05dbeU9HWi
hr62QzS4e0k01cqFRYGKZ3Y6U8yqMthiEumAkg0RN1Su0pK6miLehulXPWo8cpna
dK4XWTYRCgjJDjA7GFe7+2zB/htnRxivtwiK+DnfAzU6odfIbQ+JMsKfdoWHg3Gl
HEUAhGaJeY+MLESm94OGBJydKDZVkoCwWwVjQ6MPiZD2QWoF3OKrBCBY4FpV4JTc
1hrBxGKdjzKy6f8Sd3T7iD00CxzDlOI+MTBhe2bU3ZOeLxLRKwe78OL5d7dK0qRw
0ZUSSv35xVuU6BnTTKt+tqWmwEpu2kKklsA2pizm/JHWvL/G05BQPQcWLjtMwFsv
9g1P1+16qyHQsszx533GtvhveFLokaSHwJU+0V1RprkMHs2k4hJnHi90nwULv63x
yhX3ud/Ci1/McoztYft4PqbYQ0ORpaHGh50VpgpgGuFZkO3UKwfVaM3iOHmNHaxq
AybHz+wDXas0lhedGfVzByipMh+R13+qJFEA5BGlzuTA4w85k9FP2YGAvJ7IAE2X
6bGM4F3TBzs0jmjnA+gZbO3OCY9iyukZIrdj6yW9hMR1XUKIrwwrPjXE6p7Wn+OK
4Rp26+7PmZ9X79gVE5k0bmLu5qnb7ayohvrkBO2F5e7ihmqOLo9yHF4LzNWu9PVf
Rrn67qFF218b06PAR+0plJG1Qc/Vt1TKCwDiBFKuBPel8reuLJce6dqbaF5fAHAW
x2siZb8fiN7rxdMS/GLKRv5oW6SOw0htOuqnMy0X5dVq9F263M+JasOmeb8RcGkX
/PC/8DXR6Ou9o6RG4ZJi/yE0tHxpm9q3y4utMJDTOU+1peX2GnzlZrtduPe58GKw
GsYqXsVq8+t1/+WKNrkWQBkQB994ieCRH9MDH6TL2Jn8kwxTdJdM0V86jmKU/7/d
Huh2gNZv3XIERsc01nBO1Qo2MrOJ0MZuS1/RMLc1IyO7bTO7FPE8ew5s2HdT8ZV3
kIELN1XY08804324qlLTthM6WyVwvjL0gcOSKU4yvTDesDcQk11YOeQH6pV3NTfY
U87oCf9eVo7dWb2AgcUaeyQmM7/QaWeZYCHmlAqy1lfm1Tw0xY19t6Pklx6SOKbt
S+1HFCtEskz/+xn9oV3fAw4m7/zwylF4OtMBksgfglNq2UqvjY+9WottNMVCSuA8
UqjDN8KtGK1eveZHV8mMmDKrfOAhkaWbqpgHgyAP5dpa3I4GBMOv7UUjjTTpW5Ys
xgUVWVsZpXLTaiy90IFdO9x4s1BKi3uTKczV3CAWbiicX+nB2GWR4YWJDtB+y9hl
gnqJRWMHmMNxkMFDSDAjQIWxlb6BmhiBMcadFt4b6VesberSOeLqWevGcn1NGYMW
wyU30GVS8q7DXW0VqVxHp7HhpRBKapg3LvFEhY1+tYg2Tlhlo+LrNesaP9XMgGS+
96/2dEAEAJVxVVDNGZFmxFH3BMu5OPe49msRanXS45Q9CUeLFuKc8k0Cv7HY5BYY
bhDdR46HZeefwkxm0WD4RC/6QHVp0hnPi70lpxkPHMHSdHF9ozmT3H9YVjEu1Jiw
i/DBBRjQi1YuooYCgcPhT+j7iBSFMTfIxo/6Jmz/IS/gNcMOyUE1smPQ+9Y+PXfF
gvImcpAm2oEXhV/5qP0kN/hggnghoX0c/JKd8/fPYx3MTUq1DNeXdjnZ6JZ7OhyF
RpvDz0DBL9mEDxwX/SY691erZH4ayCMviq7mquCyWDQpjlfxG1I5OCzjyvev9KFm
e1QKvA7WrWsAiK1ki3L/+XNpm3LWHUN5KRTayl2ZsjJAlD1Y21Zf0bp9rPLohfku
PALAzDjvg9ahyj1YiU1wsyIl97F+hdIOfwcSdKw3tl7aMhWkRxU5PXYcTuS+J0Vf
N3jCMAVzLtD0ZKfD3MIfw2quqXuWBudUU28OBvwWgFyjnUJERHpvvKH0HAcSpoPS
drvuoZ9Hf6WXNA6PayijTvsQFK6wOaaPz1GBw1NovqxE8aBlbylIb3FvrGDox5z6
x0u44L/CBSK4acCX9pY4xVIuZO//3hN1w/6VNj1XhmB58mAprTdfm32Qd4bIucHb
Gs5/hs7GLM3u6cYsibBepentxMKE1T3/Pyp9JvK2pFg+oyhuwveQMvbUh0t5bLEz
Daa9QSFtCWd4LXY8N0maU6MRkn+2gN692o1SzCrX0MevrLnZHXYT+V4jYgdwDMZg
KCZ+IaFNv026qKt7qonCvCBMRy+rGPIp6E4RqP0kRlN7IxJMyWj7x4AtwcUwQ8pY
0xpydw0zU5ZA8F2kD23Ph/USG39PV+jrgRfv5OB4r9dMuTWXI+Z892l1q35J9Qdx
dBEuWvQ8k1tb8kvhnK8zrB3FKsPwOG20zvTky1SW5WBTthwpLlZ/qf0KG8VAPsPw
gUdfkmNbgX1VxV0ql2tYBPzg/hBlE16fpFJrduvx+sEsGuy8/AEKruBY03t4YXwz
afy0iVTNnvJRtdOMfAagBLZam8Y+e67Aeu6acVgZ8uaEk0S24NXshCpcxAlf8gM7
w6qkJIq8HK8z4jtJvgGHiHrDZy/sr+TmYq/S37JJZZMATOMgXmBIjUGFi/NlApmy
tRtWiyz1EGmqkluXF0u55pM1KqBMRI7/FUeqDeFKy8mrGhBvM74IcMqHdHHUfE9E
215AS/0sZ4jqjhRQ9wnnlGveJZVy1xGy8ESaWwVAoNEzwi/KtCFWG5T7Y9f9Mmhg
j8va+b3ZjFEdSzJDCZ4IQoPb5k78bPhYkVeIx35i0BLSVJ2UAnevoYzsDy3jZQ4s
kn4BZtn9+wqQe4pDUjQhTiTEuC4wgWOlvDnlY6wIBGaXXEyl+HOCq+3ipxXoLfnO
gKF0Dyr2zw6UexQ/g+/ddD9mLTgOlm5nYgFpFudD/KHyvWGrcIBFBODKcFQO7z7V
Izwk5qu3483RliQvWVZ9DgeFQFBn9yyVUtvq2j4CXSQs39Gs3c6aZnNtCgZcTZju
TL9hOEXryuez8fnPNB0QY+VSHTnJlYb/xikWemkv2YYcmVr0pqDprBNPjAG1Lche
K7YvGhijP4zUZTqnCygqEC7J3Rne6vkvZ/A/58dTlTuXNFbBPZvNwVQREUvCq6HB
dmFXI87MMhE1VVGPFA5kGKrBBWZbfc4lOKBf6hnvHcvmcFkOqTjoddgUX+kYvyaR
/dV3bdXp1tpM1QU7V5HPEqB5TDoG44i1Ywhg1R2G4KeN0ZgtQGDdpKQZznEr9/Tk
Xu3Vks60bqClIFsNeekoey3goBg2q4RXaRr58eCa2wE0i5I3w/46XLVtUw3Kwcnd
Pn47O3i9/lQNiVvDjxp7D2HXjcScRya7DdgkCaVEhtRHL4dTPgx7e6daUOJuHAcf
/uzsIzj11c+65BtzpUdLjPMeWC5ACRGPolOWz+mReSIdNBSTb9aq737+IqicseVt
3XLZd0iPy4MadnADZFp7dMQONu5folbp/43GLuzAT2SwMlMmtnDPTDmJA8cOW6/G
5t+qOxz0D6o7xr6VgUH92VK2wHC8xeGUH3D0Chcvy2fT4KM7L5bg6mQq3Bj8r+6n
nf/cNcCVYxnW3TyiTyskPfspXMMxMPkdXZPwhvpsdSf19YVJtQXjZS/PT1KJQdba
OsJ9u3/xwuu6rZsa5UCV5MIEKyRgIVK964fm/Vams5UZ2QNESFAjCDepopMHLfWR
0KZ5Tow3oIqxLqR33zoFQ586g1Bd93UdijmWnPLZkNEX2kTHSuwC/tDGshzmo+kV
G9inCjrmUdKQDuexOtYrnXlKEG+mLpLhYxBxUSNCOlcDf508OMeLFAvmYnPT9u22
hdCjpnzbyw4xvpUpRP9F6tZtkHBueXZWKr9gvtv/pFXmP07xY7QPXMFN7J6uhUlf
4Yb2iOeR12Z0+4X1gWoMntILoO/v0Qdj8Ev/9nKRzwZylwkhmof/AXbLciMtu5sM
7lfSrIFSszcupeJJlJKeV/irun/BErwbF1/CHxQ3dI9owYPJBIHP/hLqZ7t6YkRb
1wJmY0Jf8IAbQMbMt3eRoFJ9p6MpVXRNDGqPoStgiL4jmP1GZngS5b4qmQEWDzzl
iTaXTmCP9hwP7+MpnsB/+k/tHqsQAWVY9YLw3Nndja+Tg/eKscfPr85Oc3tPSmDr
ltninRz6qhIQx/m2rp0genTk5+WssCdNfw6mWxBzZt276f1mj4w9SXQNTEZhLVp8
igICiRNIw99wORjfmmb/Dp2jFN81WPA9s8yIlUEdszBGnc8RnDdt7r/qtxb86Xyd
L249KpZ8s31wgZpi7pqf+3xwVUsM8LI8ezQVETRZjWN4WTMsI4DHuUGjk3mTcQMx
PahbY+5dxmsKupKxpqkD4h9YGcLUh4wvoWl75k4tI4oMW6Nv3fmMOIrjZppNzwmL
aqBOtcSVIE2s9LnePEjvbX7w8IutbNUmSMpzAVNQ1bOqVxbs1eaPyNRWzi2v5PwR
G3LuMFThiH/dHlWCk+UTRix+nDfM6M0pap2m1Mml2RFz9ggGj14nyGxuljTrQU1q
rwufyLvsoKD8lIx7sokl3AOnHnX6jb7/zV3pH1RMjrSR+T1YzvG22Glo5duDTBlT
2oMA5EhGHPi3YhaxuDi85LuQxGWFyWTPnOHkyBLbeMdsvAZjn2QUXdofgT7uQG6w
RwPKSs10WVmCoJprTdoAdSahKmu8xgnHVEpAddEkFDGciyWUUWmy7qjuyKRPN8+3
eMvKRlLa82mPbTr3gvBU5FmiVXnyj3eFna59mXfKH/yrL3wcyZSbzgg6zoE0Zf5N
1AouFF5+oJRnEHlO9JLVObFdJIy3qMBCtlSUBnMmFHd+wWATuI3xPYGDXJf5Bq6E
ZejbKmFaMTBtu22mCNLeja2qBrwRIkIiHL5npViAEkpZZRk8Qo2iieDh0hDWI5x8
FsKzI5H8wxdMzJCEWHGtj1zDUeITAA7GD1xwOubhSV8EtYdgcxx07x6Tn/ocTrcQ
IAeBg6R0hkIPhLj2t/v6Wnl1C+bE3JO5Z4By87uqqWV25Mg6Q6PC/c9VsB2PZhxF
2gL19EG/B0wGhq+p6GYF8WFYouK6GeQJo0d3Ki2NUkwQHSqhPbPsxiHmqjyWhL/o
xGZoXoe3Os9OWp5o8b5zhVPTrQ0sq25RTjSDH3Fy91EnV/eV7ij13t8r2VcDsKnH
LweFhUwBaz6ylR2IZdg7q9Yh4xyRlQHdtK0W9euim1zCEH5MUDMAjLx0eYBXXq2Y
0KvaN4K9MlL4NDYEkRniE1I6vOtCnVFUnf/EZbGJSr8YdA6sPsDs+8+CRIDle5fN
OHI7m2c1C3pSxmzZiJcSx7554VkUfmIR7knHlB2d8hAnrwRRaKDX2jlWDGKY1RU7
08U5DCpWqU7MrETq0ob2P78iQmALfj6l6014oDorNnkRVewJmauPsWXqAbLx0ZxD
xExHV/lju0ER2n0aPTpKOPup9wIXypoH4sE3KBeiP7lOr54x4lMw/cMnaN35C8Hw
pQ4Tc25one+xYEC/0Ur72j9FfNtzd2wyTiM1MtoXbAxV4wmO5RkF47I2M0akUtzc
cm0xuvoxugi/k/Ooj3ZSDk4ZLEdg0jJB2SD2wRYggMwaWt+iwBt2OeQiWKoHnpeW
Pyp4ib2mGX41elbXBoKbo/vmKlKI46OlkKB8JZ8ndmOY1cGI+KRCR+SaWhZ57oNP
Hz/BOk++I4rKIUAlD0enPlh1DtOknqYmR5sjxeEt0boe0BCW0qS5ADtgIk2LSiaO
shdMxdHOlYTImGNbiP34FrdyCX9wMxcSi+TSikjgXtQC5xSINBP2s4Vfix2I8orf
aCGiOAXa1XR+3o95cKBTOimXbL0GUofat7J+bptOomqfb65iCW642mvAkSS95FiZ
4+MP7k+RwtrvvaksxAjzjkz8n8bXiqhbhHplY8SzXw9aI83VwDGis9IWS6uSDG7d
yzuSWZpRh5hcCMoO/MEEHa/nIbdLd7uehqxOmNZI/akfJyNe71ihBf2Vc0Y21lVn
nR4rUuuQcdEEbL6DRmushnjjEM0A1+hnte/s5MzBorptLPJ6WBDAWyjVqsgjc7hs
eSvDgQstb4xCRe2Uwh3uwQvcq/xK2MunJLMhUnvuht2Ci+8mTaXr/F8kCgiFoeDQ
uWZ+0dC43emHIyr9thBprxsjzxgSgv3MNa5f4zw6rCw1bnZ5sWxpNytMNZpLh5uQ
Z+IyI5w4JBbTCitx68+sfCMW9M/ZnUTGcDuJDMsujnQBb6r/Uq36znbZHk9Vg7zX
xeWkbpfp14i4VTOck23DyHkL9GH9eo2c6DggjpGeEcy7TBTt7jc3VOi2tadO+xgV
d1lVSRi8nReZljW7NDem6JaZVSV62oVssI1t43ghMgIOLjcB3lV/3kBK/Cbkhw3P
hu93wxSDkCXnwCzRECpvG0zBsrnTJAs2MiC0l2+rWMBqp5wsUCoTI9y+pVJo9tXf
B71TNshl4AWGRDWx7CgLd61jRpVz9qSkDtf77pwH8vFMq8FqhhLK7u/zSLjxIDkv
8RU4sFN4OQW6GzCxTWf7IWrX5n7LLiDSYnFko649ape/CCR5aALkfZLTIai8c0aH
uW6xgcYHgcD8e2HnP5Yac+HpXx+QxFcm+FDpU+qLnpHGwuKxF7sfhv4YXxWPNQcv
RWYDap7FLxHng1pU7srLNIF8GM8Sdz1Akoll1WE105VJeUgF2Br5h+0/ojaVNAlm
9imi4GmrKSkpKtLRAiy0yGHP99TGXFWCTMCKyA3c/VV0W38u3KgBFZ75atweyWZC
T/YZvwTTCfPK/9jHiZnkfo5VoWtzAH6LWmK5NDJLNPnI2QyWgwNqvusQfgyyj7mh
Q1SOMOHKaq6uo/Z30qKDlFpftW2VjNnfuAq53Lm4desDlm7KUGwNmFpz9cr2sUsk
1hBmhi9clE4r4WZy7BMlJNGdgUjQSWRsLXoE/4KDrPcXclj4XnJ1U/VKw0t/UR1L
7rLBPxR9U0Mrr2c1yGfwROZXt3iy0anMayKQujoHM6IZZMRaKO6ZlI6W4VXadnDc
gEUyT6RGN9vi5FwTpWy393kuL5eXKwH30krkBuZKsKYxvNs8C5Gm/A1iD9U0YLlh
jqBJmJkOYguV5brkbYmFLGZZZ9nlyCpkqitk+yYmhnUab3GFrUM5coLcB7yQWxXB
PGkD9o0K5FJ7kdhfAQZHVDgnle7ClYA3WVIALc20ILVMU3bd04USDOY9zQAVKwdG
8tnoJnWRXh4V7qfripmYHTd3Ms+4hp8OTdaavvDFyYiEujbnSMHQiH/RVdySYcFL
xj+JXw34jv6VzdhoxaRSBl3I3bpbIJhHexYaZAwnMrtyt6zUPRnthksuoCo1cDUM
wx2zveukipG7ClDLrNIsBixfZlDksm7gxISKfwr7PtiCyL5WrZKwpe96FTV0EMbL
x2+HgvubSGgf1ItpBLysQzXpPSGUCL3dwEVor0mesnaFVPXw/YNw98oJql213OS2
TkUz5qzmk4Uzrlb3V9yY8p2C1Cfxt//MgnzPT2Gkrvbv8gH5OKUr1DMESwulup85
uAZ+IWKnCXG1yaF+X396hYpUrgREwvEMcnLh0axHJLl7fNCKVuHtJyKKQUOwQgx2
LpZ1qgBMlXRVMi1E86sOXqwotcsvh4LuNzfVf7+z4cCKJrKql8Nj1dJK0nzTp7aA
hen9Jj4JhFkxP4deXHGOoQ9Qup5jVJ5I2t5Mh2dhlQvpR6HIJB3j99Ww5ZMMIzUP
ShLpYOLZm1H1E0CZIoauqQQWpCxm15vb7VgqP/IgDTb78wpK/I1qFARdVb3YR3db
KwJeyPAZIUfrXDNpzyqe/cONBVk0RuVrI3fdVK5kTXHjgnG+bXRgeBsMp6dEs14e
E/QfoHD00Kdvqd3JcficXifRMOQkVSOuPq8+RB9H/4rTbyXBQ9WmLEr9zR9oRPvj
eYekC+MCgvUeqLORG3GG7YmZTy8JOeEy6noFoyA/JWG9BST1ia8qD15ubdVNBMLY
k/xava3t0fFPcKFWBIs07p8Uj2QXbHvgLiuq0tachOHgse8HCCAILajAHRdHdQmm
JACOyi31lFJTsTj+QEPzsR8f/8vzg8V6sMQRHvJWDPTrz3XdK+29kkrIHEycLl7N
Mo4XOL6IkUyVdIWfTvAlZ+fD5PrQSFxa3TNVWJo0hZ/6FDO8Z2vUEnZNSaskTiNk
Wt/8e1EkijmB7JTodwlsBUJ7Z0RT9jNuIN4CFzOiUAj9Ki6VqGrbl0/mt8gXpBjm
uUbP0GC400Ig9ap9xJfrSbnWx7UeNE8u0JK6hhZJMb4CRNOi+wOFZG5HyByNoKWI
oO6d12Wj1R9fLm8g6gD4FGh1ZkX9Pk7PzLVxr/AnHzngu28T13+szadGOa1lfypu
MXtFwO+mJWaL6iTZiF2PI3pDIV8mFw1J2sswV4rpzpAHDJqA5YOH/5IyMM7GaShL
eGT4a98f7yYiPx864bba6ARJFmu1xaf7CkclLamPJ12VhZUBjrdouUAHeq2yPuZn
EKUeUOuDKAHRHjzMTr/M206NLfvER+8NU5ANENBgCrMdCunDS6lrlrnHBsaYeD9g
bIci3RzhG7m12BQ817YcMz7qm0Znfd5CZFrSf/fiO4TVJimD78mBlLUttKAWLJu3
LDiClHxFAm0CPMrzWInlC0qJ+guavz1aZPKc90Z40dtCzeewT1BWEpSFgBy/criI
xiymkcX+7l+sMcpGuPAgPQ9g6jSbYO0UvystWwuqEQKVBJrtWpOcpPAgE/LrL1Il
tvVRvd04c8K19EYPIZXX7mbCWWD4RF/9ofHghFAWhTdiaKyuwm8zPEuiZmvytUof
6PYr8BMR1rAGwmhmw07QabCBOqVrwCMiJXbWPmxq0kmV+R7LP5XUEM9Z9p0d3qrs
h1pAeMD3A9uuXJ6oaizA0KjyvNmoCY0uyCk/UPuXxJStOL66cGaLVkfZW604dJ45
rTZKb2Ik5bDubO6R87XQYA2xqdts7gtQq+jmyb/y7pAASwHA/eS0uLShV0WwMMrK
Hcvnyx7jXFQOKHcU3Iw2SH5d9dy5UV48yzsaJ961Fh6NFMWIRlcmvkJjM1+25Zkj
ipFBzu6r8cdGVCcmv9ipibE5E6DHxS20GBf3g1HrqtPCRy9vBcKChP8idoq/+8JZ
a5ta0vG5xK7M0+cxV6RR6aInaSkcAY5J7IXLxwgi6DiFCszAr9E4fVGlz9MvAkPW
zM5xkNuLaPJG25wHdKMAYhqWkY98c9x76fj0njLB1XbNVKSAB2HcwJeoQZlJYkap
8xIexknXuH5jYiGK/eQzP4za24t1THts46numu8jtsxPE4g13s/DVKfidu1wzRAz
WF0I44Qg2fneAEYYryEUoRlSs5O1oVCDGvhG+Kf5SX1Wr3S9pYNfLSffSe9M96NW
UavkgKrG0kFzEz4z+yau1qA7u9sXmEXvdVKvDkn5OctzYBsM4r9no2Q3HEjognLr
xG3ODbMCibM9UaEtYi23gZOapoe2FEtt43fdP2FYlw191k94vkOyf3jRj24uJTyr
Nc6rJaWuL8F2Q37klEFHl21JzaRQPK2QyI6ZH+61dQuc6EehnEZzu+boLCF3J1EO
LNRkA18a6raMdITiwhsKOynzMQkAQ9gPq6JwMRuqwhNGyspubv3Zv5AowBp0AXPU
vXcRaYdNG2x6zxkT3Hg7CQKQPmoljPm09IKCO2oRrsNsZXeajhVehx2G7IyONPDB
Nf9OuMjalb6qNWCVO4GO4lwq/Ljq0liMWArmeSZeQq2JvFSsTNliUn88Z0qNwneQ
GVlKe0EDB6EVHrcXonBqrIAhS9ulanmg/MoLH8w5ujKrnhCaFSmzqVzTMQwTMfhV
cKEZV9uHhRn9HEaC3jn3CRqFPk2kp27y2c3FJQfzR1Zew5I67By0QpvOGMxTZm8/
MYzuwlhjrhPFhxgErsCsBLPYi5kaWFsFcDlE0C8QEZFBFKat4J/q9mZzIeFBzGyF
Wyje4VHuZ+NcQ1FxS+NJFlhFiuPd4mqNV4R5Q/gs5kc7qjMTyGbAYBuig4TChnVD
1LxWurkVHvT2oWPkfOQrVJwIrSBkGbV8nF4IYleC+IkXd5CzSpxrYTzBC62msx5X
XCG4bWwv5F5UiFwIlENiBm8fhZeZbU73ZmAvgvA+knUI1IYwS1xKQ3p1/tuXgzQ0
MiINIJfBHdQ3fVg8dWzMtM3e4bif5zzaKw3/Eu3dGffUbu42UV1CS6Qoe3nmzRip
KSrDVsr+mQdZKDXwxNo5ue691yffi4V1YjedOKvVgIoyTBL+KU9RbqP7VZA8wENZ
P6l9GFuKeODH8u5nKaJT3QhTsX+CP36nJUBoXiBwdHLIRP8BSHFgidhbhlqSMvZH
Xji9qBez4+5/FFNymdKzgjMT05tzZzQMklkT/Mo+ZQt/5anwabeCRkuEiEjsQGYR
mvxRsVklFXVWR13I8qQe67NDL3wPO1E8nZmssD0sf9nZ18uT+OZqae24HZPiBefv
WxlRcTQQK2y3pyZu+laxl/34IV29J7QpLH5CmhPqkv6hjGWrGaNVNr1l82NE3vFE
+hJ/s/xlclczFSX2D7BKJCwVVdvs2BX3Ra2gROku6MxQkT/apzLEr3vGXCU2otD6
c+kSapxKDtqtV+7soQFrm4yyyQE4YsynYxB8Tpb6cOAwdih6hr0MbOT6jq3KY4+u
0tMaKMXvTghokxxoGWl6YxaCzbVBrYbE6ZX4K2LpHMULIvujn86ZSouF56Ag2tUk
Ni5rOOKTlK7rebp9kI/lgOk0TPEBJ5EJcGmFOigr04SAQ3CWDVzwl8BcUp7fIDA5
ZOsVb60w8ScoDvr+TKGpOGYfpsAIk11qJVDXrRmWMx2n6k1RZ0sF/u2j7JIDI9O/
r+0ituLekE6caQlVF5Wc90DTN7imwPNNTbxxLisDuie3nDFlpRmLmXYNsyM6tvpz
U9IKwyeCCILVdJC9mZzZaHO5ipsa9ckZORJfISY8Tc/O4RXcY3LYWRxYk5erw1+K
hgKyyyIM343k5SNZ21wBUfCyqX4aDbdoEYqln7oq5IZB9K9ntcMG4JLdFvFOn+zv
CFXWKiBxyd814CNmxEo18Wsgc9beVmZ2O4BMYkmKtpw67U7TnUXP6tUv4qtaJuq6
Ob8Q9w/OKevRxhzkTPhowYrzAwqp0CJwDHLB9hFy0TlxFF2qVY54c5rDVOAnvrNh
yDAq8dPbB3PBrAIr6L44Qx5GuQGlofavFpvQGQekpSnb35mpQ3U9V8EQGbUH35Xn
fJ2cSQ2YfNpYIUTK3Ds5NWzUp53MYBzarXBaLwIvNXAUq7jRK3SSY0805Az7p0UG
26boTXIRmavY/YRV62eOZpZVRwS4Bb4eX14SmeAe0p8pc+SDuzP8JQpY7FOaaXZo
ERqOc8Di7r/DNfyXPJFSEQyFbNMtiadFLMGIKDyEPacDsB7NLw+IiKiqNHmuxiyJ
U9VqZ1HTo6N21fGJ6Xa5ilRRXlksxVgi3QcZzxMIqxOfz+UDt5gpkD9WJZeDg4so
BGjQCAVEwhbhvCa0WWhgeXb+zTtsvtvjDg1Pm0osKkC2EY9O4Pse5no+hVLXrrYy
lJSk6pne5F/ugh4u97uf72rjC7ykonfzDh8QW5RnYaAxZsqLsDZGmwv7X+cPvNgX
dAY8G2rqg1A7QTbbpNeIByd8zgvrtTKoqrWXX1ExDdFWGex5n7H/l9IlImUPUbeD
pJdFX4UM7vqjMZ+uMHZPrjDvz2hRxDe7LLmrfVQs64rK5mq//O42jbB6eiVus9SY
yj6w+6yhJwImEBhM/Skm574X4OfLblLgD1y+4W7q7Jg93lTHNm292UIhEVj+DzM5
wMXK5YZsw1Z8L3cGskXydFzcqHA/+hPbzBh+5KvdU3RtDED4I5vhELtS1rkn3oN7
9AU6AFYe1L6+olO1+oWQJGK8DrQHY6A7Jvd9zei0s92TKR0WMnrAJTvuIaklBCVk
GcKWCtiwPvQErea5BqS2M/QNAvJgDRD2XdzIK/UHbVl7J6PXdR5ssgzIQtAzdH1M
vDIYsfScND1U7U2QR6PtPkRkxzegNvfi6kDg4YFiflDCHzfNYRDLnI25YRcRstiS
3zRyRfB+wroa5LmS/4qNy7bwvRvuQaIhmCMTor5aPFcZb81kSrI/Jr1doNrdkZYR
/4uueLpxm4Y5aKBi5IivonaZylZHR0PxOXbMo0P0hM405aJQjQVLDNWTbT2uwq9s
1lRwUrOzAQEkwJPuiMqBGTdsXSvFHJUZ2ikGaPXXwAXYzozhJmCbJdsummrY8/P/
AiNBNSOfepoPjtD57uuY4ucIb84toKNQ2fEuu+iiT05fc0fMev+9avT4KqawUQiI
GX8CadiC4evaznBh+FxE8NCJsA0e6PAhWorCeB81Og7igybG9hAOuQsBe6iSCl+D
1n81DtygDpPbMutPFeJrKT9f4bBv0kFcEWumAqvWGs+8wmETjx8w5gPUQAw72lI/
4j5P4JRJ5o3gT66Y6eyhjoMK/SIo5bvZ9K8zifl8N18KoPjdLuPDFPqDSKA6h7ti
1bb3+ThwVVGpvixtVMaRX8J2JmGGCeJstKnpzgkcVB2psSY0smAAcpqjg6T5267O
vTnGscWSh/VUtuuIhkLvONYrdDqqHIrhhqFsZMM55Nfyyhybe/w4QAbqDTH2fF0p
g344whGmOWAzEu++u9hTeLCFYb5FLYUZFrxoTSAS76ghFChQV38jT1TWxlQ9cYBL
VjHOOX+SW2I186RkfqbyzqrL6lHSpl792MOxpe97RI0QWX1Nz+C77sCSZgAnoulG
eIXBcyjrjCcEGIJNhMf85Km86HML1a40+6NyPcMofv/3pgxgHeOueYZjPSrMgssw
JYBqAvmwfKKMbLMGWSIRnsT+8EOToRmDG5kNCjI0EdaQH70PLhIty53jwdAPBWuk
VMYX+UMnVRhp/+qNbvxtYW+xJ0v5DO1uKDXUbVzPb8U3jd8UtAiL7lSoP9pXqHxh
OC+6lIlWFmRUZrKFxREVYjsaqO0iFdsJJ2ljQytWAuknZ4VsI4Hk0a/wlReVDxn9
LlUIUFUsjK/7aVGe1EPgoorAdViSlyxzCRI59GLvFiorDsaJO8zk6fW5oa4O/lV+
NxM7O4Zhj8rtp88IAI7IKhMzE41ABkzSUzfh3tUSJ3MTGudsiygGRWi4prhlTPyo
Cp9TveMULlNiMCu4OtWnh2IdGV4lJMwVWlkEWpl1Ignoh6GU+z7B9+d+r2W+Ipyk
7E0Va3GfS539EUWivETaDpGMYwTnaQ/skwvAM2uQUPhjPgNP8lYEmFg4nLuC9sM5
ORrfD9n3IRLisqihTFy3sblB0VJoxdAR8dbqoPhrRN1F2C2IuY2eB0jX0tY33Q23
MYCj7CyyCJ/vO+Y1y4nUYv6hjYbKoZxYn4jOuUiIiCGYma/OjWENChB0MNCb3Nae
wFmLDPdZntMH1MAPBeBgVi+zHp60JW7j2j7kwRVaUz2mFTEWYO66eSw1zTrE+Hj5
uRJrosVE1zlSqg7R9dTNNiNAk4lroxg8SHcfk00yAJiuQPdHgyoWjKzv6g+IYZ/u
4e7Q87F10a4E0CbAN9fEwYVLvmqLHtOXuPsSJNQDdY7dRm7KIf/b8+tGkUmGadw7
29S6rRoUnbtnG3qMtdSYKSUYgc9zv8u++OpI/VxMaHjzdI4wsRJnWBvOq+p3m54f
d//tFVWbAiJoEFv9y4GDpE2hzRXMtPf9jpB4Mkfu2i6f14pzv+oP0ISPRXDHOG9H
4WjqhjCmo/Szxls38xfrQRvqfVAAjqU8Yzip3V2mz1BeONRKMB052WMB84FAU5Zj
ZHNzKq7xTGKRX8Lho9EChj95tmiv2zEfHap9DUErZ8sOQuPqaYC0a1xUdHpV5BGi
HFgY+L3gqCwRSOYmfm8rPaz59nR1j+Y3kQ/cQexHTAojfcRSepZGORNGMAH3G4fJ
2cYTNEYNyPu4LxUq3f80PwNW8X3h4TE2FiWYxjXY8b2NBDVPn77pLngj5hAcbq7u
beO7dG4dO3/0qaTT2fcpk114TgXY/2YYaH7bowcqIjc+o6Jj5ds13aFWRsKIIR5i
lHQgmKmNvurJWTygSdSvyoaGsTDtcVhjjuVj+GR0wNoOz+BcGWJhRp9C/xY7iRXG
dj0b4l5K8iVOX2NQHPGIjZPwwU+ggWzHtSlPh8xIGSU+bCGkIulUGP3tWyjRTLKB
fpK+RzwK2e7VhkbfC0wfIEhib4IIiRXZQz4mrkvGW2WT7+NTaqXgO2OyWRg0w/+Q
vHBICEA51hlvsLaQCLy21zIeB8E6ZBDNd2lQdQLwutlcZ/YjnfCgU+3amO2hN8Bp
vvBW0cyVuTSmRX7YUGxhnJ/QEOI0Xq0xYj6e8+NWKwZ5kXDHrNEqHkj2y4OA9GM/
bcsK7D4lxWtUXHFCAGlSDwWxIHZkOIoPTmMvNh1c+o2DYayXuXtDKVxjg2fi21ZS
jPKGw4KH8v+dpEaj1rKg6IsOUEBKpbkWF3Y1sybe7fGk/U1JPygCbnoUkuSJTkPq
gBFAM6xZLTrQUOQk59wGpw/nXmQw8kYmf3SIHHgi4zS+ArF2+esN3WDcnHrRy7sw
3CLl/inb/BSVDXkKsIYlBpWfefLVl+9VAbmfZbFczA/Ru67a6wL1m0Bj/dZeua0X
01E5oelUGVhanLD5p4grogKxmLF9d/ttmhjM/vph3xgJijE9wfIhACCf/Ez3bKI/
ha2ilGB95hfxjmvIE+tgpFm4pbm/sQcIOz9mUVp0y2OIpiCcnBDPsPBDlLEC1QX8
iSACLwRQIb2bwXU+a26TNawLNQ3yCGIpVP9/CcvTa/F40+9yXMMzJscyI+/nfUSP
DwkALhoHYHxlAX2B+0W4axZAx+hhfIPsm/XCKzAB2i0qMrIhmhAS6F9agd4U3YSp
rKTp9w3AoJdrJcdYYacwScJgjjy5Gua1PD+n5a05Mm70AYyu2y3GP1x6Ug/EB3j4
FpEfAOLcrafOmEDoIkUyWUsFM4ekncYLCjYy3pC8C2XocryLvla0RbOAK8a7aoc4
jcMKxrzBdcDFZkeYb1HZgJUPsPJTvmb4HDoOG9hs84qe/R+XVQlhhZuRkqdO7VZT
IiGrcqBZ6lFWhcjlPtiogm2UMvZJpKOIT+QsTmD6VlYY6k7HGmP46+0hpnQsr+k1
K2xhHB1wlwOB/A+GkZQehal/RRb3gc6iEh9yLvmoH2Y3lvDFb8YNDHGT1HR/1txS
Y4Hjjz74OKhD48/ViaG8h0NZB+NVaJHsayNKbb2ZEAhHoEOB4rZOrBVTIJ0KNvoP
xZE4yxhijz+eZQujQ7pjEiXCC4jZZxbL8jnR+OOQsNBbbUa87aZtPSVOTNv7QT5J
dDEMS4rrQ3a6WSY+g+AXiKxdkZbfBS0qjCPeNuyI5TOOcgd6uQMbQjLUEJkDS0nT
ew0/dUb54dgk7MKWNLOlOOO79CtVT21gzyGuxHDjoD3RboRdGqMsGRM0rEgRDF02
IL8ZNUvsHQPTMZRtmzAbdBG8TiVqEn4Bm3om0TYocE5ObgVYOxml5yCNt5dcyvQi
Rs4hpxardBVRFIm9DLgapO7qPKIg1nPT96k5qYzVQ1VGPIL1bwz1ByScDwOvlIyY
eNISygJ0ZBSjlWQcIaFAQcyibGhIvX9/bMDqmiaoZRgX7VG6zkTyF/ieGhG/Lml/
Ui916vyZaB/UsgA4dQ3hFDTeFSjO3cuPcIKeXRKTTzguTUOXMLihM8HPlqkgTDxA
jEYv0w4Ge3ui2gmwLx4SuP7bPgQkb2B2xc4g63QYYpzeHEJBQx/5qSihdEDVSgTM
B4chiH2hsR1aH6fYcfGWrnr2y5JjDWg/K05x0wKaLwDEEhBjH0hT+cczRZY/kFwk
y783yu6klwbBCGIIgjIlhQYgezRq4AdKff9ukhJh6bJio+QpKx9iY8P3qOTlxyuL
3sTSO2mFldNAIwFQsesAKNYmQiGlS4TAYP7BNqbOgmUbXs1vAO9AQ8AhSZ5A73vi
3sw/UaB0KuTGnFeBMSBNDf2bdeKCOLAJxCrkt/OjT59yhgJtkRFjtGoA0AE9A0c6
LztItDoxwfPXCBcMx0JFAqiHFiZ8W5tZPhzL0R4lesS7HkMrFIdkzKbbIYqCphTq
5tTnOxYIHvslEe24Xj2rjg9Mng+mGoSj9Lj4xsIK9xCmA0vu42jkLIHBGNLSgoGo
LLsoE1Wh8QwuxjJxGgcLSGhqpnGstAnr/T0ANkXqfxH/0m8L5x199ieF64o1PSdR
DLYnGMfaSCabuP3+ezQcotDYE147qoROJZGIi28vKOZffbpvOt59JYUTUNe1CAqK
uShQLQSH/2qJ/nbHSakyfoIhX32co4gcn8OTkNK06515VDa7WbunX3/fNff0Yppt
GvbBF2dJE07utF7ZnmGpxTE1hyAKX7u3qRaP/QmLqMvF2qrIq/nF4P8ODK23/HtU
r3kaGcXJItNXmCv/uFI0wzh62dXaZdzqI0YN4qH0Y+K5QprPeWnpFB/+lYlu9jG8
k+OE8Oi1nQNW1XsRlYivVR3BiVE5CN8X1CaXMWMdlt/xvL5kKhVG4XxPVbuuNuNt
rqc0qLLw1ZCHKv9+RPtouq13hqs+xGdFxopmMsiFRAxJmCWWSfEFTnnUuYb1JXy9
mcTUvE0YUr7TMFc2dujhsB96/aiptnS26FW91GHgpUfYHIlhycfrkjvXgUmxJLBx
bVi6IaR1fl3Uz9dk137F/xeOEfAo5vH0kSmfUc+X51NXhhChVHW0VpZkAC3vIYHo
Gt2WCZ2SFDGuV6LUSSgRrp0F1hxOA6H/8jTU76sHPBsY+gu7EPD0TPtUGodRtJ5+
0Qse509F810rroM8HRGbSRbSVGu0ke8kaXxLF2TV3Ilnxu3IDOwxQfPXcEwdibb1
bdZKYWym5CioR5wBZ4vHIwrt7K3A/GRW+1RdH4fxa/dKQPiTwfog7z1vneYkFaws
NoF90YjoG1b3njhrPRARD4ibsx261MNVJ3hvs9E/o0b61SDy6uUddTAARe22+JET
XtgtBfdfVUYujBWzC8V3DlrB0mUAUliShwdasH+6OFOlWmMM4tokPs7sq9GNBgzC
fMDVWKP4NAxPKmRuWByPwLS3Dpv7ubQIYT7hedyvOn3ADVrl9XyKF9UETPQ4LmPO
XpiZaOTC1O2jkc2ivm3ejphPlsX+I0UMazZHa6JRzJV37k+AI4paUcdUvw5tDFn9
IrA2036KGFrBB32YI4V1yihD18/XoivKQ3yUooLbw7N2W0NVfQC7v051QeO3MKoC
AW1q8ndukGUf3eOlIfc6Peg647LiV1FK0dlglPEE+vhpWgfm11Z9R7hy9iLp3Tf4
iqDbDCkuFNLXWHt+CQWpb3eTMoZj1bz3ocpbnyFuuSb8MVracJBb3owOJs8nyLIW
jemcefFdniCsnvjYzumOvt0FEDiQkViIUYk9wOMpRXuokIbF7VfLce9xrSb51gLR
+1GJ4WVIlmAv2I5ad/tpWJFiADYPjB3fcVgJdNk0EuSBQHvLTQPU8QpUsekHPOdM
NSaXrhl81QQv5JExd+bqBQDPGZcL6g+pDeS2jhhak7veShZtnqW8a7Qi37ogm1t0
957/UwxbhX5P/muTZiLyfAcrvdfLuWbh0wfw6METPINuFygYVgJGBJj1G4ZsWCc4
GCVTGaQCTIotdxdTaarzOY/LzI1rYfEBDsG4l5UJhQKFC3i6btHX0Qi08Z1RnZRV
kwf9XKKC6Tik+h0+d2QQC25i52Mwq9x+R6jSnoCYESAXOkRNPnRJE9Dn5Yg5GKqN
VoAiZWBnr7ILCPfIHaEHgOocwTdjyFKeFwZxeFCfOMj8H19ru1sSTjfcg2z0OHxj
mLfwS9jGF1Au103TsWJdXRzsbqSI+o5gWi6BUCorMokm68aMIKUfDJwU2mPTC4O6
pNFg4itPHrRI71I/zaeqlB4Ui2lj2p4/1N0DCN1CKos3mVisFWjtndnT19H/JD4b
dUJo7txznyM8v/RtBoGzp0IOEe0He8JwY47VZAIyprrB/scJijvzWUiOo+WFrFlA
YmezUYNHh+tUH1VopamcXuXuTBLhzySHGsIUIGvZpQyICs9yOtCp1vFt8VA5fk4/
MP6/zPhbn98nJViq6pFxHij0Dx6Gn7taW6egNKoz2QIZaEcU3l0bCVGh3pizRq4U
+1f072Csg/6URUCoIfIKFq97zF73+fYzF/UIlVEYQYtBODzkrbsD6XaXqa4tmT2K
JYNzn9IX4BvgQwXH8pYtohmD3MS1rbY4u+mxmgWosenJocexiWGPM9Ip6rpBelgz
NQXFd3zP8kQl5dPhMWJzZOVS68B8hNT8+GXJb7DIsi+YUXWbHk8UVgLam5NFkjVa
6exHA7vfJJVOGUvA2DFQpVoBHKrOhbudAXXTj3xa2r3oHx0YKQMzsGyYQ/jOw1iJ
YrDBMbid+9K6Xb1s7L6ajbcAET75LRDFPhXPwRFrQ2KY1WQoI9UM21327eMduyzN
IEyVBN3kaU8ZBzKwEBfozPMfJaOPzN+91yoYBnt9poUJbisYNk5uiY0mwJtr4Wh1
DBtPBimt1YRVvlIQUVls/uxqsyTc0KjMegTprCIYj7pdaDo4raznKZpiM49Xyx5M
fdwFBDr/pBqRhTJlXD4xaKQOEhIx2SZ8QAOGuXqol5Jt3D9KQRg8ddHo4tQUvOv9
QfOdcNvRqT0qGVQfNMUc/uAaFu8Yw6JR53yMa3sGxBDUR3NbuDQk3QAfcSTgbKLl
RjicJAxjLW6H+9/TN55MTGnfX+5GTxzXxvC5DqtDIsS3461AMSIwYimPWgoViFn/
n+8p89SrdQgVkLhJ9duPRPjlZ3kNDvLAFw5wf+ha3nAxzED7vGxFVMU05zGriaSm
D2xJcKlzEleW8HH7Ylh8YTy5HlClq4XLLA2JEVoz3jC83Zaf2TQfpbngH0Wffy+5
4ksFI0gKl4U/6JOvuJZQ7ouOn9F5adaPBqE4Ruw7kNdPDPkmFXV8U89jbjlocZuq
6i4B7eb6xGiWLFvEy3PyW2Mp0kIAudgXiMnvScCGABdUY2NwjckFN83epXPQ0e/g
cnA3pR/nlfEsBXF4Li8YhMVDNVaPR54aoNHvyf58G2SdCwYlaNT0xrJ8nXTCax+r
1JCzLIJTBdKm+7wr1Ya6uBr67QYb2mO4fWlmmAk2BQd6uNSaglWUbiJzb3Ginn+Y
KbopLuIrExGHmrIy6Ne9O3xXotD2Knc4WWgO8H9UOqkwTI3u/0itPv4dZf6Rnl4D
BkN39PNrSoAXi23MDAcMcwNF0MMwrT6d84fXmJYu6IvEdZ8Cw7+16/M5H3bK921h
5aqypocekYvnrpLbCrO2KGBcqTiZ7xx3TlgfxxbbGAAVKLPYvmqsbpcau0+wAaM0
5NTZOjxAhbKdxyzI0OvtSPQO06WY09809q4XinhBkPKQAyNzgw7h2oCreHhj+qHv
Lqzgdo4y4STPhSxO1OpwNP44bOqvKYCxryiR9Tvt5LqRyYQ9uSWkMCXe3+t1Hbjn
a3QwwK5bsHJCHUH8XdLxeC6rS9bD7a+++acvPaNOfFRbmP7FMsmI0AvvLJ896UYs
UgZqVqaazwMmSz0p9vUsa3tK6K9BcGsU87Vj1BdB1jse0X6CwUnjkNsfsPWiabNS
tCathFZu1PW4mYdky6JDVmQGg7f4yVSF0819LJ3KIblGCcJWM+69N1VpmxD3/adA
q5cCJrKADpt04okw/llv3peSM8ByDQKYu6OGA4FdJtk4md/xD9hOJA9pGTISw+N1
nZ6UyVB+IRxSo0XMCZkxL1DUNxygbrisYFvn0nAmmPRAbH8fgcuGPr5ISRBcb+x0
G2pz3awx/5mpSS0nXMYkDp7YI+uu0b/ZkARNMIxBBLFBLdOcvI2A8BCSKJguDEAB
sU69XCPjchXlM3CQiAkzAaglw/MfE8zie3rDTIRCiJM+qlModXPFd0ll1YIMH9jK
PeZ64cSS/e42tp+JIbE2FaCJ4LkQuauvd/BNRVqG9CHSfVZXfXT1K2BjAVGWjV1P
X0Jb6BQ6iUIe69SqlzNNYI27/Rbs+eWxyp1FT85zqAyyVyPLe3Pt1IqRMU1wsdHk
C8Gqonv/auVdmsxxLObAo+l9ZOLaMCiVrID/nInMBl/fTdIo95ZP2BiWIoX64kAK
qdnSxPMsy+NdGWereO6xmap31tE3g6zVjNYRq+Rw8aQ63r5cW12Zq9DbiVFRaz0f
ztcw8TquccsMJQ8hP9s8wl3l/nHkBXRq3UxsIipqZG/l6mnHa7lDoAHrzgii1f+i
qfyws5Zcxk5wos8ha2Axk8KeItC5YVDmF+9mXiuS0K9oM/mDGbjAvq4zXPwvpoX3
2PW+wCMjnHbhuRBm0k1KZFhGsyvqJoWlgXIWQemIEtyK8ka5X5AU344faR7tM6Tv
1WTeoxjGwSd2/YegRlgLJB/T81Xrz6jouY1ac8GFS1b4mXip329iVp/x60lJ01hX
bldVWIMNOq5PCNeZd4VFP5d3UD3Idqre6j8AkMjPw7Yqys62ahuf/lyp5Fr7U6Mg
oK+qOvwfNOc/laxo2x7+7JLsx2og/QwobUa05lcWeFZul4IBJ+zKCCjBxkJAh1jK
VXArcMefUb4AqL76/QpRgienrHbWnM6G5sw5mE4SF70uoMMErEEBO7fW6fFmk2oO
wqe5E9ZQAHNFMtJ7eXir7W83SUWwG/zcR6P3fO3lx0HWoZTTRIcB/UGYvkRnNXQU
F4O9rZhCdcTVMhzK3GRE1ukwqfKCYbbgreAqM0twOwRCppSyMob/USSuKmf3V9iI
bVgvDN9H96L4W7rFjCMr8XFPtSH0qDHxv/Pv4RGSXhCOqxjAQ85FTkP6NYdtkcKv
mMlsbLSmKYeL7lmf0ktApuT/+HfR/ivyQ4wXrkMVc2LfasmKLsZPtcSbbhjoNcfU
Q5zKMtDdjMjmeYwjy2mU4hieN9pEk9d+BfBcNt3sr5FG5PxoVQjkwjMm0N+Vs5FD
Z5tMdzZYvKJ+tgAfJuDzPx0QKYvW6Qk/qF7C/sQ+wm+F2IV2DRzTMVe1u8mCKvhQ
WIwDjEEBr9iknWC6PDnfxR8iU/lFNVcQ0yDCnMf//FJm6o2VjIvsJq9W6o3oTsHA
CuNV8CuD6O/k3YHnf9ppDhiRfRNOCMNoTKdn71w2fWxNee/3sfoAVV5xUhlyuGxf
jkkScfndTsRQl8dXy3GmG+n1helPYNHZNhFQ3k485Ax5mbNgOIV9Bq5b56jjZN6C
kco6m6qxjTglPToRNPVgB9AAegCGvRrTHclTilb8JhIOuIBJC5x7xWx1P0ha8zVu
gQ2kYkSsQITS9XkzEMuyN7Wq62hWso3TYk6rxrRDSh3lCMiWu7fsNkApUFIWEYVj
fhDDsnTD57XqTWadV1/DkIwPUBWlUbrhU0STTYldyPvISy+yaTuBTIyaZIO5VC2P
Eu8C8TFmdykTCbGeS/RtkuyYJAN390JW0YVr1d3EBnpqsbqqvjyaEOK7c0sqB94G
KfXJXQ3kS5lYn+lyylX5bUhOn1RnxZ3doQXi/jIeGOu5UoCxHcqWfcn/+YlLeTH+
pyDHJikC8lVvbWjtSf97RUVNCBuAhXpdVDElpV3eSH6xQevXGEy6lXuHtFcrMrnN
tTKEmYG5DNKRrTA1+ja3/d5nP/abi0SNLPV4dYvF7iCziONEHp2j6OHYBmw8nP64
PtS1nQvf9WZ6UsubJMqeOiS41O/VhOevf6XUsUX+w/oUBCvLgRuOy2cyyRjOpTyS
nggeIu6wAa45mszKBaGte2lUvY+jMieXnSCX79HjFAnJku4+zVLBae26+i1WHB84
mChj1fq2QtsI9v+PrIG/1G1uCtSv+pywVduAeyYfGYOE2mkJYcIlE7nNz1b+xNjp
b237lR2cc4tVHg8EtSyKHSpouMPB8i2ISHx2eMffliQ5X1GwnQF8zqRkhpeRuq1P
ZI5yKsyDrgOzm+l3+nOnoeP6NqpRnsaN6V1dw7IBe5TqeItItXUg5RH+JKNG8VtI
gk2iew9r5HlbeVv2YSWKTwbvtE22KN4pERu1QRGQ7T+Emh0pph5+4QmFQTSkAOPP
ILKo4COCJyJxv36KeJACSYTdqCGC7HeetPhROnkVrat0vp7/wNOBcO/ircBare/p
dxiV+3xX4EdskTA3rzzwglM2pXQe8A0VrqbJ5/nm0BdKDBay+ZNhKyPcNwZY+Xnu
EymIW//21T6wOLBDjWU3Ni+nrpe1LRQSFkUkjmATPpnmPdKaqEmkVw254jtUxd5G
60/VuKW9ZaWdBkeSJ1T9Fo5tBHElULLb3ooup+1yhGVzQaVUhkojX4KQBEjMbVQP
5gFZqcBSPMF1UnLXnA2V8cKY0Ux24rx3sqXXu8th+1V45rizS001sf4rZykmBd3o
n+uyKIa/IF+oqm2B9pxkT90n3evOkJ6MmaLbFxFNt+dHBtqbIIl8S7y2l2HNogcp
+kH9Ys6ekDkZ5mbd5JXcdy/4rztr4kgQGU0yDm69DH2F+oTgm5t2+m8jTZVbLr0G
0QoR4WojRcg7NeBeVQfUss6nGaWURWZgKZaUmt/6mbpHI+D53dA9aGSaO1ny991R
PMS4ptz1Ym9pV9+StL72wggLMFbEcaXQuzqa/Uyu7yxg1TpPyCZKqZ4pAn6IDWb7
Q7pEl+oKDDN7nEADgVyriCFHoTm+wV3vdLyrkCaIqM7WfmjfMh75j44mVlbSrr4i
aenaIsvkpKFLqQVf0lBnGkSKJgRgXxojfoWSc4nHsiB1FEsT2BzAz9X6nOBXJkVh
8/7HFq5B77ddVPeT3f3NPZM9HCpdK7062oi1DQ4yHv3pw7igYmiNo4f7IjExw+xw
w9Xb6XscO+oMrGiqaWkJG3S6byxQxDx/EMosln0fc5PhfK99IfaoEOAi/jN4+DJf
X1MKmIwTdzrBh83br952vbQSQOQ3HtMU0g04rZVucENz48vrnP0yvRPqVbnpArXx
niKS5mApDQGhNagebAF6q0RYRN0PRg4+oLsO+OWbn+WjdCFyen+xvAW+EIZyTK5F
M8kVnYIpvpc8IzFuLszuAt0GPOdrFvarHhfUm2H9uaY2ClvrZxmJccsRGWrNNp53
ow30JQgqQ7DAerXygezc38MCgMWPVZrXhZCm+CHiKn2xya/xbnyvedD+YBoAJ9NT
8NKDVMUo6AH8djXm7OxPh1oLjBPygVOmS1RKKxE54o8diegqNHmdld92IGv9UVQ6
sboLnOajFiB720KclTL3bhSWUyTxAlBzYUp8dY2zTqi2h1NSqTUvEoXTa2C50bmD
ssv1sigsvy+qPHLq8qlhSvCf2PuDrmt9FeJG00bO6mqaP80vlDocFuax548ZLD8v
J67yUp1zCeHNrff6+XZsalFY2mOaFdXqjj6tj9kg2K84FeJkVzJuzfWLU6u+R89X
Qd/Di9KV4nZUjNiEf8gSIj+noFuCaTqaM2DwhLKt3n/cc/tPu0xvO0CaHRz0X/UI
zGd+v6KXhrmca94ySU2YkVnmOemHg+v9A04H6TCqpNqt1O51+bnO1knC1J+TUL7A
+CuWnsoGZ+hAYT/xtP4/q72P9EUR3+GlRwzr6N82thVZRXrSS43JvocajoK/h5j2
BCoIBeKzIFMClSAytxg3ROE6EESng7MQWXloSKjpWoNwZ/jdVixUR8aW+xwlh0yq
NlHemifcaapxYRUPU0C0HeeZbSiW+Afg5qfMpnkOtV/avaVB01wpnVD2wme1CPgr
fQtBbrsasF5mUMTIbWhKtNdndrS3krVGuu8unyc4LybzaNDsmDVBu1K6lyVMBRHQ
pJ86wEJdKW9+WSCz/dUbYkFAkZpxxe3i0OuAxJ2d89zdksrQ89YnJZzaS800qud+
zVjEvExZjbOFO1D7L87pVPSxFAnzE7+1PdWA86hJJp59rwzvfa+ExPzSHaaG8uSn
OI1aifQ6vjQOqgoyWKqJO+nr2SPY0TVZ6JbEJ1G4HU51P6QRE4lp0DgfZ4uzXp1R
fA8NRmFZ/2zqTU/RmkHZfJXaiB8yxdFNz+qgDlmYwAw/7i/UWHtSQPL0sxovnEjl
AhJpmFuU0hV7VWe8eQK0QD4z1zHpQoZacwPCzvJumsCPqGpHlop9NvILB7pKHinq
od5dByvCN+2hMjFSn8aqWtiRKSsj6TSCAjF6jqZzIcO71laUSwP/iRl+597+ugUz
hZm6ccm6e2gDtw/3Y5e6vA5hfSgiU2cd7B7Y10UxYy73Tntzz7T+OmrKpYfVztXq
0i7cUvgHSc/NFBZqxJKhcCytkFqD2Sx9SLBBXjk3e1zjg7+QTzu7T6sViRYcqWuJ
tdrrqleynv4NtmPuHMHSsp+DQVdRITcnAdl7/chIYHVku6MS/fDhH+YNj4d4QVym
pGvMvrM7CbC020dV9aEgjbvMhQHwDCHuJlSkSejkOJ/LOtMuvACghFDXZUeu1x3Z
oYea8+jLq+c+mpceWPfWwYNxneybwdQwitrnq0C9+XapYtZ0b4qD8cdv47xnAesL
Tz1gUkTJfdoJxkj57atstYD717HEYhDzp3lv618RimIagHST5SjrC5J/OYNa3vIo
q+rwvTiyxRslND6la7pDtxYeHcSWYO2db53a+7RroT2QqH1isVDK3NYzV+rHmBkD
aBzI9FgW5utrQp4Uyp4LLYh1bqZTPkqHbyLSBrlQc4FoJU5/XaXgVo0X8T9GMxs9
x1u6S2T1aIW2oSjfHpamC876jbDvlCnW8Ty6kCjgnXwuWxa2DfvPep+SvDJ4u7qP
G/cLEqmQtLSmu4X1BhyBNb4wU7Z7ESVwKKuCCRgaEt9udvNodGXwg1T5T+StLeB2
tusIh4KFI+4w2sxZXTzJ8NnF1nOvJmzjTRUvugaNOuc+th1mE9cZSGI5iBfrne2F
wiAqBn+S4MfzjUO4HV8OkPDjrfGbnX7t80pmAIJlE4sS4lvt8OcWojz9hFAoQzgD
9Xj0jtKZ1uaAYZJAm/7oH0t47h759kpk7SKgp0tzF6yBH7D2TLZNyndhKI6UbxGV
1xHrPtdpJDfncTjfuLDzLzKYjOXNgqazIr7+/Gg/tTW0Nato102E8UHmeDoRsmtq
GdfbM95BwbXnaNGOn8FOwKx4BwEKJXDI+Befvsi9CwUFUV3ot3KAwaPIpxfIoCFR
15G6iCBZ3bNS2MdveHqFh2SuN9mDSWVvc5B+3uB3nttOTS1bWdSP2BGhf41VQsNF
whQKjtO0iBuh2m/VZiPmJjGTyTy5VSXE9WDGkUIXN4dsnqwLPgPoXVzJw3fJQAGS
QEfsstaMzC/hgCzpUfItZES8vgd81U64uZf6tVCO2y5G4iBmG1zLFLNnGCFawdSN
qCozRq8fB642UIgGln6REkN5OS1a6M0XP2LtiiegdTVflpAklVUF249HRsFXx1uJ
us6X+shVuBRpzGaXAgZ7+2/iKBdTS29Rnt84lj8P5JsBOPyZGy9izOPC+9PHi1/Y
nwiDbGUTKXA/XJSoS6idqZn8qtrDxalm0+V3oNpErUMEG4kXjo7p1OTcBrcR6rCn
rdWMPfodVJILVr34N95xsaqpHQ+UBAZlJzdqn36VfrSDDR9KIbxoa0xU8b7klC+4
gWOWQxytA0fy/cqS6GSFqnX1WUk2S5yesdoraxJepri/wj0sVc+yesDvT5APD/vZ
rN+9ZzEgggiNPPhA5RdtCIH6DDK9+rr+xsZiX/GlWWapi4bhvIOWqQZjJXuu1Qsx
vTgx2jsxkcsf6Z6k0psbS7ZD8aXjhSU8lgGQQmdSXW/5Uq4jtE9QDdVfioZ9hOJd
umJGFlrrCmER9xeSJjOJmcHQ0dgA4RNVuBEz3xwCwWxVwT3aBlNf60xgt+fQrsFy
neaCCiWN3xE/s7Et8Kl0NKeIXAyrI2nFFpyuYUlMP4rkVK5duUJ5HW3aEZs+YmDy
y7gVsilhaz9557Xj3RqErQIHidf2DkyaQyHCDkMYpM9hg2mxxN5fYBrdjNqmaHft
SWyODUA8RiCWBURVMAjv0Ry5JJGcOALaV1t/Ss1AavAmPGDqME51KeXB2IQSbUgM
6STQdvVqD4ccgnlV3J3YKy1PfSwo+am6M0mhALeOV+IVJ6VZ1dqqkPjTzkTtQL/n
XT+ppr0uRUUC8b41vS5rGRnOPNY3XJdCT+ROwGIZZShoSZJiXsmkvyTB7escbXlP
XfJk9+b6lRtYcjW+bXbD8RoWzOUoQ2aiWwKGSV4LRXWjDRFm/IOrgkCPGzbA38Ze
3CghoiBr5g+u1dYsGqit7wDe9/QtGfI+ZwcvSSKj6O5iJcDvQInPiP8Wdgqez9DK
m9IpU22O1htGm3FHObZVJyoqqxdQvXfIRZWEKOyD/qjaDSicJ+5qJVdHkh987Chu
YCsONRQ8k7GVzCJoZHMhh84wE8yquWrcrtxkSMaouUhtlK/r7/uGzwLcrSy8nkO8
quP3VFzMRIlujol3DySDRnVrDwpDjreO7NzYp0CIF43xobcvSRSRGlePMXedCUNz
5t7mBpAyoeBH+fHYVums/Ed3Z0+b61QDMWrvq8oAMZUxyYdrYo7Odl/7ECa378Z/
lRDkzUWT//vkQoIalV8hRubAyeLII0u9YvAVY1KMz0l/kyNC0P0njIUVN2XwC6hy
Z+pPwI+NS81Z+CDmUSR1ThvY+Y4g4EQOD6rXXfgMLFsvdNdpDqr2pMCCU8rZQ/HO
sY6HMvQhk3wYAuDr9nhREwLUl1B/aU1cWKj8U3A22y31suLXJSVOmgbybrlBY4AN
c4f2vqquPwTAEhUO5hyApygAVmbCb32Bi4+htaH6EJVzMFFmqP/k64TN1LHJE0Gz
YInjkPfAjzN0213cPcf6nkYScmB+RNVhQEq171HWPqV8YuHeoQOROxbTxxGvb8Gk
dDjThe3IdHHxEpwKQYjriQ4kQ/Tz9DEasG/V6YynwPo4dbnMCKAfYO+7qR3VNw2n
Jmfk0zrJL2QrHJdmr1RVTOEDcd7LmyIVuBaY7byXf4hvd/7mKkLj+y5sLg4UQ0D1
7mG2HHNHbo2Bl9vuJ/svAdpCkUnJdiLhnamoIwUAL/ph712OOL1F/4luYKInvsAA
CQ1UkPD6DS81PC4+G6iwXrwBWuSUzAQx51iHXh5rQmV6OJjhdno0jpJlourMIczg
uxRDCyhAFWmEzXVg8O5dPhSQ7IVSl8Fw7NHVa0cn45swwediEkrqGHP5wGcXcTSD
n2eu9LIh8WKApipkgzUqAr4HD/VtW2xOWh/3goQ86advVmT4anxatWQHpoKc/QI7
bVydzLK7gfevzD/Mscqxd8MBnp0Hvpciu79ZR0pCzLb5AszWAqJ1wDZhPhCGTLub
S8UgkOxrgOM8K22ujxe6D9PZPCj/Fc8yyevlf8AlkzyJs26gd1N39k8mAQLI3dOf
GzbErqtrND1591sle2VW2ktbM8BrIZ+XHypVvEMTRCFSeYJoRz/3xouvcdHG2GMn
tnJuRxXZz8Fp/Wl5CixfxKaT1dj7FRgZAIRMGemmQVDYz1qa/idUcarYWWgs6YH/
M9GEbH/xr6MHEb6rNF4zb3CQ9qEgy6Vy652EOvSwMHTP5Hxl17sDZ1fXk4l+fEWw
5ZkTWeJpHeMdOSq1s1aZ/l1L+8D7sKSNanv/dsfbYanTrO4agBZitL+1zakP3qlV
ZRIRGIb/v0hLwOPFAf/v5VxDK98DdigSrtwKEPXguGBLSMveXjWofYfxfuC21tqt
PLf8bziI6KaQDIiIwJQYCzCu5YJYYHDzvmkAID4vNHPJyXw5dmSKD5BCv9ONMoMG
4t/JMGz8KZnziBEq2vs41NLBjaDJ2uUat55nH7pgErzDYk3qe1jTqxGzyEPDuSrD
vBdNzc+MhIe5tAHxU5xAuz7uet5HLKAdnLkdv+7qAZruK4x+v2eaprH9tLwiDsJc
BZivhrVKZU+P6RWM6n6GkZM9LnpjkCTkjmvqE3esjI1y2z3EE1uuGUUAPbblia9Y
xqgUL2jRaYbPgIpiVSGbMTHs+BAphuaeViIzcitFU5DZVcC+7Y2xYOtyPLbuOCJt
Um1ew0XuNnliLVt4q6DUtCZfWP8VapfJsujAjqsflmesYsjjBwax3qB98ydXFXqM
OPS+QCdcSY//ZURYUMaNqUE/fgD7QNL4iZYcwzcxwPCDkncmXlGswJcnJoqwFT5L
0oLn1QyiyrCBvhreYaIdFjBy7z1U2BCT6iHCgI9hpDIZeTTNM5PhIATDWO0UFgfq
u18wRllokBHTUBjlocKLw7FNYiYj9sI9qiND3vMXtdCwVkurQCYe+aNAEfIj+XEc
U1cpVxqqZ/GwLwH2zs4Vx+eNh5p1EN3XT/z5ZY0pzyfS50StvxPI8I6Wy0ml1UgX
BGNfYZc37aclSqa952u2XDpmkOl8S0a5wAhl+eJYziZv+MgbByXbaIiBubyQhz3a
byrFGs+7roL8+FvjAFN5TRaLRP2NW/dZSQ4EGnu8rylGG9uXyaC59GBDs+toxgQ4
Maigi2gBuCJyEUaCEvMckWQE96498jPENo+Btb1Z6xuDFYBc+Br13kmiU45wXFgB
2qHdLpbME5/RHbKLn+zrb+xTQ30zpsdQJUtERc/pIdZbnnbjtmwnre14DzDD/7Vw
2M/ly3beAMsY8kTF6V906JTzH2wSmfDY1EFapQJ6p6CxGs1LRavmFbJu/GOJSAec
b+IA60/xeapYD4zMLvtR+omAreAuqCPHRUK98Myf9cy87xO4g18OtLr+lRHQPYSA
9ALXUKjC+JOHqPIggAiW3CRy0x8akZD9w5VmpTxTx5TV9e/6m0gG7UZ25HDLFDKf
usGSR4p2CxbN2ETgG65hI1ELm4vhzkRfATl1EaL8T7U2mZB9Vs3OxVF/g4k3Z8EQ
kZttY8n7olUkj3FtMmpFnxijN8QZIn03h/UEwpYdFhmziHJVx2tW+Gq42TRlwmDM
YkC1oXMTYc1z4BHex0O4LH7TncSTDT4NBepjxl3EPDNZ4DifRPaKv+e6QK59eujO
JjVxBacvnIUxyzCkhoLaaZ9FuciaK0zX3u1+d4FAYpj3V+gHEVWOR92OVHf+NuzB
sDsALRELuhK+0iVttya7YCnLhSpUX0JQFb/WjVyxeXMJZl63gDJT0DQ7FXX6nE6y
2eAQe96s5TiL1n0AHbpznLQHn/GHUax7UHAr2YOW7sgQH3nQhQo7fls+Vdf4XPVL
+FVcO80JvARdNKdjzoMAam+FtjoT+aJ3A748jjDPvWx822veVZQ2eOgozBCLYA2W
Er5SDSQV3Na+gkeNO6iSbhSPjTVWcUWzxjJ3uBvEkQZA0A3glaBhYtIZtLQJamn2
Rytmb3xjY+innBkOe6Pv8C9mE0u/Qkkkjmsot70lGVqaUHRnxz/8t/xflHC6nk5Z
pk+7FzwJ+UkhRUoPRP2g69PFgyMlEQegWmB4RBu0cGKR1SSdnD9WbRmpa425e38Q
1/CI9s5R2c+5xyZXoHiQ65DTcQ8Cci9ozij4etFa6R0YFZviNo7g3r5tUBkXra86
bqmKd/3FuBJlBnnWv3CsMTPohzX68uaZ6rK+/jpGXa8DHmQgiW2MHgO90isCGYd/
033PuA/27NdlKBePMloDas/CWlsn1x2yF+oEkswH1zMhBRradfsIRsxO6Wa2pKke
KxuWQIQgznHwPLWfW3sHo0kT2hXUyt8EoIHuPb1hxHzYOVr3az04yt63mgr0uT4l
Wb78gWW9iKZKIZYFG2tvEGJjZDr9oPorcrCyanhWlR3mRO1JwzaFIy9e7nbwy7AE
9Ls5p3rM7Hh6ASuHCJBq9uJJWD6gePetkabfcKK1wfm8CA+t5SqFrwlCybZMgMCY
iaX2NCOc2vgvYS/53RvHlZXD0ZrJKu14upszo6+A/b+CLBUrEJwrMD1NUVkrxrP8
LC6PUQdkuREC6B6hd9ssCHuAXpdGjS3ZDPaA8NHGLrJs/wmbbtIBoHm+bL4JCJFq
zlO5nY5zu4mWQJU6w/hv8zISViDzpj5Y2ieiySl7TpDLvLwJVJnYH9Cby9dd0L1a
EpxialUFo/bErVQlpUkvMRS0GfFFIgpBwFOSvfHCFc6SihnL0WxwQA81hrBw6gWr
285kvUguqbJUEyXy06lKxFunAYN953xOB8SdyRJbOFU0pOQbvok3CPcXkwQo7slK
jgb1gU1kbspiQhCaNMTBvJ5Pc9a45uAe4kOpMBdnfHVXWE6HkwYR1WkMl3xO2jCn
d3qy0Ko5hgw9AkX04KyS1hLejoA+WXF/DXSCpX2roNcGI0JsSHUzmF84vIBX9gDM
3KY5P3ArqCfWcFvFUs/Rb3aSi3OMxfWjlfzQ9pVNemBsS9naIcRIGGVyCW3N3mwn
ximi2PEn2iJmk5vZK4vHoDlHRPMBj9ua3ZluuIY1q3mdjfyVx+OeWJm5NdabRED9
5DZlXKN+aKbiM/iOLE6KrGmECQLHOxnwDGlnJU7sM28SirorhPQREbWJxFpcho88
BIfaZjJeA48MdjCIrkdI68DWbWX69Y/g70/T+I71nf2wBa7kdUwGTRsDvRwpDYGI
hkiiqtCEuXhsGl4P2gKulACkyr7i04zm2+KjM+/HJf0qc4Rn9YjLHY5py3KbFdy1
0L1K71mJ3BSnq2QuHesgiXCLrhB6cRf6RkI6m7SdDtdIuXksYkGH7JElrViTMiQ1
2+T+fNLx8HLHQss4qrxR4rCjUEfCqAR6XqNujGq1JMax0PJma+s0AMyxMeauVCOs
gUdO183hShrcJW+HqUxdNfCp3BWedBimB620wtsWYGG0cb84lVI2w+nS0PkawU54
cwm49ShWgW0Vv/ZDN3PXaepBKiuKWPnRiByA/qkBw7bD/sSED4mXzktYWppl0Mm8
GiauKpwdgOurnxkGTuxtlTE9kSzrBsANN4ll1yZu0mVM1Ubf6/19vJgzS89wGoo2
W3Ig0p/UFfEUPJ9FP3xaREPV+erzxHkXLEDpTigKqqlDxm0mfC8LWqH8xgO/QgWJ
6nFU10Ab1yP4KO0pTwn0ttEDLt2oTN8GiAiig1TvliPpS+OvGsz+FGoIE1h280Pn
Z4e6mYAjtYKQrwWsCsG5mEMQScpkXKBQCpAnDjcJxae9whWBfva1arrVnq8ZhlXR
B32J6tqPSTlUdFv3+6+ncsghnXqaoECeDZGXuSAU/xbk7YlI0UH9BU/jodH7bOxg
c+eCw+vNxofIZL+EXISQ29oNo3wJdsWWDAbAVFkVJJlP2y9cRbiyi1Ar4yzFOLZi
b+ZkNAy8nsJ7zQpuxp7qXsVqsZ+mrWzmdnCyqFKxaex8yL1gRIz18LgulM9c6xY3
OahC0Ql/KLzWfO+vyyjxAg6AEL51XCCjg4Q/Jl1oRt5g95OYID0oaDcqNK0u378D
HHOTx7z9i8rs6ms5E59G8969YWs0h/2W1XbWB4b35jsZAlwbO/JHKbXPcTTitdzC
1B55RBbZnGIGSjbo0GhxSU/qLGsesEiuIt2WRG9OCcmJLyZKMRd2+WlIX1Ism7pB
cC+NyMXx5Uk3BzneJpcMFlwnJuiKSa1C/b0JMmNxdspi1rQ+Iflr8s+zHj8YEMQz
y0vUK6DQlXM8EYwm3Txz90+Ja8o5O/1h4b/8Ksetg+bUbMLfG23awjT0JTo0oe0A
D24S493sU3q+Wss/rzh9XwxpXa4kCNPXq7Lub7/zlcWU7IkV4/ywR71/qX86L7pY
3Y8iHAuSNZZi204j/iG88MBHoIBf6sySlbrv/RpfU8TT9HtpxPssOFC0FcI4y1Qk
XD7R0fKE86hU7So1cySML+I4AxggsImciXYk3tBtKwJg/1OhuLUJtTdd/jdyY2Qb
JfTQwgArez6JfXb5Fy/fXSA9byHPZOwkjmQr0fIhNsaTg4VZa2l+0C8/wI3EkmbM
1k1JCUEseFg5S/LR+REEcDoSyzB7UFZEQx3mhwX0k3YY09K1XdObm6PhCC6YtJmc
ef9DGuOfWRMCRmkewqJApu6a8OsLl2Q0HShXxciUEHlvOdySMnPRoZbFykl2q1A9
ej4GbDVMKk20D0BsNcdqpzDeuWcNNxWAN3GwWo95cu0wavOxxrZJaA1E+o7rcLgh
IzyC0cnClGWY4449nkZSeRMoFfgTbWvgmXildFKHMFYOfe6HRnTTge7VjkHvrDlR
OfXX3PSBk185FiJnJzGKW6Cbj+BbnhjxxMJvltGQWk5/JsVIZg/PxP2doOKkD9nB
F6Q+d13s9pFqNxigGe6eoIjkuy3AeI2Iz+I1zdnURrWSvBe+lGS9zXzqmG4ZjYEM
PNlmnpxUmhbQJYIRgZQc4Jymkx8KVB7PZNciSVV0l+6jOXdgh6N/0NIbd14IAygJ
ldOHVvURd0OHUymJ9t54mariG1lbxLrn5OedLWHUAHLDMf/K4ThqIxhXsG9xWIRh
2Z9Lm4IueE98/iOPZnF0LWRrPJv4O1aKjJ6BJmljkk8Y4CNkxMcDJhiz1N7k49EW
ekKhpZvSld7XvPgpXrKL7GU3mp0qwzz9kMDHh+ZrY02mq2BZ5GdmAMZRSuYRBsOd
qlQ6rnaHzelZ5M4vGLw65WhO8XOLYuTXGVvwwTHyQmrssI2rGTUjyl9ROHMVWP5M
YtGs6bmXLOMbZ3e9ZYzwcVw8KU6pIDNTv6bL8hRIxHE2ZrvQ/5/eUdZscV8eKw4T
egTFB87HuSCkArlKJsp+Irf4zuykRFgrgw+4nFd3iPWC5rCWEt25p4Uoj9JMNfz3
lz0gLU7FAB9gFLks25wS8Mnk5af++DNnALiz3uhiPC/IiNIyzNpIR0IuUVt9+BtK
CZ2vgeKas5aSomuIzboHTbu5194wAyM2KHfzCumPCPep7NmWVIva/kzL+tjTINGs
sR0cfqmpVX+4qaaIbSyK8ih7ufkW9LkfzLOGKnx2qQm4INi8hkHohGVFd9LYOCdu
eE0rO8mpc2LJih3ISJd4dXazFqBF6Ih5I/jP/C8B3GKrUOmfGy3lZjs+/AsE9d3I
rtBZUxYCuAThEsyUDPY6P50GLeETKpz4EgoVJiLtrP9S/ToLege6rWjYTmxFb3Kq
1hBcWn/WM/RTjKRQwcegFZR6v8gl2bB2Fz5IRU1k5OCPyk9q0QSTjQzHoO8hfy/O
Ut0PUsSwixXbeKByQ3qUXDOecNuL9NSzLZwtosBCGBXtnECQGKyuKJP23X59uW1u
b4O6sqK7YtWVp+Usq8fImZxDKzymOBbuhury41/mR7/RX99Qm0JZpnXw18+xt+Cp
SCBWJZ/sXsdaVcFBxx+IOv+x7wEhUOdUJul2Jmd9MlJsa7zYrys2etKiuwOKj/MX
LKOlC1XGeJ0LIOZjtD3F4PSj5ATrFXHG9IwvHoyiW5OXosp58O4mvU7EaE0VMjLj
d4yBtdd+i9FZpr3yN2w4PtOBtSUK6tWGMaz5lCo7jKfoxf6I07W0ytE53mjOn0pF
HaWWkktxdiKuNizc2OLDo7QatOpQq9xBFx6Zgm4LYtX7ov7yR9FyMKFUz8xwqmH8
qA1ilHSocE1GHK/BNxSdyUnJNyv7UOkDrkcvYL5e8t5pgY3ubYXc4FYqEW83Gu6K
1/vKPmqEy69ztV/QRywWrWwevxiKAN2MEjVXgODnaJ4bS/8nlgtRr7Pq5RtRl9b2
knsob/5uTEsdAGz6OZrZ/z6HbtpC7fIWA57iFc37TqG+sncTUibB2qjm4E7Z3pjn
581daYG1E20gdl0Rr9JkogTS78wJQ5zp1mpOKHIBiwyjm967CTS3GX7eGOdcD/ct
QTu1+bj3a5qP8PtR5UwDp614wjYMtVf8tWuoPfBvtCeF7yxeGGld6nZQs/edPlva
hYRe7t/d076lMo/v71nVpNUKIb3FoB70YTwo12tfrxCSjVHXY/DFAyOrOXdDNS6t
ZV/kNHOwnGRVOeDvTNx1d8hchGt/F5FaaqwUVd5S+hrzNU7lTBK2T8XY/81x9QZ+
5ddOiFITFbhhoR40xG3e2gUT63vNaTOTuI3MvdHqjkiHLl4IWtyai/2udSEEptyH
+tvMePOeX+uO2j/149RqHM5l9P4YAJIZ3Q8QU4z+HEwEuqIlLJvZ584zyxSK5ET+
zMzO9oXZ3P0ohGD6k9l3CVjlq7+qLiQQxj1W9Z++SRvhkg2Cf6fslZUr6thiP7Fl
ECmMPOsCCB9pvCkvzZ/LKNqNR6qibGyuKiKHQ7MOki3jlBcSlxK4v7BtEgzqewS6
iI1RBGoW3YvookfsSyuCkP/gPXMrbgzdbfar8jJB8z/AhxcS0Ri6YkOsi8gFvCIr
+pDXHOPZATO7XbMLlaF81QricwVv+W2TL3kHDHdEU8Jl90cBAwBVEto4mTozQkE/
mC2NWklDQNADdRHvwKxedEQU3hEFINRlAYNmYU4HxdzjwRIeY+xBNks4c2I4cljM
f/Km/KOBeIzQyfVEEPp9795UKdMvWsgCZyhD12QvS99Kd/WCsuc5iL4Wu6CxdzLD
oaEKqH0dUlUGs1BvHyrLVwIoIvXnl4HrkM4Yz5tDsX5W4BSoLu4ZLNAroIqtoDRS
DXD/iepzC8OjdkUgfl1tri6x1oZEKt3gXSsK1s6tMNg4W96LpVWgPnZL4HOFMakm
vPWweND6SkgrHwdEZBgEDX3f3lm0ulU4YgxY0Uj7xOYBJr9ibzpVoIRoudbNCK8N
VhFqZ7UtXTqfBy8eaw3h7utBajSD5dmsHvPVYNNYKYrPRF75Oe1eODecMbV4/oQX
CiR1n98Sg0719JvlzyRXl4IC94AtCWpCkyaR8nUdKpsKhKIy2NpZTVNCJBR+sqvk
AZRETd02mPWOMqJvz8q6ydWFJ284RpsE7s22dBPUAv6kTg2AEUB1zb00IX5tf8ZE
7ciklY0zERlqgB/7J+NV8W2gHL/Y1X1roRci6EcEQQdTMZo2Xq412/3L3vzXra6b
OLB/+Lqopx5XkDiYXD1yrQ+BLiX/GzZSpLcWquzfisCnjhQ77H0lwYIuXZFU5O5l
XFJSIbHo2hZHlUIa1P9gg09vrPbcWrVXyS3pMjj46ZOBO58WNkxH5WBCrPduvyeS
McAR4R3MpFODa41MxqzKF5pgxmj5xiJKuHHVxaJnGpjDN6Ii3ysEYyO/wohuIeGe
ZYPMSiiy5NSfWQ2Y8cMxIxUTQrCGxSd5fjCcx79nNEfhq3gz5bmtLaLQzyjAaWAF
KuRmf8vr1muMTiyNGXB6XbbNCzqxVuYNLzD8aaRfQ9I+pOWTg+nJpkY/djMS2jRr
k3+CwuuzYjfbSLcTRVthez4T1AkFoBS6nBZ7g7+rtpqWF/OK5dzwSP0VCwOezXlw
GXDogsgrxhGFxhH2/FgMM4oxACe6FjXEn8l0q+QEp7yGFtpp77ASXN0V+cmvGHWP
qLvvIxEaXKdoLAN/CmT4ubP+sO8RGLiFlfWnn7R6Pqfc6pebjmAa2m/d7fPrnGhs
wQfIG5v0QE5URBb07Sn2elhRSRbax9Bpx3rKqq4/9DvlJJeX52umzAVURyds+UtX
j53qoSIpnh88Z4EVyGUwT2KGmqpYy+XhlLD0Ql25eVRODUHsCHZ+rSiJADnbdAqI
TK+R+TwOtaD93RQUrk9cBhaYYqE24SD6TSucjq7MIEhmHhqjBzYU5SmVyyv/Yehx
J/dWLS+vOOVWPbi6cKskPufFHTCe+qvVYuIfTa5AoOsufOibHvqkz2ctgWeOk+qh
GfHoFE9EjamXtyCbfOSX5OeFBMHheExhR10MvtOTvpAh7Nkv9OwAn4rKzkTVCPRJ
BAtjVin7WYL3SmWmEE/2cUHtsLFYsr46+KwKt1g5Mdoujn/qMOfEX1+Hzefr6EqK
NIgDK+nMQmKGL702eEiSU4lisTpE7WP1fwwu7K+W4bdo44ywfSU2Lcl6RuqdmtTv
j0gMXivR6CKyU6QLx/91CBb6UvMn0ZZk0cSq+c/CLo0pSESfh7S1NVZ+JwrgAwN4
e/ObeilHYrO8urlmYQ1jsDDS5j3YkKwf8G+SJFBAT/QKDHJ7DPQ5M2phVS/RQr85
OF8rDWMbIa9ei6VGnRZfFmgtfPYrgBeeOEwg/XGphXHqvBbQUqF49kRAoqMGRw1e
hpObDeutYldXDJ+rE7i9EeowqTVxtfqiHoncBmyLu5hOOiJ1bxPJDlJAkZxp+LCu
44LtuG5m2fLnF0mNOO4/ZaX9MkKnUeRfXoSSGOHyDZQrgF0Jic04DPhe+2jVkZz9
ocVZpAL613WeTAbi6LtOGAAKouoOnfm9Cq5DGJmOVouGLHjuY7Lr1emTC9JE+5c9
ysEr0Zcojn+xPtmRVCv12ry9AbZndnyH1R2b0htBCDrk68QcbtUKUhBlRV1FH4rp
A91FRaSJXAfxueMzEhcVt9oKa8cuIALzxCJ6M1TOZvlOgzoePsdpUtSfEcQ+8g8O
qxgNRQ/DlBS+eKm4KuWQ4bJgQ+zgQ8jkB7Iv7F1HLKlI9Z+MoqS6IFYzSLW21Mn3
Pp6Y37O/JVGnt0sPysiKROWAME98Z1/phPHUeDbX5ErQb6qAC0TzPfTuDxJ9yr2C
PSgRQJBwq8kaEsbJlMX1H8hH4HeACLW1Y+Gxowq921/I3i1U8rv0SkFUd+kQ3mzl
+Ey+fJaxFfl54XPVX6KRhvfepe0yEGq/ji3OxNSVuVQ38Jbunk84fttKx1PtPokm
rpeMWV2lEGE4yNmpHaJWwpaAOpRIPXYx+2yJ0m9Q/EbizFKtjfhkxOor3AJ2loU3
Lq9vu6TpaxOfM/0gl0Do9csPzRk4oI8fXWUei5q71wZgAFqWgcUnFdTuaohV7XQc
x9DPnIX71AlxDXkpOdNezQVTBTfrNfG6jEzgcmEE4iL86h6pzEyGv3Va3Xbcd0yS
/XmdTqlfXBBZnERDZZ2ntBv9lEpZatkq4KjSvc5AJm6EcUtW63j9Et9AAlgtoWog
dVtcr6O55/ZryIoOkIvxgt1hX5STzV1y9suKl28Yi1EJC5iBCna1+n0cE+Uqt8kZ
WaJq6LSi/T5oEA9DuBu5nchKIpoxeQNJVicKrP0Mzme4c/SZcsvOk4MEqyXYnWJS
V327Sng59CXHkhsHrG4va2oX6UZIaziaicc70QRvTO+3xr0bqXazaXNoIEf263V1
LC5///EsYIgIDvs8bI0sH6D0SAie7r6o/SGtpeEmHCi4wS7KI4MCVzBwM61JwJjh
IPJaFldAz9RVc98TjaINgmrgWA2PQTtIbzv7AG+WT1UreU4hqK2cKRSoosZGfWBI
RVgrRSNcY0Z3L1EWssyg1BnVLiw7Uug6lZukApZ0zrY7yBn8i4iS1FD5A1Cp8nn/
kCJH+NC/Pn432Qro7YAQODnApxNI6DH3d7w5xS0Uq/NcmuKQFeAQYeTQS00T9LkL
FpknLjti+iLxqyGkSMMI50BU4G1pKIVXqTwaL6P2fUkdwrCae90iUd6Pvhq8PjDM
H7QuPNvq/s27nulht+pHQal0JPNpvfNeg8IQSnl+STjI1Du+UIwIDrU4sa3ujrG7
CRcbQbktf6rXFgMQ5MwIzRvGRiDPJNNrMIYGcb0yfiXQU8A5jgu8YaCNj3MTE25z
mXEcUlwEeHVoEuQrrWOop6u0iR/8SgWVzCtDqvlAYD3Y/Llui+p9H3C5NgrF/cU9
sXhGFABGOWwd7SD11YCGdNllhwFcX4gRvYT1ciGmjxGbFTT2CoSGBPRttVq1B6YY
sJ6xt0ucMXMCQnP3xKmsSGmFEMdTAvwcV4nnIOpLfVmCW/T0P0O+4GSG/7huN37N
Ren+D4cFG8U9uLuSPeNeAoa09AosUhzfQ9bxH/lRAQ5Jg/ihyPwN9yH0QBCkl0yu
9c6/N3UTfPwtnW1M2vIHPFf4d796LFWTvUrxO3o0SPrNgYV3ZniCvS03mAamAAwo
lVILiYGD4QTZfTxjZjUBnNdjjI+l3s7oa4eiy6EWWTz7/ADVjEWuNqVkW5eDsCE5
sQUvhnopQ0AXV6ngUURQjplsuLIZjpJzojX+V/iAubRJzx5j2YThlGY9wJLEF8B6
pE9voISIGbAms2KBWunBDz//8qFew7AbWr1ZRQVnCPfnhyWmS7UWxgr6nFlQgmc6
cwspwPO106Hd37bkRinknCeOJvAQgsQXuw2wEVx+yvh7v0yIUCbZZh2fDrQ8Dhzc
wePYsELURidQRq89XT9RbGj53FfLlxhtBjhM2dgHF6zuoHCXN5ju2eZi2/pDcvxq
3MPZxa1k0Zk6sn3W8xpzDQ+6y/rmlalHvij37KFQh63xDgSMHk1DjMnKdbGibKgJ
DzuRlRgrTTr0EE7/EoFUtd15tguJ3BakRDYkoGu88Ij+6CzskyqrQy97pFIXMrYz
OpWUf8ONnRIPLX60RlGJIziyr0MOvYVA8KnlTidaG2QgdGsH1rrQLqIJxIdoHGcq
ZTJJGPubNwBXh5efwNHyGuUOzCz7J9/HaqM7/L7T4c7inOdzd42aTBNo/lQUSDpM
6cYgh+l4B3o+pvmNUfFkGf7D8GIaye8209X3Msrhp5rSOAFPLzgEYGR2BIJTXAmz
dg8VP0kckhLrEAttTSkfyUEsoxoZDKIqTEPHE7cDdlh0lKnSHClx838ZPaTV4ZHv
UfLwZcz8ckjGzyXeAcoBLEb3iizi9D6LUnIgxUSk4opx4ZuD7jD84ukJg/+07oPr
Sag1VTboG0MpoIfADZJAcYpX91IBMnKvelyxISlUKYPTHSUIz+viM63CIM8aP6Xn
f+l9vHn+mIM6OGUhTdtEh5LOhI98eZpGPD1dieYr0nZAt9lhY7jqe4Mg2lu+EdUA
n4/mxseUfaIPGmVacFE5yHKKmdbBXIjpbnpIzNSPnkkh2tQxKbS3A7D27LVUntSV
KLKTRfLz4qd3z/aXM8HNBE4Ey2lYOT1t+JF4b3d1mgLwklIefo8SHIrSGNfQRWAp
Odln1PbOyj4Oh83YQgUQp3Jf9Ugn/rhZGWPFuZ8K1jysKjyWlFsyk1vgzXrQ4sfl
tQgpUhql+YCqaExnokMM5Q3yvffdwWeM3G8GyIGFchD4U4UflqaRURSfmC2GwJal
KF2H7HjDnXfO2WS7e8OfGyG0YA2lL9viL4v3ItnDxxvLEdPUe9h9u3eFOP5J9ZwX
e4In9B73y55XTgtoLFnAG6G0qBExf5ntKTSh71/vZ7wyVcmVvRAEB+6FuJvQexGS
kj8Tc6fHJdb83KAkwcixWELRNC7h/AiHlmyZ7+5CmIdVS1GDIq/R6QSGGLsN0UMi
sk8jN4ktgEMSwmWNgyrdid2VcmRKV53WEGJmyzAVS4qL7hYL1HWjQ/yMAeSnwDUu
yYLnjJK9MhPoGp1uhcFAcyeCUooYs2voh/U6OBXSXUw1sIHrC27idMH3MRhp8GDJ
MsmQ5MUU1HWP8c32D3vMqGulguATD0qIkSYHsGXC1JXT7zbtP+TKru2PfDxhyf4b
HT7ymfAa9XEaYvFgZdOSx+ZIkj2CrOiHjrIwkZ9SfegEkgYKqREXMBBWC/F1Dt48
QHX7v2DHOyElXPqEBTMuSSkUv7X29uzh/+lYes7TNQD+OVPR7M0IdiGPjQfc6x6K
99aosxZu/KhC/nalXNIc9FsK9mGsJ/UicnkUnqT6dxIhWntdLpRuOSgUyqpY7/Wk
ZCIedhmQsraf7YHeUQ64I7zFdNDy4tk9eBtok/S8JLS9emSpq0kULcf4svBMw0UR
OetGjerXDfNxLqxX9VKHvVRdWOu21qZ7UUeuOdRvPd+FnHCqyXSZUuaFyZ6q9Pv/
os/+f7sbobA5m3eWC3oEU9tMGgm3thKqXeuzIBmmuW6Sn63PLMPB8ZNrhAvFRijq
kjvi/kebhmF3EZSeUJkUR1jF2RBL+2x55X0pruarxuV/lDZWvxniWJvaas64PMF2
ECLnavKKTIw76AJHKh4dKuShmhkMn6Y4hsw5oLH+ozlpOMZNk826UWokb5Tqpckv
0sM9R20xayCojpnhB3VlZgsWQ9iYSIQX+Y4ZEfdJxPdB6dfdcJuS7Yz/SzGpYdGu
7HCptM5bx9+QsEej5xlKE6XrEokBE5Nxcde9RnO9EZVx4x3xTDTtfJvW+z3uvH72
26n8ieBgj4LLAYRPaYmQ6NF3GW41NepzcunOr5DvYoyZ9OcED6UDoV6YlI3cMw4H
P7dyW6+t84mJtkDueYwekhwN1++2piT4FuuFki3W8GkzVdGsOHjTai6aLqKuMhDl
dU5UkK9L4Q9ksLNOWSs+Ev98Y+EzHI5R7EhvC7Nqa422YtobTtvBRR3SsCr8Yu5s
yemqgr9uttWkVkglW8afbwO6gL4WAH8tmnuXa/hhfd+fm29B7aSv2VGkwHmDjLXo
KwS6pUXYwQQy2r9zsJ10KxtjspHE9bqN66RnHF72PMJYO27tNY5Hfx5gzFKf0f89
Gin+r2Zwi1PD+ihv9nERKMBXeo3aqZjLQhdXrIe/FAk4qc+BiMCXjq4mW2oYJVZy
As/pRdcvceO8oNoAqouCDSZFuVrs43i1/kBG4489crJzf4pGPY7oE6EcdI30kPLb
2gqAQGofwxYEFeycstcPR1vnQFeVk78qbv7bxJ1C2Dj4hDu35Nb81111Ob+emg2U
0qwikA37G71bemL4bHgY/J/rLUTERJsRuHpy/VIHtjh1n0RxKvnsFDUOnA67Ad0j
9JlPpDKH3WrEJWTQy4qqUmc0KxlBUwt3OCAYS6UToJrzUR6pHGAHJdx55E0X8TWG
OGks5AsY3PL4I1gDh4o3Nc1wwV7pohuK7Fo9mF29s4ul2vXiEcTqwgNP8G2q0XXl
XYenWQpj8/EJnXbqQQikxEkRM//u3R4bu72TvH/jFPNxNU4jzrIuY/gIwGp/bagO
v1sla0ZSB4fZpfYgq6z9s4vkiF7oaReI43u3qeN56SCzBZJ3OTRz1eXSuG+7m1/v
F2KaWGpwdjkgZij3PsGcGpadfJU0wFXFAy14DzkeM6ug7jKyv7DBEjPPIRi0GjTO
oegdS0mA3YFFXFHh+IoZsErVTPnjjAGsxqZXO+/786mfoo4VcuJZLAsFW/5iYAxR
HN7pojxs3DcJBu2QTNiKPsxw3u3HFHAM43RzIzOoQTl7+5beq7/epjQTC1gqIDvt
aEQducgwLwRDiednETdPvrSN6UL8Iyo1Prkd7wDy059/FtDOwA8/vHhhqZr5JCnR
I65e/ImWYj3cjalyKCxbhspG3BGKUGm/+ZYBZ0PysT2+iwwWz8OmEnRhLgs6U3nS
JePpOPMluzNMl2lc7tpGgml/BdDdVbS8Ys7r9WrLk1vLdYOaYYPHv+pxAz2bLf7E
VN6bmncl5yWSOltGUTi0sxKR0H6bfEtu9j9l5XA0GiIMLRzpcUWg3+1+9d4JgX0N
E43XvgGiLLDBXM80AGadbEPTYbPeKuMOSYF28AAx7KIv8n9P/KTadt3doCydrH1B
6MxOK8KOPWvOBOeA9f3GQlPq6IleZDeTYUrtG8oU13Y8hM4YaQClwoL818c5RRyV
+fPM1ei3O/svb2i0mwKhPzIyJk0DEnLwWUbbrW9CFE0N8W+YJPrVAgfONpTTFpju
3ZRBiC1hK5wQTsUsEFpuiRZbcUgkaQg/00BcfO+HXeK3Ge9XyCaEJbKYRnf7eUCc
kXxFHfzTmeUfcxe37cgHhCYX6Aiw4t9+Shqmsafm1Fd+OXWg7sTmVSm7k2qrevDj
4mrvoaRS4s0I6FKN9jpGSRkFcuphLPRO21lNKPrbkbzCXvuko+M2hsSrxaQU6FJQ
V8HyiD38x/K3XR4K4e0SVsoITvTIcHurVVvitdfz4ZfIAej+EOLIvrgHHCGUGEtO
IdrUKB2dq3tZ4fAL1MPjDvB+6ZV3S+vf8kk+cjca7JUco18WqXflyoQ7ZyfEHiRn
vdNeivIXtnRPGUN4ZevkKKoN3kxa2QLwD8j5L8uCFNsK9C08Ous4lkNxAPa1D5cM
RURNRtpFV6k00dx+CQVbbaWOobz10c8Po3C8+Et37z7+RB7dUMYFcC51RIQc+ZdC
qOaDaqwjrnNy6EcActWSI6kLaNxjTkAQJaD/Elo0Nr3wGNZkv/olfPfZO7doKGIk
MgmJ5+piDezjQBN5E0cEN3ysaoxVB+Dx0Tn6yeMzFF2j396l3Kna5ItGSvjH/JW+
U8y8UfRv8Qf73N+Wth3bv9VO4MQiGzUZ8c+joWOw0JsRNj3g3sSnESfmDH5P2ETD
4n0H0Pvigm7KYkSkYaStDAnzv5ANQJxRsDTXUuxRmklGVyADNM3tqv9tWxYlzHQu
wFZjS7AlhIBvANl05CppXecKCSmi2bfZLE5SDEpKAiLW/E63pYCa2/KQWNa+svnw
Tkap9cGe7QLqqaqG0vLGYUv+PaoNEEtuqvxppI3Tr/vJCHpcpXhLTOAoQevCZb9x
aoXIrPpP7Xnd9jDJ07o4HhuihWa+bPEf0rkg8LkNos4HCICsBRI+g07dBnkMoRRM
pso0KuQIPyEyx35G5oom/io6bVuJRC/6baGoiRSpRgvpJKRly66+AIZqYIF4I/yC
2J73S6FCbL4bZ1RGG5SIkWLvnpSD1NVMeW5gP46TA7A/tpss+M7bUlpl1m9i5p/m
6r63aALWqS3Kl4NB7262KrP+kTl3R0+RGrGan+aLRtf/WNwhtcMMMMEXebDno6nm
jvhNmouSO7xj2ExmcQTHX39bhcuNwjLElLecMoDBWzWdUVpbyg+Zh8Lhpn5vK+lG
2EPdBnJvZfCqL+iGoM0Mr++Vd9mENPLUwGipnAm45V5TYix35JCxGdhGfgXk0fOd
4KyBNZ4SsBdbbEtmbhVdAviSoO9Ohpt1Vyptdm/EJU12jPY0qbj/+TluwaC+15vx
KNcQzOuvCgCO39AADWsdRBx0QaHtUFjvmRO5YaHoIPF7bMGVKfAoru2EBoGIMd57
dIpWfycUhJNwFCK9Ihg7mDX8O7M7QN8SIhcAgeyK2VPzkzp2+R9tOAnvCjWPuo1g
oq0kI/Z0ZrjU4f6BRLLrQLkdgzqba2z6usb5D3pIyULK+ipPRWIQq6PFac0mzCfQ
msDLnecErOW3tijTNxAMrzRf0G1X++OBDNWXBXm4eM6AsnhDDNMYY0s6BXA6K0d9
UfaLV6lHJQes0vChPOKDt8kjDOJync841WA7LaF7MzXqht5+LMzIpabtDyCH+daB
5RVO7B0QAs1zqJVG/zyRatS5AXV+hiW0V0giCb04Gv+8g4YKN9b8/AcspZ3rHKH1
2ksfKmSjGmmniySdMyfi59JQdw+pkHlXWoWJJp8jfr3y1iebqb63HFucQAR4oVVK
RmHeNqTflI1ZQysqBr20t4ULuGGvWfpBIhDcRyRBkIuZnTaG6SyTLzaXVajd8HOf
o2Ashpa0aEakDFQdYP6FFehSwu8BAZJKXHoft039pYCH7rBqUvttN5XwEvfS5aqu
H77+zKAL9PNf4k63Eg+HvGy8iC4SRaVgq3mmc4jRQB7yfhiHiNpoDG8mJmast2j9
16hYz7dMQSKy7Ro8a94A6LvxNXx4g1UNfvghvHho0g+apDTcRyWqwoQ1Gr5Ro2Vr
odXZPBPuJ7xXk//i6zkpMQq4B+aZGCvwC2PxKAWFleAQTVUbr9JNEaJW6hy4Qstj
AETyn7oooUh4PSuBXzFwJcty9oRXRPWupeFaQkBSU0pu2mKXyZKjWtQk/AxLPHY4
K63tRHXdLTvPD+QXQL1mVQr4qn35K6vnxeZS0iaNXB1+QzlUTLFlY60k3KLxa1Zd
TXfVMtK4QMiEUgxFSdKe0Dok1mCK49jJPBuyzmbSr7/abwRudY7E6EKo6MHbSQhS
1Lj5RvDsue7ucUjxvPXyffDxnNbrIoc/OEiNew6YwgfcnPafMHAqpVMxVExpE/Df
9Vcs9J8EBXrRbpflXFWZdxFx9niHggkIYI88q6dOFJW6bZy2P/Od+YQK5E4m7Nz6
gM9hSHePTRKI2eXzztKMglKhwTNX7LGH5Ko0XBMMoaDbQ4ra66pzd0r0I2H63YO9
k81ZH5T2obC2GfjJf2hZI2cs3AsfqoXZ/P2dx57+SL89CT9TghFIhxkc3mv8qWse
zumdzCwqSSW89h/0vx7owQyFs7HI43AXJN+5xnGmDfCm7lOvoUbsjzRDUfmomzds
CiO/62Kj0btBQDOkNBsDsgYVhhhJ1/aleof5aBfANQK4iKLIarp2+4il6Q1/Lgh0
WtWUd6VPLOngjzffGCbZzb/tc0Cd/uhRMZSTSQodPhfkBSnUnmaLF+XkMETrGmvH
4swDj6ISOl45h8zuX0yyu7aZmaPN6J7ufXaNjWQdq9TCqASRlOESAkSea5vOTQHy
lDZXOiQmwyvis1WTAkXUH2iM5d58mtw3hE3apcTrGvtjW1+GsSHAG4PO5LCGfoDJ
lOXzvxD7h5wtQqsMT+5HcaLCG1Hc00AuqFK2m3sPWeXHCKnuBmE2VEW6haIrxEcx
AQwimeIiAkHAYD5+VBi394bEcryGtN0nn+eQvkg+2pWqNnHbWveTLA7I+TZsD3Rq
lSw0a/NZGvgTGTUwO0Z6AlE7ii7e+3TZ6HwnJcMSjWn1u6TYl0Q2pZemqvpoxknh
9Ks1uJci/U87xBuos/rFTyRC1ArfnvQve/Bc3Dh08rHWNEBDMl4hXR5AGSwIJlYY
yFN38cJJrrGc5L7K1eEBVa5Ojf8JXxrZBy3SMuXm7ik4F/zu6Hr9RDyaLoIazJ5E
Ni7t602lBDP6aq3opvKkfKugstam/RkVSf/HvTpxhE/zjpThK/zIDg3hH11NB+Fe
462s/g9oLoLwlxugcYxcfIa+crwLZft+8u2x6zuRBWpr78YfwxXYZLP+OegSq77a
3RChjBHx5N8r5J/xrM8ohFUJB1vQhhfyP/WnkcZy0ftElsHbGMlPc8LsFZAUXnzQ
UMvKMS7pb7XBCONxjbhWRKkxGKF9G3H0mJTXH0HDJwyUK5qlF1c2sVXshXj2zDAv
kCULeoR25cBqLdRIWhhf6pETPOfJ16CmownUWDjzc+1KS2JVUNEYUa/XMblS7b2H
SQFC2FTFBjjaSG/n7C+gfU2aTjKTCnoZXKMojglKPtCXydCUp1UKLx2qFz20Rswp
F7MZe7/N9WY9B7xuxEWmU7/SRhI5zbjeizmEl7vq7/pcFUmdodYM7saZKQdwDRiA
g6q1ITnpbv3AsSYXPhlDHyRkkECUWi3v2J92AI/EF04ko79Z6bFbSorub7QWjjRy
oB21J5LNV//p+/l1b4wphuEc7RJWAno2Eb7SWIpfUwK+HCckLJjZRZOv4e4JBULL
36ZziHM3deqyMxFD/YUuotnDgZkzTG4yM6GG0v8VMNGsx1Yn6Du47q1f03jSRPjg
bJfI8sWZLB/mq+MHwd7TVlnDbC9AxYYnkq95yvBtRNZ4neOv62Os07vDIku5uMhq
Ox/C3GHw6I4dTPcnmwOK2URw4Jf/3O5IiSpl7a/X7BTBsIG6OFW5HIES6eN7YfAs
ynHMzIbnL8o3i0It35IKRYOg3MPEkfxQEvjRhND4uhp0bNwUqbemHwGXoMoihesy
RLq9f1o9md+6AHoJh/9kqrXAnV8zwk9K2ciO6P7Rkc1qn7+EOjs0ulPM4yi4D2JJ
Od0Kh3EGfLuU5BuRZt/Wiw3dyG/vR7qsqTCMbO/UW7n/BbKNZ9Mnc1cMccyjKDX8
NUFfebfuHRAJNIb6EMZ9c84piSvEcEbeCeCL7AP+IYAvfCG1jytDiTy5p9Re50BQ
NT1tAiyXMIE0zA4HoqJ0FP1qf/HSzQpJDgPKlQjXSg4Knh8MBo1/suhoF4i5Hpt/
RbC3w4JS9O71XcOBMyHXy8d2CAf1sVkC7OEqTTu3aSCdQhPaGpcWVibcqoQndg39
UkAXpFGtiUPy7tIyePk9FEBWufnU2Kp6koEJVaJO6DvtS2n5syonQBZXvO3ybxW6
naCaLWhzEu6ctMcULp51jzrU6Rsat3UmFRoJaLumLHDMdHqoEGaZGNE8KMLGZYvf
Gv6XUI7ygu22FfvUSOE5zOVC6B2mt0OGvYh01vc27K07vU5Fg8U/Rb236c/VVV2p
O0z62pNdvWmsWYbUjBfXbCyFTTZ8auIbXeOGaXGayE2+c4ncHBQkP8HHQ+NbJOOv
PVXnW84R4usjN8/VHdEH81S7GdbQk3A1nSp1Gzk/6lAq5zdZy9vpoLD9vM9N2L0p
pa3cfZbRzIgpSbQ54SvpSp4wKVyM5azPrFXGNHTVOUY0Qg5JWy7cCMM5m04eriWZ
PbgBVELspmXy4gd5F2yw4GH/ygwx2FJ55Plhadip00/NywJwu78cMerTMNq/6OSr
NwGrR0fsMbsvu7P9fbH8LmiBIGIjoQfXQgwNTq71FssdtEbl7c3zpg9b9wiUw3Lf
myLvR1rkWYoH+Awe5Hhsu9ebvB5O2b+6SL75cw5klkzCQtkJPZq86MhyfqNNJYvC
Jk4pxEzd7//J+eFe3GMC6FKfLIKfiDBsr2Ra6eAXeRPoBDID5R6zmdOrh0LU5SXo
BiHOGTXnrd5UgHKqZ8nBO+6ScutwN5Dkl/kGZmczT5VhV7C/vh7cb7a52IlU8bA/
dv9175Yi8VTEQUdN8DOIBpWMoOggYI/f4mEUxRjbzbJYSpKXZhoyzvOsfGqPnlBz
A/tSiZhBavBZfth6MU1oEgG+01cId83/Q7PPXhyt268xZAqqv3ttG5+9PHCTdYDx
ALi7jZNd5pYuuIGXiwzJ2c6/c8m8L2yxrWIwhfbenhhcmOsIcpuXj8hp1PJ4rR0x
T3x9I5XPBnR2tPga3mHeRRr31le/CIUgzW0o8V1p6jk4iBmdsF6rprxHeGpeKcGi
lk5cu018FjRVvaoiIPopfoewth7unoqa1yW0KQR6nczHCvgzWM4HR9V168nDGXw1
h5Mg6MwdkzanDu8dVjJmA7i8hA9TPd/siUGDnDuDtKSJZwDrbPmH9/Z0QmOsr9gc
ETzxGc+JGNND6aR9JKsPh3jRAzclkzheAceYGRUdYuDI9CiIZR/QYb1tw2p5IoFI
E1Lnsc8maN6kMK9tO2YOj1K+LAHitaWmrTe0ajdTKtDrDQ9JRRS4pLBLygNv1aNZ
mVnuL7KzJPFBqneYS0sAsM4eBrVgu9uAKODFZXHvrrHLWY0rHTO6RCFCljm9OqaO
dGQOi++Kh0ij6DGNQmb/Sbfqb+38hbqKkEm9Lrl5VtKTEDrPTeP2yIiGJiI5YYNE
5C5dLGbEbojZqs5cx2zaeY4ETUQQLHZk0Xs49KB7n0x5Tbg9lDn8LjhBINsDx1zU
9M/O2WUlIPVTSg2FSjo8sV4PX/3yQBjBBX5ffpqYRbwXAZupSXsvdgGgeuYz0FLm
EHMzrHP7d4lVMEwuxAZ82KhDIEJIAhtPz1/e9da+xfoNXJrx36X2/Mx+esGoAhbm
D+495+6OyViy7TQS9IDYl14u4VEd0HBVUQOBVqBJypKkPN5BI7tuVlLBq3dlTjBM
3n34Md2VVtu9OyTm/pN1IOkjkmlRQGc8Rb8w2AmN9tDX/V385H8rZ6QwQOKMoUNK
F3ATFYWFDS1cPCaOu+v+tEJ1Sf8FkcL8Ndyj81pjeN6ngZ7rUYrTPn3xMmqfR17m
aXIz/kQAJmX4wcqUztsbBXLiMnM9z+qi/XI+Aue0oeM0IDfHPHUQAXuiZgKf08z+
n3DiDlPEpAyvQJSbeBFSvlu8jKeW3l5+SkoHaQNUT7rTREUP3SA5wikc0QkGXp9m
/tHsKaJ6LHINu8Y4MBcPnb4Cj6eLFMmInYJs3InM3wtwi3OblNKyCHrOi6NWdeJj
2ZEQmDdlSsuDR8fGuq9wzak8NtuwsTMal3XtyGEox7HpVmGbWioa0vnyyyT8PFNj
wQQHJ2ydBuWsDqxoIUNspaFkVf55AaA5NP4qC0I7NRj22bB8eASxwt97eYtjl65P
rJlRWA00syKtoN2GlvvH2U4zd361KfNoPMHWkJEduL3Sc/X2+6zXReW+trcv4EYA
i5DTqZEbm3zDzvzCBbIm7Fs7gfxTC1u3DWIWftqVka1YkpbC6i2KGUrUp4tiCMLS
zw5OoB/CNardHQa6YY2mwXCjXqpQkSIIHc/3m14Buaov/OscvtL1bmfmK2gmabU5
c3j+AwQiOA+1NltDODxBPMvyyjJDqyR0bo4yQKk0w8TYs6p9ykGkFZiqMjz1NKxv
72SOk3Rc13SQ+xVnBxM7T6WbzNfIy6TwteHA75Yih4sdJCbY3nA3po1AtaXjL+/j
nAqHEdE3XcN6tq+BHQTBxK2xzT8IJkeVQfsBvv2/VqNsURFGZGwyvdGtxqfcDVGG
v8nLzbZdKYTBooHQ9TU9pvsvC6celZCqbE169Fwha3yletNqk+rFPRqXUQEQwPhL
hH2BhZxQi1FvdAUzxaQIADaaFSxK7UGdppalGp2C2MFasWEOx6jCekTEw18M0sbr
iejDopKCGkLjaI1MY55uhOFqQsCLW5Y1hC5PGBikwr0yrtllcUYNwGjP6bbtofIQ
87zP2la8xDn8Mf0WL9pdu1cqpXpwrUZknR1Hst/FYPZOSuBLkm4dxnZ18/TgGaCG
NgN9zkZkhCmRCuBLZ2mYhHR6OPaOFwO7NKx45rlsdYUMjONmr+Z5Im22m0JKeGWa
OfLqW85mvfTw348RQJ5+nYhErswM3YcVB9efCSvlvCJhM/UrRVxIfOnDlvABJSRV
f+lE7QxWRBZguHIKPeLsTl3J31NNVPXor/rr0sO/QdpEcZEG7tDfAIw6LWNXUvT/
725c2qcF1ORSj2NETV82vfalS0/QlmvPHOZmiplxyohLlMZG6kDljSKMAj/jJrTU
9moss7pjjnd7y3pOTVWwoW+/0g7jH8mrniO5rgBgi3e0Jf+A3pOoQMn22kdbz99B
fVLz32mZ8QzeZexmLJ2dwYrnhjvtHru+BFSAuLA1Lw2JBK54kcef4Z7DA0LMrSW/
Y7zypHo/FkDVsz/V6hlh6rNa7Xw0a0YGWDeGQ5JsNE5IWbXdo3muOAzeHEjuA0PY
2X0KpIy+Y/BclQWwLJnumYTu2XkJqMxbwXM2OZLXLXwq16zGpuEmiR7ndO8zdic7
0xhfGtQGMcQPCAhi6mnJ9rXwutpgFJXvqQ+Q00eOsCew/R6XJG2+WmaN+ftU0YdD
Hb+dLumCe92cBE+4TecZmKC9MN6TJ+zGhGkcx88auk5intR5HfeHwNRIsAj39h/9
xR4zizgM92hZX4Jt8bvW18iURINlqrWfD8FQe+575E6ZFYqFYU6Zq+saAFRMtAMx
/0LPgSkGUtXuuUsILKMBkKZGxcU7nkInk2w30pEcxsX+h9T2LG6IEaOJfh3VvVlI
+kI3/QSqv9Ao/YWAOCyuLQqkswJaX+jA905voJOXvrwv+jwtFTJWirh1QCEI/MJA
+XT4Gj5pVn7brtlt2+NxD8HqBS23+RF4eYaChfhrLmEVJuZmi7ExNIjTBfk8kQqG
f8+OEKz+vYpzJDlc80L6E+KD9/QLlex8TcfGNBIqO+zGzKyTgRQutuVgcCLHeLoG
9CRd0tah5LDXiJ3zb3vFQNmP0SeL9vsX3r5ivG/yDaRkQSLFf6OsHPctSJgxj4Kg
EkwrRXK5olGt/R/nMx2zlsxZBXMDnaqpohBDjoAYLjJOtQxyzTlO3VtqEp9GvWhS
gUUSuCyDQzdRAr4Lh+lJvC+vH4mGIm7eYdmoCObrDDLm5yc1IzR6Qjn+/DFGBRqw
TP/xAzj9DbUSUvozv98rMvHfk7inHl9ngz3Oz5twZRIq82o0i9gp4Qox6D3OFhjf
mx8x+vGWC16zhW8J443+Fbk+wN8evtjrqr30wcsoUmsJxvlNOShAGPxpw9ChFYV+
qvzaN9sZCpVDmD/kIklMJ7QJHo0k2hXiu9Zq3+TEq7WEtQH4Tnu8nIMeuD99QhI7
E7f49GwwRx3soDbM2xuMgUywMTwuCj2s2iGKWPX9agbzCulihrrYvUx3Fez4BvYA
W2QX9oQavdy0Q0WgWQX9dRtF0GCGiCYctznF9kjt2a1kWZNwo+NBaD871LaznIKr
1Vv9mHGbLKZ2FSv16pRvl2pke57L5SNnO4ySHK++ezEG37Te8gMiAcNbS9NgU5bg
UcmrwX30gRpXBs3XJOsgWv2kTdppuGagseqb5H7mmRpwgaIfI9vnSpDyCrV7lyek
9evXeGQy6eGxROCaoucMFiielfZRHMzA3YuxgFFzA4yTR+wPHWfIVFUuao+6u5P2
NeYEBf6vjZHhXiQ7nHLR5VHLHFnzrhDm+KAxMJGvkv33FbvZ4e9F0CQpcDpoMsTq
zeu3ApgfxQ8HpPj8KWfOglUO+r+EGD7DflTsHuoz0smr0sv3bOpwGEQWzHEJyHn1
gQ8w6sU51CAmovUhmOTLMTQnb13KBf/s+dYwKb8usX9WkdH12fO4B9edjWH3DlJF
epTCv3uf8X1BbnvfAZV8BYjnmoz2tz4i/mUrti4DYgeikXjBBXHyxqq37J1RU6Eu
r5iJvdoIav/HUnQpERbXPumG3oMRPKUA+mukW66Yz+IMKPhXGNJjpgBeH3zGQWJr
ib1kO/WISpKdfXbDQrTpoj6f3ZtrzOtniKpaNJL9GSMkZnRETQIa8kGNbjBQmleG
uXWIWYSG0AI/85gvQPSkyKcaOl+6UQzozQLXxXFEcuf+QX9/8wGR57BpsiZyFvXO
GdUSFJiqz1nCXsjR3P2K2M2xJSSsagSy2ja5ZkM6vXfYFEwOo4ERb6UuLFtUt73e
UDt8RFEyMt7ceTE0fx3bUD56buOdVPMJU7+VgCreejnWRhbW6Bev1V5JRN1eUOs9
cCnbQWzFOrpJkWtwLLSzKakp271M+rgOSK6EUJ4v1Pkm1GYprrKU1jltvnjkVu6H
fFibUg0dihvXBDBupveXwNGvONrce/VWXcKP8oR7PVDaJWtiDXJlHQa2SUuylTuO
Rrgh+4FgyiUbJVKhho1sAmMSd5+EqoDD7n0aUyGgCgbXPAS4/ztVjTlzXS7XvRGt
n5d8Z1vZ3ltFDKQASg5WhZOYHchG25PbS+JWZ1pKLQuAmZ+y15xlWdhvVMs73FkF
iv8BAIBb6XcWzOmJM/XHpfybe67Dmds4tUt6xYXtgPVW0D3cnmHqHOjYM0SKDS3j
RNzPiQS1LXPR2yw3SOUn3uDIkQnVWGZpbRUhKb0dLbdB8R+ociDdgU+TiYa7En6/
WmQ9De/LoW2+aF2JzMG5wmK/wQnGy0PFrJBPIdyk56MAdcTKPUKGAsKJuawV2i+9
Mysae3JZt3rGvjZr/cWqMJQpX7BSPSxt1WukLbSLxhgGambQfI1lQVGUnXMBJgif
7pf11KB0+HXZq4VOQTsqZcEFcIvU/hny7xcQCx49StqznpwvEJIRDzdbk/hA3h2y
IP5Y/txwsfWQ/Qtl1zHUnfcdOwjyaPjZh3N6AcRBZ2FphhdlNay6A6yIjvmVMSvg
LEXwNEcWWpyo86tA5ICADTUnCPcE0Io30cZyJhv5Qw7hWsqkNB/P/BRJc8o3PV8X
Ww9x5P9ebd3nnCo3VP6qNvWJTp5HisSYh/GoLkCV4oGJoOK/cJggwS7eag14riUo
knJjblYmh0b0ngJScfc6KhakWiEz9lVsd0qheUflC5FhiVPSxjB8uULIPVjg8oM1
Mqjf9X136r/txb3TWPqSp3zhPEwJAsN9IsBnLraFixk7Xc3Lb4IHRtt6dgewNgcT
SLl3DJZ3bEjaBJiHhO8vuejKakR8bvnuF7Ljj/S3NHyJXNQ4TECVTOHTNebtD9/V
/HYl7OeTH0z95XZFZCjEpvVc5aa3Knvh8W5a7e7SVfcrXe35ASOMdOH0KmxXFf85
l3fA0fVLAuIKlZlIo++gt3U3CNcQCSjEfyVYiu2ynYkXP6HfYbs/zBQy4JDaRZs7
R3zNITA9mekzWs/33+M/klC7qwcRDpCvc/dEe7V6GQN8gPcrHjlN4Qq8HUam+r1O
lL00mfgFnyBYLqOw5YPnKeUC3cRoaSz3BV2yOTH1B1ZJWumrc6JnbY1WcglSSirX
bqOdWhYR17DQJnPcejohMQ8caZqhgfj0yOakfkhb9Yo27mfF1GsNtKOWWO6CWy4k
W4px66MAFNmvfTsPKWCq7g5ToZ/GblvQ9J5K6KdCqxV/PlecFw0ILHIczwQZcrXz
mbhozLbbYOmidGWHtkilr5E96jNzRryAxptQR3LnPK/U0iBse3KNEiuW+nZuFvbQ
TubAzzi6AhFRyAz/ZyQ1zM2YRYRbZQMzIvxEmjK+YZgbrlYNM7pVZdqR7kPs6y67
W5mp54PXnvK2E6O0I6e9+KPydIaJpLIAOzjdei2gT27SQIq3Y+XkjC8WUtnQlcDb
Iz8I3gR4tGyrMuLy+hIGabWuU6W1mzEX421WIFNmZo7cl6RlQHKNpZq07ncijtrB
TjyJK6+ArgxcRlxXBwUApTvo+vZYBT09K8TJ049BeIiNypJG7e03xiNO8QZKDY/T
xfxwxkOQKmMFJ53sNbeppjtrvtHL9p535ce7oxpFdO1IYspNLuC2vyajbaJsviRE
oboRafjvs69xfyHDpSg8qxxCeZEPCAlNBF4OPH+Bw/nsQfBrYLxcOmQygPKEc3Ek
bDDUebKhKsJrQs2Fp+EOBwi4SLjOU/keMRCL9bEp1zfIzLLoGh6aktazuTmlt7te
B+RqDnPl6ju6zMvaF+vKX93CDY5QHDK61qmnYmLopzU129TV/MgkkrrlNsLZwCVR
+OHbZsONly6RpHzajWDqpg1QaInyo0oOXHg/sllzjGmn4LoO8fa0JSd05g7osw+b
ssNr17nZPH4JXPBsCAPhhPNobHTkvz6ObBWz012R/+nIwmfzrU3Ov8ItfF3Jduv6
ENMCKBxKwT5PAkO3P5EbjDbP8yq+XnONPCfOC4l9xfTq52z3ZDHypemxhqRUOaMV
pbE6wiYFgqtP3IDK59+9FhkLhqE04C02yOhV6XK6BMyQ3v/gxuehSwzWZekg23dO
T0HMbqE07sO5gjSu7+8KRUtWPHbCBHd8I1GCEx0K4isjGXWo9/j9UfI9H3fKJcvp
c12uioE7X3MXi7Y+g9QQaQW9Nm7mMeb4yiVtr6hszl16ZwXednhm2zyfWIO13YIa
flMkkT/ypsCokuMdghpr57zLFcVq4UmOTEcB2jFgewwbyDSmJu7uyYzpPdWorT4g
kQqeDd31AdmuK2EekVDjfpmO8dJ9k38PkUVtiFVWPQKBcyRG3zdZf2fmDF4Relrj
p27aUDfWtcbx5oEh1q8Cx4LUKmMnHWfutjEKJI5wLhRr1o/W0o+RTS5Eca749xuf
nwh7iiwOS8w4OiF/8ElA5PP4frm3jnNydTcOgNdqw0XLg+4ZzajGvxz2fVf8SnTu
iVSOxvJOdJLw22nj9pijdq/wHQZDY4XRLObv0SVBbeJBSE+Lk3zfavGs6rL0/kie
3WUWxiOX/fSxlTCoGQXcnkT2p/Zqdfdpb2ecVglqIPiMmvD6bklm+vPsPZmwkqFy
xkNE8yjpMlfBZ/EkScrKAB1byygAhT5rB1zBlcs/8TC5fezIHpMbqttbGki43kIq
unLIN5BBEkYm1tL9BSQCE0lDx4N1ZpwdQdtDNGAoEYP5t0Hch8h/7xQ7eNNbhXF5
MDohAgD+eOfCrGS9qyAvEMmCdl735r1ObhYzV7TTU7ZrKZy3MRWs3Ncou+Fwk37G
xYS/TQ0rcAmYxbYtZ75wn9WhkkyfER7XqyUxkAv9vmdbTCg5gdJvBSmB2MSHOnUk
t7A7zY+YVr3c0mfJfcvlsvRNEKb2Cwj3a2+dMi5bAEzclda5CB54fdAWUATr845e
JD3XZQr61/v436Q/XrWFvwjRqzouuj/uGezI7YnadVWXUNzcp/GoBvvRqX4/i5oX
f6I6wKwnnWDl9PpqQ3xvEvkUGQjCkt3AJHhGDeMvRv4+hRHz0IeBu3ZDVid4Uw+b
1tmA+A2i1F/D6Tp4/DXduOVB66tMWKKvRh8v6TW/sGppUvvWZaI9/lhWSdI0vNL/
9zqYKIFKq+YbdnjkA/z+fQ4AeKtJKT3Orn7RN9RERu404F6aeO5oOt6uZOs8UoJq
XX31Q+Eb4EEreB3559iv0iLFttK3rwMTdvxQFL72DHHjlVDirEpePTIeMNKqqo9K
8xobN+cDWs45FmbdWOBdHI8Dgq+U4/EUkF6xMc4BX2KDj4X+wHM6OeUyi1l41+5T
vyuvb3uDQfCpb3fXIDv5/V8APW7MFxg9PSO+EA8GOakgOrwVXS3pNt9YJ986YcGP
06OBWbOeI33MsfhMKeR8a7ZXdpCbdUZJJ954o75pk+1FxLwe9sVi2eN9bhMhjZXu
5sqPdht0CQ0ZuHA1BU6Kz6MnpRzvfDNv11RBa//CIiNLQ8LQkuKT6dku6YWFT2ZH
eGBuLbRwPb5IVFiMDWpwvPAtwhMhmCihukQzweIqI4QOhF8tJJ9I6LkRMQgrWxmT
gT98y80to5/rSw5SdxDHrONGFWveFaLCCBuGKjh1YelKamB3IIk86f4033mT3yHk
/Gv2f7NebVp9F4YZvUbol/zlaGcgJLbVB0Bko4uHRsCHPrEC2i/MGhYAy5kK8QJu
6h/Jtqd22PaGQwgPlgHIU68Tbi+fFN1c2/k0A0jAGFeb05BN9OVvmPUXnS1wU3tI
AhS23bM9nEDKKvdW+4GxkUdiTwozeb1SQe25D2T9TeULnofPR9YLCdbjtqhDnI2x
DLUDqWfURrcXnfdwlujEMhBydeXh5+Jimc2VqEbgjiirdrc4CD3tsxey2sgjQTGj
xfe6rbN+pFBzr0bnaj/awDNl2vBLfA23EodtkbGzptq+6L2q6wiNqi1co6RRQHQf
oB9Yo+coyiM8V4/sXs2+1GGj/sIpAnVemaMftpogY4847RrAMAVMTId3kM6tzzWn
NEV+i+TJwozQ0Y/Te8XLjPtt7eYIwwQgsg/XdErmj2WchgCmQrpMOR9SNbKzl277
PUuA2diM9nYMW++xEK9gJzRflzpmiSAcnr7BCvxg1YHmVIFgFqeCmfZnX9zZzCWF
76WlEbWXKYVADYx2qJOsFRWU0MUowcgQmFd/xPRnK67WSi7Bf7r2tvxD2zXrCJQw
YQUWI8rZnqtmAMBDTbqDxME7G9O7+9PB/qYFdCszGWEaaKjINk03cCm2W5wI5BnC
q94yq/SVxqI6JIR3/OXM+bllkIjD8FpZECv3mcEirQwN2mIiFltdXvzOx4+exi0X
3snEtCoF3N0RDWA+XARNAL/1mqUTRpwizq6Gy/nfJuVSFJ5e8OEhou6Pwwnn+fiu
0ghIeP5339CG4z5ctSZgXiZFJmlg5j1LNolBS9Fxv5Gqc9w7hNN/4tVD6wnqos7G
xj3e7bpLNuPkfjMAH3s3ZRF1OVO2qdfqcHHcqcVJ49oBcccNIKJxOgg3Mqm+3puh
1uFAyzOenMXOi/uftPA+3mIrvsn4PYudicCSVfS9YBbTHGWE6feTuyapH9yikt2v
TMr2x9PVLbpe9E5R233wZmXdoOPZBhQ1fA5VLGMQegDc/TPTUkSPfCLtvDh7m+hn
6wtJEZ4LW/K9Ht5IDndEG1mDMSig/XCDgZr7/PiMs4EuRUPsw+UOSQHz3sJSJ6xr
FO8f0wttQDSjb+ZjSO55k1oh4Gx6hH34KzWzSA7StSReGrZT6Hf94HdxJiDRv/yr
84lGVoZ2TuPNXPDPqxl5Zi5XUV0Qk+v8QshiJCR1b9A0CWLTZaalR5Re0g/eENBb
93sQP2FmsiGMKOuMIQh6CBhPbPxhUiWMkwLa7Ypm2KXD15TiAzdH9ijSISHWPIOW
ibgco+CNLP5Pntk2fmvLPONI5ocesghdGVGpvYMcH2WgoHfQNEpObnanzetOJfs+
q1iTcyuzPeqVEqK4pBOgeLsJMfBMEEus5b2BchJE8e6BTU5E5OuLbdRd8yAbq9Re
sQVfoKdFh/Gi6NapBiUeG2ImmMi5ZfFGXYl/DMQPIF0e5qq0LHkfutpqJ6ZUrhLb
N8GeeZpm0sTb7E24M9JMt4YBoAiotRkdAWHxBr7EZ2AO2F7PLgExzWYMXoSKeLxZ
csS70iukVtixR2s89k0H0qA6RnjWK1GDOcyN2f2nraPFD24e5bSBrBz9hIIJuHlL
AImWxsv/b3I9HweutshvMGznk6cx0COcq7PGJBMQ4hwkbiBTivbiTKeqmLcJjkzH
4/BE66ZbjntnCH7i5KiREpYT+msQoihA1qrpNuRYOa77P0gdbsG90GmEkIyKfE2q
EJi5YDRJPeuLl1A28g6fPWsLJbTaSqwKjm5IogV3bvehxdT6HglOW9cPq4eV+E7X
s0Aza1vUlPk6Jqs/MHmBwxQl+YcLLyucgcoKYNr63gq3M2sCRQ+XSwCHR8ZkeJE6
NITLGFxclktEGRzm+1S1pLR6YNbnxXIuWFNejq65yFb0qzlwOg9Q1oJ7QtcqgK5C
4rtPhW9tt0zgEnscHHC6Y3fdBM7GJo7pXaOFh+j+8uRmBNQ2BWoeGkUeiegpV+7E
1MRjvapjb8PZdvHzuW7rRbO7kZkpOl8InCGDLkTjZmwoQAuQXDfJvqvXxHlaaNPN
LyBuX3jbeAkTJKXt77V7zPp2XVaLsLB1OrhsyaBIilWkOorkcP2pntOIlxRErILI
yrcM5xN+oNVaOYsutNtlbDuoovDqEKM1QnkQyDrv90tP9WYlLGzqSkQtWTid4nIQ
VVnSJRo0F6psNqX5H2SRrzPPmEznOK4VJlu9rKdwbjHh5oFo6X6P6OhJa+R1qXSD
WZU0X42eCbqzE+XQXEBEZLONDOxZylTRH5S2I7yBn/LxuwTt78oJ1Ig3ucoIY7L3
LrIVXand1KDCQcoJKXPMzzviqKWy3HyEj8LvkPPvWOqLRqpCgBs1lzx3A5nXmV4c
8vN8aFrayiiQGkxAahj85xX9+QgZbNhNXunD3lf8m4lt0MBM++/4eHwH0Hcw2ucN
R6IOMseJ6zM34z3Z5AbzjasBZ+q9ffvbDzTve+jcytuvFgzSof5prJNe7O6yk59p
RC99PxK7EXeyHqh3flQmxamr9WMaDtQhYQXFRGmfDY8LxQmcwk3rz2WFF4w8iGCX
Dj09iwC6m9100Ev0eP78Eff8K/570fjz/pR5ZCcaysf7mUv0l9J6YvQgoitQRG8t
Dq00BDpK1MZJzCrKtOyTosHtc4kX4QB0darr1cg+arKyLRfYnQ3zMx1GxUWEbDzS
ltWMchbrKtIwj+Ge1A0ebNYJcnRzf8Q45IPMHWfb/PfFxIcexDAgD0q8BKvAbMjh
NnJHMfpFA3AO51PrsetHzvIzy0HJPTMAQjn2y0sEUWBctHse74pIkxE+M1I83yjo
MsgvCXWXEWdQYHvrCytKt4PhZwCGcv+MNHK3HN/MkT1kdNhXCmd3f0frcrUIsPkx
V7nYWm56pSAHwzZLJuHiboKA4S3qEfRFgV9FCatr4/fxLPslOAUES166HmUsDJ6S
hMWhqrt0rUsBvtF6dsrdkJZ1OEMcuR+LJNH1FL8ijlxh0tMyMX8IIda7pPvIDK5L
q0vcbgz8ASXBF1Rnbbp9hOjhTjF/zmbQlSsIxEP4PQwhknQcXkLmUPpKWEd1dxQv
gN24MeL+YlsmGKW5MkR6nLS2hyiP/o/xxpTLqdQhvG44RbdXycA+LZqC/gkhJg8s
tNSA6xl9VuQ1GlBiAY0hPbF27+bqr+HhwrTiAClOrpNry42uCzhybajge1DuU/3s
QoPy10j8qUAYyBeZrc++bYAwLNEaRRSKVl+0FjqrxAA1bIAKqdHkMPFi+BIHA0Dm
b5QCr/bxnXj0MRmpSB8HGamcfRFvt12Uh3OaP7B6igAe1PXgkeltsZ5SqoNbr30v
l14q6gNChaMb8wnm4u2VnrgsHp0kZBahCQx/7WNWmE9aNebfZJrTV8G8z+JklQ8U
B6UnzBTIZD/TlBzdGVZ/mcC/LlbU/cnYHDCmQbRNk/pTrBlCb77v8aOLGhExmKz0
7r7xmsmdHZtwitZa5P6rYd+xPEqmYNUeU73zQxgRuXl28wLp83XdXF9KfueNo9DJ
hZh+I/N+erR7n1rHu630jf/+8bGyLKv1Q/KCMRufUr6tvEx0xmyt5yyhtr9wiQTE
rmtVTmbuUAj+bLPlAgx0NgaD3YTHs8gbidD1Q3iDKuko0wKemhXr8MwSK/D9k/VT
6BwbRfUA2OEC3lHLXcQeAT5L/XMLGVhlj1bZg6G9DeW9DtIdLbRLCXUEV19FjxSo
++jFAmssG6LT6q1dOI6VZ+R7gZY9FyU5ZEFerhr8tA+yN6R+Wv+5rnUPHsaLTvQo
3Dl4ZIE7JJI+0OoAORDKdAxrwkRks7Vmo4lptk5w1HDW0i0apGqzwvdk5oWdyaLO
V6KdOlMa13kqy9O/NiFANGCcNAzAMTjTNTRC2g/dm47EuheyQSQIYA8ZKYUTgLl0
O1Y1eT6hNVLn10dn99AeG7Mi7U8Db8AodvEtXOSxXTECF4ZIZqF0E0k/XLhHGiXq
`pragma protect end_protected
