// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Vme/xv53NES7IHZVfyrD+Iopmm9Wgg9J1JZqFZq7vFrzO5g3x6UxhuLvfcVF1BuzcrtBCiWASl2e
wwyu+xf7UDO8hi+5vM8f1i/4FBNuqV/gwai/PsFgtUSsbHmuU0/9ZWD8eHU51OZ8A6YQj6TqUKcH
IEfM50hxsHhfkKch9zgOMtDngWLKyXxwYKH9xoq6fofwP3PWnssq7AfhBT8N/x7Yqnpka2wn8RW6
4P2vKhLlJUMHWHLMFP1cMRiaJ3pqz/gb512v9RcSG0jl/d1BkNIkN3vgEUoRzxZhnvvZ/SbtmBHj
hxRqnKy+3cTGNLKvoxQjj5xAeDst6a3Hr0WAPg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
2T+tAL3+bMFDOfxly4OpXkPdmp77+cp6R02zOXLfKt62Z79tpieq35HGYzwu9nzH1TN1l59Qu5wM
m40AsIF905Raea62Gyvta/CYqFq4NngUAN2g/arSai3y0Js+lU1OpIOtbbeK1JUOXQnZSblFi4GT
/g/4n3n6Nkhm+lmnEte5ytiFW4okvF6FESPRrNrOvWRCS8UfXsi7tQ0KQFD9zv/nqy7g3l7iro+S
GNqiwKn5Qmz9bS7mw5Ln7J/AdGx4/5ts1TniP3B3R6+9IdSqbOVjZVzcEdiqfGTPC6AMOJrv5qvM
ZKOzKXB2lSbI6K2sSliWpx+1YeGJGTJ/qct20ESHtY9q8nfzkUi8aaG44AIiR6Gi0R+cXbtKPuxA
Z6yYBrsEkHJEwuVz0dqvBxvApHe3WFfWm944krkaptVT1M/KoevVv/j8xLPU+nUrZfDWb5Y4Yit+
4H8ieReu6e2XPnuhzKUK4j5Wz4+alcBqhgB20f8FS4eM1B2s6gT3FXWG7F9L/ciTMs7VglI/xPuc
WWhb9DNW9/PCZaUxgwKBoUBcZvjvOWQhVi25euZiodUIbJ1bWeeiQa8eim/m1Ics0MBPPKb6rWdn
u9xGJvn0zAc/qomX2G/hoSx+LDQ11aDjputdE0kEG2eob9AEndk3gfjFyFI9n9NBGuwi3MVvFLCq
Y8hmpGsFyl+9hFj2C8EdeN3/7vZ1uQDbpIDwuabOV7lNKFpMR3dj96T5vFIl96CHsMzHR3m8ehqT
59/TwlvjsxNSrisNfO9nfSZarZ+clD2rG5skX1iHphGHaBcTikxh4TdjnPnfcayHn5F4pFt9MSSH
vwr4V2vEjNE3NQiDOCwRrkn26CzObvRTZsED1jaoNWoVx2Klwrg9OVaDH47O/OYVwXr8uyaeZO2K
LOBzz05rMThZcV+hbm04V/AmUUnseh8UjLCj8y/QwIexUqDZOlmZwZGUO6OThBJRDtJMn3U/uoAx
GSITR5j+pX/gcJvAtt+fWbiEe9LFp333vAAguhMjBYtincomP+C26MpLG1Eiomdmbce5jalzPAxc
6oPM/AphOX++y5yW0527v0Lo6wKbpCmTH8v4jjTVgcVUq7hgZ5vW9luZ5ALU5xw6HTuCVV/Jyshm
wA95IlAEO2BcU7SzL7ReicX4gO8i1JXRgX4Ps+9XzMTxTnhIxKUzMpUwcIv28M+ibNkQ8wZj4bXK
w2iQS45Czf8Nh4LTFThATpfBM/bPLaZHz0IjUcK/rlukg4ZaMRh/YgQsVeLV8gIu8I1be93wRWMa
uLwEuwJCuYObSvqNvhAYM7zyJ0FpdrlK+GQ7+GknXAaXuTarKgZMKoXrOubMVcX/NOrVK2n6BPKt
U6PrQQtzbMbTdeBxwxHsnJt31+o1UNKYhX5maLHUPOLA+9SL/gvvsKfGsdquZGFYkpaPty6FOyqx
bulCtXaMf21grPzFQY9WXPkjEAUsPw991odVxTJQNw0Smu3jwIPFumsVNTyb61memGYelaWepxO2
1iuB8aEBkQGKa/ETy3xvQNita2jJVda6UsDMIp9uhL0sFDFxjVub8KfkFuGcBvKpg8tFjFKOsGe6
Qg4AhM60mhPrv1I/ekVgb8nyOwWxSM39rtIwb/0n6FP255KhwLsS9nv4nt8LKFcLGDxpK6ymjV+j
zoWfRW35loanp3DTWvDI91zgXf9iFb1JrhPqPeIRBAB7Qn/VU745AemhMu5ReY4jLFVbxbRBc13P
u4s+Ulh327M4ZulvEm/FUt0BEBRSrzSZkrU35a8hnOvVqOcayTroNMlS49NE7vjYF5IxSeE2fV6m
TbPXOWXfqqjW3/HJBZ+VatP9jIc4B0t5FJXgAPBzQ7kymoAMKWUvWaYLKh4NmbcOulyKQztNP/nr
PrhqcbaBqPSJbCtmu+BdbV4sZJUIgSHHM3G+HJ62IVekb1f+cXoIaFbPaDbGA6AIUrPQWCCdr1UE
VzmkbPTt/NRgvx22qUCOni6012G7RffqfzN0yD9f8DMM+wAUFQPHTZhYmsV+Ho+/QqnJI7V+1sdA
aKs8WTuJIbL7nZehwEMLgoiqqQSjITR8RV4DOpSnCGf8MQqYz48qUj330QgRK5R5Bk2MqUwaBjiR
VmAwkEpqvLSmD+XnBzdkICBugw3Sh//mGx59D21oWVkELyC+jqyMEGD2KIwNo4bY0iR1kCpe/raC
gwXyXhhqr2klZ3t9dzAGcxarzu3v41jbV/kGPtInOF5nTmPsNa2S7PedUcsesJZFhvtkopuQKEJO
5rt7WRd7gUqD1MEMUncQWjXXfQSpizVCUHaqgjd2/zHrywQE7TCndRO/XlzetdJ5wwA2Q1a9arSz
DQcMoEJHuZTqLPnl6I+CjIW4Rz1YroY/dBBLMIk6frIJ/hZnD349Ui6V0mcjmY8lAUohpuc7bc/W
2JGt+QCfY/rmT+LexFfgCsxYcjutFRpzcKiFz7qo3DjZH+abwUoJh/kKvDCeFT0nmILHocD56wfK
0LbK5fSltQOcDSvmvg8pXkmR6rnbQtu5MhKyVsoWRreUa71IiayNlLVONmY/83+bkhaH3G+Wnr3g
YBMyk9iCOOU3k5iwDuHWIXJaaV4+5Ple0ylsmJVj7Kc69mkhJBcY+98/7P/BjjwtFHhKsBLBAQeJ
NQQRwTJKEyFW1eeqv5f7JnrsDKvGvwlPAJhdn3aO6BjMzNBQ0xKu/roKSjrOSTltyrRn5GnWzz4k
E4t8AohRBbiAUJBq6jplAAZ6zHVUAtkd1X1bP8l7r/8U153LyzyMNceciCQZ5xenEi6UeapbpuvF
uzxND8OdBfyJvAR22XuibtJcfoOROPtu2nET6yL3EnaMZODu0CeAt8Hz7J4nnveO4mHpt3lv7oCA
7aO2RgUius1kI6nBTAJwvWdSROMbXdS56O0A60kMDUsV0SP43npRbvLYQk+pzB3CpN6NEXKoktOK
FKxqDU0RzoUsMxn1jx96mAiq/BkgGHodRbcAtfxxeBV0wgT3GjkKUQN9LghGbvzNSXHr7x5SQySA
T9W6AzyjEEYapkW45UcPAKihVz2RsigQ7ZxeKpSQTvI+sQ/kYgTU2Bt/GivqfPsOFyUCYQgB9JL0
iuyoK0KaNeSaXRsLh3RszUNV9ubLtgRZZW689Kah4zYgD5Za9RoWvirNKsfUMaAKJMATy2kS37/q
n0fcT6+kIYotgrwK86TjTC/rwo5v9H3nBxcD24gE42vbT9WcTnwlAmAvLUL5UY2lzzjLJAByGivP
wKDmg+XCevK5dF3FB7IDZyK82Ib0+7Qi012LF/eS4XBU7XAlgRW9WlpRr2CYD134I5ZSiX7ONOAT
Vsgjp8qnuQM3Rk5TnlgeIqVj0SiHzZ62PzzkKwfNsnpQm/hhlSdcwufqDRj6Vb5cIKhzmp5AVIZn
4rFwe94iZITwIzvvmCuFj8TaGAnjpqvpE2BLKYArZQjIHhdKNowk1NhY10pPUcWuR+HMzD9YMAek
YBWIQgtgmTsWDXSJxmlFIyg4qu1maKlYaZOFe+/io9ukwZAX7vGwe/o3jyMoa39+le2BghyhE4MP
5+R2XlSrbMvq/EHebYbUzCdnTa1Fi1x8C3HEAO2ijOfluF5ZaimZN4R1yRKBhMKTN7CTXwxe11Ti
hWw89/bEeZGbaj/b0U+ep0obn2FkyAVpfIDOB6Hh+IYSkwO5TRbhKVeAmu2qui+h6LIZm83HYJEf
nS04CwQiCP1qzuJiLi/j5fi2K7CU6riSyXN2as1YntTPqwJCDkz3FNh//ijoillFgPrMuEr1PaS/
wXgEIbmt6UpAaZbtdCQx1r6sjGGdcBXSVYYwWZFpLm90rViu+vP8D+IOTdXm2vByzkSo49fk5qdO
LFdTYezVlHBvamKSTqi+ip/kfF5Ouk2/084KCGMF9iE0Lb9nCenVZlxlFd7h9zk5FkFdeY43ANL+
sJAak+ni2EuOljGDBxOfFfcrVDkGsTbTeHyh65uKxxiiHTl2V1P4gPIh+ad5c1PZIG6cZDsULzvZ
zKtREab/yO2UA6k+L9nqAZho9+Qe1pw1Ae+f/hBXmJ1Cje+bQR/054l128B7vpSUJzf35tGjIUwN
7WmrA3b4IuifwDUoFhFpRsedA40/P7NL2M3feArogG/N8IaTbyaUTqMITL4dabKBTwLWBV/RtNfS
EYN9td7GQc6/iNYhMijYTMJVJ5sh7w9s7G5jopZDZ78p1+3GDrBe4jEH3SFInYsCp6mQ9zKJaxsP
cRfBj2+F0Q+VNogGUKlffdRQfMgFh8HuwxaQ+Q6LCvBvxrUoBIOW9ZJLiIOTZyOoQYdLXefuoOUj
a7s6nJWqZV4UKnje1tAvG5OuO5NMDLAQ8Zl1NOFrKJtqQjkLSA7RbJhR+CHxdTt+/6OAhWfLbE05
b3RxiwnYmiSLKKZStazDvBzyjmGQLsEJALyoB6l/UvHEFNBnFKzcFePIuMcuNhp6XHrT4QpfxuHD
ss3ePMELEU8Wicr+Hj8H4/RBHbpUyqKkpC7MYI3zhVljMTI0WDup3oo2DcsuBtEo6wO+hXQtjDNx
tW7Thacazy3vZqqbgeAa1XWLZf1RNo0UhDC6oSgjCADm182Fz0kMF8N3B1S2Yw1akgEYib09ZvkN
8K69lzdavM3PVuRenvEmNINvt7Q/G6yG2udhVSnEK4M9NFEpMLBzaPm6S/8Tu0NfX3lHNOY78Rfp
c6c99md4+3iX6NDBcvVP5RAwyHum85jxKb7At6wUYH7eIakJDV18QvSUTw1JiaKXUuUchXEnnXNx
uYc0368Cyk/awP3mr3cK+ZK/r+V4v5NBXKhA4+HnlmjQ2L1H9zD1+3xwWjVHYHrYcx9NMi/AXTXJ
f69xawa+V1Kb2c3VrDPMHMvy+tt8Se89fjhceSaYROtfM+xVICkOJUiEw4eWLv+DcNzQMbUW9Nqy
gvxtaM9PbYDNjFc3PT7/51aMhkFnGJhx0F1/TSR1sChYArFoR8jv+rA2TiBEnCTNXyhkisnTkAMi
7eBZdKeaBBFmEdrhnzHKCfQa5MFmMhEZBmy5Y1OjCwZkm9OL3hWbgwQYmw/+KFwcp5IQRG7BLdor
Vuz7vmZXjFKMIM+7yAPqhys/qvG2S+nyAnutvsnoyRCJ85XBdqmf++2BdMINFtf2VMnVeKiNZmmv
4d7L9Hmc3u3Obn6Fxu+l9cMHgwYWLHq6Ny+y/LcsCAr+MIi9DHqo2wPBoLmax8gicnOXB6hxgHr8
/NWibXgE9BceJEZJQs2MHBQxYH2f1x9fxORcsCayUbiuSzVMkNmfvHzA00mgufRB3ATjxM2bSrlS
sZN9ycnWT+lcp/SPfhESVPDOQ6bueXnBSJF3fOD8ZDTwF0MyDiCbCjQwSrjEWc3eyTRPm9GLdM0W
wNssHnd/otI5/3wZz485fKHjgUZrteTZkzmjgp8ivunS+6q420A4ceKdLcReGOVe5ybP63BuIqt1
T0d61u42eGmmrnUfQ27l1Lka3YDPmftFfLRG/VUCA+Dps5cNSjN3LX7pE/lKya+4DDGQ2Y8QoJNO
oZ1Ng7pX3DLgSQjefYkB1lOvA4gbqbzxWUn6dMjcMqUcT9KoWi0LEMJPhyIRE7bWXlUs5eQ+2ZIz
RnOoaa/oxSzX0S+LiZNYDJmiLHJ9BOr7axgY4mgxHIfoDrNbWAfrFhHoYM/MjlTQP0Vf2n/25QM7
C9QNY4INZ9egWv0ZGKfCzQDtH7WbCbtdUfRJ+BK8ELIUZN6xKWYzzTBwgx6gb/StYcdlBOo2doz7
J2y11BWhcUZFbDeTcVVsVd9VWofEcGHUhH1XVcN3sULuaziQuT5vyB3RgyVKapiwONyEU6JoDurG
NWECXNtgYZE71It39Lw67LefO+dfQ3m2msTHcqjwVHTO16wjLmcE1rytF5tKho2PTMqMYIws9LyW
/guuVLnXbQUPE/y6WHwx5B9KgWwIZyuBIdreq86vyrzmhog9De0ibIM6TbEb3v3ePqBHAoOKwmQ5
JEyHJfIv5jxUc0iTMsB7x2J3/bNEKCKWUUC3PJI7h3eNlzof8OZM14/p8PUCPsCT1GU2kosXEAdH
AvhV55q9rIPEEvf27t5NY/vsPVTKpJwusb0lu30ERF+iU83eNFkxUR1ZvHYAvfEo5xfLtKme+8dO
nRJQE91LzHJEBSE38mwicHe88ZQeTnceFPaJWa2RudxUon9S3QTLHWMIMAn58sUQcrhrOAsyfhAS
krJxirhufK/zVjy7Rv9/NkAgXGkaYqh828x/+OcGp2o9tN0Gw+W4gQDd85j5WvNKhFK1VSr3upD0
lFS5f/YzZBbV2a1sb6idO8gLPBAY+dhRNEsVJ4L8ohjHonwMBYLsMqK/ZBGC5TvLLVef1hRKnIZ4
qSJzo3YrLYCMnNh0AQeGGrfNPpGvHUCey++wCCDxgCjs0jvkIAKUce+GSSeBr7C8bHRqrXcJO1bo
1YLdYgyJmh9fB6TDnnFFLlIFD1Dem/GQHaWgVAifjUmxMAgrKLZuuJ6tRZfqFbcPJJwZfHy1ZmEt
tfMfY+6ZRp90gy9Xd1MsY5I0PIgyCz3Jf6hvammuQ3P5Giy+zjj6kHngVw5pYvdl53/XlrCHbAi5
cuBUNp5fWxmHZ3C2omPX5W2C7I7Ul20PaQvAzVdkbpWCNt0LZp96BtwvD8sfpPtkznqIBxGCr3X3
mJmFLRCCZHixEWkpxVMI3iH+KMieax3PJbGWJSwzaEdV4dxKRAj4Rg9/OikGTJ3643ceCc+ZNB8y
xOVJ7v4RLIbpWo7zsYY1Hvga5mlwQV0B6D7OUjfNA9o6N+Q1pRdQvJPbEZ0fYfL9a0wSYcAU3PuH
mnw1XrHUYtSE0eFVILhrYtfgHhMOypKvVny1NrHv5H8IPYnNCgtkVkL0csH8rXMD+5jMqKMWgLWg
E2MdytFHcerqwhhtu7GaGiyBuG3v8U6siVHhRAWRMMWbAW3MGupVtj9bhkFxGjHmgxvGV0PHX4vk
dhXhE5dUloqiesNUKgPNCj6dxpFKmi/lvszLVxdJEVDFUxoWq91a0KLYc3giiBxNftf00VWRmtU8
6wetWsr6pKMqWyJlJlEXOp5t525adrGGPc79zTg6fb4zAn6/3wwOAjkqpg7vdv2j5ArjaRaU6smE
/t0PNw7XbohfIw5cFqXUY7ki1pAx7///K3GWbn+5U/SdgkxHEtwe4QXd/yB2U4wwoLZIV+gYplLr
ERO5XiZfEKogocUZfPqhYsNveCYuw73j8Cyfkxds42RjwzO9SrP06Lk2VLtfUUZAsrjAJEq8H+no
JNU4K3dtB32GKUJ5r6Wz+TQYfa7BLnuK6f0u7CKQ77oGRLJvn5q3hQaq7GLy8HpC3HrbA0by5bSs
B3ZMVZFXLzUEg9jK3ewVJdnIyjXNhgmm+3xFsR8B7/E9mMVkAbErw1rSB93Wg9JgpAZG7bSkYEDe
7tYN1TKY0DGTMVf2Jkulvk5xst2vUOUpI+1MUxZyhDGa5rGXmisRa9bnh4d7oBG7Yvef6xaWPZrf
U1p/oJTlPjJfru2fFrL33zOIe1xUTot2KrwLrGefo+yUbbdN7FpEhtktusqkWeJ6s3q5ZRGuDiV/
mL+EQpuotqzk1vxaqZndU81dMtFHUjzbgL7ksjq/Ob9ANC/yI7vxesASCPgRljAW/uhfcB5nxCo4
IElB9HlS/AYafNwIQB3wbVXAY/xCGuUxD1F5FoOvk1M2M6RP3fRH2EjrLZx10mbLvJlhyvm9Dh7L
fKPVvUEXpAcMF64GlBrUg+7JxWyfjhEeQNaMueAARRZcr6g4oJWjh6snMs2frIpPz6f3qM93FE73
TF2cdzWG58fgOJZtzWydczzj1/LJVd6wDOngV9Qw//CI/79m/nedUmrpOif0b9orI+5g8dr9wRLr
4nmRWoloG2wWTeYoeF4oaTna0jrS71AXvGIFjrjkyuokZUI/O78j7hAnbzqX4Oduoysqd6SwnLhu
MHqMe/tI8aZysD7a1+ZS4KUJo8HqkgHu1dptPYacL/QGDwZuVsrg0fPhVseLQPeeo07utPrR3PLP
L091N3J4d+oDWGvX8vpPtM25QIDQVziJv6pXaU7Eoj6ePBlzG6rWccVr+lGZmKt6yeWPifaTYtCz
Iv4b2PLUow0sl3I2J2Dm/egjkA2+CVTlTG43mD3yAAYsrOTNiGJI0aJYrOpzeIweBhJ4OPqllwoC
WnGexegswq0CDqA40RUj+Kua3Qlza3VQpBZvdt9j++wFGgrSTOptTlC+ZM7CM+DZ4+9Lxd7bMvxY
6iO4RHAt5iALU3oZI78DYLJT46pntc9jNIaox3j3FjPvimnb5iLiJzw481cVQitwUERyr+yWE3yR
6222SeDB9AiktkU5vTZoRu/yjsH6RTw/AB+g0UcEdezPnYHwtcz3UdxCUs7HQMma4C2rPMjvqhxY
Uy756kGGQ8MSUisR1eD64B44NhtB+VNP3Tmu1Lb6GB51AtS+PiiQ8M76LAkCDpU2gbXws+ZUpEkh
mfFNS3/w0iROzqFkHiMFALGcnQujHRwdMZ6A/IbhitKwcvl+aM7XIjRK97vEFh/VGT4oe8vhPo4U
irs6P01VGyKCCc6j4lWiaXJlBShnA0viqwsxARBWVNSbsCkggk0duG/v8Y3TC7umc9Z3tgRrGryG
AOvbkkxecM4TskGF3Gh6onJMq+n8joAfbnKAlNqdU4M3H9EQwbAFlPvWBx+BgyDrmAfbJX9pxd3k
0fm4xmSoMdIMj0Vt7hpEel0Qzr7q5RGx3coRthmfRgUC2Z/PkenGOh+CvJH3LDTxYMZ7sBWfKfSu
KUOZdXQ7N/yncoVuf1kD1xF0CuZdWuJxZGaoKBUiPbil2N1yOlB2Mc79WbM4IeNOKLTFARfWsPxZ
5mVLX/npIrvUSYsNB2o0MKxCM3ySmIcuxjfm+z4lehexrB8TpWisoerlB27vcom0I7+/HwBiySXv
HMX0PLw+bu66JobhFmzQK+Or8qfsz6mfVrDOW5NyevTWMFdQ3GjOIm4T8JF7JR1Oyr4Lf/0WT/kc
CKtBzXlJxSQIC4ZwA51fxbCDVjM7kdEY2WjzIHNGlCkd9/Db224rYMO+58rLJDCnyO7sxPcQVVkR
6RjL+UXDLf2Qcf60eLFJbYnATyI7xdtAVMwvRhvL9cniLFgHN2RXbbfL+cX7oIvIs/SNRwTTQwu/
n4HJuNrIeVtjZ7hzCG/PIpFODjMWdcd2RkYe98r+LMIGxPkqkK+H01o+E7bVj20svofqoAiWxben
VkXxpMXNpSAiMKnWBhlewquY+Pw4vm5s2KCWP6A5XFpHsf7I2QYKJ2fKiVgAlz7mlSh12sWjcw/z
+SXOdmH1HCtu1BHYLOiyPDYpI2NEEqWLj2vu7A1YBZh3FshT69GUALsyKgYRMo/f3VqdcxcxsncE
uk2ZgH5bDTwPm2RkzAEEnhBsVXmBODNVWf/bs0nOm9HzX6ZeOdjjbxIvYZjSCbytzGqd2/9TzhbO
e0mQeVuxwbEdtE4ZKVVKIKobp/U2FFoK5JMX6k4784PMxbQPq3J/lI4bTUNGLSrkIPUkW1V08hmq
6DvcNwHz/qgsLJJgW/9jHxNo+c/BvNonbPhuV3ow0m5jGIlm/p4QEUB6fVgeQy+zVIlVIDvVN5T2
XjQ1pAxfM4Srq0qEyEJqNXnoJUBz1TQn1z73spuUCqUdn715krqLAgQsCC3b7LOJZnelwwAI3WNf
sX/gQippNHEKmEQr+yxnzvGSQt11xv35mqJLrxgL+qJmiVvFAJw03OP6iXZZCTR5BN67yt5zHvd2
S8UixgUBRJzEKaW+vA3SvpeD6y0dCntHLXZGzMljf7UfK2l/G8XA7ge7ek8mH0Hqm7vT3Q2DzQPW
plGZgoqY8ygP4QsK040ooSn+6gX2sNQ2DxpaVyq2yd++R1OmbYNYQ1PbBmmALwo39HUNsP9vVQGo
liwmNkDuL+REhJbxRAUQPt14drm80lU+P9RkwkXdkeTT/PS9BaMfG7HsmF3+XkksLL9/dcW0PO2B
HukJS6A39rpOf5SelENKXlc04XQFAoBbHrWzN4K1X70mVh1YwXfsqzI9diDzjS0MwvZNdFU7ZRQR
tlqojlC1kmd2n6s3wmMMgLPQJDgNwypU0/vCUfnwRruvCUkdDLJRtjRS35nLest+TitbwTh/ptw9
IC9YM7rXeECQUnq3ttzGVtHjd4oSePVv0n3V54IQ574zolngC66jcqRGo3MC9Fj+x6OtUxcL2xyt
PgogrRFDbbTCe05XR2/9tYFhgnsgMCAY/aSPIVSTyWziMB8vD1ZbZB05NeDKuB0ktmek3qgYLwZj
gOxRfSYnJq4xST7jfg+sPJvRiPOEPCheUHNzzot8S52s67p4OaMi4u9DDGFjMB4EQZ7ZU/ViKFB7
WR62J5ZmWBbnXDkF7FqAJTl7T2VWSed+hDRUHxACxWshxyhorczkq0XyCBlfhAnmTFPyXpEE0v6e
XBxp2oJC61LPrpUVs7ygjNG7hw5QonF+pHe3uj/FvXqlS4ST/eVt3HlQcbYVRoIEAz2YmwTUgRRV
XhFLMke6ImuWn9wSArn3vp0xf2DKftYbhhiobW8poQF3lMGBdcAvwBMme78s88BzugRQV2LHKgWJ
S46NLTvUmX9yQzk9S13BD9UzCNU/sJvGcYIZZms6y7lcOApJ39LG1T1JpN6KADusJ0Ft6NFt0W38
/JWTHwsumddRYthU9TmBpZcrTUbuE9OTi+l1Yl+Jxy3T8d3UZb9brRytihiXMmP9cboPl33uZcon
a4ehNyMFxb64SD/VRTD6OM78zMbjSVh0ZPKPw3J31xuHYqO6G0H2BPYVGifmoCmj/fGVYY50F6Cj
M6MaxkCRoXLeltb15iJWgSfMy1bSJ71ejpb9yUBEF5HlEzRhBN0J8yavNE7L4V/FComYSG8MRZIi
FVICxAGrOxb8tg3UZMiW3vrVhvSVtJkjVgRfXNY/6WuyLmyK/jSj36Cj72gN490CGe+PyPbwVfZs
aTjka8LHrAO7ZYyc7wEYiNASlzS2Q1UqHHMxZs5iHoXwjvoOcsDW5z/A5MX98eknfjnll189ygol
01chcOEAtMPq6B9rzFeFzZ+++080rmd/Rg2jPD91aERIpZNOkWXOatn+eyI8/zRbXCgT9VvdH3ZE
/nMjOWMuZRAEVazcCKN553unFcfCeh3Bb5YBpgFktKBqhyu4/rzJqOVqrgNnxK2YjLvxBDKKY9nj
ja5Gpdkw4zUT7V1UeedIrTVh2KGNUMEXoPxtWZt47gLAyErpRlTqi7ERHfMdE4q0UYSpDyzWF4bG
dZTOtE2NympkZ9nT9mEbCQH3K7662JIA6nwp6lBgeIpvSmzv00C13CY3d5dnYeENJo/yM+xEN59o
6arWyU5RdG41LtbMRMHkHAEWH/6UDnHRzB3889qKSUFw2jnsn5RM+x+vOdTkuNTaXNxXkxTAmRWm
SRNQOBzK5HyIKCUFmURn/FfAYvSBNt1KOQBpFksF4pECwSQjMhZVDJHEct32+hJ0JgufVsTcoNAr
c5dncXmja3KMFn3sUr/dKKL4fCcI5DAEfQBNSpoIe3Be8Clxc8pY4OYfw+zaiRnAHrfteoXQW7Ay
rvetCnByWPcYzIhFn8qI0ddA1LR3ckiNrqCDkntBipkr9KwOZE4DDajrxePKdNQa0IP17t0xPkPu
l+gGrkj4jdfJfXGfHV6a4Xmqagx2mdYvpQ0NsQREt1VPqGRL2SrlBO7cPls3uq68/l8fAB9Pn1m2
A2+NhgNJ43DhF2HhBBEWNzT1358gs+uKxbdeXPGaymThJ7DbsfqwQwW/WBfgscnNBBVuCd3gcjfI
IP0/l2W9KsHXLwFej9rkIp1BAYpFMXouyXjzUpqKOpRXejwpPqi5Dr3uOOqFh4fW7G0llUkOKSBp
V3vObHq1IvpbjjqIKFGHpCySolI/O69EoFNORmdpPWQc+lPtsgM/QAUao64KtQV746jLfbuXHL9z
p62ohRzsgEzki18LKd+qiY0IG5Bt/hlJK37GTH7gnd5Qt/kmUAJJbeH0/x9GZweOMa80lyPue9+h
D2q/SxMCo+TroydWOKlyHoGP1Fmz9p8kK8im+jdQ8S4f07T0zVf0iNAcjD58tADD9/O4dnDMcwKx
Rw4UPNX34N6f+fF61/rf7R/UhM0T/Lem9jDQzqKWYYd0gvpkQ8X8E7ShXo4HCZ1plHOZL8e15Unp
txousDmjXCkYqsSo0mec2Q4erj2qzlPGZ85/M4wX9dF2DfiYoWn/MD5NgfLo/Tu1JlN6PPfPncUJ
MN5HzMlG8Y8J8rBMLmXfCxUwYZ3DyYP8U2Y/x2r6YGgxYFNhbyMsv8XAZhPNuq9FmMBjR5cm+fhT
6y/h7GPLtPOlmgxTTx1CIuHunBom2aM+LI3hEUdjaJwRyHbo/7k6XrNu+AlKUVzxcu4Z3HWZzBZi
navX8pBfF0EElW2z2VZHwjmz/iKxfOCSGHcI86xpOIzRV+qMXZsQt+wM6B1xaZZxIdVQAY1f0R+p
fhoNplLZuuyOiMQOfrlRp9PJbn68wtCvwb35rNHdotdsbsErFi5Tcrce4ZrTHcQdaY/ir87BjUlb
9lJb3VlAOkUksbiRcA1GpoMsXes+n8STxw0AwTEixof1Tje4h83N84VqoPvf9hADrLqsQPYO8vc2
tleqRd5xY/gFoeYsj/Bj8xTgeGNlNQ/2YTH+OvjYHef2WbrqA7xHyV/cBHk2QZGrU8L4/J4+Wmsz
AgIsKUSD6G/e4dGRzWNh/eu1imA8sgPjlK6BtnJ4HCFiKOPR2b7+a7uCQc68ysLUjh699Yw/NrD8
3S6ll+eWy+WiO++gFRiJh3pPMvMlpBUz2gEINUSfCtL2xZOtYcqrZE60u8vbyFjBqJ1crVmf65+o
Asc/VBsy2MiCBOeqOCPIOJ2QCG0eZJor2/cQIevgbTi/GnCnrqumH7eUV0DQ8KCB2W6JUlg4xm0U
bFMpTKBeQ7fwBGqRc5YefwMjb/bhWMGM9qSwoaoI3LVt41NgqLIvO2h2OxZo1y8TooDDwLnK/6Fl
8yLOXz5VxuSBAbJsZ+5MtyppCrW/OhyECV9AKqeAFAARw9FtPwHZTiPZ/IzSvCwCWa0STqVpRuDz
hackSkhKVuVoNsWnn/qmDNszw8R+0XSJvitvQFMGuhjd6bBZegRhOogjvvNDkE4AiNOhohKUjZIQ
ryb7oTYut9Q4RXNDJaBiOhIaC1c7SQtipg0pZWhibohfX4KboAtG/U5raG8alYjscj6Oc2JU4VXX
vBVZ7W3y6zgyrSkp6viHPTrYmYwCEWn2iXAYY2coGpc1oR32JH7rD6N9PJFTYyJM2FXSDb0mrkM8
zp1MlTYNeZdGpLBfDo6hOiwGoTU/mLQBZUtNW0IZagSqgbHHQqQ3oiz73CB652WLH4j/xjsrmYus
5QTvXETLVWDesHJToXUUS5MDioqJC7VfRFPOphQhVVoxouypXGLcfmMPOKTtl+tO1nm7SvWwizze
UZr4mEvk91rr+FtMipPwdNz99X+BS0eUq4K8LWXNQZHlQ8MeAIVnpDEI8w0LZO5YeXDNj2uj3+Nz
2qm8Wdr4Cc6Wb/al176YU6BJSvv72v49/J/iJtY+z4mxItM4xEOvQsrvpbPiYJVVAJsf3Ma1nbjn
DNmE5tkiQf40R1OVZSNfzp82B2NHm7NVPm3cHkzg7Tf4EE7SVlJuBJOC7BPQlwT59SZM8HQ2kNcB
Jw50daR7slhpJMoBHWFUVb4thlteuYt9FUG+ugnYBoN/vhT00zwqVpgXBVgHislaMjgkkBwHAA0V
BkGftdPv49lEkJLa+tUS5eBeaQRgKLDhd8t8yEiuodW9SIqrALxtx0eEDkMH/wFIMLROcW1SNsN2
i+kbPqgvYlz0hPiKgnPB7JSB016HSMA1Mja/Er/jPmnpwauxk3XWIpdEgdbKbVK01/eUi3OACkgZ
N1wreJyRel+i7kc6BNBRhxO56vRrpho6ByTsVapARhD7cIC8444L26tNp/jGwL7W5+7R73Gw8d5H
7yw9KwpVH40HDPydT6lJEpuVxuRss9v/DUD5ysiIw71TSpx90I+NOlBc9R53UaoLKpjX/S98vDE5
mUmA2Muvm0q0DOWqZV8qsA4xlvwUGzLDOwIxJ+clHP8GipHpt12MfNHlq0PQoEC2BINg+Iq4wMkl
hp5JV4+BiI/zk0qZQRNAIOGiA8TIGOhWoqmquXcmarX7tCGa4emzimdHo0BCni8GckbxKG3UPVNa
Prl4mABPQDryjg9IAinIBl7QdXHzSIO8k9DYgHoCr1AflcKCHgOVvvPGkOJY2oIkX815PgvjdESI
YPgLM6utOiERtw6hNU8sqzZGixsmAWUCfrxsqN1PA6lFW9Vug5Ec5rKt1E0UY4SYMIXH8QX78UoK
u7UcS+4j+1X2Vp2Ahfsc/PSQuZHxFcAWaN5lYtw5/MqR+wDgIsC91kvp7/B5eoIFWUsjklbN56t/
OwmQASOlSmsY37vkpHQw9fEJ2Q9aGr1iOZLc2/Lh2s3WFfS1QPZvMVXmaIJYg9lD4LW7RjxeZZ4S
Hrx4cNlI/NR1hagaM5ddOXvAzQ2siylMZdBSLFUk30n69nkweQGW8gxZsGS3eh+Xx/CMwHHuZWF7
pTD4sCsqICuJAhK0i//yZMzTMIVyJLq14FVkIdDywhAp+xBVbgQ3BSm6/gcRVn1YIa4BXiR/30iK
wHzZYf0WpBBU6Ic9dGMgx8j4e8m5t9rNuzmtSNxWGwHpx9LIVvnQdzGPfbcwXsnbArrca00jFUrE
z06yeGjoH7X2ydmQTeiPN42KAKHv3hM5aYuwIOUZv7+PjrtZ2qjJjngQN61YQbdxRRpcggUMCepE
qmp3lIilXDShNisvOiY5O2lt4Wh7Wq9nvhqN20T8q4FQc5aOqb2aRaupyzEoBezMEOUDExnS+KSh
TPOKPn/LwudXAhrkxayr559bw65rHo0hvQKMGLwpAeLJJ0idoTpl/ITqupLRgcEfNUV1zitpbAsx
rkQoLUudJjzUW7h1kNH9JDeAzeJCTF/yfIGQxrRS3n67gyxtBHA4DeHuj0HJ1dJe1Ua17HjL/+Po
m1cI5CFWvby/5VQ4nXWvQa7o0IHovoj4r3KVlI4GBiEzM2WIbuKSkn+gDqUV6S5Pkdpk6ZS21pys
KQx8beMkln8S9NT8fzgcL9LxdliF1QRHoJf4AhJurW2/OWEREYiaObkdC7S3mSOVPEfjdkYW6/+R
PEjvMUmNpXlmSst+4fGBBHwB5zCEwo9BFnvDNIAJ93M/88H7Nfi4tCxRtE/5G1wAxCE7Bf+4eRPT
920r8NVGiGkzIRDMHe7JGR7jfoxe4+0dh19r/lPPnKUeH0GIJZ7RRFfHPcXMbLbz7woQkPA2OJbA
qD3sUZgdvqU3rvBsbFDy7kWQxsiSkDeneJVbKOuizpd68aHmQq+rWY3wOuw6Ug+t2KUbKcvjXE6h
5FTtUpVdAS9F3bLdwl9O95g+1Yd5Dvs4PQzmc3yF3HtP9+pEwbPlFfyGJiiC8c2KD7IcpDfzXxTh
ZXtkCbbEWHdnYllwyYgpID3b1y7ewDG4FCJDRnI/KzhSPW/OYZAqCAuIi76TmOMGvaz207+bvdxY
irvBwzTViJeRIViMMSLFNjYFWW2xWJpQtRS76ytLZMwJmDQtSxB0CC4MncrlNoBcKtGKhksvZTRw
3jntlj3y9pBqBgsjjs1Fpz9WOVjMV9ukmNL68Pv4ENePFArrkMNmf20wLYXSiycIPpmMumr5P+4w
4cKP7J9EjWYo6wgRV22jyFEmnqnbXPCRGSmJgTvavizgi3ZJpNWX1yxjRw5/xgYSoMItWHi338CL
oiy9vmOCrWemvf1oSwNvKVlfDMdsZxY6iVzce5g5vbHwPBuHn7l26qLDt2FgkBpg5ZOPSV93UnZz
rx1CAHm2SNITcGY19+pbtVvaAly1k2lkx8B6b5mD5vXlLLrQ5812tT199Eh5QfehctKstEX79fHa
JWeBqIPep6wpsn6Kpbj7z+nRncmdhmCjUOC1OJ45s9XIP/LXoqOquG0gy/ZBYAD+ybSYkaCQp09D
osj7miNtSxFwGtGav0ickU4Nu2Xqt4WQ4Y2ULq7XwfA9PqcpeJfv43hC0O7VssYZ2AvKmrcGwdP9
8igw4X5AQQKNA8eblGNOTYJ7N0x5QIpuTXw7eo3fb+eb8dDxSGW/aLA56DhXZTZ7q7tvWsH4a/0u
+FA7aZBJqbhgEkVd7irUGv8EZ+JhWoKbjM7GT5Zoa9dQdRw8fQpZhX8I2Aab+jMhEJ+2kGcR1KDu
ZkPLN7qjaNDEyMonSktSPmiM2FKPXPhlAlC4SSF3dcE1Zh3C13GBjU3g0yyxhHKjoOoIjkKHHNY+
FuiPpC8ZyvkKQtDKMlsalzSptTuddhAnjsHahf3vUbkq3QSlEBTscH0MhQRTaQXqzIgicumzUpqF
6Qj6tYLWaY8LNrOTAf4dCcRPVZn8jw5phPMIzNugxJ18ChRieFgktG+g84CpZ/2aanWbfBWiBlZc
8bMmWnxUuFYzKu2bn68rEo/jJzFSUmL0pbNilJpdG8HFplZmB1YkwLfIRohmeCt1d/ZgsG+1oX7R
drmqlDzVkJdMaIGtESEhqZrdRKjl06LGfeXz6iJZkhicPVg6S4PFpXj22MtsnRR3B1kMaCA07iJj
h1nyHcz6W9+Ex8Y+q6+qb/ogPc506ZqCyyyE1IEB0J3hntFH7d0dwxfDwwU4C59XGcojmuFj02OQ
e75hG2E2lwrVSgthV09cae2g2ajcWOBr5Gw3k+aeESZByfzEVMJvJrT2oqhEEi9HrwlyqRnzJguH
D+yS4ZXKXJxKaNOcir36/24CG41pHFs4W12F6mD/D2TYFr/bcn/XUUhttIaegAV9pRpoFl/jdL5E
oe1QZsAuskk9njwHbpbNaJVookue3KLY6pAzikEZXU1VnBOjh2+/lAbPPdQ//RWHeb7/mOpkHBOW
+2Pg3mRhBgVdzGyuIUtc1HoxTYz8J7+kAjRHu/Veq35mvxgKJu9Y5Pi5zUyEvf80MHqyftv6CbkD
qmOI0SlbkM8rqudnfK3wcMadtvd9tY2I+3jKhktPOYDwZudX7WpQyFFuvjDyWmedQrpCiqQnIknF
NR/tB8wmVxk7fUAk3jOX6ViQY+yzLiFPwuRgEEbxqV1qkOhCyUuW7IFrLUnYosSGaQvBAsnF7L0Y
IJo3FNdLpj4A1ZfWFYAxS+3g22Fl7byEkSplkuDG1LgcqXelgsAk5cSNvnymbYrbF5J13caNh4Vg
PoZH6BisZlayQ1PRGU5kkMc5ycoldq6+n7UFzGLT8NDpA5w6mFgVx5VDD3j6cBR+4C1UNMk9jRD/
0bxA+d+qYdap254UiJq3n01FrwyZs+IYVTsirwGXHBxp7mWzyKEJF00nHjNHH8t2ZoIJyterzdz6
ovRaoXrJWFEnOv9l9LKrDr75WkixYEMtqcsY1XZbeaiMWfzN8hXcOklOg9wBpqkcRSM/bVNUQul5
1KDQ4P6NcyZxodG7SpSTM6jtOFFlJFrT0XcMsH9nP7FDYXScmieMO8XcPR3C/rvz+NOCE3SjDGLS
4qsVqguYAOrGNK0zqCHT9Zk8bfVg74YKV6g1sv22Ax8iEGIoW4Powrw0RsbznTO1uAO5Dz8U84Hs
rxxtX4hWszOeXzudhijFflmGKT5NY4S/H/mh3pFiLjXvcfDhNDVJSXCt6qwVFDrpa2aYDuqlEiqS
XQ4kznjseBBi5TgWK7hUhD8CTG815QoKJN3thu5RwC1y74xrdRC8F/4ak6Is2yUVf6xop4NSVBbL
kHv68naRvlKQBCcZY4wQI9sxiBvF/CRW2alid9XsslWx9A4AUaxDjLOUAz6/zIE1tZKjroHg3RnG
SQFHYGmFi+HZW/xnvWwy1IxCmAzlNQOeOrX157Yd59ERAfbh6rS2NfzE5yhcsQMcjdKW63JLhifu
nt41OgdeG5HwBRikWk0ry71VlkZyYs79YGgT8l+NYh67i67qlsUeG1O5HJ9ri2MrXoHYkMBV11Ou
mYfmhHNuaU18xUA839V60Ioxhmle6zj89Yaw1YD1IyuHhmf6sTyBKL5mRchq2Cl17lM384iu2Lm5
JV4MpVxPEHGXHLiHusQgppwYAwG2ysof1e5JzkYLqChs5A43Ju9KUODf/VAYFWKDYCm/uxuacE+3
7bw+0xIegX45Hkht0UOW0CFW2HPLfYQ5JlVnXr6TInrS73e3H8b9vldM9NUnq/RAB8UDBog4AmiF
i6NpLImP/oSfgLFBHckSiiz+dRXViwW/05iTogL0KpESWIjRiMYO1y0k/t2M98osa4Pwp5l+1v4h
w/4MFoy1Z1L5AD6Gqx/4unc1GzOkReq6Ymw6g2BUryvUJ9ed1debJj7sSS7bcvpLeuTRz5oUHjP8
iAc0EvSTo9gml3v+s/PbOO4nBeyAztJ4POkvrbqbmzl4JwPJL4BEBsm3+8wYfsZU8VBwkGCcvvwz
vUfZ+BuPRsRsm8K2wTNIDx+5U/jOY3jMWnM2dBTxPmLz+8mM6D90n4g9M22ac+pXh8hyXYIZOVSq
qSc4kqqcIkDPSegloqzeaT8EusZnxpNlrrkrqQFpA7q9Z/DfKHO0nRwvbpOuZGQfvREyRCpOCdYy
Hyl4no+7oQiH+VJG82mg5smhEWP4z4b09EGeDc47XMFK0DnvNPfuGgE4UVloy4ABC2rKpT7oHnAJ
pLzBYlDfoFlgEaRp97/NsQEFsxW8S6Oe47pipL+q4Z/UYq/zZpk05K+0oY1KPCh+4LiXnYq4tqID
f+Tjw3kQgble25h35ukLKh0maCOrz7VxWEn7mT0mSeMZkaoIJXa9JhgLpIkWUBhf+xAZESWvzutw
fxINplcHwpAMa2AVis2gbVweDGBy+ckTn9w9M85sk42/1prhGM4nIeZgMWhUqwNMWFJSf3XlbjbN
FbNjTMEhoFfz90i6CT1gqcXRX2yVE7k3sy1VxI65WqLUyt/7Fj1I10RzxiKCNCwPav6KKVbHmcH8
olsCmXq/6DvzmDA0uRPhn/vQkMeDP+QYyzLBOSAAWO5XKS2pVKjzp4+AxXebTEUiQXOj9SfuJUJ3
9dLodZn3U+q8RssCReOgpJdDBcMrnDg3VJgIrZhyYJtSd6IJEbZXMA86dZeW5abbWc4y4mOQyfFr
w/J7xB0jS3Jq2Ieqz4PPrgIc3eRkW5J7pCrHbPJ5GCIBRQlfo1E0rYlGdYxAL//mMLrmfP185rK5
n6ldW3DSNTWHW4Sls9+r0KPG+yIXStXBBKVhFDErtbTxI4XXHgqynbLeUPMu8rqfTV2bCtUPIAQM
HdoRosS0q7AWFPdZej2HX4yQEXL5xF+Bju3MRXWXkeSlSwD2nCZ8ZlHSZQt6tBg3U/xTmCD6tC8a
OMcaMGUNw4pMgo0AjrdGO7cuIKNS4Pz310kQW3KE47o70f9L7wx7z7699/2o2e0wEjCajCvFXTtC
BmbPdlaYhPpS1Jqr/QKpGLYEFqHOxVNJ2zzx0TZPf/1n6BT3NGP6XHq8eWnIjhNwqRRrgsfYSUJC
0qQFsm5vFrwssiyL5s2CW5SfjMbW5YfaWvOlBcGnKiEECJi6Z1sdgv86ZdMlVAuJcnm3yQ8yFua/
0uHBXh5b9ce43o4bujIsn3lweUzpJpoDsXShNFMKH1sbKyaKCyLDZY0fX2cIG1gN4dIE5ukBG/fe
7KHWZhWN60jcBiHjqoGjJH1W6DJDE0uVBI5E1UeaHRa6RR8c2CqiQw8ztToRwNU4K+EPvI+uUZqT
LXLdVHFP2lL2DcoEGX6L4GNILHLd2bBA79R+fywPWMKEhjIC4nRkeneZOx88Q8F1fdfMBi5MhdXL
zMxMmRGe8nyTQbj+hnNjXFeUgp1Td+gnAhHs1Bj7ue93hCg1+zbpJBPOmcBCi1sqMeWash+5GJjP
PwT73t5Njw272/22bJEmbsLHQYCQy8zR6uy1cTpt4c5Hi5eYyl9JrOd0JgsC46P3IuDOtkYJDLai
gGRBbiz8QMuJzMdVhKzDl30AHNQ/p+265C6oWo1txkkYsIjBWohFZNGakyvnIBqGKBo4XQy+XHkw
uNLA1tK87FKVbdFQp7CHGpE0JcMJxG98Nw03zDcbupDjOFwPeHbvMAXA3S1oRK6wI0F/u/hc8ryn
rgO/ol/XR/S4p8IIXTaQFrLakEl4JcJlY7PlgpWVOjPxUPvmc8i4Pmdjf7CVkxcaapFMqMbjYsxS
+UAwKJ8wqZs7vhR2q0DsVnFc3B+Bi8qJrwhd4M66Hk7aR9a3nnbH2txAWVOCfkNNt5J1CIjG5Ko6
NYfKElWrTshtVzWl6sKYqg2l+Up3u7Kxqmb/sSzNhprTqVIYg+lk6LfjWvunhY0Or3S/Y/K2SNbb
gUwfwhS7ee+VHEbJUtIkp/pBhY6OWd4M18BClU9PEbZW7iNr7BXjAZaJ66+KLQF1EC1PBVgjS83w
O6Q2DvrebsHhGL95FWhRQnJZ2GKQ857YUICuinuMd95ffWqU2gAiMXpZPqhcAEZVJ36U8l78AfcW
fDOfLiBrmAcvdq6C2nQcCJdZ3W6HUAKqV5WUln7ou+5ZjBtBkL3PNRvZYWNknvaFFngDdz6OdpfY
WgylDjy8EwXvgsugroOpeDDmaEug+mxILnVYz3nOx2pbLdYnz1hnbi4oB5Q7Cl0K/jb1Hi//f4H9
PvzNfUqbypt65hEUzWRIqhbJIGOaWMAu8Ifk1kN09m6+2YLZ4/SjW561b4eu1fv3UC0b4s/NHOOi
/seMAw4vCNsRCDEnqImsP+kmFw1Vw+2jOMxSBY/n82WPHvyXT/gzbZcyarM32/a4yIjAX79+G3MS
99VlbST0xV40qd8cz5OxDCe9o792BfsySOL8ov+SCM6E3s1wH/BR3kQbXhKVVIYgDCEH9FZmdiaV
nLbIhLuD4rcdEtSk1GjU/MA1zGdKKuwokGN+Dz+TQCl37Azy4kQQ3Aj4tLLUKyv4guIPIcXPyR6b
3zyLcqGeHYiTsChnjR0jQhDMITpRB8azkB2Pyoc2I2kIHZIpMDG6/ZjjtJXJAkLg5yIH8UeSQjUy
FnMloOLIoc20p2gqjQ7Nf3KxKMSaEhykhNJNmpj8JqagyQ+NG4vkAND6v/HxeI8Hk/FP0qsHypes
0fDgMwdd0hjufcsW2n0qyG1Axuea2sYKsa79WnBPkO2buroYBj63Bew7ozL6ACMdDM7y7+KKxWmj
fpafKvo7nDwUqK36N5SVPrC/ToNrAgO5uYvRABeLBo3zng8MXHelskBSWUOTY/S0AiFA81JFU+Y7
88ByGdeaZTXN41sEtjFRn1zjkTphuZchevRTQhM3l/t+cr5Wk5l123cltN8gUqNZ+ETcx7Y7ISk5
tnQPW4hhlZMI2jnUpITwmLuVAcMTxVJyN7CfFhFJ/aWrz922hPNRX9RJ2yf8sUZ7rAcAQWeCxcDa
emnWgQF9LaWGOnwehQpUz5z0lkdtcPzPbLjm8cq5o4aqA4+cpA7+h0Nl1kZi56KiOJkp9ThvxeVs
gn6f+MHIj/UqjKpgyW9ANwN9EhAimoO71k/1JCDJ8lLtH6jlGIl5l1W2FlttUf1hNyXHrZS5Ywp+
iF6NW/YYEUXFvb19lwr28D/aT2gE+xqSlOiaRjtDPW9QKc/44sTnL4wZaTwIQsHI4dRoBiOpHQQk
SQ3pZm6s4A9kZjZh1E47EWafAaNQn5jZ17+31P+9EKuCAe47tIU10CMQZ4ho7MonRiqk9d4ARNK9
dbav1rqhhyK/FbAbH08UoH13nw6WWTOhne9BQROAgmFJatr0RDSGGocYTJiyZOq93EDnwi4Zzagq
eRQJuYjnqyxZKWz6P5bw5ecrt+Mhbrq6KUCs74eVNWXXCqaUJwrqXpaXBF7s/wPy2TzoD6etBvjA
DmJJkEDRpw3w5koEOoB01YPjoOuogZnYMb34ijIv3Qtr4G6LhR3X9GBbMfRi0gyX1LCDSSsumUTo
pFyRyMsF/xk2MypZW3fvliVYuytM/dMrj6ebtMt/IH9cEkkg/c5GklJ3nW7axOA11i0lTt/nIe1r
A2JNvZ+ddOKETjAD/6YUIu8NDq187NW1ce+LHKfPgy/Hh9QDEUihOnw4UpoHR4ytl+bIrlATh4Yc
6LCObYAVPFDNCtA9nRZj2SAJDs/KLd0/W3WRCw4fhOyU93QS9c8l8cPBMn1pAI68vqbl3ZOePtsp
Om0dC05bJSOkCUPlhNqEiPnd2RQ0ZFUFVushifmAYV3Jb13HX15sKNzajuPCM4+GVUG7gZ7ybOYu
egWKG40Ya10F9RJRwoLW0DyqIlSLvCdZ/sAdc7ztzmfl6JDEc89k+K/DXmt0o/wGF/9N1K+V88L+
yl0j3QBgkR5fmzuiBlNauchytPbHLqI9owyf/vV8d7ysof3BW98z1lSO5N2cs4duSJkpNHqHgAUN
eIn1QfYZTwXiAailu/NqxyuSXPku6bb2c5HwM+uRYnw9xz2dGCJ49MSAw/wBzrx1jU+lJ3fBoEDv
HqcD3NoGhizaVtiqlIhO8KoGChz/qyyBxiUxwSmzbd24sCFzzf5q7mwIBT4/mGaLggfT2jiWrgsO
uieIcgKzFU2/ODVc+dnQhwomp04tnsIh1YKnU+qTfA9/ibiYhN6/cghWKnUWe4+OEQl1qGl2FckO
nA/epZ9jwgy8XYzDq+pBLd6be3lycxS5igl9Yai95pPscEztfvlV6R23OMHLt+hXclU/ez0hEoW6
dfxEcTPAeQOriMAwn4SRpatS34EK8/1Zvnvnq2sotbWfX20FiZQMURXKxnwDSayVM3FMfphBIFP6
OXokzGHO6Vhhuc1BPX6rfIv68MS1w6+OKu6WKPAijqnIzxyLf3GxnNRKeuLsEZHgeDbedaomDSZG
Br0Zc6ueEhWTT87J5dg5kJF8hr9zvyEoS4ZwrApuKDj849bO6qzeRTl5K+ViFLQcntHS3hSiGIHd
3D/mv64KkyRWSr052qYrxNNN10xEYXw99x2AiEVUVhsCSHromWFnY8UGFm5rFe83teKKQr57HKUL
4ZhVSsLuAQKKF8BdNEuXQE3lWRQJ/rwG6BjLWM4GB3g7rAf2ojPU0+oVKjNeW6lOsHeAQfEoaKyK
bjOrbYCUaYotZMUoFMSdyCIQBGameM7R3FInIWPJwR63Emj3f4I/Zsy7sVjkFrV4bahQnmN9sfQS
HNIzTMl26jbSvm82LpNXvnQZatzYgIWOEqi91QIk3v3m9XwbnVYasqk78Ph857gik9PQ2sl0Y1zf
Ou0G24nNVZHJ/0v5DH2/VtvUvTvnj/FTK228O3RAVaWPrYhQ41sg2DezUSTPHSlmz+T6TX6Dcmep
74EBAmBPIIWrs/Q/hnXnBuG/YUCPNPEDjCO5WvxOkmCXGNHL2FjS4RqE7vtWII2VAGYzLH6Xa+17
SahyGm7SNp7jNO8a7I+mYJqvIolYNhAnPDqoWFApAZqHco/5aDfQ4DtwxcyrPvkr0nHQ2RtiK94J
JO5ESHpKtgD2Ge9wcmR8gLTw6UX+GzlFb2uQv/HyP4xxy++LLCBZiwQ0vb+CiDOfM1uoPMGg+w+p
Xz9rePnLL8tirVhGlnYE+EcO0/bPh/TH/x8xbrniUjpR1pf20RI9dkm7wyZOWGXKiSCBGUqBJxB4
koYKc9I++vUymrR61RKUvBqtS7sSeX3yQFa30RIFEn16S88tQKUxXcLd9OLhTk7JV8djhrsG9Ubh
+91Qr0DdKjfl9fnfki7iSUei85AysOsynRohP9ffEBxegDuIxqJpkkh7pgXjorbu3H6XvG9wAfSH
MAglabwO+2/Tn1GjbHanAip4fXGekO/7to187R65s+velrYnD6qtPZU3Pova1NNzYsAWjLw4vb9g
XbKUL10vi5Q925jygFHOYO1xoidcuFGW6rk9pJiHef6e6urNF0/xth36Aul91kPT9Bhc+aKAjayM
iLSoj1/+u0cpnjj22FK6MnnzRAzjNUBAkEyP8V2NP7kMSlzzeZ/zV84HhNQUbnXkfQP9ZkZnhOYB
lceoacVWaZj8Q1jXg+wZtTUvXv7YuMsUkdJOY7tPB8D4OYBM6uE98F7vK6OmQPx0E+bXV/zjzhon
iE67pWWHsXrhkpiBYbDhURIcEVjSWUN0MjJ6WUChxQTzskZpus3g6vUYD4FGbW2CXIWtl1qJsO9u
0gcG/ZQ5qKbLtchnsDuE4oaoJ3syJBTjKHnCFU04SZownOgGcZG9i0wPMSB5V32bRtptIRRd14HD
9zATtYWxjjb8mqUwTaDvJNSjJzayzDqawA39z6FMDvaLiJya96dlkaG2puVwrJmQoUQ/pyoh52yh
cBL+oDXuHAMTl3/+UHfHgCmujtMUxa84k9ToPaqnDeGcTqjtgAH8yKNaB0UXvQgdmcMq+jbtBTyN
2SFimgVWWx4Vg5NAlwp+wkmkDxLMKfteqk84DBHP+8drMbp6OQ5/t08RbcuWyueAZask6JI1Cjtk
CuhzCz6QtrXUe1DKhuUmllAqC3Et2c5R6xLrPV66tHEPiG/CuvD8kU2oBdwuaO+TO4uAg6qovKhH
rU3fA/jMWZdGkwIbSDGaU2mbpbQeDvH90fdMiZic/7vVRKGYFq9BP37FosBVmr84nTybUCQaEr0b
BaDXkh0ypsuzyh7fs9NTZIDhlbfNlkcF4opYCb+zgWXnvKLY1tmUu8NcwFMZrHigK/ah066Z3OR3
ysmZaYmDeulOcNQ5+b8b76iXgr8sOoymfmJ62lmbYtbvVrD65gFfsuIkEPFf9nFTSLkRNUpkLZjd
CJX3DphRUhq7i4u3iGPMoIYu9Ql2VdpyQAFIdhG0dM1oW4yUD32x9MQXwfcMr2K5AbyPKCz/hKr5
5dil09XBCnapw3v/3w9VidwmkfThIq+zEbFUmZQP550WbRFzvzIfzr47OsZuhT4J7JP/AnTHaVav
+MQY1rmYOQ/kgsKCBAgPMUQcVDcgpZBJRlHYaLZsHaZlJ6ptaq75g53ywpM0XqDk1R64Si8zufnk
wtUi9CQmsnThw9CBBfS1OrMQ1bK0dnspFGJ24T6Tw58Sm4xiCdC4lqE0ovMWmmG4ifNn5Fhs4aI7
KLTvaMSMXgf2tewnam+dzxb78hvR24PuBqJdMTio3BpuccOOgY5KdaK34kglrCCKQhyBrjkprIFf
FBovtxZALlYVGzV2hAnVzP01Zgei5mTacAwCGlvIof4qaf2mbm0mZvqywkslEM4ERANsaRN5f+S/
3IJV4yZMALH246fdO3hfp5rwzrKPQgcEmWU1YO7jtudq7gMORKXc1/wSz0CKrPw0r+DrsEVlaWs1
NC5vhtQC8mw9yirkkEhamRFHF0q9eh38kb+y3rRqLPc+Alc57SpZCdM+Vx5/H0aBEEvQWocIAtaa
y8d5YfGtGjvLGiJREimcyJDnZwxoUqG5qU4uoX+eQWsKbEF6PrkVS6I71GVBe4mCVnzTzdRzOORg
wT0iMDGxu8urdcQzd4OyzgGJJ9+d2ZVhhYeaViu5B5R8EM0m1i8ZiGNMBR76p87gxIwxb+nFNnYi
+u5p/vG9XcltFmcrQqA+3DMmMRaqWQjPxtyLJGK1Uuh6pbInp63WXJYnQX+Aauc/fnIWU0QM2UbH
2acd5aMlvXvs0q6Sic2gZbP28NeaPndNmG1oJCvvJI9EnUsDx4cjy3MegQYAGzUbJrWTIQnL4O7o
5CIOthAmF6ZzD9F7oL71iFZHZBQx23gKrviK5g9aAekxdS0t0Wf1qFoMpIigcEQqXHiRPMPGhNgt
n//Byf2VJCyOB18OeOjuJzHObt6X8enlbn5i+ew6Qlqg44xKkoSyB64cqEjwRT4QgIqpTqZVCmt9
V9HtrjkhsZoaCZmpOp9sQ5PUkwJKciFIdnl6VsEPBkWKp5MowVMSsOGrz8w0wOtzcmVSRFMZ1dr7
CPPfPslYigU9lRCRTLymnO899j6H3v6aFLhK1jLVxa8a3VcpO8Zo5vtr6gZ1NrMug2OIr6Ua9Hgl
ukDw9lj2blhjEPCMa2fH16o6Z1AdY/587+iu/mUg+DdV+DE9lH/MKhMpqOMbQ3xV9opKFktmIv3W
kLckPP7bv9kV2muXQAedc2Uxh6+CeshIh5MvYZzysLt6a4d6GDPfYXu/gMQEsFZOlmrHE7vHs1KY
46i/ldnBNYJ2fRzZ9yoahCw4mBHWnI+q/UtMiFCJ2nFM1e+7xbwb42I6EaHKsGY6xbSiu0IIcNAV
CFu5ngQim60BFKtlR2foYVvUnRmxYA3QmzFUy8P1A08c32IDGbliHMe3y7bYB8aJdEdBPDETkdly
5XkrDjjfvonZeYLTJUfTEWYbuFvW9WIP1JmXbxLFoqdqQVkysyOEMaPm7z6b7n6AJH6IlFTNrXKA
erQYbRVggH46ASAs12+quMbmUB6OgKMHwxZQDnqyqfrF46eeOQFpdgZWCfzXiLTJBoTRMVdiv6Po
iKtptwDi9ZW5Qc0TQgNkCkRLCwJfwJOVu2rpy9+QSejCVU97nJ/SeiLynLlZCRsA1OgYfbrerclN
OpCMcH2TbjuWOl6k+seTmPWSqg6jm+e+exAC+56mdMBZUyxJvuSWdnGNTHmN2b9QUq25JEMcuHC/
CqIN94Dk0Qc04fHWb3FM4mUh+Nhm7nJwSzJlPhmc9fDJLaqdhtkcEpQ+pFqsuRPKQ3djfrjbCXWj
8ZZR3ev3VbuufReOao4qpKJ3HeijF7Qs8wLDi6s8SvPn1CK8PkWujrXqK0WBgGdXZpMppv4A14wF
uYibHgpysADuWGS3kKqe7mpuzYv7W7Mc1Y7+tVPNN9oGhvQqkp7od+M3aQ4VwiR9WW88gCIOuLXy
+cccjoVHgbDXe3z3xuefrJOQJt9aGQs0VyCG/vAcJ9cUIlvIUl5X8+aIImUeFJFs8IbvBZARgF8z
zF6GGYJbBkH8NGm3UBJLYorGTlnVaPmwSSE10TqKb+wm5LuXkj2C/egUs+pfzKy4HH1a2Kud6cNk
+GVP3yRq8lZ98giqiWU4pFKV0TZmMGaNENimJt8qX5PmhGqddmr8vVhdlF1A7Ebuq7CEWsDmTsTr
jVGBtbXnSkdDpVOFRxzopRPWHstdILR4KOLuHN5Ezndh/02I7TSoeD+splO8C4IY7Tu71OIzXi2E
WgCaktZ2n4Wkg+ShhiwHQdzbhJ48ZJbqq3sC0Nqz2L0Ovyj6dRna0lPr/TmnIt0YeyA6i/hwn4cX
PRDHpr1eNMAvuZkEMrp3Q6uayUYZUT0lg0G7WwYoks7NyK/EP/k+JsXKyVBFURIwXe8kupHzMoVm
QWj+U7jWoW/3t6dEJZZwkUqVERHzfUaEdLBIei1tYP5u0/jSF/9gRmuCmR2jXxz01FTqzIi4IGUu
ScHaY8pWynroqpSdu7jTazumVte9YKNpbzKz8OGJpBSKjQaX4P9tMz44Peuy1HUn6PU1GC3loAK+
2OixuMp6ydVLX22rYSwHNOin9MIHLh23/BiYK2e5+r4x+i4Q9R03FY3/PEcJdaLcqdJP92bCYQJn
PG8DFSxUCzWLRyaw1KYPCOGK+KHlB+mcqGpQRLFM4AXR1cmQYEMicRzuK3ANUcNKgmnfrppVlXnK
1rpBci1hS4kNzQJIrtdy3smQ4AL/fN1fHIbo+BNgAVfpz3XQeoKNNfwKmVrya3rugwsGeX84L1e7
b/f9RwWbzJ8M9npM+WBD1K4dBoz/Xz9i0YVpEpqCLgBrVau56hAT5MyDPTgKFYg5Cs9pBhsClUHj
U8z9fICgbazgyc6oIeVGuxHy1Tytv2Dv77FXUJ96wAm5UgrKnIEOImVo6ZRG5UpE0LTk+XLNYMYJ
r8Hvat/qEWWJ/BlW+/A1O/Rgn+8J9Gr25o/mBSS8jKsfl7FFpt3BM3CR4cXHR+qO0+ZxMn2as2SC
AFjwzhbmNKAFP/7lqVmk7qPDryg+iMFF+Amuyhqd+ayCAWNdNbj22j08wLVEU/9KBRSYrztbD6yW
bfoJ2rdMQ5tIOl1c3474GLbaAMVgpgPSRi6dfdbxsgJqRTffvbBuhMoq2NWn1q0mgE79Zvhv8h9/
a87y3MUdb7tWCf57ic4Rs4hHhCCqr/q0x7MqKkmKwuXbWhNhzsmDMaUmMPe6aqrCiNoRsl1aMFG1
6ippvIQbHPYaW6q8Mdwv+603GgG2POT3pvTm2UB7mxQqhDqIf+SajwLYrsqgyGR7j0I8wOCkgLxI
iCdqEg8hnU9ZLFQS0br+PgC3AqWz8pIJoROgUXY0RX+o9rTufGeabQ+tPkgrQsuwZ8KL0A6UbnsW
v7L86lxdRc2KMQLBZK1QZZr0l8e3aOdLUQ8bGGNo4xLtUBmy9dn4nX0SskYVF3FC8j6OC5G2CASo
DcF2fu+vN/5zFmYS/aZEBiuSFtEfjjNHLkKXCxwBwiAKkureENvjECnSEcVqZs7C/ZdMnSOdVjHe
9rDlVZaLbQd/ZGRRA7ai1rnlP08CWAj65W6CQeimjYCiqZR2ljsxiOZnet4ZmQuYsmCH1Bpup8Nj
mZiVn8Nt4ckNiBb3b/pToGLVKF7C1kDJDasILW3EyrE4T9DSWOFVDmy25rUjXKqFwKosGXDTXQ9c
x1fKiPvsH+ilVfc7+I4tf1eLag9K7+Lw63UuAp7kxsha/v/EwUxp50Unppc4mcD3WfMvo7dv7da7
wHXs2wCjh/p5sF/OsKqwMas9dE6hXRgeVFD3n3JvrIqwKw03sOIyFpZoc2u3lpTXJ5OFzrz6aJK/
9oBaMouAhmDuVr2y8sBRC6vkBB9FmY2peXUYTKT4LJLQtxe1AsQZsRMCzckJxWzxQcgCYWgy0lyM
944Lf0sPL6l5txU8qUgo/9laE0XJmwowXWpNC4MsmrKRSfnQNSM93pabEFc16fiKTkpNcxwjG3bJ
YgH1rIhFzuH+GWVO47KlAQzeHebRNFq9WiZ5VrN1/CDYWXZejiNvRs5Fl5qCLMThtzH2TyGbwkys
QcWmYrF2G3fPSNO/F5jxnYeagRFP+qz52ZCHliFy7PtsSiwke6wJY8As3/qsFs6bTsCh/Hjmpskc
to+BDqjFFwg/9AxWcT1vArbGKDsX6UB4Hpks1trlem3x5tx+FLjAMNnKnjNvgfBG51s61d4ciOQE
oZ/zPOgIrD1kek2RiQtxu+7y0H9vzE7Eu8F+uShiNTGRp+Eo0aa5KtPFcIH9+WPJRfWS7N1puWW0
/ffv7XE3PG00wOh72GWkiWPqcB2yAQWjv/DLzV/iD/cjix3AntxhaPnkGl+6lE/FmJ19p2qZsGRE
AkjmrWsMy6+FgFocLgCSxXogfW8OKlUrKOVQk+IrRkLUMc3q0jwDfw76y3NsaC28sDG69NZw2ynO
/wxo82l0MYoikbz/hxBEZSDYC17Uxl7U31BBthpX5AbAGI7zELsch2IbQlfImU7FE68FTSuzTK7+
PPcVGs3O1G3C2ih+/lcXgJuTuMZG6l9+/zPW6orWgof/rhRM/LLgR1LFq5Z/L65sXrKYiUtLjO90
OvHu3G8lcIWCcYT2bzSuOxOJvsUQ/NOtn8vpxC6SeDjaOFrVwC736Pdwh1WIHJBdsJ2pWsmAFh2K
OMeW1T8Kd6bPyNKQ5VeqqziD4R1sHvq3VwjRkDO8sAJLg0uiyHiJR0cSQCKM0Y6dfi5IxVd48pdd
2HWHKXzXhtnJ0vl5dgh3BKbFEjzpwyMCZYwPysVBJkmA20a+XZXQukowfxvB/DByUF24tnlUIyTI
BzjP08aEbZTjwhIJHT52VdKKg+71zLTXJZ1d5GWYkJBeRZ+885Rl97xsPxaJ+umLCQfZhMrftE0m
/mvUvAV0xy7ONZ8FhGGc69SLVaHhz66uWb2AONhLToxrYNk5mEC4CHs2Oo7IeeZ6PlyMGCBTiy5i
xrFd2Nkc7iKQKsB/gCTktoMN9qGkSBknfZxl0i2E03aePFBcAxTihzJaFPBzCRz9PlR2ivprbnRh
RL5teonhEj61kai7u3UYBOGvSid2TxaZ/xXwmL4WgY2lEmonMoLSSu2EOaZqTCNNekLwRZ6G+Vr3
Q91kV2ZiWzzcAsUXYn8DjxdCu84DTe7YwhHRU638ma15//bnkzkIxSq+GrY6z4YSQT/LLnrVVkfZ
QXcwCqGYkFkthWA3pl6ElU3uM0VslBPsaTyQGm5Iv3braaLajfxWuKQuMJ/7/tQutwyudfNnpkHL
SYm4s+2rKVmsZK3MBGuETIoiwgT5AqQCA49aEPj4eQXtB4uiV9iqwu6J2JlHVoev8Ifz0zYLl4Us
VtbFa9r/7UjM9xaoGqBiEz3HOHXD1zdhuK5HwAIxXeZP4n/MFsrMWdOwUwC5rm7wTg+yfwI6bNpL
SglnLApIWD2y77RjC5U0e98u2Ca3PjuhaGKbnqkJ7xnu9gtIZpvFcZRRPfaP0+lptPJPxrP+NFnd
glKftI5iqXK/xfiVOVIaZsacct2TfjW+1fUBHPH2GW6/oguEX5d/P+1p/BCUUY6kNiinVOk9Sqna
5Gt5HjfXjmKS2D2HnHR/ZYN27MhdWebdq0JNBtnSAABXRia6in4ROGxNhri87KdhHsBr+JA3vZFT
UVhQ32wB3mEUSOeOg6/HXCcPHtAgzBuo91bpv7VbGGORe6TEACb4FiQr+SsD6OAmlk5xLn+TvujO
tkCtKpQVx38bq152VqeAjInQ7hOWJO+FBzV/4/M59YGmrNgJCdhf9iX3ijzfuWqPb7c3fce1oyLz
TP1T4Ak9bm56Iwm8ovUyY7SQPEiyolrQryp/0LvFZ/DkFyiNCpUIYBvjvQKjvbGIdvQcItRCMIX8
rV+REcvPJixvULdt9pVsEMP7B6O8DnG6ngVY5zmW4Wh2JJyrxI0881baIAvg/yNA/nYq6ohlAk/z
aR+NiFNvDrR9JfXxS7T10nmlSvJd2m5y560rrRcnvCeTM79zyVtAevY1Jf7x4Ye/DjWpWuGUtkyM
5ZclpCzXDhAmJd77l+w3gbOfj0AvY+uMDzDf/i5kQIgkBWwSkbw5MAoD1ZZc3TeSs3+4Egs3UAjs
B7FegU5vpebWAZz+juk0zaWU/pZMLFDW72qIiQtRkf7C5cAjZuDkFOtTm/MWX61ZKJ38eVLhnph1
Pk0Kv76q7ozUCRPeHa3KjmOmhrQbNQDP9UEKM5UnjDfvzayl+pJwcIOxeRC+rhpCUaXjbWZ3lybn
RrymUhxZYXWsjJYT3fCYqnVlUfXtzdlmi4iPvjd7iZr1YUhdsNUGDPpJ3e91qLa9ux20CplAbJsm
7OuAb7m9ReW+kz11z13rHgRfkMiKRXzb7kmyvps/oLJq+M5G2/s2gLBtY93m08fjwX14tvBtuSt0
rmXW3SaJl0XYeFDVSqN1QR4fKx85m4ISlUCDeaLbhFH3Fp+tqRhDusywPq31HvNqHo10oaxhaNf1
YjytSRQ/SjfFqKLDta2WHN1ksVDHAJsLONpScSGLhyq2gZn/MdYnt67YkxbhSZO5f7bwEkAVY55j
qZhzMdQFHQ420uJa1lUv5pIZ5xpcIxwHBvm6vFoTi/aD+NxqfWEyWPX8S9Dxho3kRdrc5PPhcrjr
2PS47PiRFW2QgbHpKBMmKI2hn3r/b73KdQ3W/9Bxa2hl63Jx7xfUyptVUS4aL8xZYIdfH2RgylET
1CXeIsxLLHw30dDFkOe8+YF3SJpFgYohuLMdRCcc/uJeEVxSkjtR2jO1ukRDrS5fPpdczAbQG01U
/dBybqS0SQ3o6ARv9bxLxgJmOU2AbZ0TJvqwuz59kKiDgXxiRh3uJBkv2y/8vgTnI1DqHT1jVbQ/
YA2V12/FupcutT70iwDhfBuE7I6jmMb+ROt1DIAsygXAdZHYcQxbY83Z6qpHVUVxXP9ToX2u3aQJ
QsygUVmsWy93M/OC5gECKwOQNeMJUwFFPOCvuw91lveqGY2QHCKlvzS5XboT3zJSLgil6maGYiSG
9t/W/BSa9/IZAxx8RDOwngVy60CWHg3nN3SyTqLhhLHC7DPtQfzhOiXy5XHpO20SbQ1AKfv9BOhT
cuAgEgsHUwYnCgdWAkGXO7yAMWShVWdf1nxtOslC5jlRcJPDZWhjfytKT06uBIYsvGDXiCA4j7nE
X1vSDkYaHx4n5gctMDzHGH0IDYWd6ZHfyra6auT8fMu0kMjCn9L1nKujuRI52aoz0wlY9CLOPOQ6
pp+HDnJGvgOcBrBXK9LHgt+5XtpFp3Yi72i85rXE6GpgIeOQG/YqGcPcAZurJRpOfyyraVg/zo7m
K2Y+A+e8W4G03w5StKJGXYRht17ktzQL0zvgGj8vwkm1SMw30JZTdJy70zEnFNEB7CdEDfx7+K7w
jhJtGatP52EEkRKSA+9rf02lUzlNTnx7fC7Y0BU3SrEWkKQP6z8f9mcQZ3ZRhnJoEZe8W1ynhWSM
plQu++PDVU9rwbFpq7YHhhGLVaG6iPvegz1ZhAUbnmnu/8+uIlkqTBBchmx0TZfXJaGbdGsC46pX
5V8f9KbhRVgoX8ZrpCnflQG5aQCxL05CvTPMbqKKp29N26XoZX1v3T2g6J4/v2UlOPcG5vpcVWMn
FxarNjY+VsHjCD1GaB23kiTLLBKyTqonhv/btkK6a3Rf8BlW3P1VFcB4T8WmtSwZms2pjlQJ0vPA
vIzIdqLd6E7/dobc/wgK6kwo3OCmbOHITr9i+rWxdPnzYb/44LKNStCECfw5QwoBu3UiPy7Yhj2o
epfHYTm3fXU/2SlGRfDRC03tdqYuNZy4Ncq14FHLFD/OF2odscu/yRTq9DINu6jJe4bEFfLzqRqD
9O3/T1S5SRgfIqdXWTXnW0vPYLypGQi+A9QLGCGHf7is3PiJbWl7MD9LeU4Uhrn3CsB22B25CMbz
0ALCQdIUFFtwnte19ENzcLwIlNEBSGKdm2KkER/PdvgF7LdN4anBSeGHoT8L9oKmRQO8LZuAvTIT
P+7n1cWkCHIhtqFJd7LfCFcTTkOh9OTBldlXLYoFGjO8jANA7MHYiCEFXW0eApjSUtiGgCpUTyBv
QKMfSWVuxBhDG0VwcTKUatRzguMGQV0yDTKM1sc2ZdPDKd4E4xSykjJfMHi1Z5XQhmwXgHuIPnfk
iqCQSJZ5dabuC4Ue2cGZyLvLKxFsxdiHV+531OGYF7o9lOqAdVzsomReGwczn5oBUMZy/erShiYH
leJ5705CLSqoarTm6Jx8bnYnx/wBFKI/mPx85C12tIS+M+QuWgwL5jzDcZjz2RVvA2/xSakqPJ2s
QADT9+Vmo0a7ENNG1GUWGk05E2deY8o3xl/cPQnE9vXclsqLzZP/2UBjJT8R5e6EZ9jb8J9sEEHA
ES8kE60T1OZ+BIXWqt2dpDwdum1UV/99AAA7/nACoPocA+erhzQSl48welRhTTkDzPwUi6MWQgaF
NQApewr0D/o1qQ9Nty7SBnHIQ4E4DyVdLr+q5Vzku22AEvr37jDp4k/h/5u1VFpbMNd7F51bR0Yb
540BkyE0MZdByWyCnkLjaAROsPA8JVnOBdSjAGcpn1wQGPrUnWqY7bJSTu0msRV/8X+TK3FPeGY5
LjuW4ehQ+QRiPth7RJ+spKJh54zOcCNHPxhboGJRSqVUaXgS7hS53+zbJufXhZO5GflNnUP/rgKf
+OqVMbCVFH3AQCJZF2GLGO0c/a7hqXT9MAVKlMlLmErABmm3yKpfvRPtKjyJ/7v4DnHZdPtV/RYX
/T1/0lgBpAFC5J5Vufw3qElGOP2E/dBRKPAWNkESv0RwaU7t1m3sIKbewb7XdfsCXJBO06Yq71sh
11xBRnPvA1/wzJAydxkEbCgKxaGI26BHqJuvJamrFcGcSA8lk/knVguatV1UhoE5Rrd78KixFc3G
BC3+TcP8QRwPlngTA+j1cd6vG/YBtOd6yN2D/eU/eN8KB+NMxurUdhmXKgZOsKsnMFNIKVEa//Zu
fvLWicbF/h8CSWdt7YUDWsTb/iWgdA7/qWHl6LjuV89IiEfPRGcvwzwvnFLcbwGNB5b8D61KyIgJ
EXQVsj2LE1Vc68d1Wo4IK3/fHFykT6nos//Jpco6MPsYmGurO0/rig+JZ9x5SUQ6uYq4FPNXDo5T
jAQz2GbfUjUCiSv6bhNYofoGG/DjnCTtDtRO2pRKCBeRDRf9kvFnGyq20DHDL/Z1SrRRi3Z9ucV2
k+aJmBYsiOFsw2yf56M1i7osJZdP82NS2/8RC2a4QtcRLj2umdMNJPnpxmBEdwodgOF1GOeE85iT
GDQ21NBUTCipgj4fz4+p6DW/vl8ZbCq5oFQ5dEIUuA7QCzScwr8qSP//Iz2Eqkk/MGh3vh05ChEr
kykiapay/n4LtTIz1DOaH7+VdOtX0rZTa7uEBf6Du5vMMZj1teYUlWDqvVtpLRkPutg8ODpExwo7
3EvgvBWfaGyrRfJfVLnL0M5n2Ah+D1M6RBrnDgZj66kAODqb/4OmaRsXbp0UQDSFW01stjJn5Y4+
CNIdADlUke9Fia70tJ685qpnKCV7wkojcENIoDMesX9bhAV61u1hXxchaN/m9jkeJojaaUsfa0k5
Xq1+ibKAVFDTyPF7TyuV8a7l7gljMlgwYCoH1VIJxA2GoYC8Tks97EiFSo2l0jeOZIdSOMB2T3qM
Ho6ThQv7GGv4vROagIEiD52m8+r5o2MOCUL3Kp91S3thJjDLFVQHAyCL9lEyVMN5KceQbFqvPgEG
+AerSxXtanssLCUlDNMEtK6JdaDj9McU1I5M/Z36zVxRmQnqbhvErXRzqv5Y6m9YpT8UIS9Vj9FP
7V6IpLtMhzTueCWbOgDTqMVt4iQcjrGO4Z2vnQ2aCQM2uR528RyyiwchkxAOrh2nMCQUHNJbnu5P
MmSGZ4ehKDVsrP/TdL+GiLvgP6H3HRr02WGLb5lzHhMpxxQH4NvXtRQA06zi0iMCzYdZ5ww6SHdS
aMrSRLGSSXh77h3mjYyFBXKSWmXZGnUi5/BL8s2l1bdK7tASfggyFs6Y1YwfHhuXY5wxHuIkcZi8
B+xjaPppNvX2UK0o5/6UfsTyx4si4UtZEuKKbbqU/ZcTb7jtmVeQEjrEcOI12h6yiRcWbU6O1VDr
YJJGh1RNBDrCsLeTAGHTQHgJ43WWz0JTHCffhQGIkw5IXTBjRlB0fkHW7tUkXAJ1vLWuulNYePJM
5AK0pUMK2mrPaOg60DDFWpvAdqkrt7cwgvRn1MjRpqYHTXOu/1UtpLstp6zFb0Q48r/NN85UJixT
IR9+nSxAxEhzDLiyB+7RX9QglQPcrk5hY1R4ot61m7X6UpLQ6NGTkYjBzYwRbrSvHByZMrf/EjJ8
kQkxRKTyEAo992bgnf79x2A0nEMvxYhW9HtuwcmmBjZdtg9Q2Ez5+sXFDtOkyse+qc14YGyi3RX7
bmKSEz52Map9Gzi3grNjGt3I9DSb58p8gqwZAEf+HDrnpq5sSOEIqqiQ4CpTTL+1FCUU98CgseHl
WLaLQWdqQ9WHhWr4fPe/2tA8tK4xaxB7UWD35njX07Sp698X6l+uiFB+ZGBXl4atvZpDXkhGDv0o
cpyx2VXCzrhNfut6hMu2GtHEGio2XoFI0zs2QA1kYYHJIswAXXDbd/JxqNpqtWCWNcMOzloxEIgJ
kh9aaRyaQk05wPZ9upVPk2uOAiGw/Tb/7blOSWsyXdUTr9DbJqYKunF5qv/OJQWkQ8pXVXQoqhKd
h8W0ZYnIzP38CjYuuoLRzd7NrY/p9kOJ9ce1HyM2r0pmKnOpHZgxPw2NRA/z4dETtAgJTEbSGWBK
HoMwCXi4QqJW8gK4YDMWp9kgztW2/bGQ/rgZ/tv7Rp+wnxd7wroyfRT+Z6liYzTS5UsMc1lVQRaJ
b8Hv3m+/OfkyYDgLUwFQufC7PZikCIoWaniyyrk97zo0P6PO4yXb4jpwdQc2OpPUvTMLOJP7Ni/v
UtCy6ZZAJkqBqMpUDeo3w+CS7zhIIn3IPkYaN9G7g+ReCvWf/9IvIV5Vpz5KqsMiWceVuENgABwC
1Gbt/XxI9spCKC5RNagxVrHdSLUl9D4oZcDC2CflZmRHSZEYNcdyHFHHh9e2w65qItpcqPUrqM3Q
QnBOk+dpz5QMRCUx0O7ZaplPSe2Oi8ft65pqjAUpci6CpVJf5k/xiGRI/9b9l0Gsz8bDpE06ZG/8
5rW2vWI0FhIGYAXJyEx7vgYujaSPUTuParWnHfeKvVxmG/N4StKdeJz88QOqA7t6S7G3rFnPH4OZ
9Dz2484Q0llPugLFcI09CFEFSJYVv0r222uB+8AwKOb2FSXCuYQOtCqUCBcYre8eF2TUplLxdPGh
6wtS2JcDTn0OCWKjLBDNNTTo1+Ti/KSUTTW8QttcujBJhDnJQuvV+6jQ7aHGdsDZbGzFPCVdJr14
U3tR296mr4pPPnZztpfQdBOsjsL2JVPVUX97hUJ9/c/6HzsU2DuEU3ejmkSc7k9KIDvU7qGSidPr
ZWQyOlOObMbDH6fR4k10+08Ezrw66hqN7KBB1IR/AMqun29lTQImpq72qS6glwaoxIN57XnHMo5z
bzIMCS3hJD4G2R6ha4QSsEhWCI/i2v9XxTAZy89vYIrzsgLZPJ7EZm18tnKPmcNAXF+jq4BryoUE
cRPwKDB6vqRYd8BszsTUyEKBQKjVlNdURFh2Njjt75avdbv6k6U8vWRNNChTNVJFE2vtgLee4rh+
PtULyQ2+/O40Ai0QW33udZeXxGjXVvJe7IosaesOC8Mlbx5ZtlVnx+jnNvyA38J9/fAELllEwJSR
r/IJ7tIv4e64c9AeruLB9A/209mdkcj+VI83D3o3FqjY2P45LhK5WumnsrWmI7nAbT4yPLzLVNld
ibatfBatV0aNmg9Y9M1uwKoVbyLxyiNgwbWDm2lyvc4bvWn4WSO0VJEuezNXa6zX5lD/EynlD0xL
7hLctRmqeiSHTye47zb0t+ogfoamLTpGAXoSrpDplVHYuJxOrH0Sp1Uw3N7oMCs2Kv+KoHqa/voD
EtqgJM65S6prNAnUQADZwO+Cuu8C3Y9E5LRYH8ppYDGJJSGs4B8pge3xDI4ssNjt4XUgoYrn8hnI
2EifovE9wLVcl7rkaCg1PlM8nyvmALRLoFmr2o9fyPeBRYP5gXoy9LDehOKCEkOcxpln6u6hPrLS
p4AVBxnqmY50Xnc6aQWjpl3q8OYnwNZ+ZC5JhmJnQpcUwiF6I9ZlJMhESaND/0nFxxgXDQgZBPCe
rptSexmT2mhxud+iiANnWDK9nZUl+2WfReuX7uT0k0r6wKpbVG7wFA2aB0fji803fHUl0OfpRiNc
QqUH8g5lpwn7oB8rl8rsShrmMGBw1zQ2v4JT1LBBgionck6pLPSkmyqXPlH78r3IWP0LAjN1kCqC
cgX0MmVQSdemun+elMx4c79bQXO711OkITiVhPx8l8dFxS8BAb4Cl9Z7aE7Z8/nEoj/LunMcyTsN
bkWigr5aGhTTHBwdqL+ylnLkspThp6STbntPCBYbwvTnEqX3VNNhIr1agj96Cyeqq7wzPI4IdSUh
61ztLML+cQyZJuZ+Du1qwwm0uu9MYzKiwgnQnZiRsRlDjJStq9hAnnbMYegEVUON5Tf+f1G1tuyq
xhh6z3kqL1LFmIJ8jSEwqS7FcGfzLdft9iaJayU/7mw+ZhgoRUndm0n2+UZbiwi5G8BpXvmtM0XM
lTAXjICTBgOmw5jATuKaoCZLomT9pK/1MOWXCWc8B2QVOaX436H4ebm1kz2u0Uvz1Mt1HGvn/7oU
zFPoCgC2f/S7yIhgZ3moTnzEIBjo/OIfYRwJ84tYjIJep/sXkHXl7/a1/ruBsV7lb1dqHgnmc6Ze
0tn/O+sr1M8QwvW1moMUZSJZLJ1eetniFRr3KXJOIDS12UkMApf1i1SGGhSqWa4AkYYEJBGk6sbS
Qy/C0hOEHQPYzMgBbV+GlAIPfWwt/QJoS2sSHb0CJa/884+D8OJZ872hAHhwMop1GtbiNf3FMJyR
fboosw7j1VKvmSiyQtmRDM9sbjL37ceJ9j+lJJ+qPSa06hAMcuHZHRXJpeA/KK+Rnwo8q8c1wQxk
aAyeIoXefiNquTopkOZJauZ++R0MCybUxa7vDUfXpnKLkjFQSIQ3BO9xOD/huDPWY0H87645Zleo
B2qHanglQcRC+cXHpm+Kht1Hh6u1l4Tt31+8danof5AL0a6BLEYGZL3Fp/H2B6IPASp7E9zVdyxv
cL/up2oAywJLtEAS5wi3msEYYBbuihcURa15jutuEtuK0snNdJN9ifNAi9myAChUphAxFBQTWuKx
XT1lmof6xbixLKSIgraX93fI9NeTdn3TJN7YqTqx0dslDgQhUW6nhOaTwjGGIB8zufLNVLBSVBBX
KlDPPHJprg4KvW+/XKUbGAAkARH4l822w0QHYZfdHgzf4HZS9ukxgA5VYF1QKmvZGzPuermPRPow
IgOKy4qkxtVIqLamTJgYv//KMDfgYv2YIITjCCS6uQyTnyS5OJZ+EXLun2aDIoFtdwon7uFRSisU
MiOQAQV5mHwd9yGZOBEAaedudQaZR9xTPtF6sGT4OMLMXzEZjd3H1W8aAeO5R8ibG1CE8rTsp7eU
EbeVaZfsUrbmMvA7fT3D7SWHXF1GUIbfCc0jkqrCZ996BocGtEugoBArPiqQ5WNoXumxQ/uhJDtl
zPUq+wxvEXHEbt2ZVMMZcp1Ahi00B6vRLHm/IV3TcF8+b0Xl7dusF7bkPaOXdEvb663jSpv5+R8U
uBy3LJMIGc08qjhnDM7/wif9mtZ8RYxZypF56Dfr/sqWisu0dXgT8o0JMeRcg/zjXU5sKnumsZ1O
Myafcrqsm0HqPFea5fqnz7dAH1vY9CPkBMr3PcEj+cO533AQVE8tmqQwezUj+UIZmH6hTkgrcfwe
N8G4Q1g1eKO3MMSsUkzfV1mpSeTezhh0GPQKSqfcuXDHAh4D70rxnXeeYdUoZVop5BEPZrHPLwAO
kFNE5cptVSoC5H2VagzLcfd7KXP/nvfpIfOgn74LxtyBl7MnPylBcrlc/l5ZcLCJO9JWRCCSpvAI
X1jKxgoPgvPJvy1y5cKmOWm7+LvPaBiAz/PGvP6/U9xvpWpzw+1SekVsd/V9bBiXiWsE4rusxjTG
Luwz9eNY7JNm61F5J1tuhajRQi6uU0TVmq/KtAqix10TgHk7U9Hh9/Gza97AXeuPxsqLDocOWv1d
PBi8egam3mVYbw0yM8HdfNiYRLIjmzVLbTQd7TlsfDd3vCOnV0qcTy3oPNCPxYMZL5/EUGXysp20
1x+r1Q4p7RZ/38EEfhPD9ABaVcNlmWoFiwe0VfzAcFHa8ymF+gszyOVnxoon3Zs4i25FzuDjwIiU
Td2V00N4H8T9EDI2/o9pyrY5qU9g1NTw/uSjh76y9q/io6g1QdyOBm5FY7A1vvHchMUhm34ByXF6
UXHMTRoIHeYgHGgCBEG2mma9PmJEZFS1GqxUTdTtOVL/4Sd6ZZaW1iXaasL1Oq0laSs7vokTjMe7
8hmnZB1QcjL99EHAuMra6exDkxiziPBkzJWXQ3wyA1I9lYTR9CHoY54Y5MkDn0eVWuuIP5kM65N2
LPxTfTxJfg8Tnz8UrKQV5Z0/ITxs4EGM7VB1lQ780ym7uZsfAq5A9xxZNq6SBR9UbEHqho/vf3Rz
tHwENBLffYM732B0aJUB4UEgoJ03xEsIRIJH9ysKavcjWpJdrRFD8VZLQcPHJFy4TeU1uxbwYumP
b679caSF0acjpLITJWKB0KtmInEFevNoLZC4frh6QuVmSu2+U4LdbK9rjjjBE7EqC0Te/SwtTpDd
tgCxnQjoA0wmffp9W274ufQdaxiHBLRFmL0eUIthKzj6mrUHZtXGFW7XXmiLgdTOnqniapy2Vxkk
6MWNd5M+48eZFLieH0Ux12RTJjxX5kxIDyfO0mitLiiiO8CZ9xbZClrQiidmkQZaeTakyt5o/ymg
Ouoc2KQ0Jjulvip5bmstyz0mR22hHFTkI3A3x5QKBtg+lHWHQZ/vW0C69C3RB2tb2ccxD5JTC0os
xE8q9s745hkweNHQLElOgwtG3X2ugAgQV7KYk1exU2rSDAw3k6RF4yJaCq48SRt5Il4EYbSZDWex
h/dSLHQyfwSYG9MEzdFUAuj042RLQ8tJ1G4BzZ8vucZK5sAy/qdPxkJ0NvTnRpK/HFUdTqn1hrO0
YAOBUeZZGPEfrmi95pLM0H6mu93nYGHnqUSfUtKoxh5iCLslA/IZS2+JEQwhGRvoxlIESYRoor7U
HrRsuX8qx26htm2En6OqcvLOsaYuQonsngIYlWllOjKw9aSX9HygHIxIdaiHSqa3nyZEFYSMXdqN
vG0Q+ZTYTGnwynS3dmk1pvsv8bMQy2m1uMtocmIi1EHsLX3zVOATT7eS59xGSSxjTVgzh35QkcLU
HxA6FnB2MF1uVUuN+RKCVjpgO3DLiuqRhCyQ423pS3g3Wz+/3sfNnHFdE8tQbtzuG5kIr5TcG8+r
kMcU/oZZtaJU1705mX1K/TvyKf0YEaiIpuD9YEvtK+/ugMpzAD0ezIoHKzvk1U6M/SF6PESGFpzD
fMe3CtsmpgoO3+u3sJgXwcVbo75SNHX+gF6cfH7uYUkLsvJqzZGjqiqBN5g4Rfky6lUF0YyLB6W9
B8QNCQH1IFZBUF4Go7d6kRr1dOAUz+tqXTEE7G9eTHKK3UR0tyZJiR7chWe6/WeRqnzyG1CRsZg6
v/JPLfA+VEef5r8YnoSjPZtR2FtRKqnC008Y8S/4+YHmm7AaMQFFsnCduKZn8RM+HlYlvcwZVyyJ
Lj5WwmkhyD8QCQ2Za0hMVnJdjQg8+MRhXOira+qTK9m2ZWUXaauL+OrqTioDbBUGFIjzMfCNi8hC
MfmFAbfsGnzDY0S2Ngvmn/2vEtl5jr6Iw2NfG96iGbANXWJnCNra9BhOacbdkHfjBeqh/f6eJ1vY
kVwhVZ133vp3pHxU/oboKUOW4Dtea3++flClJIIZ/dYYPAgJWMhJokjIWIll11G7Q8qHhez/VXTK
DKa09ukTnKTqm1MibtQAWGg2o5vsdrrwgtF/YYvsDVlDFIhmclNj7+vCIFZ5EF8ccE9t9+4Y+XIK
Pe5gxLzBeWFzCp9rbES16LWuYdoF+jmRPvYAjYyRlSQ7v12KD4s3BfcEdRwdHUYS7Ck+kWqE71Xl
q2FXnsZMaYaiOl3Ft+Xfpzkddr6YTio4F+3vMeGC7QLpWyKBrlpnD39OoM6pQXEcquyxpdXFGwxj
WM2wjzOVo3gmaILqhR+HkxqDRBzSoKAczyeoKcrG054TTTm13b0se90Y4S7E+a4xrcUMej2wvfNO
u49Ck6KfCkn1WNXGQj1loXa8Y2TcoK94+qmhphNFFLIcBBffNP6kPEYLuJkqM4Q6UyBtMQoZjx9A
SFZ8KZg+6m62pFmHsxye5pOJBpgxoyHCsoSPDW5FFCNncOadYg14LwhHIk18QTaDur2wG0JV2uVp
y9eFriMvwhDiulhQo+o5Wt9pCFhHP9T/Lzqsl91NGQQM4AfMDIpMqiYk6DjlyU4y5vfdmJDnElgt
GnG74y3b3m3t/h5h93GUFKWgu0vPk5yAINZnEidLLkVtpCMJ3jLiVvVFVksFb/buibyr/7g88CZW
5RJVM0h64/eTK3MVPsEyez9/VPinJgXOK40KLcKCuBH1OvHs4Pxv1OifMvldrfvS5b6DmNv8rBps
zWImVc9s4RB4mjGJR36L++r1Uhl1ysLWm/GUQHYtL642k1BqWYWBFdHDdykv7KReFofTs/0b6ovy
V/uMCUfA/zWECg1b04XW9LRLCrXnFj+qkVEgavvJtmKRLU7U1vnc5ZwbE03muhWjKQN8bGNHsfgM
3Qbg2W7zgmveW0cn6pqevKqvro84FgFpkbkCO4Vn2cLrLxKffU3EmauJj6EiBg2bYGTAB/YheVnq
y9GVT6lvXMklRBqAPeqiOmHpp+GzUg01iQ9UMCN46Q+3LrCi/fofRdfMcz1e6Xz8WMNDYohnrSTy
H9KtBm2wt/THKRWUz/H/KaOfjOzFj/X4Y1paD/3NEDbWEQBoaUFNfDz7p9VoByO/jYaWQ4RpngV7
NgpkM7JiVXhTr0fjaXlgxojTszXv/kz3PsLpnVfBNjdCXbYS4IPuxPfdBMHOREFQ1JyDkUNQSyXs
iHmQ4SJ2y7Jl0pyNX8BJ2/1pHwm+qqasQnuxENjdPO8UGUoDEIsyPeghmUn16SIJqLK7QxkRBZ9/
1mRccy8E+frNGgcKA03DBLab6aVDkofisZ2FC1R4uuHah6cZxEh3BmR1ORrzI9V91WWMAeDj/nPX
NN9xFxhKxeMlhvnOCFjirFgfDF4Ej4jprDAoDS3ph81vgNNKqKNGVPeoBSnNcyQLTZ/RelXSry4b
OXcjnY6UMsqH43oaVyXzaMtzVhTaELsRUUF0gFJ17EAd/l4fTeHolmtoy8VCbcOT8rgCwzBLbjpx
XgeME8/t6bsV5LxBdo00SuaEhKJRtA9CuVXIal19K1Cnxoz2irzR2t9ERbLSLQcCyRxiFxDDef4G
991xhFokIYomfMsG3E1HUQzUFdXdEGKgiBgcd514CEfMeimBwmMnu8mgIhDt2OzFaWRAaJezQZUg
I0aquanSbj5PChL6RP3r2OuOpF/+3XrsqzdTAIGKJBISSSfN+3rcif83UtA8l+a8iZQIdpKy5FoM
ViKrP1C5iHyAutdq9Tbx5LwSD337U8ryc1JS7QsC8w/egIlBZSFaFrZm2bE5BWxYv6XEqU59uVO0
0wIqqEu0PXULO1c8f+uuYZKoIV3R6qmH2AlLhWwazAhfC9wHwX4xwEmKDep0kBnTqL5TLQRtOBZO
7K/SekSMVdLkvpb6u6DCwvNEM0E31qyOgCa5WwOIDid+EqyGLHpN/5gbQqHbivALAn1NgAYmjdhQ
o9o3BvwbTGlrDAFyrqI4M9mKhNtoZuPDOd00rELu+xRqZjFKyPoCAZ0/KO7nf55pJyI52DX6vtly
s/HZpxuaAAltYpgaGLorJPAXLgkGX0nd/s4Thvi3NgiGg4VNQG7/3D6LztUoJAPCTmrZI2/UKOey
vry/EP6vzUGnvqQPqiVxBIHgRxjIlOw2Cs1KeYaki00qSea60ACRffYZxC1GgLGc0C0cJEdNG7ZW
J6dxsvYJvXdB/7+MM58PvYSkLs/QzOcRrbA/kk9B0oKFv/rHLtLCCmBiuzmymXDaM24ryvNIqcuE
vDOxzbduiC+6WHoHsGlmm6OafPng9o9nmviCmRW7UMoz99IH4pSaHY4hJbAnMli3zC2GGkqQli+M
+ht55ZK/qhLG5FF1fI5lcDi9szXpsDYPcMwMcougqEYV1WxyrhnfvRs1dMikO5VD13cT1CpTlB7r
nWu/qKgMflM9hmN2NOvXyfAO2DdTVoWV9NeMA0h/cMagqDxUlOivvhMwPvNGmGE9bo3HChdQTXft
PqeKBjG/7gxeGkuSKOsz2dPvvNBLhHS89YQTiLS6LNTo1M9e+ZUkV6diRGhh6lrIuNTC7WAbRY1w
lPBIoL/G06YbXJnSRFwN23u3IHSO0IIKy36vh4kRAvY1OWbCPSQimY/wAwRllBbTaZ1/ffFGCFim
QRzZKpLivRizxYFK+XjFKXFbOFMLn02PtrflB6MyRMotJw/1ZVgBFphINetUjTl8qPXUBR11XWAI
mq2OTcFj0Ky9iaFbXbcCAlooEkRhOw7tk6Ie0nuH7qz1krvVtD6ZaPDmv5fMi+c+t1V2Sv2Kpr76
MQq2OVRSni5/0YUCLt8lbNcxcDfeUfeVOxeBiyMY3qHv8uDPFybVOT5ElyrMhLbdUhobNCNDmedr
YW53kRYkYiteMGCgp2mAhRVVedUZr9aNa/JAR2owZdctlhLMx8H8OpEKNmahgPBTzPVMiD8pTrFb
6locQo3cqb/jfmc3oo2EtDVNd7SnMFOn0uIljKs4bFFSX21cdugxvDslQ6BqBCO3f52Ce1NvU+vL
pk9trQ4+JiKhEMlG94EO/XfK0EifGZ3TZ6HtWqnu8JYBEf70zi9c4vp0WY9vfWEbiyeguZvPp3f1
NwJKVs1wHm5nUA13UGCjTk5yQQkx5Sdj7+9xSlXeEzhvvLs0borZlDROqamIqPLCNKiojqZxAvpX
0ezZiuxdOmxR/SbHkNNtdpvQVrvYe4kSVFCSWe4JGreigSpwpSgkU92TFBp2ZLtAai/JvkLg+ROe
vb694QORAp264za1mzIgTwYjnZAJmFx3ErsygE4sg1zqmob1twqOgjNSvAyypFQl/s8NoSgy+4/H
HmYx1V9iEzOZ9ErQM8TnHrMIXeiyr6fOjo5zVNz9KlZyEv4YZXlyMNzli5rmX9zwt+sqkICHE73H
j6vxOqw+of25hobw+fB/jXjFvz4qG4hMqNx87dks6/f7n1YxkS5oo/a+1zEWTfBFpQQC2qQuRSMb
r+/LB/9gadxjAlQVC6mkQ+DTnMP2Yq0OkGiVPBIn3NMm5aDaqb6P6mM488TLn/wBJDEF+GCNfU+z
SXcdrboFqOBCt1lh7G1mnWuqXjZnoeNlWP0qhhqkKpoO3I1TK4NrTBy+Xb9C8DTgq3SUIva2IwZM
3q25b046OYEokJR7QNOoOGjbwKEDwFsATP63gO80LR8SZpRcFVHYXiyl/uR2OdGIPFaRan58wjjf
03Bwf7tK4NwkzYF5mmFLQ1IHAIq6Oer1YYpj6nDqSENpzqWHXnokupZ6RzbbCyajz+QHu9sRBxwx
2LdaDMh+aHejj9fjl9oND/JHm8I7bQpPKJg+0FVwZy//LpFazX1SYS/JgFvw7B40cYea+ZTo+j4n
oD1by2KawxOknBZpdmkjXO9pE0iMhc+9ZusPrNVXnEb7x0iOrV7tbIaUeJvczQCGGVg6s3XhxumF
/YUqxD4rC3HvZhyCe6sPK47o0NEQj1dQl45QbK24pczxLCnVZg1s0DqALi6f3rJWE59UiJh/OfJI
N0shAcaGdP0l/aw+r7duRO8vyPsAMekJ3/3cv1+calkWDTG8GKdlBhrrAhAFhbnGjADTimacdPB1
Szy/rIylxQVK2lhJYx5kVnSckToZpYkCF1hLVVWurIr/yb6fxSLvrCVyZ3BrFEIN9uCLCEkviXRD
QhzdhFmm+sHVsfx5v+jFd+0kFoc5sec884gOVoCfgy624pFj7CDWpN1haigBlVugvv2DTcgfqrZu
QfSrKx1UJ2EmxDJcPu6BegUEjGeiootJjT/z1qRYeyYAv9n3eqMnJEoMOh8DR8m8TfY6Ocx3myPK
q/7asBduiOFyQjgvDRRuPJ16QAVC683d9qDwAFzPz+cFuWIramvauiXVJEe+YxKUI+vee9OGK+XJ
LCBZJwmp08fIwnqPKO1RRzo6pd6aiIWTOpkHOaax1Rd5jyw8eOdBacGw8NXkUB5Aj9gouNLYjBEf
4CVGxMwU0/0orO1u0Jw/MHEKsMpWuyajrrJUoMo9n7tVpp1H2er8fsse4DpQEMSx8E79XQrQMXIz
08gV4WDPp8NgUVqnOnPqUlsDKvey+f9krjD1EUmn1ETkw6cZTpa6ixDv+M7DY1mtokIvYIG9da0K
7hiydn+U5x015oEkyxVdPkeITfC92NRsQa8zUAZl6PZmcJhuo4gWp4AITWvN/A2HZfChDpkU1SpP
z9hSFGfpzvWuVz+zSCfLaXPhgD6av0POp2OTR6JgjojsuBkQnM4vr0laNaWJDcHftb4CT43YHl6q
Mrag6twgeM/iWm9V9deiD1XBxzTPkAuecgsYOMmbS1G+GStd4t9S9ebK8xlNMKMv7S2K3SDQ0PaR
XXCucAS7Z9U6TVfo7iPjauyINEqHc9VRFai5qPZxLUxbcK6Vul90Pcq5eq/tPMKSy4DxUASc4QlR
gIFYnnWBu7NvWUcSh64JXPYAFReFnuVEFoabXA0uek37JFdH0uwUYYDY4qDmZtbeZoCYOJgjuAxY
p2RzKhM1cAIUJtS0kH2cucp+TLxjTq3KzSiDQsrUYbNY2l0n+XkpwVkTh7sxA2y7Nfz4bzr/YYIZ
OZ69d683698dzeCq074cRa5f5YbVxJPCa45fhHm0pand9zN+KWxhdPByfuYX8E1GPBNukf/gXzH9
L3jlbz0ZHdqD6lPXva1EOXZDSLk6+Jg9e9btaa1P8Y4Ig+JxLX6VCT8XppdDEoxf4pTNpGugRoNJ
DxOss8vgwQtRAR71gCwkHqj6SbnTjb1m1pToomULcefUCpmfdOsVwDdmwN2FyP2HKNe2IYvYySEv
bsicL65W8b9dyPBZ8kooeDI98TheS6HI9o+Ol0bthcO/fbwk3dFNt5dnwDHKNM5wx9fLK2uSKkJb
lKlx8+BWeK8j1/+hAHgK51o7LGnfNrPRnGZ1USTGT/xgBPNWhz3iI0HMClt2yOYO12XThQhrWTuo
p5ylNAzmhgz1cJD/AVmzr47K8qBTfmej8Ae284XgpQ54OwZqHzdb+Ke/pKD+4ql8UWuIWcoZBMIh
9VccKmMWsrZq3qxAUYD/l7Ypx6h1rkHRLGu/TaHHrVs+TWs6HJW8f387ZLbUaqbV7BmQIhKBZVYB
NvTZW+25jDo6nULLAFtp/y4200l9iLTi5GWXkooDoek2OPh38Kx9reJeKLkhaW4ugfB2Qgii7t2f
txP7wj1qRxiPuveE6GtDmwMkiNamd+gKzteJ3aAx9zXd6miPhN5WuhVQTQRpzxR73GM7Npixkqw5
o/89uka1GRHe2fg3d9ORgd6dJ64QC2tAKnIsQ6gM3GqMakfCM11JeAnyaf8SPuQ7GjrqdYJsTGPP
BoWYETSdgGvBgtRZhuXWoVjgHHAYkUCT31NSRJPiZ/0BgrKfBFm0nmj6EA9yzbCSoLBKVtVplEyU
bi/tj8UMS9lDS8jVORoTibIugPdIFjAw3EnoGWMzEA+mQz7jecLqfrl78WkHHAE1GVe5yLEih6m5
/jxNvGASO3bLrxdghmRBymsuB3Upb3NP/k1fqkq7X5QMSEbLDfy2v3AiXKnKlcezggQ21DPbmi7u
3wwZ9eMFk65AyVDo6YYXCToriiXp53O58e3P6mf5NRhBPpPFcQeABEFHwhLYVPOrhuyt0YMIlZoj
ZZ+FmgxAh7PVpz+aqzgl537qLpWRdx1Hn82wHDMvH1ke8a3eqwDiL3rmpp8/tlAOuT4zNuwgJNX1
tMLRb9uzCEt4qNfMdQ6Q1NeUrBRMTlF5abaSBoR/gLzsLmB3wbghxB/PPcvfewLDbVL2WFEONF2Z
03uPC0pDltQVenZaL+5HXJU2lDdrv9a6GWJSIh59qsJdNxgnFfJnXkKTwwo35AdO727KwqZZcaDd
/obMfniQh0AZJcCpoMk/9IpdAYAqpPkL2d5aa4xSXUH51vpZ4s6CW3NzzdqYJIDkwqToYN9dmTBP
F6hIpw+7MsZrIAEayXnFbGD7cs8b/vP43v2WpTneaFV2uBkHOWrAEm2O3QnG9msClACmWIAd+J6U
TLtC1ZGKOH0jvyDYIWyZthom5v9ye5Y1G/VyE8OYzBaCnULTJxejelaeV9bI5R+YbbKRsjx2XfEq
6amd9N22VK4iL9QP4SyDE3Cyqpz6ZJZ8qx52RO6m9Emh4i7dRSdouwtS7tNTeQrFHcUvu39FAtrc
r1U7Qda+RifsedduK1o22UcUMwBcOngfukSsmmY5q/u/KLS5spu+ThrIWbj234mZ/p6GzG1+1TQi
6czaOCxalJk46eTJmMQAoBc9ft0sKv3QiKhvvrRGbUhuDllXCbtwAFehc8Hy2MMIWuhVUQd635pV
XyCEi90ObQgk6OsL9zRrvO+8PfHM39gWM0xC8MtOSI/cO/RSMvWLntP7Nc0FK4ikEIVF8zIQK6Fb
Qmw70ZcGf8+57VbKYboWn603DH8F2PVbRSBk8AyN9c5d1+Z51iXBAYqUV1UnfAvGWGp9fCT1t9KL
zQHmAuxUJ9gNf0lFu6usGSm7JB9RUJ3O9nAgRM7o0dN5eWJwREnsEhO8l2vse5mfYEvmCmUpakLV
t523gcv+fnN9RD26zjz6lvUO1q4gKl2ThLz0FOnjNY51kM/mMIB2yalejblFBamKQ+3aBycJ9MJq
q2dxYG6ZN3PLUQjgb9M3amh9EHDbpBVGsL9aZFgY8qPDf73Zlt2yT8nZkkbBBykeav51YYbt1DVM
/TycRBHelPltXm2+tw/iF+FaCyrHtgxcE7N1QKtJaOKvW2POEeHcphrvfJpufzVDTlpP1CCVlfrs
prOmeivFYALsrWVlr3MbGiV009vKSeFkm5U8GQqB0Jx4jp/Vwls4rFVeIbDtnCl94r6U+bEvwnlL
TIuIHktZO+3l3DJKy4Js2C5QJtTWasJawhx0FIWnIbd5RtGThxfbM8PYqWfOteQwGL6TyFumrivk
u2Q+QxAO6yLl2PWTcw/zv3YiftW8VcaqwynnBVYd637sWk21piThWS/132BHSfqAa2HgaqI0Kdfi
+eVNNWaUdRjZUSQoNyf49MYtASFhdNX2fWHOM2me6+UOwztc7GGGQrtbvV2IBE8yUsmo7+A6NZwD
fYGtrE5kwd7ZcoBRzQEbwsNSejleg41NTfrfm++NGHwNS1E9a8QotBgAmUeliRIkr04f716LQt/9
+u4cEnowebKETZ7EdlqzkIE9Lz7a2Ac/evNjS3gQ7tDaDF8IiIIHiKiLiCscVND37sgQRbsxsfRQ
oqEAAIcFZZCSYPLFuD5Oi1kcuWS6lv7Oji02Cji/Cav3zXhaScvU8I76rcxVKo8LBMUbifiwXyYI
2MkbY08C/1D3s9Au4xEjCn81YU0bC1j4MFoNRmpBl1NUwqXf925o9nXMoh2WvNMSyJ4NCwtkWAbY
k6cyLiSyX62SJVd/3jRvatptfL2nNm5KkVHnggAzyMA++LmFusr8k3H45pUcuYDIZ8MfW9DkKINS
qsjcdd06UjaaQhhcRU/uoBT6QQTHFgbHcJK0VX94RIBe441Tmgr0rbrayj+SBZBLpsTqNrPFSCo5
1PGn0c+tzAWQoGPdK5BzruAs/2U9cUkXY2+KFTsYiie/WorLPJsEwyaxECBHB/sZd/jHfRaZ/tX1
mNPwpMLc1x0SS/viUHgSC25ezbKc+b7WAJpF5c9exASmhXubLCDSETidsVfDZzO4c5ZHYIPBOFUF
9yrrrNJM4D08nCOrAJTFhyaMIF3gW5TsL+MWduyoOD5mPv4nMbmtPVGHwF1LiTZ0O05eWeZxyIj+
NNvTI/NMVH7Ogid9B3bSYKh+p8CTBxceMTy0kBt22pvRuy5zRAxGJ6iCwwCf0BDQ8YWwxunaiE0U
9O71Hd+lbL7RcEyu4Lc70LPZEyCRrFzFbixA7Fkl/1d8Zi8I30Erh9DQDTQod0AUk8WBsEr3rTfr
RB3tPcTyHYRYd7vxQYrj4UrF5lGE3KY74cEXocrlUlnjegBjK+UfgH0XWvOVK/CpGRi62VNrHvI6
OruuXth0QOqGcGjoAVWkhNHPUvxdIdOxEywGC6dsWt7n01Dtod3FKPTNt6bta488so0T/vS6uyTP
qONZC8/v+viu4dFb255NkJnawD5Ur7ficJmVHOj7+mq6WJ/ak4/JO0Qk3QoZ7127S/IBceV4VqnB
HNqZZU+QGB1lvY5pWoA25ntQAfERn8gm35xiFJg5Itx7wP5YAznsvGNeYEl2bxJ2vZ5u4Jx+9CIq
LrlKY9iYVHAHjnorhXzWmcO3QK2kqcigixICxA1qwNWsAf09HAdEaAqlA9VoCtGvKmTQQ38N85bF
xjYrcpvDfiJ6ixi2AvDSfdbWM7BwRbPPBnqU9ZPPHfBm3biqOGNghuSRBq6/RKE0Jv3RrqeFv4Iv
0MIt0u+KcDgQKmjfY24vCy41XEv5z7rAQ7tc/1prMBE+aIoAEtYkYoCLqNwNNf09R5WRNGXYu+7J
lSxRBm43+MwYQQush0xc9i8ioA4mqmjgXNiU68M4bnK4H8/q1bW0vz6Bpq5562dcHYOwNl47pBJb
p6gvZ9OMrCnHFyYtEGIhZnn7sCbJPOa3iFILJ6qpHpL7riO/x0Zcjvz5w9PrG+ceue/LKQSqMClj
REqWOrGxED/soKYzLZ1oLHr10OHdvpTI2oMAjTUqcm2EP8Kypp8pM1s/iTpzTHC4wNoD1ug5EeL5
WEUvpaiwau0HJZ+0wtd36WTbAsJCEI6uyWRyOqI1PP8YDYOT+9/cJ4kcX3JvgXGy2//efs2wXWjg
0g6aDMgpsuidGABs89m6MwjS2nwMRgy3zrfAArQPZ5lHGt2VOGTIyoyK3HlqsLJw4bhLNZFkd6GC
HImE0YpE5aFnVGYR5eKR8UH8mmT6OVFFWcyr2xiXJGsVGaBe8wfe6NxiwpzJ/mQ4UjvA6I6xNwSj
TKS9giThS2rjelG6q8sZYB76C+57FCVv9VCrqMXo9Xd1e6tRrjwpQMc60QfUTRZoA1etsqcXcYWn
DVmk0GLYZ8+w6KUacBgwz3t011P7wwv5g0s7WD7Qt8662eqB4xrWv1uTNgvxs2yJpcuIDbL7ha5J
dfS6aDQgbPHi7JFovyY+bPFw8EK4he3fZdQrwSshqEzX9coZo+SpUq27PuG0rJOv/hKFHTDQSRQR
P78/MoiqMRn9zNQJMICPgb+3Ucvx4zKK3BnhHFKRlkDcRR9NGDwYsvMr65sNqvcfGcRHSt1SpC5n
3ztnx2FZoO7JLNwXULzQynsBpXOQnrzprnXt97NxpYuEYqDW0B1/9akOThPMV2O0dCHfjOuG0Ghr
qVOiwKuAdgYJSxYr6Ji0VjOscDKrK0W2MVT+ELGIm+GfaI3OPmiU+ZE+w7B3CyTP0pVTon0+yS0X
zkdOKdiAmPSyc17G/HNA57T8LyoH4omqoXfUgYTEID7kJXDQUhkSufr2bEiTs16VJ9RTScuY7CHa
9J+2olTDVtLIxzjvxh7TqiY8gWUUhbaCUiiIXFk4a8NJKpwQrlls9XqBaEujvaLDTn6zMjo3nu8R
M3WVh9cYAZAyVTIeRiboeLW/X2WhBmARQ+/g9uIdZTPxXgSr1TLbL+UTGe2C3bDVqpFGDrrjC4aK
1z0Jiar2LWyx9vVGRtzfKyrD4bgu+EGZd52WOMKbxa5am9CDdKUgbNtVzUf9bCUgj9hzw984k3p1
YGePauZ+Zbe4V6lO/F3fWtO70sIkRylo5VwDiNms+mVQFQe6aex0MTFARK2dVxYMnU2SzV61/iAk
ZOxGSXyul3M8BqfeQe/UXnw8TjpXSUvB3Lp8neLPrcqv+BBEW1ZwxgLII4bxtnkr1RNGC0z6CFMS
uy1bOgFgEi+lZRQvN4dTmfB9ihkAUn6+DDb/GxyIC55ycUtwRGGCrs4473z9WFGcH8C/C2gcRUHl
sz35U7hGmMyqe/+hGVX7zCl+R7B7x1LcTTow9amHrFv1cxcw6oeFb94N85dNvdgitOrGxr2pFkvC
XtR9bUb3MVaVEE+Kda/mMN4gNlFRFDLe8A5JLVMgPski2Dg1JtSiQx77nqftruNPqMvhPi4QJv3f
Iv+UVCnTUHA7YsUdxbAYWpZVfO+LmwSaHXTXfSRGbPJ7SKNEWI9ly/lkI2/aY5FWi0+06f2DO7CI
LLbmBWyzn6HHGsJMm4/vrIAQl0ojXKlr1ykAjfMZzYK5rFN9lcuY30VyREaa4Y0WuagJF4PFE3dv
+zHoNhe/RWmla9umZwHYye4kQXAHXiyCHT58j+DsfXC7e5a+kUY/sJrRFeoBYufplvWOdUF02EP3
jpYXxQhzb9ziBneITUnrZTBNvC9CiAzMYtgWGCFI8IzSBQHbVGhYnDeDC91Aha5JEeChWiB3xufB
kTyZTIaL7O5mbBZOfJgb4GV5lFEfHo7DcOI5RNIKT9zIPUkbhhVol8nLxbn9SzhnKiLcmwpQzFZI
GA8b/xKtCihMovkasgV72aMMcQjs9qUMIje9YjdzhYimtawfqyBtPh3GztFyVBZQtFbJcseVWuZA
BPrjgVSJ5rxrLq5WqraAt6TM/rFTpuAvRasOem/UBZifcHkWzI9TQdb1AvDWH4JukjxSXURl/IBu
7ipbKvP6ZHplNVQ6OFl78il3wTyvqOlI+OBJQN5WcnaHwg4lAbDRl4LWmBXiflB2SHQpkFGbQ+jN
qa8qqb7RQbszxKmaxVznV5cmi5NQAXKOkPG5D+ammdoGTq3b4IMznKDBeuo+ga0TdW+JAwnIvq2W
6XGg+9hsxw51T86/UK9em2he4JS7wjQshScBijHmYqXqyTELKW48rVAJmBMlnz5YeQqDRTR+ilTY
V1fPfawxS1sp0mtHJObQN57gks2Ua5cKKDpErKPJVM0+numGSgYOsa7FqaAtz8W7jkTvPoPigaw6
lE0wIA6Ln996L+4fwf3kV6RK5Y2ou3+tO7VXCCOEKkO8BY13Sjyi7WolECQrTybUWgtLPm1i1ABj
QERpEln8ADKAmFpbeibO8ees8OKi4CCXZICgWrz7WY4C2jEgKsbreNf1EQgvaszhRenEM1HkE7In
7dDaH9bXBGKsTkPpfpGsYzfE+gyHMILksCWxLX0bDScAsitQ7vdOtrBmLzxlhQwDLqQSk33ivK7n
KkE7zJuvECLrcv8A3dAzNC43lmtUGW3DX7x43AXIBjYrPKvskPaKg0T+Z42FO5uuVfQAJQc9ypuI
qEblT6k2fyP2WByXTj8g+9tvR+77AZhlXQkiJ3Yfsm4+DW5AEMIem4Uw6z6r8ebrCzcsKD5Nx0Qq
XKEMwB/Hn+sipIJsXXMKzMSU1uQvTqKn4CSNrdehMV3j1jmedQIJp6prcS8LeP1DZpOR8fQYxyRC
Q/hXlSzI/VIxxeXgmcxIKtvCRrrbdQNdAiZie8nQ6takwvnk74QFEie4hhhMfUvAVMm0ipwpkI4c
Y52Rt/mmBYacLCsZTybYbArhltDV3a6WLqAqhfG3292LoSqrc3C7Wbh9Qw/qiQkova7jCemnBgXA
EBau5sppMU+U/p303nSuZdANUpbT6rQwULlWd75uPvZTwW6Wx7qQO92duHVTCZHaCwQ5mirbf2H6
lE9u9a0hAPYPMYbDPDsgX5QEKcRXLnlAdpenfo9eMevpjNS3Th9ZMNzka1Dzwk+fgxCqylZANdIW
lAlrSkPKzPqNGYfaEDMemKoGlXSefbHMbrMvRWy6oSQEUeThhoulOqGgHZqDdp4BASMpRf+BwNNc
Q4uJg+M+vGIs9uOxnxdrSkGNxpWtScGYOLlH15rTbqhFJZOu3T12h50zqMdz+36pqtByyjKgKhUC
JvmAC4EuN7+GS0zl/kdPYZaMmtBuxTJ4aOt0Vz33ib16dGkDAWdAIVjqKkAo89sOTfTJw74dsN5g
oAHOXj9BO0QlT/mzQQeI+PFRKpAM7wUWYTwU+w8tQI9gP06rnY6q44LAD5pTcX0LedscpdofSCoN
IxSYNW2Ncj8Upqrtf/6Ay/+oaWLGHVvYsHqraYJoChZzWjsiKrSGO1JzQVtG159braBJdLyUEGUV
Op+1DjinXM946uqS4aaNbor5/6Y+ZXop9qaEbjYoaknCgqkdgPfcvNATsrF9DZ0elJP7vrJTa8N2
y9SbVjdl//SMcNcKWgHIecHj3cAhV6k6UtXXwDfMtWkRunRRoEmDiyy47N4Mvn4Q3XzTB7DvJygn
gWBERZh1WZRpbtQGptpNJ3fecdM9cde6vU/IwyrkzbI+cG3KGDcxK4/wrJY4mutHcysa74PCvZLc
jMbsIcGsGicMJSt9B+pwARMk3mbl5dn3gJemwa+WWCfbNPyGV/nor/m5TqTEqFcnyFLxdN++s8+z
HIzP6HL/hBKBDtO3asvV8hZSp/EfzwxA478nenndLz1JLKkkd4mCj5muxTmqs46u5qoTMNoBRlVB
oqQ5bgjwaO7D7rvpGTD5dllpR8N3qcRATY1UHIGlaPNBdJOUyk0f+JOPNjfb2OLyfoADhWYORp4V
HdGKstns065CYdailT+p6SN0W91mZAUoFHEFHTHeMFNxHhe9stDsS8UkVM5pJOW2apRMV52wUInE
CvgtZFkfopChk1ibL8jDOs+4+EBq/Bp+fktItLpf+9RAzeOUgblq731PJZL85dUKPviZ58zRgzSl
BavJIFpxYXCIhDIUwW7Sf9ALdzBgQmJ1iFs79adRAJUWrheEPJla04p8vhfraN5w+uHJRcjr49V5
TGEmYiV4KrDF5utz9gIBCiy6KhTVK6yX+89oqi3JqjHT0ddF/beR8XJKHY4Rl7P5QD4gkZE/d3z7
z+estwIV71O+cKst0jI4hJjkMWQtaFwbuNOz41Q5Ed6I4eOoYkqu+1AwTqq/NX6W8mJLGCBpuEkI
ovlhVw1sZGb0Rkk2/offLmSmUXyau5mq0s0w3huvP6FiWF/koEchtLzqXFQS4wpS6+cYSsNMNj9J
66Jsz+XSTPWoNrqV0EVEba0peRo5g/gkOpS68jddQOCiyKm0wWK1wEtfjY1kACM0HXfEW6NF7Lb1
JqSryI+6WJ+JPDTjlaLzzr+ZgUQaLe13uA1MPGOsFz6l9Auv47lkKxIF5MzLffrdm8XJYBGJqpy5
1lnm6k77TGcmXfTLuVNpHSVswgPbXvDIcl6DOP4M7nq2mXfYNE0S9xvWLnOUYmbp5aMgx7FhEEMR
fd2oBLjrxOM/Fk70ubcCr3iiTaFcHAMZZsHZ13OP5NLuT0W2ZzkqVj1//hGvhHZZmti0lVI8Pdp6
bL8/mW+NVH+qUfwwinl54sR2Ya4Typ+qgWG77wCOMYd+NmHI8z2omP6WLlccJ5DNwtjhOs3BlRo7
psnbkG23qxqna4pRLD6Mvu7kyglBaeJaxaR77GaqX4Ni5187m0xZl8BTpF/SIxik6UCxuaCCQAbV
r/9JUe5K+Kcm2bhsN6WHCBpB/3tyo7zYWeKkHATlc+nWActiPHC5d0k4vzXx7VV3fK2eeqtrCTVs
ReVNbJmfRneeVxQ4JGs5c1swTzoURRPY+VFKOW7eCu52YAKhOJ5NcS3hJ8wHm3zvkJe6Zv6Pb9ep
hKSHRwxtUlgKFrmR0k1kC2fCQClZDmoVCjCGdZZBqqM030p/tVK7mUl0quydqVmR9pKSG1/UjuS4
QPdycV4r2nY+03X5JqNFYmI5pkurkf+o6cpZk5aXtxMxiXiTTFLQchTFfFzBO+WhuYwXYPj3E/O4
G79zWwQOXIp2jmEy32QsQlp8++lmOLnD+33N9kbHAl4kTRn0YTblvyEEimthkL3rVv77/5x3JZl9
6UraUN2/rXNus/Lt1kuv1aVgP5fwGqc+iMnx3ehlzkjJEGy/oCOgtzuDTwIRXRDyox7kZvQ2Is9x
AI4foq8XHvtRMP/jqQfvjUUeO3jdhovLN4EmqwwtCfAaQcMk+y+1VZ0RAYPt+Zm4Ih8pSMxsUM6I
s4yVtQPtj/WOUUeXmVHYOwNlxf7/DqGdlloOK+6fs7XAmjGSTzvmM/7t4PKxJ/eB9kl3oA5CUfxV
QTMn5ouDDZ14S1p1iu+Wgs0xjcLpA6LAn6oXOJdR45DPy77fauSns9MLEhC1OFMuAbi17GPhe/Kh
pRecJdabfD5Kqwowu+T56TXBEcCHgCiJdSShPx/mJZkVVTZFBRfVCqnRhQgu9pR/sOyek+FGCcIc
En2EGsQKPDRp+WJ4BHaR64YyQf/pDu0guMHcFbc795wNGduTUeYK1FyyFrPkBFHFHup8enduXfe9
AHZJfc0cvQ3WufzIDnD6vWFWsxe4Up0PKqTybZ50Jwr+uIxTNdO8YVXJXIs92GDG8kK/rua5oPLe
HJzvXPTudfv5JpTZI+xhHdA4LtgqiyFSZoO1iGKu7Z4zsWyHAGbZgLZ5Od27g1jm/48r24OGlVbi
ITJ8rYCr2EgJWhsOAXSstAD1pTysiHY4gUv6IFDqlsxOA23Ch8GlTNZ00rgCzsHDruISNWrXMCJQ
e3Qzf0DSdW1rJUKbGwEyeagqmc1SsnLmR1mYBhliCAqgh9nYyZsgHNX9UAwr6/iVppZPeKdCvKL1
9F0DOrGpWD324XSWDc3lWhCOdW1b3eWPMy2KDBE+Z3cbs/QWV3+4pUlOp1s4YxHPyx0aQC+A0GjO
YIVpmZeZCKdzX3IEomrg3O/qcZR3/yg1ajoNt/p806rGXLxVlsB8FbjxMn0a8AlGJl5eST+teZHA
zMYzIPpWRY61VgKLkY6H9VJYx/goakmK04u3FHHSf1Qu6e/hTks6C6HBTKcn4uBzR1Gnds7va9QJ
i35R107kvmQIMhTlezOF6+gFnrpHbCqHW/wyDkxBghxgcbhLLc6Rj/3LHU6odgSm8wKqz2MU9mei
t9tAgQHS6rCPZewZh8A86McfGe5T8nyMbnuMXaw11LMn0JZn9u/fDMkOqkPj9+qZLwg8vKskWJ5b
RxIEDZhWm9Sdd+08UTRHIiOtPokc0qYvL8cAuF1zMAOAqw3dh8FChpaGqkQgeTGO39unPwXEWfwl
/IHOwHf0/Qu9tod1Zlg/nRAXP0LXHT9dUxhvJMvbdTvJPpgSSUd5tPVPC13g3P4jnl8LA2Kaq42/
NLdZ9XF7WY7zsLNIQo9pCANdK1WLuAJ1qji4foBMtu+3JYs9MTjIw2kc+2Cj7oYvrvNTB707+6se
ceUkW/UK6CkRMvn04yXu2WURstyaB3PBOwZSEhiAD+KoaRvcR/ltysXcvsTUHAlVdqWF/OGwl5sW
2xFkpMNXD1k66juVFMtLh6+8Yp++bMsnf6djZgYKix0edYPED2Z/s05ACMKAwh27C1Lfu0IArMrc
nD1xDGTAPloAbabY1UyNj9UTPaT0NQ1V5XbhXBN7dqfCN2ukVx2/5qkiAhzw3LT1fqsultFsyKvU
sSONDM+7UVvm59ohJYFjdw0Lq/4ME51wskEUTg8JBgOWWKppn7LYa0HqIbwflv1mkey8MEv0Iv9x
leEjc6DCk11/BTjY08OzFeUPS0VuPzCU4oRveUduGa+wNtfoQIJPwCgClKIsHJC5zIGBUQ4X5CLA
bDhgwC8E0LjPZcDrUbCXphQiqiFHIpDXsO5OY6ZKLTl2ZEygMby7cXi/YTyNH9ANJaiJTJVbCDjN
ORhxDxhWG6ue+afOzDvq007c1jLMLtGlswjG5jKe1g6nRiqyGRS0Km0hbJbSf3vHyI6wSIGYPLEq
ssbxuK7pUJ/rPrRg63acT5XOVJSbU4PTvUtpwPL8Ew/4hz3iWxoa0vAmIcHOtjZg6mPzyLN6If/2
2ZexhnF3QmKUq9gKiX7IrvGWwnVmIaDNU+T/6aXcllQ/unQLvDWlf+9fMkzg1jp/L9bKUQGYF0Rn
aYrtcBei+Q/BWhJ0x3UpWX5Zlqm4jNsx+4GbFW5MroQTRNk2XNyYEJy1S2n3kEIfx5pNXerbLjQt
lTVOrQVOMdu5kQdWZKgrXdb1H0G0SdpTDk82AKDlTH8XvJDWNDK+zJpDDDzPykDVvZ0+gW0P6fcE
/88m4UJa22aoqpI2eNLxvD1uVn2HXF+SszafnR2esVLiS8gboXkY5u84jxC0FLZ1557KDZ0wlKt7
ek98xOgSRwkcv/QjSejrRfEry+jKbtJalJzMy5RZ2hpYbs6RGu3Vma6GtcCFzwYMTKhxYuq5D0i6
wwVDh5fYKrOgIKsN9s0Qx2TCIqN02JYyFWXgrEiMBPF7YMIkMyCR1VFVoUvybFBTCju0j97mJ7bB
JCXQjHoCxgtClPEkk1DRowE1IpRs90cW9gTEiHCVBWfOPqLoCI3E80zf/JoUZcxxP+gdO9zSK1v6
5gkDaoqKCcEqJvPOv0Z6sDU7cGZNW7tFvZZMOUI2bOt5tXjCwG4hFJap3kBa1RAOtgS3MqxAyZ2F
+h5Sd/MmiMsyDxQekOpMfTFpACaLdDruPO+4TpycrESs00uDavjKomzit7BJ4rjxVkr8LjJoCtL0
hG8+dmtH8YF3stBh90GpdAzsynEjoh7o0Zlq66LRodevVrh6l03hooioWbq57yBTDOWfSnDG8d8g
XvSAaTVF8lecNHBmETXWrdEQM2Un7ezmA4djciAwBfNi78Kbkx+cv54xYltSZT2AmiQ8CFCXUqvi
QlgkSpb6fF6BQQvH1AXsb6VI7el6NmXEvOyb+GDkUdPent7NncQD4gNtd/uCYC/WBNfDUZlNc2ea
0GbvSoycJwU2f+rQsRUbbCwMJr0CoZSQcOdtJ7kKCpMvjHz+Q1S0yBYxB7r475ogcQk0gsU4BRD4
LkrseQ92yeHeSNV1afmsZTjKv7+ZKUgDWDz3j40rV0OYiZvNuhTxeTkHlwd99YFgDS8+7SsHtGz9
T06ZF8Jho7vPBLN6Le075NKOimmkul2/FeP02cNcZsTBJ4Bh9K2eh9VKGC7PYCzkP5V+eE2Psp5S
5dLluuqQ1TrZSZy/sQ/pTDQUU5UQIJ+b8XH5bq6/nfKegcbUF2X+3+NfPaR5rnL99PIeeWX86gFN
iZAbxF8fz1GERS5JRs8W/OoD5yn7sL+Zjm9RxfTzzZvS580nxwnLro2jlMy5KLL4QkH+sZ/moEN+
t/LkVqJ9QEZSHBjYx0hUN8O3eBoazZNQWk7moQod/02tGxgAdn3SUA2Xm1mTsSJIaeuEcC5fRxty
ShT1V/bQxh/Nc/CG626PvRBTAohHqn3dV1gmowhT0fEHaOX8T6vv06X7o2IZXA8VVDVC57YojDos
uLfZ5Bz+DM/yVB3hLEHZv1YI6Y1rgzzRe//8QX0k46im/T5FkKwBkISiKVWJK/Sf+z0xaD9cvouk
wEtFhkJ6BFEsVq+7J0utBPUfNJHfq49r8hQto9ECqIbO0lo7fGRSgC5gC2yWjPXYsM1L5VhRyZes
C2moK6yYykGbAWu98FLnA3tWgewPAfZDgJxlssazgE4A253cdF+a0wvaMdedBOXXGiDfWsq6gq9v
/3IUzaE5sCjMff2tpKMeW5UtRMMvwxljcj2E1XudQQNgI7ZNrn2qorXOm1NVslP/svNP4FEOW4ey
08BFQ33WFCbY6S/LZh7BSHlvbIo8Af3YBVOYdF4XJlESd5MGvKPt1gNPjpQVCSJCXu3+XhX59rPh
6gAhDRrYGqePhNyj4j3Ton23WKv8b7g9mAsscyrt9+q1jTCgFPvf/M8cqyythn4grwSTTL83akqN
LsvzfPGzwJUTpNk1ffOE9fuCsOEjS43GZBiUaZ1/zVmXouvq5KP59uhsyaYJ+tcl9xlDPCTEFFLj
8+jFh5YwRKjRtjbE6ylYe3eknbzT4sKJgWYe8w3K8Y4pFZx4yzVBOIO9ubuGyEOWsUL/pvn2R+nT
XFnbGD0pMWuGN4hRywG8Oetx2qVKY1M+YR88UqMYOZbuF07ypeaQ8DN+RAP2tpDdxkc4ayXgYuxV
hHVQL36nQNCNJN2eOYMkdXxc0hep76dOH5f/dWIQGtjkqirsLUZHXorTOrAaHhM6mmbbrV78LW/m
wwCfPjUQB2aRHdIJsAw1sG4gBDfh1BXlnQ2xH/8EXHYo94k4F8c4IXy8gy1dVUctsBSm8CnT+6aM
zCHnPN0gUQC/HNbhWswBogke3EFZnjBNRbVJoCbPUj/KA6JIbkUPPSUIgg4cb/tjRKQGMWFvwjDl
SYXYRzgpSfSErL4Ao7L18u+C+UWmWmpKzJSuR1RpWmWJSfV+u7t+HWv5LBEInhXhIwHiPuIm2RIf
PxJjRheDN+pYhoRpLQRfWyYwLJ2aqRRCAeBJM9BmqpE67OAs7zwanCVOqLlnOD4ZzTQvDPpQOMMS
wqEzFb5gtj5SHUZM6GxNDgvxWqqnouThaaqGOPvmv36VyqssdBbVt6Vwy/CZDNzn4TrIKH+/jLpS
THUZPGfhgRc3NQDZbig1Y8GdDuOGYoT7CU7fdUAek+l+rORhtL0f+EUqFT0DzU+mFpBJ3dBWhE6x
lZM0QlfRTTPFBThwmAkPRPGnSFOej7aQ2J3Iv8dfmlsWgBpKnXSfSMJSO0o97TH4LNj3Zddqg4la
Mw+2oMo+MlWzgCqb3eY+vREIGkSDrFAkOxnpQG0BF9LGSCPuRAwhL8WIQDkk8pNgyq+UdmroHVPU
1jWouAJ0zhYwadu2l4iT00g8yS9JQNQUvjbijYi9uiUE1iaLzg8EWn3Wh8Q2kvwt6U5uGuHkddRZ
h1/6G8zCHkyb6rPZrtoFeAoJiX8t6iohIbC4BRL1j0/xSByfmjd555Ydey9usrPgrN32bHrxsV7s
vTbnMCvc5mnPuTaw/Uol7Nv/C+ltQo7F+Pcmy8hR2gMPDFTsS3OChhpOG1yqKVeltoGUsxhVUMwS
fFUkwQoU8PX5CfMmsAQrj5X1AvPHgZ5laQJoUJB3XnPpsI4o+CuY4yWXB3l10V5PWoIaYtqu2b7Q
zHX3C8bRFz/yGbWLqR044wBiZRuArCV/cET7Dlaq5N7UBGNzx9wI5P21WeG7TRQtSZASJ6saQNnp
CyQPCpxviJxCnuauCAZ7PvCsBSpiPH/P+a3daco20yKlS+JAgBDlSXX61PNbotKPGMwoGJamCwGp
xq8Qt1uavHARoAuggdR7p/ykBI7bzh/lGYXczrwq+zyj1hgsTNfU03i7RnCOgscg74BXoNof6Ki3
aIy09hsKEqN6SjE4rblmrtN7RuJR0R1YMLK63T+YGeVe1TNor1Tr5BrB886fUzhNeeGM1NycZ4w2
6SMjxwSBWjdaTIwGFBWE6u7yBZDQfsMdyp0ikUkddnZgWiass+W8bfqN8zq3++5/m6Ot/hJojPpW
PgWe7+851xkfXWY5plsdyYKf9gK+xWTsj69hJrIU6GPwC+E3OMpxYiYf7ilZd3q9ZD5yewlvD0c7
K3iZLgNHiNIM60ZUSoEgI1JgZ9RC4dcm5xZ3jT50j6arvUcdHDx0NL0v0xhWFn8dSgYm9A36/LTU
1aerf2cfiMxnPQzcMjLyMsyoJBnRpIer8lF1RyVbAwwQnJEtvLZ7mKrG/ZuS/Rjt/ckUtIlQ6+pn
TCzPGSkjYpcqQWEW1oTVYO/eDi7XYbNzotJcg3dyeTypyuyL7iG8AxBSBbiIcbkEEGKd48QPJma9
pYSni9dN5ElGN5qpNGSZ9n6bZlqRCYSxW8u0TxUMloMY/rbRZZINDpNYNum/1ol/5bX2WnCREZmK
e2kDvX2hxFBRzWwspi3Cv9zMHpIViAlv3yOAN68NuEsnDlgHChpHo47417iYik31IlRywuOYCRSX
fknHwiGooyYQW8FPb04SlInz6sg+MrOHVYT+oxXJJ4tP1ErwaVAOKq+CMWdK9zBwphqKvSQaWZvA
HjTSNoaA6iSwaoUddFTfimgjLK7Rk52bmDji4zqLwOxa9VFdPrXtpLmZJ0NT6Q9Oqm10xNWpyC3y
dbeHn4nI0Cen3z5Lt/zma24r4dw7hZUfsOARXpAhYU9m9W0469eEcswZFt/s+M/VHBLc8ZWYGcmF
MxqAibhTxRIWBge0zrsxtXbUNJnWbFRjcRWM6sPUBEqaqITsTlXY8JDuwMa35Lyodm/5+PB5D0VB
JjJeKLVFRRTW83JIeWu/RCsKXkXmFc/kgWoIqEU+HwFbCKSUuvMEMyADpnzhDuCdBBC8Oahvtmy+
dqdKMtU9eu9fh14zkic+rr11jisg3aFXVSmFyE/SMQcsLfUNv8A5adc4quJzsMZTLv6SqpbijrVr
vdPfJ5loC6U3iba9wjmOd4/Ko5UzO/1786niz3gP1cxkX5nBi14TgtxbWWBt0xw4ajp10xvsLUkd
2pwkaY+erbTZrvJ9XYNAaNzjwwwVAnnIHeOrv4T1s+WoX98kBhZ82Bv350X77pbz/qEkwR0mIp4U
Gi3P324LtRzDBcKlelUhqWMiv5bJWI10IyW+6f1tjqL65WutmBZXZZCFjrYutEwSonaPSqx2Qzmn
Zh2XaAFBf4dl7ymbyHHlryXmajB9bWHnn/ccTEoeH5XxqcFJB+Z3pecnND9dEIGNI+UEaNQggwuM
jJReBcX0N9WH+3pUnNQGoWNO7SA26kA+jusfS7l1yJyEU0rBFRB7jiN2PGuQFQ68EPUI1EVmtJCk
JtHmh5Mn803xDxM5wtxSxnIGT3UavdQwCkO2YxHfhmDrGvg1tp78B9FFS+VfsnW7EucbcPcliWbh
PbwIOua3QGF7TZ0VTivCIhpd2KcrwSi9+2fRMOnH5HYRJmxLybYsunfxh1Z+7KkijOLpwVNROjDu
gPaWZYjc6qlHtVFTh7mmbl1J0uMRDhnPbdpIBvCeo6SWtiD6GisT1Balek10jleA9McuJFmB3fAy
WTDKhgxF2VBlHi0JaAnW6OBvEiSEVYhmaxgf1T+OV5OyDeAwU//LQAJPhSXUYG74et0CgJtCv3kv
Ms1tbjg0NMtVrh0ZqHr/dzXmp4yViDOICNTQvoH+Rz4s/+BoTcm8OHKw9UBIS6YO6J3/HPFDorDL
b31QHp9eBWh8owQOpu0uMV7qvrwHy8KL9JLPtH9qtEmzqQ9F50hsb6TVsoHFZkkAs1Z5UyxAeHoO
zS/rQ+Bbp3zPgR2mIJ+OBIms/rogcNfn4JYu9O7DRL9zEoOVf3Fr3LH8/lIASmiVzTRHHZni4jnF
rjFLEwnYv/BQYGNLBiZMrL5bPEB3huarC7YnMySvlDFXQAEwOD9vvRUbw4T8BNdjwPWfMXlmrq+C
/SdIhVorSfBoaKqkRO9Fw0quxnqQbYLtPvNcrRRzdENCTjwaS7lwQwAUwGTeKXXkP1ypMTC3cM+I
qH83e+k/X7xUOXtRQu0gDGPKWW3syui1ER+zx6+ayan+umqSe4Db+owJdStH7R9//Ng27a7gHFip
EfLpNJWH5sEegryu/AywnDsIQEJyFeCDvIz2kQ0tNbV4/qs3AWweGvIYllrt6C7SytNcJsLGC9DJ
1+Xl8eldq+klDhv6yENNoUAxjtm6omzVLKWhmdQCCWwLOMdk5IYWjpDgD1a0E1OGqn9ZG0mYJ9sT
GW8OR1HikNQpcVQ7BrBXYH/M+EPvj+quEYq3y02ifARt7GDgPrfAjfYPqUtj9vNU2Ntctf1Kam5H
pP3iwz32w6s/+B7BL58g3Bl0qTm8c6EtDJKt/doo3YzO8k+SlIaf8nu2Um4mUs9qsTpa/WxET8XT
ILz4O0uocQGbaor2mbujuGXl7IPrpRejRZxsTxFhF3qTrsLX0o210yO39M8nk7ZvpI2AfdNctzRJ
PUntYesNnUN8qj6DlqzFiuzt13FwoXvcgP0OidlMZQ/AEiTdXs+NwWFFy+yGrNemthp18L4OU5PJ
8FTkGa0Bj1LKdEYtBZX0WMljI0L2k3i5z2xO1rATj8gZ57bAySjPnZPMjUCv/9bLFryU8Biszxtg
pW0kDVEj2uIYc4J/9ZnJyaU6Pteh40QmXxNA3zAIkyO1bK9w6Xm8AcKkQQtICoDvGFLdNnaZ5q+M
wS/a0BynJ069PjHDfL8RUxT+1ALFSTExIvuSgFMAUQwxEZHx0xnlp54DpXI6KXJvRrutayZUUmqL
nDzOTSanoEEhJNfSTXpN4hKTzJSK4vTigGEOe6xODT2BlS7I0MNcibhBBcQS47R7Ur0DdcNXwprD
J3OBOEQXaILoNDnzWbGh7Z17r7RBdJob6sntRu8rNHMoCR1wCEUCSMmd5jidhcqoGAuwvTzEB6Qc
5gr4vrMBaEtaRLd+/hqBui+Uy+VB+oRK4ChLVuK8HNB9SlAOCvH/e+eAtvyUqGpuywHO33dgFlAy
Jk7hSdJhrN6FX+hTGtcbbf1L5LT7DZg+7WSSevRaFbX5waJiK8Xhu/nCKNYAymNCROyVCeXASziY
AhuViXYgOpivkN9nYDw4LeEZOqSabe9TD+SZls5B7J2NOY71qbvyxdqHjPiRMKXCigkkzWd7ZLfy
T0fyD86aNIFWy8ar+/aW0wPb6/ke9XXRTH0rB8mtfH+sXLcDvsqaYLbbfmSqW4SY1JOP2PVmcELx
HYkjrjQ9UFNMRc2vKjvhscRFJy+Ygd1wVYaSQDLB0H0SXywHgOJwtlosGwxJor5BS6CdIsF139Eg
/zB0i8BUVP//PDU89fSAPONSWfNMY7jeAL5SLOrmonbhicCQairWvS4W0iXhPeTGUt4ppjxb3yJH
/FQk+d16tDhvLCRjlQOZwQ0XHwlydWVseG6E15bxcyRDEXCPbTttyQnPSwRVJw7vLuUoqcxFLwv3
rTJgLI/KjN/+LXq+sg3XA3COdXqV+8kz3SXQWb8WASgUGI4wZ1I//v+MX0PxXfFdbk18oow0C0tR
hCVgQtNBgm0wpe1wI5SurrbIVHYSSuRD+kvJOuw3ugrpD5N5T7DcRv2UZrLp8CE6seaOePJFLbkH
KkQXEU59PpXqSWebjts+nUMCZOvtvVjoepW7w9vPe6vczd7HrvxdWmjzBUQ1XpZrFKMw0zfWWxq/
FKUbzb8XmoGQ12UFSwIJ8ntbqiTpATG5gJSwKVCBOTvfrfJ/O+zX55bPHavHDKMh1ZACc7Dj42i1
AwJ+rrwjgAHhRyZjcc620/v6ro4QvtMSdPeko+020yLY7Xsr6E4foNCtxncTSp7OZIms2p4F15CV
QQ45rZ3mTs6lR5LPyvhVrgcXyDYFNjGOIR+AB7sCkxnPNHeTa9xX89LkH3IAB/qXla798wi0cRZY
DOL5jwhr6ntoZMujFw0cesMwPsN1n1bNZTiHXe2tg016m01nQloxbp5awl6pJFY7LlgBCHd+PM2m
xP50A3/u1SYIW0ztOIfj5BM6NuwcxssnYn4IG/fdkwTecBUo66kgRwHcjD0R4QzyCMGoSle2y+mV
W4edmmepe9od+6UhD531Tz1FkhQbLc/BjjZYB7jh8J9lFgR0j9XvBDY7QbF3vTmqCzUyl8x/o6P0
q2XyQzesE1cp2JtBTAPEZuIptgxEIB2WenmoPU0WP/uzkG47cO3qQWv3TxI7BWJDEsAl/cfcH66W
eXxht5x0+IPy1VX9wCrIghcqhVXU5YgTe8QEeyOpKxrAaB5I+2naMe2tkmcaPzEaVGBhHyhpXEcY
PVyz5GUCBit90jExjD5S/cPONqg+B7W6HzJ7OFSGGUqqNloC0zKnpAj/4sMfBL31G4x5rxc0020W
kEoUxgtTMxjz6tdqYLNBcmM4RURnIE4WKhDm1cqLNFxUgxl0ZfJjN7K9k/LzwUx+oE/Pe2jSpfUT
5ApTfIvZSBrPsIM9ZhDKZVBReHN1js5KFkKyHIvlBmKZ5C8Lk9nE3eA5/ZKAw6BJkIl0LwXit1ac
Fd0p734SIdIClN+L1MnxlrjW0Nl3zEPnIfIaSd7w6rBYdUGqDnrQstJV0eP3/azJAf1HhTm7VBDq
rtPY09dZ6G7Ru6QKuhyiztXoKU7UgF8Jh2ICktBtg5QaRQmh9QldDimzl+m7NdpDVelJRQfpngNq
G1s2BgKdeJBetQh00g4Jz7jcNlYs4kEMzBMJuB6dI+SarBNZBRAAlby7GosAFBDmAIZ6Y4+6dpoM
bhLH/YDnQfAotiIm6pQtobVMiznRRQYdQhZ0KN0GVkMoD4Kod/Pi7MMA2PAYVoG11CVFF7XANT4O
gMAW/JMWG4pHEaAHMwVsc4uIv9kHPXj/XbJMJchlBfZEi1TFQYHPAdOe4NY8PXYP7mMioeQeZn1Y
APm1b4eVF68Yc+2/40ZpgcLwRbQwrqWbhxFZ5BHVVjj3fIfLUV95xB2cgdMWV9XfTCIjRATPRFnJ
myBWjbydeFiYq5qijUDBswj4yhVUEBH+em5DkrOwNc5Px1ikFrQpFK2sVsofy4EDfKOHpwlUE+2n
WBijsMaFHRmNMHd31ouHc8onIFj7lSq0gd4ujPfsh8ceOdNPlyJi9uq4hSWA7gngWUgdDQXT1UtI
IOWnSTUP+xuK+BP8fHayVto9vPgh/RiHbmbC1OVHJHx2/d+T5hj0RA2aSXIIK74bnuYlnK58JSD3
cYAJPK86nolU2r3yHNBT1I6Gj2eqrfBOycL/wyvegXv0mEr2qInTGgh0I2meQo6EzBHahvHgr3BZ
KnHPu0cIEiKhfVhyZwtQww/ZbUbyqEPmnyLEsCVLeYqi33FL8LunBJK7sRFKhWSGMXzUadVTXGIQ
nV+6VgVka6ue5JUkEQ27/enK/RROu1/nenAEzyUaY/HytyMvSx3DAya+7l4d0d9HC4X4UMRyzAtu
EEcXn9F1V3Z9rfhBngaoOqkT4GGwoa34t+26mRzNp/yaUxuhpD9mlIGu7FZrINw4FTPCOjbPCi+Z
V6HwRhKwn7JR3qasrF/StpEzimE5TQDLq33GgC92B7MYyeBwrQjz/y0tpmoy9slpewh4bY1qcUsd
L0zCgSHaBElaGea+XXys4HrUlSTz6HsCDXJ8YAE7NV22QiL0KC5R1UZovxQYHhcTcP9fbZIrJpyt
ZPCt3KK4S6AWVyUSlFeQO+4Dh/mybifyxXRGq/jvkmTwIvtSYIdpZgSQ6sgL+sj61vc4PFkuI1wy
8a5czhBKlUlqcutEtdHzoYvgGx0+pB7C5P5uWOqdTpAvQNnPkmtFOhADN2Ey44AFZEqcBWwEI++x
oVn/cVW9jcw9PpuG5unIYNY4mz8mqGfzIbqFPb2rInit3X4f6TIPuPCbRDcsncUOBhdKmiId/rPf
26NBFWSIt6U0ButR/jtTtOVSAR50wbXAchEfCSISXZC3J4nqg8K0xQkcdfqGvetljDSnzgsGNzdE
w/27xXEEHUgMXuhMdLgyWuGcqq9dg+r/0qDaHQg0GSmYjUcnPJUDl0FD4JoQk4ZDi+rC7vatD57B
O7p0meuQU+c7Ky3+VT13z4de5/0I9fZ3rqk3/2Nq8vdzl9Wc28NGrmQ8ed1tj4At4n2nriCKs6b/
DMvs2qNU17RExP1WailST7nZYY/LWfmQK+ypI2bnuEHIWu8PR5Kyp0rhOng5AOfuAgNzqa036uuq
tiJNMgzBkk310SGzB03UyAssEtfq+pZY2sq+wfIOL7s1LUmVqP9Ml0yEzov/UzN4xAcvX71pxtYs
4c3GLmztb7SUWz7HUauTOACCwUgbz1hok4fNX31SmXzE0tfY0POe8RN/RSGkJ5emFdfFLJ9rNNog
A397g5hPb6+SC+m8RfM5EdYG1xV7JaAetc0JsCjOf0/EWxZvpV2ZFd6zjYrHiaXHiN6hf67PJbQR
JO/MWuRjrz8qaBfVP7ePEmV/Kc8F8gCdJ3Rk5ieo40STO3eP6NZ4D7JKv0AsrZJ7W3DZqndwIeV2
WBvw9M6GPV6sPn8ycem3181Nq9IxnaIPCQN7SAgfs1B1bh2S6dbupKUbU5MufzGtnx8+T407MEy8
olbHwDJJpgZc3cMk0If4g5okmiSLXgM3/YfsBE5W1ZjJN5vC7th5cx0HbaUfVrx2iFedqmtmx3AB
ZMGOpeatknpPYTVBomRDn6ftKJyMV4gw67tEmAVXDUjOrSY+67eZutdKViTI5AHfvE37hD3D9UPv
6RcuZgR5qKJIdRDQATvHZF0oGytKzVwGHsjwKDxkYq5oMaql5eEXItmaay3EpFKaCF+VnS7Q8Cuc
AboUfDTVHdniOJ5UfnI0huNmWT4ocwcgpSiOBrkiCYB4qZ1u+0ZEcMlHC3EDReHkXMPUpyBQ+6c3
UrU2N2PX5lHnh1/wda6YLfcp3Q/OUOA+6UwShjXg+2kPLGAtRcVmypXzgoLhugaCXNnd/GLe0yOu
P5HYvQ1egQL/JBQKaKnlNskcmXeFeYtQzKsidLvVkSYJ+HGxNlABc9YYWH1lm32g9JidO4JVjSDk
4vxvfTZU5zF9QAbwMEETk8DGc6TRMu9JT6h7EPSsORJnZqCGuymalEDf0rdqTeH1qtCllbQ4u/vt
NHyin136k/UCF5X/8TI0sYlgXu2HgwQV1LdjCQ4POEI0ddWSeBWbQhfTA2svNGQUKyh0Uy4rKC6L
RfdoQaEiAzL4FkhTmg4/7hPKHo5i2lQUxEU9VeNtCcJDdaXgUB2BzPWSJcuVdiZedazPUuX/GDLi
sGyf+HQOEpGBbUwQo1ictE/84eLBkINNZEL9dDVO5wcPPcUpI9RhzBbaAaNNJMETtEW7GH4+7N73
ug84ARs5ZBm5JFinMvui4Z4TY71azsWrSzQfG4Hn2k4RCo0auhL9BImw8w6KoDd2MljPIyvqiMbX
jpbaFd9e9RyDn2kBq0WnAU6qiVOC+PRT+9Udv595EhFXHnUouoHHxomEpQku6mp5Fmy5sY6JUU0X
54OaJFAGi7grs+Wpf6Nth0pQmmhVGbbF2s5Yi/+a5hdibEKxkS/Yu5pJBklWsi/N0rtgXO0+2gNY
c+3ihC+ds0SwS8JVvI+kzPdHRq7tjVUyoTfHD8FCr6MHWbcWt8fSZrsHY1gW4md3zelK2uM2uhjC
AJm93DdgK21iWpaoJjCB8aL4sf8H81MIXdxZSOIC3MpAXfjBmbxqp8QaN17oonC3U3BwQPm/YbcX
hPRo27NBa4oZScw72PcNTsQ50GfhexefO/wGdmS5kTaZi+3tkxm1cmKeO3oRsi0FQdti0JKweri9
aydXv9ooGfOypOQTAjuXRlK/C6bJuVQl4DYe1+glZ6VdyRoGn78Vv8/ZcZ1tBC3DALznm5Ml4c9q
VnoNlhNgXSzDWnh2PRLhD9zJ2ereDo3Zamk367b532qe1H8bekImgX+LVUx04v1BfGgsX2ZSPCPB
mGQRTHPW8XmbnrB8S0DYUBBjxJusxOIp2Fnb60i26KXwidRfEGcfWXCGt9iTH7gmCuLrn2v3eIis
LYGEyi/yYEQrR808KY1aL+KLken/uRiIsNTeQtQ/elSa/m1offGv/cUsyxgvsj5ztkzKAhKG6DC8
dBonRgddMZkJioQwhWCX3n/J/kIF0pdtCg9dP1KtAzScjDXVvtO3WNNruQpcLgrMKQ44mqlkz9UR
hAVGRrscgrMtC4KUAjSLhtZMn3hPVtLE0L2B/ms65EQk1NI5qHDv8M3gNYKSLLH8IQ9kvRAhJ9wU
2giToQDjBG5H+IfBAEJDwbxf56CMvoJYkUXBitqn6RbUO0zAfgNEiByykGP38PaGWiPL4OtivwRa
BIgM0yhn8qHl+EEMxsIW2XFkvM7d7JZCk7SDMX6ApdFajBpN4TmfbpN1pDGVnWbp9CvlYBhuzlsc
8b0E7mI0V64hc5bfytcAR5KDqdMHDESUSi3AkTU8uGYj35/aKIAKcVmVlAEIX1//F8RBOtJlxVk3
rCz/p/RuUdbsL3IHOfqM5oDhw73d8rkAe09kk52wZ5BZjEtFiVusPqs82ymCQLMvw325p0vW5U1C
08iZoCMa2f2czveodK1SmCUtIq/x/Fd//7Ym6eczImyrX6ZlSBIqna3LAFp7jJeO25mO/hMyL/Kq
lV6LYGjMRs0jhZB3KBclw+WfIplFGlJuZjnIVdd9/JWXVt7bjrXJLI58b4ZVafQE3yoosOKl+w82
PByrrFByQQam/mEu0RwJxZn05vzzBaRirGbV8w73Y4NtUozTmWapG6EY+6KJ7Tc5h/kWE0/6keZI
ugx1A6n4+vxdnGS+NRTm3zb4LBzn1rJh/1zrNyAQVpCOsPKhJIjEc1YjI5vaYuyMi2DOL2dnE5Io
wGsYaIEyZBPUW+apHxkZR+U30tFVdruVeF4GJ+XCjRutboHp5Ac5Gfv/pseP+Pc2bYoXiBohRlFE
MkRyeRnRakXrxut/Jz5bhgKDVv+/pUKmCkgh9RtOvgEq90U+oUbWzgqYJINREzkFjpzOYCvvV7IE
sgGlQvCx2cIYEmoovxs5ZznZuH054iSo+GNfXxwQCPJKrq6bP10WZ2UkbKnlLoOcl5BvNDpFf6Vp
J6J5jNDBe8zbvld8/fnZ+M3ec/qUiD+2Mbi8zCE8MsNtFdRhVrjwgUemAG8WlT8YEX8Lc5IcfjM5
TRWp1WTWA7CbHNX+KlmU4MRKBJqq4iE64J1a7ZPqTrSjX2ytBrpBznWTxiOEIBYF0lr5y2TCrooq
xgPlycT1Pp64GZYAwnymT3rA48/JfUg7G0WyDhG8k+NpqjcOzAQv/OT0YTp0ugjWZWA8Y0M+Mrnk
C7MYz7San9tx6ZwP9XLgyndb9psf12AZbfI1B1F1hjkw+78s0e0sDMlKGUSLiJsxETmBl6CLNuiW
RQIFSoHnR/DCq7NbMzpcNpsHxLeJXTpIFLDMOYZ6pkS4pZpt3d4gOwRbADaabDtGm5AKGhNmtOKu
KXTu0/djA+nH3jivgC3kPNLvm5udd0aKDkJRAzIukC1WAZ72S+tcjoL6Q+UCa0oJM+NqQrxT6t8w
f9XyxIoBgOu0/5W4solIvdsz/8mgkHwolN8Yb66k9MF/9lJr2iDPE7vqjYAGmeagmRub/XTgQ4/S
IN/rGu7LKqu67C0/meWz3uvHb+RXyOJm0rPVo3ER0cq56NG11ru2QBQMuyUEKU+VCmk95xWYtGYu
HbpSDCvo6YtYv8cpM/EqwA3AReuVj7pncNUqEaL2om0icZwRLT3rDBgqwF6x4rEsfLOCIA4xeyy6
W+w0vmpLRrKhDeVAMC992Kam3y+9w4W6E6HgCl5vQ8zMkgpYaBsdJNmcgibxeAUEAcgNwYI53OaY
NZkGs4ity42n0mWiQjn+qNVpsEdOJFi58KRzfOtlue5CF5hqH5UuRhTYyjLymHWQO5dQ1zA657As
yLhoIvM7vbMypVSWtylDs5en7hCfDobSww2cen8SKQg7Gt/Ub0ayUNjf3L1L9OErnuxdiYD8ixqN
POxknNj9n9rOWnnBzXN9i1TiZ3VTTFeUMFNQKLFwYmXDvW+9IrH1nIp7OdAavdrIc9EapoAG/LFV
Ovad3uEZgBkgBLqj5N0tzVWylSnXNwahb8tEHV3BCBi+QfBfv4HBZ/rhtQ9UAsmIAzH4jic1ZBCn
+pOU2RLtxZlY1UvGO3NZN1OJ0j75Xp+uFUYcZeTEmdYwe9Shd7VXqblGSkk80qe0cp8cR1wHQuzO
JrXd1NT1aH0JgpFlqdYNout2gMtxdkWw1T3I2eKqzEU96fha+ppIfpItwJDA9xrZaW6xsCGsjG+H
Bw2sWxAmqsGr2Asvle5OUApVGv0nkPNKbO6z2q1zd2o881lkEn/37zCRhakqY8lJdaPhjsm/aUku
BTl+i1l0pht7Ge9P+20LXIxt/esdbC/xisWTFRO+oiwO0eU7g3B3eAcG/tKQJYBa/g8Zpv74SX4b
Us7RD2y/GE4rXfIdOmcg5akFp9IIW1cevm72zsDerRyfmzyN1qr2xjL/sg1bm10X6cEU2zPey8ge
FG+BoXHrsDds/EsJ/jX+XVHOK3WkPwhNvVPrGrwC9KphLIsNfQkuxYgLGEEulzg35tn+LHBk1Xm0
qNgR+AnX4PZlc33rCENOkDTmFUOPBbJo7leDfrd/NZeNIj91yQBAPP//DtgsdYlT7vcLhKPOqCZl
4nsBISeetBJDm8tkNvhW3XO1Bn3ghlSVPfwWnyKZwA+wv5FdrbnAbo3v7l5ou0l2efZB7eP41cu7
szg5ftDI1z1vuzc0+rGYjWm+7B+dihQqi9XZXOyyuOC3nzlgVVnQ1ymFtDf32ijq+ujJ70+XbT7H
++LPSzSCY4kgy6Fot+Y1pCWiA1UmpvwsW3tKlgZ7uQHtEG+doEvPMykh53AfALBu2TfAqmkQjtoG
/E2YZLjjTKINmilIidvdrgsYZtM8MOvQKybiA8oKrRzSEQQJSxfJNJJgnvOOl9cwA3eGhsCACacd
4oR0sGDS+QuUbreFoFcJE6KlLRx6nSFV9CjeU+LtxmmRk+p217ufJ8a7nYCWYhwguFGDw9UVnTMW
yZu7Ly+ClrqH5SCx65ewN4NW6z6CwyOxxByIqQWzFTegS0r16NjVuIBDrLwTQz2gxvLmccQUznis
R55u28e8xNbJmAZGqds83GSl0ZPgceONbqSJWK8GlpkiRgMDD4n6k+6+zWKaNcZd3Ym4RarYKZkG
EP+Weg4FZNee3J/13Y3az3OlIsZN/mxuKHwaH2cKuZw2FKTzTUGdJBTlTeV6mUAlEYf49RNW2OjM
3MDPgoq8pKe2OW9cvHBQxrYDqUd7lnzf6yoC3dHLpcKNIIyxJC3OpSQd+NCnJPtWD9duGv+Gg4iU
me8DegY6psJvbbmJ5UJn168tJsBCa50XlBPMVbtB7cQ3bMt4Rk9v+TeGuN5L+crkjnxeOlBRtswg
wUJAppr5ZJLLXc6XOI0XPhQqKOcj+Mg0oWJu+wFlLcp3cARKzqxg41s33nQApSIKFmuX+08+Ehf6
0sYvmmUqWUkGdjsPJQTv+n5FpBh4rfvWziYGs29cwhGHFlPq+uM8/GSvEYHCURQZP8YZjV+YvZsu
2nYU531B/rpyxIHkhULhIbLAkw4qTJc2elQ3nxwl+ipdwhVcueEp9RMCjAAIGbFXw/WGTzQojVFa
TRse4NW25QH2CbmljdUBMt/31cTkasIWowEtEBykEtITnnKzjxedtymXe6bVHQvVdBV9CAHeXniZ
3TaT/es4ocsg519auQPfgncWU2ZkXT4BsOZQSaz0mG13CdqlmRD5m2YShVErst4graWYRImN62yj
tuMN/l/dS8xAqQmTC4VxCxxrr0rYsazquTip+//Ah/UFM+QQEyww8eMcL22J/HeIh5Q9ZrQlPGlB
oM2A3edSq15kaidiU4R0JWcs+C3tN3mbEw2YaBsLw8WH2XpZTgyggq6jbvt+WyBYeVlZ1DipTT4v
cF9H/e1HyyJO7b/m+AqTjJKdwVYP4xZOOuoF103ujr59oOJIDvTpLbjxUhxkQEC+WW/ySPw7cbC5
4dGabHHhscZjAjS03DMbg+sQzC9N0KBGalmc65nQc8ZlNCe4K5TmTYMZWoLK80/nKOBUPUTUaK0x
KJVe14dEp6Ay6PZ8aI5MLxn95gF+rAvJ4uI2jXPH9fiwIX5yhOz9Aw5V5ayVIkgoJ3nziX1p1kD7
sOqaJMdlaRokwcYmYcEI3iZu5GTw8fONIzBW1hHiVSSgXZy5TsrN4R/ap0VcGJ4j6MwG1pnLuFqn
ZSi4wjryC7FayDKWSyP2IwQoLm1n3+5wqhGXGiPSNFrAIHe786o1LKzMqaj0EkFniMLjo37qdzYM
Spbj3A+eAaDtPaVurY53Di+49bqWk5H6W5aoDkF607cZnim24Kak4SfwXVFqca/EDYjkRU799jZ6
o5TWuPvKBIYWBOUU3ImK74c8UoxMYkqRTE5vSD+uDXnfJFwcQBJa1teozhhJMEdzWU/b7DPGSBnK
IYTKnH9f+m+in/SBa1jVBGw0nujmDfI5Ygn03Wg4ak8xdD+sS5pJHqtGzFfSlBXH+wp77y3PYS7s
jJ0p83F8F2esUhxBtXsSioj+w8otTl8CTkkZg5wQVDlYrRDp6C/ajQdejmiOXVb5WIUVY0C+rXj1
rNzxGwBvQmlpn2e8vtirKwpHL0msGt94GQovDHTFyZ9pC37QaIJLRsvmQForITnzX5vKoDpR6um5
nJv1ZYFs3cL/38oOoYxLdZCO7wX0RezYRMoXzTP5v20ielhEyiL8f+R7jslg2hfJq1qvPiG7Qezt
bYKZ35gleEOgSHKZoPeS+pqF9TZyItM1ZofWSDIg3N51yloNvk6GS2opj0NtUO337aBSahOgJKVj
9zUpTRJmJbyM52QfT/G/svAP9u+U0ghiJshE06/R6lp6b1qHSwDUEaElaOa6UgTlW+LpUjv2byRF
XdLFjNiYVogCmwwAYR0xsKtBy+qJKVXkqxY0RSFESCWU9BgTp7yRQf3VnJJvC8p9OChLop+f/7SM
NXAamgMzWhfWv5HsMW3aG19JjOPXB8/qfMNW5KJyTgXCWBITGcd7GMXaKYqcbE2t+11f/Ujyswdd
UHiDw2r/okB+wmCpukzDKmfpPKScmKvSNoJe63SptxUcNBDsfJ3rrCIFzVZVZKf5Gouv3Mwd/pGD
FwA21vquNUiG5P028zKIb4aksgI698iz9P1r1qlKP5EnkFhwIQ8vuyim6utJ4hqCMlmfQX3Y7PC9
j7MuVsjdsjB1updGBzbi02p5YwsbR94YezTiQxHuUC1UoJU7+Jc0wN9WZ3JwqVj4XnLxoXtWAPdp
15nCPOM8Lw+VrzR7WjkbrwyfM89kCgW7FRELEPC1OvekCEXcb/SBzqzQeQjFtacXZnsS5HOKaCG0
nooSFjUAz9qiSKE048zMcjOiY0GL7dEXs5TqvP4AXRNIPE58Hien7roqgc4kHajEO4DMBcYb1H07
15MIlEeYpJNsemHy9FhBiMY0L+ndD5kB5EDYwXi1A2e9IFXh8AL1araYoSu3oeAnkzcGc26p+4Et
wOhtGt7oNhON1dPAxe6rRsEkT9IeY1tGPyD4HU541yEmLDzKstiimp/qSPHGdEK074J0w9FaCbyX
S+B6XJm2x/aLUiF2e50tJSV3dCK6KB3terJEW6Fahu+d3A21TXzoh5QIwGEOg4UnhQ8T0D4b/36n
3AGqvWYzsVRkXKSXwxi86+VLnWszY+Y1853Cc7Kyl08Lf/cChjpST95w0i2sYv9BdLgIyEEUhWJe
ltFTTNrm3qNAHwCGw8hpLENSZqs24KOY6rKL3tfdb3Cz4J76eBEUPxIuIBT+rzcXoel5NkPM9BDw
pCG57zCofIkoI4569Knon9zll2/yz1H9HI70zddQJN961BWPJUXikheiB56b01A1Us5jS1AzPqGD
g7iF5JfyuvceDs967L7tugm5qC68u+v7hzV+bT5F/5xYgAE4htxCqOZ/MvzWmaRKkF+8EJnOcqXM
ACYFRT4xS1m7zznMunvjrZfhXLsaoJx1mp6DceUt9xAGZHybVdfuZ04QzS9rvvHouGhsIEIpKCiF
tPDFNM2/hcrQGOUTNDIMwELUHapGiXIA8zGlNbTvzWO54mKs2b+gWugTYVKIyvksDO1ebA85kYcu
BMkcv7g2FjAm5qPoy2pr0PzyY3MHubhNQeZgwpcZUGOUaAE42Y7ph/NN2QAX1CGj28FEJ9/foQtc
RZBQ0q/+Q/1+9PGBhR9NlXizKrwnNxzguGgvtSYQMYEaoBzcWbr+KRNEAwQPQyAil9XQNnntg8gL
PNsquNFq07/NDw/0B8klKyXxhvMg/pHOcdVJDUUBr04loEglCTeIeQ9ODD0VADbBRIprJShtyIyg
HfQiNztDWI/TOugY4Lqd4t5/5YVH2YcaRFnzJXpJpMuqWdrKzyLbz3zplF1Id/t3BECPzP4nGq22
x2EPrkRxgZo+ufm1RX8JQXRwiEuONsQ+UCQyP2g7XI0XraOABtYqhrscGPhr4d0dS5TUCgEsSh5i
dol12TslRoJhzNKA0e87MhNabfevIcZbwA3CVmypH5vrK4rc0Afig2VmhxlmUsXWjj5VJJ13ciU8
BOG3/jF/6amX0mCXYGuCWyUTVrhGahY2fbxa5cXMFMk8ZN9SYWz9uYF2RXGohf7PWzPZAs/Npgfl
lO12HZJTEaasHgtAHyDWY1oV8G6ohoj55uk//xR/RjsasroT3cap63T3wGYz0YBvMaUQF1PCS/sZ
sYpyetR3ersNjD4cRHjUh7MCIUkgeRSAEKRkFlm9R4oo/+rZyxjSxyAKaoWENQOP0TrF2GK6T96L
7VeWxd9ZkqrR08g+n73trIPU+mgeUQFU9k8zq5FR6earUuItAIoohKsAYQm3U5i+4I7iHvgTKGNG
zY1KufFs7mnKgMGIINfZXEesK+crEukML0NKvr0hMT33+zWEXrqqufzrtC2Q3eBzs+GO5MpygfHl
iPHM1PUQAxsxdVOaANFIM4Wj2wtF5iPyLKIjbQqgDECeJ7lWRYcVUagfUl533XMemFWYvp3Y2hEb
tfMSqR1C3n8t2SX1amUFqRpvrz5ErsMOeq0BmApHUDmb0CU2t/kdKl3FaHGrZq/Wprzaqmzi2I5a
Xp7MXNslx7njLflSSW9Eag7nWQP2cV8J6RlQgQnTSxY+1/THZCOJUwR1WiYWZyIMKYhaLZWz6Ywq
d5bhZWiDQu/SKPw70a1vG5cdAvjHNaVPduV8yyVtPN8Ogqb/n2CA4sZHrYa3klFb3B6OLJ8MxJwg
kvLedaQBcuBtn6FReduPcVYAFWg/u9LIq6fC5qKxETPG5vvPcQ3m91AwcvmPd7Jl/1Sp624iFytL
/7O4+xDrPqC4domClMSUnb2IJjtLt+hG+uHLvhQbS6snTMCP0/YB4Uf201DCBs3X3YpVx2R20MOS
IpH6CYUEdCu+q3yYM9/AEYlM/1q0mYsgKYjMGsMLyvcfVovy8QeorGdvHIi8AvIDC9PNh4okHhc6
tprtF8/w0HAVCxBsQB2e724HHjK5W5JcNCwYS+v0cNw+rffptQ+TKIPAp8Nc0bWHb4+M8WRgo2Da
Q10H2hfHbqgu47OZDJj73R5jmMV92Djbp28CKM4XZfDvEuwb+pZ311/khRqzo2epSeFCKcfnPesz
nTHfe0vB6X9q+yr2OqcWFViKjRlwMrDHa+OELQJWmLUurAzvl1BEjILWPcOzKBnY7zoxJtDq4Q3c
kkUSAFQOdHdV7Hwgsa5l2rE5GO5zS/bFs6MGDrJz4unGpuVvqBEqQFKWjulWyzlxjcseu7wAIG10
Vf0X74s8L2ClfH+DSYErIRO1itsv6ELosZIbwvLBaOEavT87Udl4JTdX5i9y1dgBbkduNtf+6z76
93EAPH5fZOXiyotWZCYGII18NesNoJcwfSwLA0Lz4p9wN1qROlcWYyZtrUGYd/boGFGFomXP6En3
SS3dBDt/1Vau2qqA13YBtreADxvR3n1o33DMnjMwN6ofPkZb83eYthBNQ0Eb4QdC7GBXhnXLTb8V
cNZSagsYYit8pXtLzefpYby4Ppxi2++coDSZ3V5m+PCFOK3matNk9IPy8t4fT7fs2vvT3LzfLqVt
jKAFDIudUqzTshea7P2GLL/DvtEPDEjGPric7tbb3O0l5aXVZAKpzFR1+PdEkumoSrSL4MC/0vfy
nCa8H++9sKp0+ISmZp9hUo4IisS1lW/R/GT/kKQqk1vjYOf8dJa4d7xb5w0lEti7bSd8X6aA3MnK
J3wF8kxTUX6xzerrJJN74SU4eKdyutCg1GwWPR9C0i5QUrgMS+LIKB7tmj2szQkiHyIsEcwbqPur
6Uy2VZSGO+WOxmPq3SzX80ZnRDEPSMlvipHv9ShKb14pd6qgBmgovvdn5Ye99xRQ7qrSH3x8XETy
9h+AHQSOjsUC6YM3CZRUGTHepQFxwkOpOnMiVNMa6dSxupgIoktzdhHThpk8ZfEM2C2Vy4UNa3x2
W41m/YW453Q9EjOdLPixQw4g0KkGBodtQB81z2BDgj5UOp/BJCdwdUrtGxi9lPN1xbJgobUpknkK
Cxmcqp3C8Q7kj22DtDeUx5shFoTDTP7S4T6AHy3JV4/Yoajw7oPMk2UGDvh/rSRkvIK9a6RUnAix
CJIacc12YtTpT55JAg1TcxmOJtYaDb570cE1Lj/ADKJdvC4vQdncDK2MTY46hccoQpKBWnq9ubtW
c+NwAbDnm5Uk4mosFPKWMnhtyT/SQopq0Y/LIZIexxVG+NCHSeRxqLI0jmucb8M5EdqK1sfyrIAO
bfwsEqnMjHQ0Mtfwe9NUpIsrM1pfzaBlsTgAaFwa2i0HnuW+d9WbVh2imJgVvyTXnhgSo1KBYYkQ
k5onbfx2cdmSn7NR4E3znlx94eLtK0YNoT8SHd2Gbbwkt95eOSjnmtKT8mztoVIyJXCby0ouGTEZ
UEhf0ehq3RpkHlMOuPbVFJ8nWF/viPM0IAu2PmKYoZxVQJ7YPF0+NbX9xzIdaOEIpJlAqWtnVIks
wNLjbaDvsdXF/qo9+r8xAxKVkJbIhUyI/Cqsii4X8VjM9B2dueniu72b0LCjvAC7gKk1FIwWlcRU
PiQ1H7UHthx0i4SWSp2lYqF/1HIrVjDM03/WBoiomBlao8Ml64XFMReGNe7iGzOGiMWLV8KnnZA2
gCbXrzFiKrZZIvzI65ZbOprDC0mlQ84IZyDAcjGWLp7PQReo0WQjVs/BXxyErqbHetx+0VsvnTEZ
kAIAElkXyMF7D+UNSH4Se9xaa6vriLWYI/BxOM781+BY8Pw8gDGQnn7mH9WdnF1xi9gTPTdm1iII
0No6Ygctna5UfPAAIzpfSndVkLzp7D/m0qOEpejflQKedBzBSE0pbMqtwh3mJULi13ksYoM+YCqD
P3dJFtzvmM14XsxlaaHeHr4b+XMTGP51j48CCLcDahe7EYtU1+lNHDpQEx3CH6anOcR7iUYuNB+J
V/RXpC/n0LDMoVcglo3L6QMWhCvSNk4ONZ0TSk7/NUEoIOINiBXKQy+tQQeKZa1TG3aCcpQNQpj4
4TNwynHBiLHeDREeozDZwpQ7jNjAdOJwuyyhmDWkFrqf1t32i5liIcpiIuvbG1ixVhvOVzmP0amo
tQejZxo+tv8p5Z2w9nJpoeqy8ghQG/4U5jfgr0qYARXgCJs5UpEHVGA3021V+eWtXmIMPnL7f2F3
b+UhM7QKUDFzVdj1P9JIBqyTzcvk0L5g/WJFMRhNEJ4XnGr+KHfSa2taBFrDieT73PTgHoQ6No05
2V2iPqec/Rmcp3cVat8wa5NgTCXB1Dy4bpCcA6JajhfUl1/jAxY4hNY3AfUs3TyBCPG7MnhVVd4a
Sk9QkA8Ab/f4ZYsVSg4QdAH3MoUwl5td1Mi2EzizX1IID5Bt1TvrDtXD4MYXx4XRQ6TD7dhRE+5y
ZMLh00c2tzu9IkYX8bbgieZd6QStXa4VRnZflw0qZV/zs2zjgPpMqua7NgAl3nrYnlU+kR35nYw9
Cno25PXi75nNuiXKkoRtakyP4ugYaOIPg+dNrkDSDH2zQtJ7zdi48TQGS2wQGGutFMrAHX1zkD6b
w7z1sry/Qjx5UDioKvM/LENbNkZ+VUgFsNdIj2ZY4RKmrSL1xsAjTNG+V09oQbzJCT/Xbp519yP4
+nlzRsGPZ0rs97MP9HuXGZtW3fYuRGCQ4u5JNlubaXS71717ValZ70ImUc5Dkjj8W4FiFx1ruT22
moAnvwBT9YeYxtV4AO+mVwzpEevi1y1Ayy6kPzkt5DBnRu6mpPn4l7Aa8zvGVORiKrx28eAqzrY8
wE+gcWiHgMWUjgSec8CYnc3N9LQ3r/c0Ht9d1CA89ulbPPlEV63V//7l9/aV35HByWLm2at8U2Bh
kVuDupq62mIeirWoaiLarGyDxp6Y2WKnQ8GbWzpnF+HQ8HMuWj1KRilP1uhYJVPKb5j+WKRlZjL9
YoYMkvPkgFNOYlZbkPqKw2mMANDf1XyMnCGFUeTTz15gXZje3xZmUtEwfGSja2m7CsSRUK/gAXUj
n1pHpBNt75r7PONiCMchtvR1TpRtHFANljMzBL5lTt5oOjw0y3wQVX78MBwSM20c/1f0a+8eVNfv
pdSBJQBqk57cd3to4AW+M64ooq04838Q7eiULnJwmSlPqkQ8tQetXitu09e6/Ob2+0re+4e4kJUK
+t+o5XkPBOY848qxzF4zcAvDXeuDAplT+j2rIVD61hR3u1u3bopEk7OODWDY54dOd8tZHeBxFlY4
UO6jAA0DBpVfh8vVzne/ii/7wftN+dPCHuCZ0Q2Ru16skmh3hDfaTdnzDoVtGZq1ntGZKCjaNEAo
25v7T/+5K5t6sNEO6wLwT7HFRb4YBYh5/6tmLxp+/hGFhd2qoLyMN58+7nNXLivgKPsaleUOb4Rf
75nCH2tYG6r6UN7+Xv0g3pX9XUeh+YfRxEVju4cqOVlT4zhivzJjzseMzYyEvQU+dz0jI9f1rOwc
grhK4IaxN1o+/4yuNwDN65FFgaUDegOk/PKEzvqbQi5aaUnq8/J3B0WvtFI3lBrXYtog5v4j13uX
Yp4nb66AqXTx1y3Xmg4r0XlLIj7j4jx0lVeKTGrmJkWT/9tX3f8T2ie6j76xq7YvcH2xHQg360ZZ
lI3aVK70tK/Crjf/ia5Jjb2RWLMJ/FUuc351efziL24Udbgz7Kt+dJQLEi8U0YgJIvonuZrH8fRC
KSntmEU44DGt73bnC9tKuEdtX1KHcgiwahBXarbK9qUNByTzuql+WsgH6OXD/gurUOeyxZlNrcuG
Hamg+12eGxewYE8ycWUxYKslEYiLE8bmJrjIqIKXsuOq77A+FIoaAM086BtahNPXqnTemIiKr2fN
8EDgHWdJLWdq+/72VuNXx1HtjM4IT+aa+WNPIoiLf0K5LBtCw+gn3qcHu0JRyLLtOJiPGh9BoBgf
v2fkwZPfcMGxSDujn6KAqRe+sPlOr/Y0o96vmmGBb6SFJ/GB1TYV7j8OAPwo1CjZ5VRUEBJGGU21
r26OQItqOzJEtrEcupvP28cs8PNO1X/uSjc4mXxyqF9X5+4Bmyznixl4HW4VRguBOkoIVPxc7vB1
0ocKPpMa5chjgiQg0p3Rw5rfAFPlz8FLQi1e9V8iOpgNNA5z56OZr0aIo+ickHxvmMAh3eYwfRB1
FXVtrFKMh9qZRuqG3bk7Obe1NZv3ikQ6FDl1rVVfT7c9V7NhYzV7NfEMC1vZNP0ikWtPXuqdpy71
4CKkR89pXekXipBnEbGdoNv6BxrmKLbaf7+q7ujAWkW8cRNZBstNOwmx7zyvOWVVAm9e74Rgq/id
DlwgNEU/PbuiiJOPAvQjIoaRJIzpKkyFeEdIofDGqLOlA25iicAzlmYXPI0UhzByVh9tthU11hiy
2o5l0YGGFgBpPASpZb3945i2PZ3uxwpVNQXeslhyTejqzoGiF2ofSeuyk6knSZvKvBtM4Y2Gc62C
1VZa+dWkCcf68pEg2WihnVRUcZ/WiJBP8Q7ZFpmxmT0UQotNYgQKaSUPXtBfHd/eQ7/sOGiURx5v
LVl8+0wnmqKGjXPGKu9aLp6oIsv4U4sJOmgB+6XbWzmH0DP19PmWWYPZpJ3dh/hipQHsnwyohTz8
2QWI+AiOjyP59iSySTJlzvLfTDU3M4WTv3g2gley0swWlBEKcbWcLhoy0tAeYTayNVIUEmQ97e8i
Ywhp3w8S/IJo2QprAnnCJvR9EuSFYq9igOZN6LkDJ2AqmGH4eElDWNNhV+snFJS2DvBhBMSLKSHo
wdvLWcdnHoSpw6DzafIuv79mIeFqsLyXSG6p3fAq+iHeNmR0oiknrUVIQ3/p8eSPtNlBS5GWzO0X
761s97T2XL4O6be6dMYPeSmzp2XIIUQrvmoHK4zIbe9ZrgoEl+Ot0Vc/cXit6Dof3eu2VLt2iAvE
Sd9JZ7+NXRhU3XVCYIEb7edrc0ygVDAFguDby7GX5XJ6fDL28hFFHTHkrwnhfg2FWV9qEIYnnpJX
qJbV/knLGAZZYc9WR4L7SKv3b+FtbCrmyfd3O2LNb4VvpVWgQTwRIooZrxxSDpjtvdbK+MMwiERH
8Ejwu6WbdKQARiN/t8o1g21nxAsprTTpWNyS/Jm5wxref5ixXnZ4a3bCfo2wMB1KXa0i9ZUSe4Bl
b+xsdyOoDoX6Gxy9SrrZ/eX1HA+2LUmFAttWMc9E4IxQV3L9WSBbtqaGyk6zE1PUt4oo6+pdFwgt
4tUG1devQTJKh7WuoL4kFMJFfyyy4+blohwBUERVuCT/SAefWOYz+0oFY5wJC5WX9MkilUbo+z+J
Ktej2N24SAv76wT9plhOk8htpG0DszZ6DxdfeXQ1wA8EDWcd35w0MRwAj2WqiSEN7/+mx78t5FFL
u7phXnPFSg2QkAJwMEq87UhMwtWM1gfxBTE91YKvH8jb5Qsg2wwrKBwYDVVcjrZM1Gc4U5ieKv9M
TUQMRkcQfFs0337MZK9zY2Dp2vgGRpJDf7tuHKVLWmFJkUb89IJPcDmYYCyqmuRLrHq4mnasXXxK
MGRqThyFWcpaFzUjZZ4sMJx9zYHQygJaRhAtX8N5xS5iFCo73FfKbyjaTquk/MYgK6wJkh5GhhrP
2Kz96BOLwH12YkJyPvmSsqWn1G63mSlyLSXOWIVEcj1S9jLfjOcDY3Ee2jYJmKwjjc/DorMQIE/g
E+0Ai2zycpJkp4/C5kB3ljsUoEIpKMWXEXl4qCEusK9puaxUWMOGSOwpXbuw6e3X/PutSR7UFTBc
M6/YVgCdfbFtuPz8R+ncfzM8OYkmMYlV/o4LjAV6cjo2c1wBSb4Midh0xLbuDew9nsuz817YX4sA
b9uEnGgm7N3aImtaqAb6jw9Ttb5AOqi5yRUKsTHq4RaZcglWK8eMBnHYqwwCrj1mARZ9SjwLDNi3
AIw1cbUW3CwtiBWmg/DHSh8FyCJXNv0aJjx2FtGXmZumdaugVgD7vhOFnxZGDRGHhpU3RNYLLFm9
VJ1TBRIX/Q47JXCgFbmXFwXRONUj0NU+TIDgj9/D07uRWB3+56jpNFsh4c1QUDjjEvUqMje/qoSs
ssx+xVYqQH3vWB7RR8Be7PBK64BHX4vGTKK1gmFS4O58LLoP2DnIMrRyW37YJRsXzC6VgAgk697S
A5NlxAq8EKQlpPqBABANfwcY1LMM+n/c45ybTa8Bj7201PEyUNFo0Z14HhRtuF6NhD5Cmnhxzx7r
75Sy9/wCk6yfLQWqOCJ9WNGsaQj/0SzoPxs8xDVtuURZh5TheZSmx5Ey72/W8g1EYZ/S5/yAs1jP
BWZVe96yatjBUKYzVE5/3PBadTgxBpFTPhmJvNEVXYWW482E4HF/C7knPmJqsSwtOK+eahfPTbq3
AxJsZSaVWAna5ncKshW1FsnBDAz7qXu+Y1DX68UD5yXxMTPaiu4oBwZQZscLckBuovG0LCR9Kun5
o0qyZ5HkTHJXgLRUQrfL1k3gGruCQLNVl5ld3XF335VTmXjtfhhuiuEagErWx+M6Ej/tXQ1tzeWS
5TIgvMOA6WkPPkU2R0tyd1IwfohVsQXVvIxPM+C3yWmqlxIGfjFhjuTa+15hT6KIrieOaSuL9Ga5
Ns3S0BXXX/DD3sTRzsFJcui7ihQv+TyLYVaryIbAFFXvW9gKnIBi3u3WXWI53gQyKrkbBnBqztRe
Hzh8aaywc/wzmcTkAmHH59R+pnsVk7qwBn7n8cnkAjwwVoIXF3bhu+7YkVqXWd4J3O3MxdtccP9W
wwav1aXEv090PORDz0T32KZsYb90wfOC7ZXoV9PxUXaNqzUPs+ueDtF8cEY7iykzwgC5peQ3ngpX
XqKutQJP4+ipcm233lw3Q/OyKvx7HCgLtqqBXpvl3zNeFikfUvObU+qyLgvnoTTz6rLvaklkj4/v
g2ZfNxz14fc63erRE9lgXX+o1G4uonU5iDYm+RQ+a8Toa7SwgEQatYrdF/5JB48/MY9iejT+rnlv
INbZsIF9kd8no9yTzL2qydr5HYMxMictrOWRgERiUaHwxAqq/QzNIlwRdhZkmvpyf7kkUaEW7/CV
cK+7H6gc1mrehpyPD8U6cfCCKhwN1OH77QeVlz5kfOxV9W++J0jUps77pAapgsNpHVmi1v5hFMS/
FrEdPOwIHADYSVz59x1WHrltobKA+aaSddxH87CsEQyQIFNibdVaKCuT5feUXbyVO1wQuupxcagc
7kjUlASaDxv/HbZFboaVo3ayBAdCD9Qcq+fcQzdswU7nT/HEupbT90Ijn8rFTA7LLrYHECc88q+9
pVlEQHwZpQNoX5ZvuBbSXRVKCzYEKSHpF27h8iGcOirFTykJLYtcDGerm+0Lv81VMyQQyjbw105Q
mWZ9+x8y9pjpLzeAKUbKMPytU7eX/xxh+FZwpXn4kL81MfMUZOOe/TwWIl7ro6IHhY9RhazGZLh9
ao+isBOOkceUdy/Skx/wIOoTc/p7onCu32uN0BBPXnL5xyhVoHu8A/ruq4bvMoBSs51y5yD6vjfq
Cp10W/45wdmtWeVod69R1Bgk4An5Uf/qN+KC9f4I0C01GK0vTHR44+SVPeQXsydNiHbMNhZaJvmQ
i9zqZHTg/gi9p/HIsZ0unJ/QqX7lOPEEfukPEht4FC95y8m2Dix76kwO52Tj7V7f+Ety3s9CXY92
kAKTGGTxGZ7GQqtt0Ob583dpGnCZPDo6I5bMYR0m8c00J8eXAeSmEucwcKGuSWuHAanoMdf138Mj
NNVfQpv3klbNwpF2/uMmXourRaxVdgsKjP6nHwmysvgtxLrmsTZ1NhsRIV+wEhpiqpDgQKSSqBuQ
bzqpMR9t6LcOsFcip44/afbXFveU6YWbcwjRU+PhvkWH6IZHnwXmr046vIXrF9lBLgccnfVEx336
/tsoxDbQDtcJVVWAqutbmVc24N0ciLTQ3S4GhSW7kT6lqNp8PXqrfIYYrhQXqrskqqChHolcE4Hp
n0g1Ueam2t+3uuzImm1s9wk0cUY2WlSpCosBYi2THnYDsv7XdY+VDxgQndWrKDPer03+6UsqjH5Y
4/YVdTtQhLeiy+AaFhKZwYZSZbMLIpwYT7MYnL815hP8UV+ZhI2AkzBpTf6THiXBrHUkhr+hHs3Q
X6ytzbvqcg6R0LXrfwxS/HeiOVaZ99OMrIruN95qQFKF2kbZLkt4MH9GQoXi1Duv0xX0Wo9AkiXa
echxxDJFEoxWepw5/0AIhzeyD/5DGpPSC8tOWYtPaeD3pgxzdPIoNNnIPgdg1GU+l3kEsiqF3jby
pd+kfn3oByxId51b9WX3YlyPVLO/lN5Dw/Dyd8VjplKSvCVKYGFzQVKbVuTr2wDmCTMtQDo6zJ5B
8FdcbzWIObqzTFl73METCqT8sswcXWRf+/+JnlQ0Hddml1E/jTluXGorM+FTQh6+jIfngNIRUiXv
aRLMR6RFs6mDVw+xJWNvWY3s9rx4vdMqsMMKu3OsTRnBimCjk7VhFmGQ+tvurQPcYu/CEpu5pxKv
vQIHxAQ8BeRdL24lxY8V1fU5GzreLbiQQlQzRgi1QE+Fb7DSw1Q2vp5BmjPRWWAk+OHsMY1rRT6u
SZ3DyH/10zX83ug9yQAZny4Ot/sz9azex6HtGsJza7tzMyZiDDc0bvwDAKvpop6f1Kix84YhxOcI
2VXHL1EvpNnFuW6a4UK6PYa7AxBXxe+YP/oEBNlwX/qMeM829JoA2rcO29exgDPfOpomP/b/LCVF
7kaAq+KO/XYP/ty8FC3CPcgnOFeFjZ839jI/0//nI6aMKJ6dak62DxKlIR9+IUB3pDv2mYvRTs1O
w/3rCv8i0FViyCtdmDYMhjSPNEBnz5O7jk+jvd17vsoTpNLbYEZ6wW1IbCMzbwPotNCwSUWShkZ2
v70Y8hkmYfnpaYLLiIPM8dWUiI0zP5uSUyMbHY8xmfa+sXyRhn3BoUsjkVOI94g+Ki4mx8DwvUSq
mWHYXF35gQPGYJGYTO3HgGiuugsePgExuP0+5i4ZrnHdYTYLF9Amv1NguxRGpDw6y/7EYg1I9TB8
aoLMKEqs9NSA9vNhUGCZ0shlGiOaxsPVIUWwX20SOa9eT7ZAG3aADb7MnqcTxtFyu0so0A0zUiIG
xcbg2pUaTkt27C8l1varMk5lyabPvuV4dMuWviACF3lwKx+A9jwWMp6VTSgzmuYNcgD0Rbj1nF/E
eYn6JrYYS6epUkRf3Aw7HaL7pc0AzHQU5/AHn5Mu+G2KyQVw253+PlprNxlnG9OKKrrMLQvZWfut
2sSuG6DSnoTOiHyw/vJEchWGdpbr3KaLCLyEIp+exMArxXtIjRBaKJEKcRg5HuZ3y6T35Ep2HRuo
vDQauGqr+u0ZNbAY+78sCtkBCpd0dYGIYkF1L4kyweJP0vKnF6FFCfQznVx1qCITXYmyvM0xiA42
CR3ngLcwPUyX5F+JwqRQTPyhMgV7W9pr/1VAYQkJvQ/S2WO129rUmtxPhmJKTJfTE5nnoWR/kPag
xcg0tnIuQEBux9XunGvWiUEtIV04BlctnAy1wteUEuqPTfTWao/Uzs3ZplVRzvu91C90ziCFQYSi
GwvnyjC0GiJx3tMCcd0YJ0ncfAfqEKgmYjB9q1i/YlRv74MXZqrECltL9wDfTnLGnHftKyI4jcZF
PC9njzl+IGEAu0VAydJP/dvLkR1C/9jeNUhGte9jkam83jfemIdX2bEuqZIWSJBqlbrlbf1xBGGu
vJ/1aCSb+ANBYRaaFFmf0Jk25eLlIK9u/oGoVvHFdDqOcrmvix54dMxn6JnOvZshfatzvkWIJom9
f3Uj2r8ddwuO9koa8dbnJHbvVnzDzqZJGcNTtUGV1b+zC6sfVK64dzqe87yX8LCxi0VSRs6Sy/Tt
2UvsenBGsa7OUWByLDF4pwHXge7Klnt9cA0++kQxEcQSl1eyN9viOhql2v7HMYaZJW/LQLs42pXG
syRK0lrwloiT7Ty21+3DvQk7IJ5bAwja7yV7Kof4tb6G/ekpYgeKWsg333WuIF/G6a+ujG4gneL8
vl8ntO9KodKOq1hN8xhLipHtA8isBKvV1SzDdUR8zkeJooTvEND2wXrR/l4wPkUrAht1VCem/qLZ
gAM3r9g8Fe8H8K1/YcIsu2WdVicPtSqsrdocsnWZouqChk7mq6T342/SFhO4Fa8WZZr24t0cQiWY
2Ada2veqEsn83619myT8u2Ad0lGN+PyfZCpEHTc09SYCKjJChzvnkj7lZVhyxWZU+iSPrYH7hx6M
ibCfdvEQ/niszkT8F8OqYnnDTpyIFRHLXZOXrtTQw8kJ7pfcXmo0OD1Lj5LU5b42c9vjhZq5WA7n
UbovE/2DvN141VWF4d9D89UaWPQwWxyUx7OA1DF2wFrW7AJZCdKxQSokNcZS7KGcBakYd1+qKXDM
Ny3fghn0xjg6iIyM3muHQteFx9XFcIRpqumHQRktoRzxXu1KTUZChp77uVIb9+wtvCLv1s2pJGBq
u9JaidtzwVOLMwS2VXdfxiTctFgjJhAgj8jtvilswEe1lxzbsN2DPJ2gP3XSk+e3XkvOCc3m2hI4
DuztTwPwkudNC7jX2GO3l9mBp7I28rqzg5chi1EoBg9oG45n8vuuw44S/a2jxJq6ONGms55LKQO4
TSsfVtxARrYPYDmrtqhUvZB3Rhw8RWfiA3OzkxdhtZ3mpEssTllWmKo+RBGBUHsYQsAKj6r9Ffva
lhjUM0f0BBLu32KgNy7NnyvsqI1ftGkWNduyslXZ4N0Dj5K4nshb70FvJQB7/CTDSCkpsUhyN+X5
+5me7M+u/CbSSQsCvMwibLZkGaiZljgvWN4YArPGcYXQll1KKZPl7Ln6WJrftdl5eUZKduoEQAfY
RnrWKsG14fNec67FnFZvS3t/SIW2NQhcTP4YYPcrMB5Jtso9cWlsJVQVCfZV5Jj9l8ZcL8yXGb9A
1AyohelCN+nCAI9PpSeWSLRlveTubCcFaVonyDJkubWppUlXA9MAxDp21iY9Sk9HPcpaJpotV6+c
oBMsBBPDtL3Kn0A9ysJaCFypO5j5vVLmuCPc5G6MdtO3K3kIhLB2T+l85R4zlfntI1rJzUAbeLvR
Z7XDYjVyWXlj9b2cxz4mOSFznb98iaCLhHdK2pIiqMYl8oXOzEldRBKxi1jzWl1ghWTdEiY4hQcf
XY717IAYJv04U3xAT827eHx3uq6q+TmH+zGxnNmpF7Uy3+Df7fSFrKLCtICs3AD3wNk8lHSz6/4M
L7IqdoSKL057oAno0f0bSYyz51sckxhXZ1/iVAbawB6fTJ879oYJuD49l8VpLxR1TKlvaIErerrl
Xi9afwnCUw2c37eESOrqj7OcvNIC5ehdmMHeNtLiTK8VbuJPpFwDLikhLH4fqJ0hjBHuZWNq6sKa
p+1ZlNSmu3u6BGIahyhz/LRBhyIa7/QnntDCJcYprF7FSon7aFNixvEVcmGbUA9r1wavozZ0LbxT
XtN9qgnQiFAVipAKKlvpXH2XAToOxbMJeY0SsBy25mGjoPPu/HJ+azCqwHphRAXEml/p8q9pG7cs
IB2FBl/P7AYGUV2e/EyDBtRBl3uTz8gczUWSLvyixocJ+d3Wa8l5My4MDTASBBBJwI9NX4D0EGyo
S3XfwLEnfqUyFvQIDrl1GMdiPTZCsvU+2dN3xsGzGLDhpTjCiNln0CSPGKGcJ/ZoEpG3pEEMfVRu
L+b4d8iUpg9DOB7SS1TsctOzjmSDBpl111Y3gTGIDMwt1t6FYsdrxkGvGmEsryvFJo4Idd6i4ByT
qf3rM447e2HpXY/oerSjefdK9iWRBT/lBXy2nS854qSvGYcP37bA8uuqSwrFqF1MyFFHjXknA8Wa
gz6d3C6zG43SQ394KDH+8l0iaC4PQKQ09tWp+9MKGeGIJi41XlGQKe9bCyw10O3I56jMfDRTpQHx
2w3SmiszfylwgOIh4INO3Z1S9C0ESlXZvxa8Vk1XnTksrh6hPx3bEUuMVj6mYkyK8RfhkQFh4wv0
JF1+rL3RpcedMgmfCEz+R/GgkYLgzh+ZJDsql2cJhRfY6eR97Ktgk6JuKBpS4bMQlTEisHmhWCUT
5dFBGr8Zc3PQLcBO0FLRjwOqvwfZQKP6z37DEDkbiFhOUImSna4jcHZKwhZXhj6d7XknKUjQpojY
gg5FZPVzfeaCd2uSt7g/Hj+3tWiSG3qY5LlibsughpLZaJTIpAdmpEd4xqrdoUHP1GcnxidKCRT4
KTlfJVTpAfVWpSq0ZxnqqaUjNxAqvAB5/w//Glb1Pi14nEgQiLNso1eXF4cFeDoTbP7ED+iJMFeC
4iOCXajwQj7rq9iilY58GV8oi9AMm5M2dmZQq5nsEgxsjT4MPIHFztHtl63tEc5XMGX1jhVTQcfs
grp4x9NPZTWnLvHUTDJ7IhG9llukXJLGh45/j0eFRjNL6pMg35nraWXsyRc+ME4bclR1Rb0izL1b
Cu/PRxjbzUl5JItTJ8KQA3nutyMdT5k1xjv8Yy/QczOzwtklVAaKPfry/SPaDJBVwaU1mVcnSZAA
RYZdobFBcNcBepvjzNiCPcINhCId+RYxNvgSesAJCUTlIqyNxL3RXloI4RBHsKNFV4H4YSiiAsZx
UBrjABUJbhv9QZe3ZIaNrQf0vBvEM6JDKD3OPGQq0KrpgNvtCX1HzvkVRri6ADoDwrGQjT8EMXqD
8Y/aUqIU7ZQuwVEJQhabDLr9UKw6vSBAzHrady/Iw5Gh7C3wwzTD9COnCuqK74KewTClpzMV/yMG
M4GsLfPIbHLGWmucbVkPJjKlSoLSTWR0KIXUiohoR4pQTFUxwlFGcAB5Gp06hNuDyyXRRcDGATGj
6P0udi5Eoh035OARbjl3mkqlb9qibruR6pBjR3/vOF2ZCkVVosMqrfiQhAjI7lDONQt9GBHMTt3s
Y38F0/3hLNTbW+GFf8zj9CrgQE/uJPhbiRKwE8zo74fPVxjCSrJ6GfjGHjBnmr6FknApfiKD4B24
uwrAan6HLs210j2tEBLhE66mfqhcZTDcpz43q7dx6UVv59J6tHIW7Q+TKYs8kar2DEho/J9ohDJc
1VGhMAII4ZMKq3xpchsXQ4W127IqMWz/7CkbIBRvm3nJqQYxB8swxAF6oeqLMkJIgq4J1NZLQW7Q
B/oo68QRz3No+SNvWIlrZB5l0xh2oUc7ZBGw+Bf10ei4sRM8C00tg2e3mMyypOcouhV6xrmwUQ9O
rJ8taxJzbF+Ia8ySehpxawDuLOOGqk6C5P0V/2qEEVkrMHLQjHwUKLL41NVhQ9O3/NVKNZMdJN0p
gXA7u1AWeNn7TFBXqC/n3L6+niGzgQ3YrzdHDOksYENTowt84sIugVZfoc2YsPXDUUDR58oU4192
Y7OQKpYUhfIZwpm3npCO51Z5MVFGf4Rj5tM+4NJif8BKuzwt40Ufo6QsrRUnplUi1NsFb0yOU/3t
P9XT70pXPGS8BaBJNIPp2TQJOzuN/4z4YwdQ97gkNnwiANDK2Syhes0XcY7s/RAhgfiGcyz+PAIu
Di4MYInm0p4a5F//SOPSehZAfaciXavBcUSP1KDMBVVpbFsmzjtJWefGdZe/g8PcclMunbHapRcW
eGz2KdC36pqsYsIw6dADXhlPCm0Gv05qqEnhDW/mC5wWw4T5SCFLs4TionS0Bdc6BGUnBG4Kor2L
GgXECY/4MVj52RJaJswM6VjAFiTCkMliZOb1C+NDb9LAQHH69h5Lp8mRjno6UMhyHCm6CG0QoeEZ
fO0jENRDimSYIup9G5QCwzBA1GcO34e2KJR+4xdJHV38QrRo5skmY5bhXvrv5nEJrbntLlJBqH/G
mBhNCR/0zuw+ePwlwx5t48yW+nLccDxXLZqW5JRpPrdhSvcdo3fh0/HQKsKshkDckIDTOVZSgzXD
R0xi5MphT5H8CDgrHnfwF04KMvTBFzEemyFEYg74WAkU0RL7LHua007qhC0XXf5kSqATvAXPLcX2
yLmX31hHXahyMLg2YvOJAvNmiBmFgQYVx9u5FurYnDgi8VbUPaTMEo/Iqd+pwho8AKzXHFnLObJ5
Vi9y/WWdPmjAPIB4AZuHFxf5+6BSfS+/+Y9i32WLureU6u0NpiwFP/5CQByj/Vna0mSqM+OZG81G
0kaTulprndnzuaCnP9yKuGoE+/27wze9c4P5knfZFfX8C6p0t0xxLe/wUZ0WZBzsbfzEqs0nYvn5
J9Une7nF6wamuS/RKPvO7J5ysHdq9LDvweRbrjWyDE5Wdo8b6qt0t+OonPA7CKPQk8oPdMO/Hney
ocA5Nm4cC5ZIz5YvclWgqsfcMZ+YXbvBuphRM2jd6nWnCS/2hc6ptetDitaIC/Yka5EF41Hp427M
JJ7bck41EiQRGuNnk0AqvJLwFROLxFtfUcMr+t3YfAJQhPXTeLbtxjnxJlUIZsfoi1Vr2su6Wadw
OKSlLHjD21tGXW0EzU8sAOCn8KuO6Xc2m4YGmr7b9Qi+navfxkd3qBNRQ4J2TkBuGzDEf5256CRL
Y5pmobjjUKNJI0RS1XmBwTAs48b9ZT45ZlpmILlQf0+eTM52ybO+nGS2hDn7XtxvMulrvCtmV8Bl
/T4sMW8rXTn64bdjWOB+3YgmEAy/7EykimdES+s4a/07BbUXeAFWkumoriPdyszn6TyRXCscL9pZ
7KCssM32Bgk8xDGzI8VL48b49emJKKq4yYZGu4YSJXqm0Ww9Tsb3rg/AWUrc7R3RWt2HVBYj4ZeC
h2ve3KgwmuCLU1Soof4hJ1LMlksp1RCrZpdJjhGmFI/z3NxS+FoXfjLE0dbqG/0Zz6QWdbtUtNCB
0GtNXftw4DGT6iz/Z6i3i7zF0Fon+43+p3vlcEXgTI+UBYLBiK2EQon3cXzdCPqFs57pmkqHBjKN
KikTGAnbs2bLdnoK5tae0aHihHqO94bc/DdRVDpN+XBh2hT+GpAVuOgNr2Xn9Ag0miKr4jgxhPBJ
9Gji9BEYUmQD0vHHBpVCf+o/tvrMuFqT7mUqmPv88JC2DNCHRq/Fys7aT7fa1oHPaofe8J2GwBCL
YUFeKGp5damywk6yjOlmBR4GsY16pLUTDwMcHIE3RhwDmEX7/usXzsYZ6eBnRo0ZX+HXkQkXjDCL
9sFKfb3sGnIok1VWjaJbQMxFDVMMa1jE2e1HvXaTq/vwqPudv+8o9SNa06ilB0n+XghmyKdQ/mxS
Vg/EBUu5zRUQ7xDfs7fDSTcjE4iZuotVcieWGgA8zquXlT+/ZNtaDaXxx3cyMDP3KiFSVu2pyrAc
8khlKZSDrMcbQ73wqu+t4InqOHv/KzMTRlkmfD5Boswb3qFijqbltU2bhgGd5S1vBfgPi9s37oUU
d9tiBx9rje59wvjQiKU9qCgp04nx20FXoCMBCwoxDMagKg9UIifZ3ic+caX3j3FvAyg/xu6EcwCa
eanzFksW89jFYQK75pnseCH+RsrG+kjjOxfJjBShX2A1rGM5NWmNoeEsUtE+hMiTDP7FNH5PKfgK
eyPPLEDSWFPVXxoqDstnalkfz6q8KVTt8tTlwae0jwuhkszKgkWQfdEQ8I/TjVN2XwGUEK9hBOkG
J4DPTGbrydoSNv3hq09CxDRrmosN+tg/Htin+ugC1Zki/ImM4R5xCGZVCjWfpa3AdvFLlZwD7TCq
Ky87O18c7V7AiwasaDI1yURw+RF2eI2pxTIQtt2Ev9EzbNibXwNbAQ1X37LkcFlIcbDQ8zwax6AI
DwGLlxGhAIk1BPTJOrzsdI2DucjqnruTuTQAuPZx9lsIcJhHI50FPqpB2TdvZH42aBkXRPeHlnaN
CUyV/C73piWFsy87BIobiacIVqCk9KopOp8Fv1W2TyqWh0WD6tPXmXQKfB2FMHb1PZCC980a11Gk
ihWvdjSoVq1BHGa4OLcLpMCJD5jEUStJepheXDsCqUxUDYXuNK1WvYKzQVQ1dpOcJMy9eGQWNcHk
pxfkavPhRqvq2K9A8l615u6XBLvLznvj2RZUmz/GIaXSoV5P9MGG5H8wkdz7Q86ogJUxI4kuRnAz
FZpBS2KNkFgu0j5NEqSPcQkqT7nF5qsRrD95GD8kMjS+WZ8rLcSPDhb6B5hL4uIapTL/GwfxTy+i
MBsHPPlweYQOUUDUVy3Yac5s/30fTRPPiHluxF6GJFOhc0Vp0qS1DM44w2QNWCuSfCXPM8H2z5jh
cPTPZSKF504N+Yh6m2oRi2ZGuOKrSMsPzbI5B+ATY988Tuqk7JFvK7SfIg2vvVcxtT32BX7uFiR6
aYaMq/Sy2nx8F6892e8Nh0pNqzQULl9mSCcGr7jmx3YtAe20ZZfcGKmDPkD6WHi4gwWhtNJcFlz6
TRIOc+P03m8+hKcY32BXIWYBGawI5mUhQWVMuvfuJIQk3I4z3uss5QZvedpcThoGug+pHFycgzyE
q7AdH8jCVZLOQqPOzOB/OlIFgx5yMEgOZ4nvDdb4URBOlBo+aSpOpcywr1HpLxxTBFLoZRs3Av12
pThVpXZQOkmyaLJ5mirxqqPDwMsVJlkimp+V7SMco4aTO3ZRh/CPbgYVwEiGV1TUFPCaWuj6iV/S
6h4xKREwkf6Cx2IicQworqSt3y3CD/nqacebsZgGcrPNiC2/lQslMvuAVBwQJcpCtFRpjSbUbl3Y
WgvEwI/TFj1FOBm9dNil3lBCklmXNdviurDCkO4ug/qUh1qZZ2iXJw4hWKLoY/0EK+eBSM65ogcS
uLby3Z8Vpvq65aMa8Bt9g1zhPtLMIJgCcihlWlNJ+LRrA9RSnd7hcJ+FgBlnNktWlkbLkrK2fxnJ
eMdrJBjDNrG1SGjpw4Z5HPyIW5eangpoTzg3S+W3Zod03wvpuvehqYMEfT8mRw0Fy26Bm8UtP4B9
OqmgOkWfF8caCn7cBrUgEZR1rlAgTIedMOjF+KWmM5uMqGe3O3KxnMEV0k9RLAEZl5iQsVtNImfv
mMbrv5vb6e6SfdMmijP9KKx6tnAz6NrRmw67DOK9r7zvJO1gXFvCL5gviS/s/09D5vhP0wz2X2XP
PAFlfEASOl+dem6MPfUpWmW5vDe5NOjn/V3cQXecXxkeh/by/v3g8aX/c4WUXBwqydNaKSDGL+/S
ga/3/JtXHQWg+AX3phyDDZef2l5bVigqCRz6lhdvsWLzZXf9NrASXyrYfMusFVUdWvgTKuTFaJ4O
mGHn88Q8TvOtyHGvWtAJs4oo+qBxu1DL8uVcCqwxL1uQVnS8Naa4S+eEEHWd8UmIjobZod/s0bfP
uccFz4SPPE5gZESf5FNEcGX+SbECuICzru2PSigcxlYZ+iK5gQA8g8Y8+LK6PCH5qGloAmiR2P1L
+tB5ZM4kNlCBesjZgctRyGm9Jk1Ww3almEBotA7lPK8eSRkPFkP/dlPa2H2ukyJYFygIwRhg6qSM
EwK5EFP4XKWT2RTrm89hTTFaEzaWQRVkMmpEWeQuh0tz5dHJg69pCUpdixUxHWXZOSmpZp00X4Tl
KV427fhZLDMHVYbaI7tPeAYdu5AtJyotvTOtcBaHq7S6jtyyg8Q2nYCZTsSAaeqvbMAT3E+BQXtq
UoVbz6mUUzf2+GeEoQd1G0lsm38KFf8aSfUIZ2IfiQkzbmt9VMz7lYlXznyoJyv2SrUPKhYxerlK
J2amMYvcO45ikhXHpRuqf6W/V53QWs79AL8lsGU+uWVkIFjkRUldeiTZ5WZRODMKCYYOmObP4Dok
k2Cn6bagrP5O6C5CvB2VrVnAntEeZvKvoslF1npluS4Azbx5OzxBHZ/2ublyamSnkeuI2P7+Ivwa
2QFZAngWbf6FxJGWbFDepTVnNgi31ocl81xT0Gil5arkiBH2cCSFCzXtilJ3yWVXoslBeCfeGvdg
gA+QdS6Y6rWaYRdT8LJZhdndmnqXAAhzeER+C9urLwUOtAygj2UclXMHFuJ6sUiuUQEtFk9UI0JN
h0QcrLI/H9VLpilqPHMviGqbmCwrthDc/W7rV9MLsfSqpZRj7cyuqKV4jWC+5LJrIBjvX0EoIcF9
7a8Tzh6VQs0sUjF6rDd2Jw1xzsnQBXCn4RAo8qYZbQEj+KAPtmOQp8aSqEhTob+hujq5WZjbMzo3
IcPSV+Hu2Mzt5+JbUA386s3MgY6otXtteXhsXgqVuiMZDE81564Anp99LGBztAwo1ImoYDozdxui
gARFMxjb+WnpK1f0eU3+anF4hAg35ElCUGLoyMq1J4W0kZM/AvoAAk8kxIi98/DMhHpx5ygmC3Et
Wl6fl/W1ncV120jPkzfEde/arSFRa7o7230be4GdfdQcqW2A6tL8Kbe0DPwe/he66+tqJzm153Tq
JVx3DnYZ8g7H6GGH6rnUgpZaI9WUKBZion7f67czqGJeZfaaUp5tyzQF7bZLzBsGxVFH7e5N04Vb
93O/a7CarMr4H8TC3lcRK6o90fjthBwONCU+ryNHMfj1gCR5Aa72NnQGbYKFSa1SMjtDSWDA+CFX
uN4hrwCrToKfBNnelPj73nRVQxxrECC4YERdyIzE5EIcWdDJcaCwAEOGo4OI+85LUySmvk4tG4Ad
iwwLtwUhlXDkFg7Wzd3tJZHlPRnwqJQM+f1s1gaxOThDl11+0B+rMoNy70I9CYBOR0/sgEkVVZXi
BAFADfiWPwnjkyZ43upojU0CNN9hGE5IV93b3YoRRkGAXzisKqDAZpIz2Ou90Coh1F0QAyPGIrOi
CqtbjS9wKylmhLkEiam9Fp8/Z5PVDYT2rLgjhEIngNoI0KP4hEsnYQcBQphvD9uTCR69IKDF0Igk
DGRxvUcx1fNzo6UdYHfrRk+WQAaf6J0WY7Et2GK/XejxUDtMFQfT+hZRV1Q8Cno6QgfKWInaqOqE
2mIrFCSXodOye+bTwtwoKPaNsqAMst8S0/HhUDj6JchjnCU0RpcppnHfY6/EwXauEUApmMtiQKS6
NH4Pgd8paNMYf3EO+ym80rIcuIhkFSjfh5B74tHW+OwkRD2GFAyQ6PY9CN3W7eVfGP6tTtP9XR1T
2JbXSUubHB6a7Bp63LjiLHQINlNCPA7LECYPNMK4IWO9bxa940uZ6yIcadQMHJuc0U9K1U9Orics
nN5lKg33//piWVNAUmXZ7NbDxvN+zqGm9S8yMsavc9V49KYEtm9OJOm6hEt+r/tsj7LQpTdy+4ZZ
JKTvpLosR/QOaoLvpF+2JnyCyRWvWhbFteb1JARdqFZKVdG0axLAfr15vFb4NUTXe2F3mFqlIwig
T0bqenzl6BK7iRpxsZUcUzc0gQepfK5K0bPmfk5GTOxdxSyDh/3YSjUQ5qaxfoXztUf6/5r7iymM
VXdUTOgNNA12y6YHRk3PQcpZr3Yq2AGvatdjOAy1uN1gBU0gAISvUgPAzlm3ZqsyXb8ZpUJtGyFm
B+O1e5zUxIOnmL2r0ISPCEPNBawJ5K1MWteOdddtqq3NbxfmqBqrFYVfLKl9bqUwXuyWCiBS1ih0
OeTa9u9C6dkxTOMR4SsBj1Em5kKvwvr5FEXKhBiy+JmPMLRG6dR+S+CuYjAY3cowQopYmss4RAZ6
Suh/aT+8kXiwp8E9wp9yxT7sWA+G0mHVsdZmZ/1kEdlSMl0vQZEjesCPrGoCIAgW9LxaKBWtLa6u
PoznN4Q7U40vEKkidwhkQKGaNqqpoQ1fupllVxthRgjkVrQSr2CgymjRuUTai4fBzrO34LjJ2osQ
z5mbzUJaIX3O7NF5Eyb7Pn5bkoYKCzY07X0TTqiHfhuRXmxTozMJvpr68oEqi/DfUW4Ii6YSmxez
4MUsxjNaOKGMjYoU8nsTL+YHAbE40zGTXBFvYNNqLj418Ezeh8lr1wt1rCPVSm01es9MorEIZzbW
INplI+pREYHC3km//4CFezuhMTcMCAd/0OqphX5Pi+JICWjDQBs9VNZK3GY5ChiyhvACzZZDe9Vo
79birrVupcfQ5EH+aTlhRphk+V+iHmolq1KiiFCUIJ5W1NZXeCwROfHi+ufFA6SZOsks8I7+uS7y
NsP2L0W3W/L3sIFPDpt7ZfMPeh2RjxAQ5fLFojv2wE2szTHd7Xu3RgjBJiQHKefgrQRnGnQjYtTo
ddRcVo9GUAlNcIv4wGZ1z7I0/qAea6iGehj2zqkqrAyytaLkedcaLenodRDPeVcoLfI0zE2hXZBO
CuAZ/Ae/5lsTNXXAqH769HsfOsaxVurteSfwvoDC+uTZoBBjhfro7rlVuThZYwfo3VkjccwL21dH
4jdWdExM6VLU8ivQc6Xohs1JVmq88+7VgEUjWnIQnc9inIt4bHxHmXyIteQyJQo9dMZZCWphyDva
O0mvj+sEy4QLNXnI8OXWxFRXodyYCrPToBPvUr4lv9s9zh87DusQgetWhoUCsmx276yXOqTTsAwq
AQNi/0AAULuvQD/5suxFtmtkl2jqCdwFuXdMvskHqhUXr1vHc5VYDpAtdRpC3dtb/Mq2lEsUeYTV
xGOlmMZ05uE/IUmuCsIgWpS+8Dw+Lq/lE7U1rLAg1M1CCuUWLnplsm7KU/cv2eSXbkbsZTN1IAje
ulfg+ojyvWS/NTHEneuL70nS6pCbvMtmtOXI/AFvR8gZi6uFu1QzQiIwnLlXJT314Ij/VIAGyK1+
W2qqbma3l0dEX/vkRc/xJ/++LUGpiWOxJ++twcmGgxumoFeTEtc8+nqA1fjHSpOHxZh+rccr4fHJ
04eEP+pkhUVy8TPYUrWNdxHfY6czJ7URcI+eRFfOe6KrbVRzLAqD05rpMACbmY8RxkLKiWdmj2Lx
ToAchWVV28p/bisPRMa+Qa2AXI8pbwGUFaZBXfp0AnMLG2mOcwYmnqnJM1MnmUHwdQUscwAkD5pO
ePLlyjqYAnixcJ9MdU+61uGWJayXB1CxMxJN2tanz00uc7wXKJ2ztklezN6mty3D/sQ8SKOLQl/U
XfcYYzn2cCJly5sswCilExh/vh3DUgnuTOfWL9HZ5Hvff9juxUqzV/WxjSK9HCI78suX4+DTXVnJ
1G3B0mmRPYDZDm05g5rOZGdo9E/kZOTHTQvU/SMGFXC2w5Kr36AQ94f5NNL91uNL3Jf9kGRPGHgD
NJj8ypj3uEqBqPHJTWw5Vib6L0W0xw8/KSsJbAukc8GlAHEAO1IxWvj0Anpize/Xs4MExJbdTGfj
UTWFX/EuaP0RgKhy3Xo14VGC68y9AAya4AHmNJSvg5WsBk4nnt04hswYsV9lY+7o6WpAjdHvpjXP
BJNYxRKu9H5gzv5lhb4W/gaglft+dqAzokAhvVBKZ+OFdVrXMyBxfwCs2/yjKCZV7LEmyGY7mNEd
tG7IY3aB34fE25Maz3pzqjmzDD18yBdA+PgmU2yOQRUx9V3XE30sKNT2TGbVMVisQrzO+rgOvnTx
ye0jgb/xZiPyaPyEkorj4jiFdFUFRoQKS+KaNZf2v1lrY0/I2t8ZgZY9Q3QainAMAosK7qe4lUy4
aOsa4f4liBGbQ7dWDKyyIy0SmJ4IRQi1CovV3keKAyXbOO6K6VcW5iQR/UY4xlUu0ZsYRvNqJeEF
nfABm2Ft6jFEKYwyzmw+weNbMzo8CO80WTqj510kph9SMe1cnXL+iG3Tn5eM8QUnc3TuUaFc83Nz
kegIHOJI8lxJSjezAQuYBKh/aIPBX4lMcLaFVipayrufkuo6aA3Z7lgHijgo4vHzF0u4mC59drG0
4AnRepsgP721VlRvIv5TUjYCESS/IEU6H4AJYFuzgJxrWGG7jLOVVLpLg63kyMP1qMTRsfsNaVfc
YjpquOgMJskI4zYUSMaTfAXr2VKvt/lM5BRZEWUHUW5AzbV3TPjTpVedNHETVVJEjTIVzOJn9v84
UGvSPthUEP5bmp0u03/pGamVU7LlrHLLB4zfv3xhvejomTgkMbdyUYpQ+nVgWUa2XrF1KkaM2IwB
+3tmh2orXZS6MaqJiEyXwfVezSBMLXn4+iQBe7Dzy52hcNM/EE6L4PZHOQOj/nwV7QfJQ1sQo5DE
FG1aVeyAloxm6Gp+GueEzUSqhIDF2yjcA7nMAX9pWWL2ovmJ3YuSL8Ar7ORwnwApcZjwpO3kLTCi
x9CB0+MqnpV/mx9mOXxRDPP0JRQASg8cI6zTFdYylrJQfrTXKhUDlXLTAYtreMnpm2WWUIdOtFxF
1JzmDRSg96QwE1sKBQZhrAPqWa9LxjmFBbBIgsLqg4+ScgeddyhxegqQjSLRVrcFa5p/voHPOrWf
kmen9ZykoGV3omxTjApA7IWujTbffjmxQnD1SVO1kZVYdWpmMq/Bu5ZmRCT6Uw5FrrPtEZo93xYh
WYsSW4NVYlZwvjShzFa6xuxytlwE2tNpln1kw9X4bHbxuSWWeOGL253/nju6A09gtPIMU6F/wnPC
hzpIAvyPQo2WH0c976xGOCJDpsKU582ORb8zViwSuFkuA2NZv03puhef4CxDwJfxpDbUwrdZhtS+
cCGnb27X733B0bxfna8/FdbD8IPfCvNQJ0KGCFxvHGtpKFUYUSASF1YZtMJLQuPLzNWAOumtut28
yEPhDKb6+LfaGYIHhH9k3VM/49IvAVHkG+8LDR575CqpORacrmMvNJknDkkN6JTeX4TdzhXqZ3Ea
iCCMyA02527b2xiLaWokKGWB3PmOT3EzqsswKjnqWVyEIUq1SCmHtYMuMPoQ261U7LpbPLhiSlGM
DFfWDtrvjEXaVaSi3AFVgA73kqoKtvc3VxNbhr/Ui9bZwnTOXrZQIGYe+ULtOTCIA1vXR9hwfX7M
wYKwBE/NOPY2fNrcyKxi3uDGzZd95TFansHf0YAmNh/lD45oH+X930x4J4B3DVJ6LlPvYhkKxzTu
HKralOQGBfMk5/cekcyv8ppaCxzH7kWbdUksNqTv9mjbEafOrNqT2dYm032KYwWeLdDuR6R0ABGC
A7vuUvdfJp6eeQkZYo2Z/AMoUQM0xCQ4/CEc4UBiNYFNpuQh3DE0jnKBsyxtBhSoDuUqGtnQOyoO
/kTdNf2WGcsgDALdUEgc+oG7VgLt76j+9XFIE+OC4G86x5abzsKD7FWDvZYZJieDaahJSZlhprBd
klofUXjSKyPVzqEyL+MpEnay7SYfI4URaTHTLzrNshjoB1pVE3SoVN9h1TA4POiblMgO6lAIVocf
zTzf1kWJDVqCatygSxjMJpSuDBY3fNikhpIQsAhCpAx/LeGxCLs21D6lVloumj+2DsjBj3aNOJ5j
r0PtTLFPx4Up3MOZ+ExdwsNIK1r7oQeyyYraRQR0gxOP6noie0QJaRPvJNs1Uiiv/ZdlzuvcENSr
ddE87N8E/LNOqabD/NvZGQpr0aNZyZRmLFRrFb5fXsim1HZqkOaRHuwshqXBWCEfv/Xg/vs2jk0o
I0BoDS8FwMjsSz+HVpR6MwZOZlBq6CukzJ4pZoYLn8tbTpx7elLPaFkVdl0AKqBJ7zFBhFsJl+DV
XDMNYFHootM0K9Uh6I3eEEJ9DQzckJr5kminX1llJZdO/IH1BFNP7NztK1xgRF7pazIqGFoQKM2W
MDkdVmuY+FCjwDopC5FRrWANqnDgKrBC/RU0Bxz2CivoEjQCZUHArvZEs7cFlsaMUnM+dqXj6bOa
s2Aiw4/YVyVM1ZqXL25b7cyi+5UsMNyG3FFDrRo1rOcgq1Nfb9b0vcCbdlkiSAECftVxP5PIwilI
9W+PKjvLtBkF2vuIW3Tipr41Ijn6X37vTtnc1STTYxgf5sSmQ5+Xm7qA0zeUmKNyhHLU9TppuwJ7
Tpaxc/YZAWafG3ea+ZyqyNoVXofEXgwkvAD89vSMRkWZ6gWuNnelX3hebA9iePU3nUX/Q4dhnysQ
MWK7JLp1i5noXr4NvE+TcO4ImsqBXdwXlCPmzKE4GPq7JxE16Bnw3/GcwP/ejHQZ55LqANKGCwxz
1ujti3+VC+/MVxNIJuDiI7FJsn9uj7nJTXkFURHxJdtF0s9jFqZ6AGWm9AXdDT/kCJ0Ct59k3PoT
NWiZMLBn7QwVhRc52nfP0VSTpx+urHg5p/vRrQeoH1mclKnix0KNb6HjxbvwuN/kUlNxIGw8J6Cm
TcLMfs2Kw2Mqr2m1lRFiXTklLe82Tr/TtbyfQRc/Z+IoaoqJuTQmzap2Df6IewpXb6IhX8yoKIQt
JxHB9qycSGGq7mqye4gjZDC/5X/zyMO9jCbjEixFw5vkyvMIxnJdkrZNvGr4OLD05sBHTXVPPjYs
Avg4iqUMeKRT4icUkd0846v2aiKGZQgUOlndCnUVAaoEZ79UjuVx81g7BnWpDhcU4wSxKC14erEZ
pwiHBTPr48Ycsi/wMdKyuR6oW32M0AdcnXiJMMKIcebELE9QXr8M4cgy0ZcHdZf28zEUUpJ8511u
26W5PNbc64Nuk9kJ0e7551RfJnt11PlWsWujZLjouppY7vrzbYHsxfuxCX92PjHyUWLS1PLdV3xC
4C9L2DiLI+iCCem2R7vDHs2gButvVQO7oXrjCm6XwZRHr8CVf1kTapPD5Q7pCwMZgYllz1XXgP+n
PjET+jDMUIH3vp2yVqWiZjYksFlyB1PDlDWNUz42jYbZ5wiKfDvxIwFaUFKPXW2rz1e5xfREpfKf
1QWtvqqM/8bepSvI3G/1j09YrdRxir3B1/A60W7xSDotQ5SmdQyrs/tkis4cHLejUc3HoQ1e9HDv
wTMot+Ndqdh4mUIgy0uFaUWvATrCz0yBZrAJyVpt4xMs3Y2R1Nktda2U3A7elNDRBvfqSflmZSa4
EDv0v7rGTe06SSKgdYx7SPN9w8yyOZVXOMVMlKAi5endMwefRgPI2BbMGAgNqONRM+TbwDHb1OM3
4d1+SHeSqhw0u0auMKXGR/5ueY6+PJvp3WLisuO1hAwGbH8RDHML3UvOgnR3/as+6n2fxV2RU4F8
SrPDzTaMVxx9Rnw2elhqsPaHeabAlQGyz94nsuvo20jZ1K/D1TIBbfGrn0Wo9+Z66tWpXclLzggc
H4z3DsDdInAQSoWcpA5AjLibiPxEG56JB17wgWKVWk4Pj3xSgElKdNSHM0/5nFHtSON8l49WPm34
ODdSuW5sJbpxYp1UIM2vopzupIsM6i5K0qreqwtTFsej9MWFXc35pnsguTryNmuTdTPxYP9+crOM
4NwWPvUV6hicBhbPUNoeEG4TvP+RIQK/M3hb/FS2ZfBqlHD4hZqjfTFh6sTapXHHEcEgBkrsMp2h
V/EB10C5WkcOaI8tz2k3VdccGIhKxUk/E1TK87Ak0Lqez2dXvfZ+o/EJt849sWSxa9g9s+pOl2bp
9R+XKOI6cmayoHEuWBSxBt75xsBsZpVg088IJjTDDnSMFXCWEmUZbxOVhNUGVq6TKwnwGwjxsgDl
29uJOvy37FiEOsmYJwTmnaIlHcRfSb+x+G3yTOz2n1KPemOt732KyLlF3vtiOqAgV07I0fAp2aw/
xQ3drTOyIEG/m+pwAO31ErfG2vhHGqeyVwVogc/eJ52/lhUNZiP9LV3VbEXgeEdjFmlAbXJ5eNJO
TyOICW007NF/F+WrJ8HxZ1YaakFzdWuhUVMoKjYDTSwa+XRsdn9l3zmg3SdEQ9KoC+qFZO9jpksz
x60GTMYQhVRz62Vf+E62VPnQUEldGfrMubKDMd2ei8HO4B9LZHyj9ORdq2bgz3m7nRiWn+mQQYtb
76pJaH1B1jH0B2onH5eEG64uE2Xy9ZCCKZ7Vn5BEGp+felip0TNwfc0UCQ/eHROn4W2zukoRwpYA
fWp2fpfCbq0l2+tyKU9PNh/4iSsAlaiy+TXwO24rgabdmKGjt/sopYqyi4NmegjQmOu5mbL0cEKs
302DrXXqwyGjvtrb92izOo775ukIty+Wso0TeRMG2n7v/hv+kfir5GC2RFdADi6o0zh0Z+G8m/Sc
hgz2OqDs6M0HmC04pevJ/Y9veRv2kehn/rk0FbupvnTPLXwoPjbZH1LaHYOh/LhoxjdSZipdWxcX
l6vxyoKsx860EqHs6HflwQlrxQ/gzwIr3Qps4smI/van1iTto7kf2ZmKdSxP9EckEA/F25yRhVsM
bZKiWCergTn3yCAnhSV5EoRmvxeKrxcJZAQV7wS23sD2hRERBrLmCRKelnBaDJfjwQ9tWQGz+RcL
rlXMf2hVsFjcMemVIwCp9S4P3hzWPZ6kAsaNafYDHf6CIKkeHQP6/jrJSU+BbYRXKSiuznGfFzzO
MBBLm4wR0QnHsp3g8rlBWzwTJG+LngWi32n3fgsRnfr9dB1rC1+FJNO0yzYU9uFSpUmmdmpmDCyh
LWFly8kA64yVTWr+Cz/6/7M+DBLTogyrco8PvevipKV+Jrr391m+16h1EToAA9ObjljnVpRQtS++
MWQebpWYB1u0blFHqBURhTb+rM52/Ml356VEwlg8nFVOoTIqr+J0N96XqDL1uktEGnN1nkbRLewh
kHGiAdZhLouOZpTZKdypTB+syGxnBhN00pFFTrNqNy7JQyzOBxa4fGwJBlffeNjTTT/9KtLSi09E
KFbpnOKuPQgoRDL7U2yriAzuHKtrkauUKZuCmN2BrPLd8r1s/5WlMjsZl0AvorKTfTxFARL9VqLp
biOlcoc1uPHBbuSGTOrU/QzpMSgedTWrREOm1sW9aTUVqTVFCQRCqWourBmrM5Wjs6pGuXOaNPI3
417uvrPmF6VSUXNhY/LkoBBzKIwAyeAVjI9N07/FJ0pXY4OwkRShTDSbsHOs9Ie7wxvRn1p9lucX
2XzP1YIoPvYcplcQu6SEL+z+AYFJDnbcrCcbkniz3cdXpZbHEw8AfqaYLHzScHBTDafAYRVFUWev
H/gqJ0e2FvR0L1EdicZwdLOVYoJjh4xTPbfd9adE8ScYBLi8zbyvrd7+VhDhrjzE6HlNiVj9lwvf
aA6oRxTm2r2iRb8Su8vP981FRimmWcXdmkJNnw3FOf9G8ODJD6Cqx782torf04GYugjlnK4A4vnK
WXg1Ii271Nc+pN+rRekbNyt5/8OEuU31XUTyYykA1oYKJuPgHwJW5zSTXmefo4g+XmeeRjZIA3Md
Tmnn6ZQLM+2Qla2YmG4cYO0zfYnY5vErr5zKqjjsVa5VWpCvaUHBzo80tsD87Q0fsQ1Y8HwD2dhY
U2CsTIB15RwW8HpyL2umjGT6Wt5VPrhfhvMV4ULqG3XIV4LG2a8ymAmsW1KxtwiH9afmUCX/HClo
V726qlCDOO6aAq4hWyEWNmx+iuwi+nbGWo6nonnNpn+Db9Y8/N8YIPi7R/C3lcxesppf8RoMqTns
MEiFhM4Y+ruCXIeWQ1eHCcJGHrD8/ndhKvndkvKzCcwTx/+5X9n2p4c9Vo3VPBh7iHzqSB73RhrU
df7rqsupGPiBMNB/4ZtkbWiZiw4l4phlM5vUlLO6i/IwQ6VEPikEuxamJEhW3jATWFCZGR3sgDEf
2JUlsrMeb9cckDl+ARspUxu//JWMDKzebDDs3OjKiMT1cdirAUKb7g/O5Bq2Z/6LD4276W9y/njG
IKnvGOwTGqQInBnR2UdZ4lcGNMI6kYOV81Te9y4reGwHVejX3WhDSeC0AWfpY54mkexBrKiwzIi5
sxaqpaR8Vy+v3HZw+LqNaYaf308wGCZ8Far7f9DkUEJ5gRtnEcjbo3iWItiSqAuULWL9+IE5FqzK
cad+UUpPWQ33OIX6/tWs7gn7Pk82Kkpr8I4/+YJVvjivnICMo8fXDziLdIG7P+MRK1gKtHY7vCr6
LW9JhfqY2DpmJ0A2IKXxwKTkPyWzGtAtlQdLbZfH8N/Zi/Y089MmQqnr6/KtsBPsEIRep6IVFDyj
4BfTH0wzWM1jUUpT7aau5SUtTrADwJ18DxnDPvK8qtPMbyUe9n2VmAGzK+jKM3GgMjeNBvd9yhEu
1KCXFhy8zASiBMD1UJlJK7OjSXD3olWJ9YJczfbJQD4ZCHzDqSO/Ijb30hrGQr4bbmrnFgBm89JP
2PCKGueD2bVqRDbG33skVFD/1ZL37FoYqLD8ADGR2rq4ACv7rI6BmWGhyZGJCGkrUheLOpFYSEWQ
cKoCh/iIn8e4P0JqiP7K0+SklOLzhZdD47FS4dsn32ByyMrDyiZmlUfxknh/78d0UrAQgiWJJ+9H
UQUbAmEjqAEtd3TMbtHPGykew7WlulGLYUH19ZaZuLO9gEjOL3MiCcSeEpL4q76c3Id1SxGfOojP
xk/Of2kF5rXYN1XP5VjBDBTjC+NFBxHU1RxGDz2rAHabHEDBeMX5uS/e3s9qWUbsjRJswv2R0VtT
Uw+jRN7ymXx9koCUIHO9ItcY7AiUr+NqGIn7Ms3ah8wp5VfrONgArhSKigAXFBaYtsSbPcJQPDMB
MFrwCm8twNmjO6LHoPqr6LB82b/DyGXDJT0uG36W3d0DYuvq8SDeCpFX+VOJdcLqUAgH2IiRBSpq
xeq+m5P4nnEpN96d7cMeneNyTZibAQk2Z+eLvwzWTOev7v5LgKd6vx6euxraz6ZiIbbBLif8cAbJ
VyqQxavfZc6dnijkQHoUBqGcmLPdNdGGQyfP7iL+p2jN18DyTxwtwqC8+Dxv+m5pvD8ftIgkF1YT
T0ND6yIHeLkHsYTbWHiRuNAMbJokATCjQOz+M9pGH7d8KoxwRJCCdl19vxf39vncAEfntBkSHuZO
cM76P7utnqnAVJJ2SK7TuY33zOYOzHIt27Y+oY5YE+kh7vE5rSlxWw1WaU7eHm4NmX6mVqDpoBTM
DNFDTLnj3Nbo+KtgZt3iDE3LvWIJ6Hthf2Ts+z3nJfF0vPIkDcGLz55ISP4D7yOoWAC2PmNPQpOX
7Don5h6w4xTcb9rMaDAY7Xdx0OijvEtPD01fVfj0OsvPYtKS0zhwD97R9DvC+9Pbf6SOAcAZwKWU
7rk0kk/nbVNmMcY2l7DTk3ZNso3QwDmlGgdSg4QAZAIhaP4ehO8a/B9g2QyAV8JkJLkh6/Kp7KV7
jO2T3dUtnbY6rIL/FTMpyNfRPyJTwJJ+M3tX7JOgzVEKsAaWYivCVeT6LxRP/n+aO1INM7H0KezE
KxmhHQLej5q2FIAy8M3mBoHqi+NxvN9P6BgAVSkPWIS3gHVWjHKj7NHbXSU4TqL6t0iRsq+VuESe
risHXqYeCEEz0l3ucn75chfDhgUaSyM49wiqs0lcXBdvNR0mCCrYOz50HQq1w0ujqM4L3S+ONeKG
okvEnqKp7dj2BZ1tVCOnDwBBqqs5CUiMVCej7/ar2D666B02sLGN7yc8k6xBkY5nJC+t7dUm6w/a
j2SbqnN1YAJavRmSGIKPbdvjC4pogvSCbM38sHWR3Ty1ayhmJHkEgsY1sozy8ucENoBi33YGEDQ+
ukAYpzdMFPG0wQBuFCq/h5Bfy/xdB2lLkC6h1GIwp0vFZ3SM6JqhAHFYncIvQ8xcJS5uYgnzFzZ2
xQMLjbb27Rt6JTHNyMkDA1NDQL1VrvtDjP2Mmay5nRkFRSJC83OMdQkUwN/Yruwy6VzkzuqoY8GN
RDn9i+SaAZNN0JVdI9zrDm5ZIMv/6HDkEsYzi4QI764r/KSlqufW9TVbVZ1Mp0ypnGZ65lWjxUTM
6/vvRY0SVClq7N7Qgo+NtIm6+b/SSwc0SIiI3dnUu1UJGiTDrNbGKFEFBsMKUjX4UM3C1GeFDBSG
KR11o3o8wp9/eKIvmIPdmOVI3ZYisFTPA8+3DFT+1IND6WdmBl+wGbTONSjWyW4GEJ442eSeyBFD
wqvV6dpbUeDd2zyFJ55lvDccTY9fTAflsWwLb1Lo1CE1MUjdiuP77IGHVqI2/ePW2pVlHJ5p7S75
YZR40vv4R/6dBNl5RLXf6uLg8DCmHL/L7DcYdxysTw/q+EHFW0G4ABjAMGjpBV1j6aiZdtghQjv4
REvtEIWPseigaymmat0isB6F6sbZY9fDxp5n+XX5dqZkPefzo9VxgRbHxL55VU1KGt0cyP4edHC5
fRjPx4y8twPPdCNr7RIGTBeph3toVYFvd3uHSmV2tkQGhS5gFBOKOi3zDYtVuHlFL9nJHzrpUTQ5
NiIY/glwit2uxBa2sqbuz++bcFeinCidNZC0yKVXgnFGQ2JCIKJj1Lo87OEpfUqHs1R/SnHaOpqz
r2JXs86txmdy0to656UKnFGhsrV5AQBaXegjQSPBr1tGQVCLu2ed5Lzr8qvt2FH5sTbuzKufprei
WKep5Z+SEGH9lRHc40J1C9S37YXSU9fbZnyI7N1+RM7+BBan8uulMra3+S5Gm1S9oizkVsFZBA91
P6RgRRrqpO33wxVhkwo1dg5Q6/ngjYWjKyPGYxXTyfW3Oyb5ZowzHSAfVe7SG45qJQ9uBKlYv9CL
EkD6Z+yfPO+fj5+6X7WpQuWeCusPOAFymJR18o2D29IE0VYMNxFvcRUj7LRHVfwN2cwryFVImmuz
8TPLjLYntTM54DaoevapJntJNQAggEKdJP/OY3PKBWkzsOjmw+hdhyiMDFCXCnGqZLZKrxY/Io5K
1ZB81AOGYlO3d1k9RV5rwZGxSo3BwjClI7M8zlUHNlJWQsrL/30suQQD44xBtzqy6l0TC+MMiBvw
R29X7FVwsL7+6E7G8i69fr0dy/P8B+ow6gqfWMxvXmSMir2CscSdvSA+WtqafH90VAdRjdwcOnuZ
JmXICkL17U/18+LZES65FmD00/Skiih8zKxx1/xjQlCCfDqxNu6pgjG0B14eeHQdzdcHgCzJlpLF
8pDGd6ooNzw8b1S7ziRnOzjKGMNaAg/AzVwKnDK8yr9YW73IxofpCBEtGnwtjVUVQDRTxhzykC7/
xyCxMnPTjmYMNAUW9TcK8nBVn/GV8FOqN1GSYRFDkatOp+vuDanMdG4kxYwbHLsCqeW+SnanJgkC
DmMZpvzjD1CAX8wi3fU5gcI0P29/cHwPKzp/xUHBKiwDwDmhIMSmfG9HKfQI0vTW4cDNyr5FfBsj
3A9Gs+7FFJJkPQD7XNS4uV6g8GTWIYRfQOlFg+oAcMzakqKG4+VzJkidIyRwBrTO37RX/MpoYxGr
aCrvn07LEAGM5EI05kokqMp8ewpuCQdSvIvgrJkvTBjYeXgZ5iFwsYqtwzf3QpW5R/36SfVkW5ZR
BS/Lz/ebEXQLHb/oz1rCs9SLAnhXvgdQEP/NCH018lslWYQS5mOvnW/sKaAxiJQd7ad/63Cxssvp
MFsxepBQim3y2DtGl35SfJxlWLDziKRoEBha5Cpt/NaW3cf0eAnj6pBvXqavP53xNtMXrV7UK4EL
eSn3Amcv6QU/aVpd1+CJJ1pDsHTVXY3Pk7quCZGOgOABh4H+gSP/UkKiyP0hoTONs63VaAgBRd1m
yXzGgLH4N4SvGHgiXjq3G0d71BiwPMLEfn8/FBktfYsV2Mm8T305axJM++F/uvR+zkmMhGH2FP5e
7+vtXQKDKklAi75HG2W+BYSK3uAxOmG56Tm33wnE2fGoB3aNVny3MLpPYELX2EkLyQG3zs1Z3QDz
f+4wzTcP/53VD0+xiuymfqnPyUnMkJSegwPvSRcaqZ6rsCKF9tuMnuTdV78yBgXl9XeNFhgJ/Glw
szZtED66xThbzCUAYFM6nrpXmbLf+uVNpkw6CS72EZvLEaZLluJpfhtcLtQH2NRsrEmlTR+B4cXv
2LiwTGfUH5I1MQqHjardg6Q59VqPb3IpYWOJDf+cpjQb4H2/FSmkksdb5p2fQNisOy5VpnM9yHVa
xStKK8E9hg1pBMTSc2mdDL4+CzMCMwFe2Rz5ju52nlWEivRrmnhsOXH411sVjybFoqkmRuTrtb35
pI2PBqp4QqCAVfgOdcIttZ+Iad+3Wp0VQVU7JfW1cPRZ+ycwwO0L724ULoIQ/9Xkjc+wAuMT7CJW
QaXB8Ebqip/5jBKp9HE4Hq7b6L1A/IlIY3DrDgRE7AwBY9PwAW98LwpUZE8KCbn+qs/3CzkPrvLy
BR8ZCw8cDit/VXAZ49socMRQwPm4ddRiB5N3KqErSgkLZVVUv873q0Ua4ZRTC6av0Xb7u1Q1E3r+
r3dJRBWh6o0a4oflyx5Osb6q+j3FyhGqsZSH8kYGFl24nNh5/pz6m1p5ciL8mUMtff7PNqAyUVju
fpgDBeB8180nSBWrf/AUe4ZfQMaHMXZfsuPRBchq8zB4vOBRPg+492fK67FPYE8C8rzXyECEgMP9
pgaGq+OYKuB1DSN841XzPPvDnZhYs24gRl5cr8mMjI6k2YxvVBwTvVb2OPYw+5phHpaU/W7PD4nG
q3PFrP4hcLzUrVKdP+TI8PQyvHib4EXKUJnuebm7Y7s/2yIAdSBPuJUhzLqiBxeeDOBYHgAPKOeV
kTYsKqXrCIp3pt0Om2nOiy0q3L7BEBx2nizohYw1bxabR8GycI5nBi2lnYPeFbBpcNQVagUITvV3
SDR7EBm0xJAduxB6mRS1izhtdGlABgWk4cHKTdgPTrE8gc1h3RybfzJgS70FcAJ/KeUEd1p6E8v/
eP1hXdwhVFJFXL9/XnUzI10iX/lzTJaIlWjmaj3adl3NYBeMcuVyB2+bHZAoF/Nkw6uJFxswxqdD
fOMjpX66QVfj0DQotj6o8cBveyTHJpHWKM6ezBq1vhNl3EE6XQDscutpvX4DtLrSlqfC3HwHDekG
iFQoCfiUTKkzL7K8ue/nhNaXyF+kG8FUukGX3gTFd0dt3uhpq5ivVNYZifI/fXJrTjX63Aof5HEC
mAcFTKfEXQA1YAHqxBDlg6ZKaI5xDX2Asw7PJUvuAgQMEvSHZBElBGuQYBVBSJWNJAlpdsMbprwd
H0Q5ytnYmq7nb1S0Dut2ATPRbPDZY/jdqOzIdF5Y3IpKgkiErb9e/gXgfFTfKRHqVXsaAGj69Oe6
/6GDIenSP9iTKCMcNCDAOaD88pads/Zf6/qftb3/pfXSOHsMZz/7P5KpeuWsZaHk67j1r+S0E3yy
RU2kblPLua4qPjW+iUD2MLOLGb+SOK1avzyVphBT+UGkjdm2d6ngTj3aVOMd77Yd8WfgSH84shpZ
N1ikkxBL7f2sf6zFC3Ex+526ZHfRVty2vol4cbge5Qs0rMD3DUvbOur3Eb5bO/3X/kVrzAhgfEZ/
GTYpCVMS2Q9oZiB50Tx3uy9d2VMC3zq0hTIq+u0zn/VR+kKQOxp3TUCexBGk8RWJH0elpag7LQ5A
DGtgv2L3jHJoDvEMF/AG951lcyBGiyuNaIpGCZRk1Azw+DQyQszRnYXC8/1bDy28cCeRmJIHrh7s
YqedcZ3LnOKfA0zrxn18+pQ/o5U7wN+ch5+avjgPXnf2OgAB4Fk4A8fgptvQwoiTMhrTeTJcD5or
TfsCwH1gsIzQzxxlbfaelc9mm1iwQgMHFD6l0BKORtQC1U3JEiV13LYWplmwSxGrXpsgYtDKA0s+
UaxpB5bxtOe9TLvBN1kki1lfTghYJSj4RP5lUQpOSsmaeox0O/TsIRX1Kj3+7g9IOZKfG3VyXhJq
qLGN/o7gEBA/uzZmr26QmJATevE9xJSPRGs5wR0+eOYAifNBnCY60K5QU6lDhx4bsAOJNUbnQN0S
aFQYxCl/kpXg4vjRZwZQ1+Mpgl05xpbvQ1UTDrNSmen/EKdp5aDeQR0BLqmh6xcgXK/NV5Hce9HF
zUSJE312eQcis/mBYpRttC+NoOmw9L9XvFNc5H06sDfXpe8oqObDWFeTkC+YtBEvzpxXcOS4EL/A
Sh4E0LWHnQ/fZsR/lVkm071IFuVcBfQjY3qa1jpsR7+GZ3M071CbBn+PGud9Yaa5ONckYeUpLPin
BVnAW+SrMx9jjb8NfVKLISweQhmw6yOvOdATH3+9eU+pDG5Lr3+OR3udnEjMpIxhJh68Dt4bGQfb
4HlZX4ZBnleQUWc4fKpjefyXVUTPQd1hB7BfuLvFLP3PnpEU8yjbFpjjWnSNS+F2DtxDyHQE5TUn
4j2MG3Rr8Q3+kQZQIAKaIVmko8GAzMpvH5PPXrxoPNLeZWJ4l0uAE/Y9rojfWXp6QHRa7gGap0Of
yzTPRZstYvHSQh3raqI1ZAV4fMtD88cOpBbZ1qREbQyobBi7E11QqtV47KA9cWxU7Qg3ORyycB3r
cbm+9W5+0V+wOoA8wmAqEZoyNzyB/Bdh0BbkH85IlfN4aMu5M9S4NRyrNqJml/ijafUrTLmzipbR
SHnnBHXRUJ3HdIhwOaIZcFd+WAzKP6RsRC5ZsFPiGuTmRMfMaUydXHDbE+Bdf177yTSE72Uvc4MN
h8653i2ZH1Qc7SjF/wbX2P+EJXV+mEDgMfG0lP4jry0nL81jZ1M/0ebeR6OB59qidkXRuDWgHLKT
2quqKhMHu93Zd0NEVVOuiNNnsY/AqCkOF1/M5uTDdLAsh/rN1/f5XXPsfcbrXgm3iySOm5quUoMB
uneJCTkqEKvhz/iQLzuSR0Tofd8gMm0oY+Oq7QnLFu9L9k5Vf3VCzVY3XWJpR3jPwtamW0E9esHE
tub2bcN7rsdA94GWeCve989gcILvLTMf/NspuWaRssZXdUOaVdgGdU9YeOa+4f0zJoYUNhoePqme
3mYz7UGmiyMyJdIvGjy8/sJ0qHTqPdiSON/hZ9qjWJQxcBWiO3ChRIyiD/OE4XkeGyUHLcjLINXL
iVrCrtZQyWFnizUjzLmo+MxX/gAIEoIRH/OjWDIX3KBK64a+jYWznMX/kW/C7nfj3R2F5nPuu2/q
LQq0WmzWq7XgM6d0MacQrVrgOoQI/IVrty9ojLZTd2CvOpUYS1PDRPTlj48Js+l4krIaxYjDKFTH
SUV5jPJkLKNPhS5Po057ycgDWSFrkuMUPGzrVqiU+NudqCkzLSPPDzPindIS1BnLHZP/RE8PZt5E
QwCv2lAvM/QPBMZiizjTWmKHdy+mY3MmlQXEw6QlxzX62Fj0BiPQRO7Cx+JrZAsT94sx1L2QrTEx
5aD+GXTJD9AUjoaI3rurHFSixP1Gdt/AXjg4UbqYuNOsv8A4+XZJ1SRiwju/DPzvGHiCBuA2Nuhs
dl98kHMzBMdEogbEss+jq2mGHSV+FdLIDgvoabzh63TWLgWE3Z+BxXa7FmmNJVTFt0teLGKnNJ8V
kUbqL0p7KcOzpG69a89TcGeglKzNftyQRzuqdUFdhtF3fmn2Cj4h/mx6bCiTJWTKF0+tEqM6nLUi
htWe3ZmsjaGi0PMJf5GabBanO3Pe5A01HUXKGisnOPSvywXc8QXqAcX8gX+QIGc5KdTmIXda7lgP
/kGTYfmmTVS2pUCyr9dxw6eopaABSb/2ta/ELIndzaBQWUFGkI+m8bJEo8WqtGpVHGfWXAythOPN
DQn8Bs8nKk5az6wQrv/TmmWL7Jq1xBReoTRQXkAA8K3Vzl0w9i+P7hVqfK5Rl4SBo0NEHp3P9LxW
TBaVuUemVGoxy6NzLbjrKrwPkeMHY7BGWuqBmVgw2urcgKfAOJBr9D5iUuCxx4NFg5zre+ppxmCb
2Ou0nDQ9n0FO2wmEjLf9VP9EZ0wzrHqMxh3fcKXcQP2U8UTMJM+BvWfM5V79C7ihOOHXO5mRC9al
X/JSw52M7rKQgtS9KPNWS/v/9grOP4DOvFEcC/g5CmGlX2jDWrVjNj6ai/cHVGYQjOBYD1GemCeO
K4xndZgrQHqOSz151/db1KUEcJLF+sYHwr+R3k7+DTRNf3fhWFnYtZkrwjCTQE7K/WjXva/asePi
oHDBPkxW31W4qbDKRt8jLY+sU4TgGwpcrayJpDTokeHJ1qHpTxUdilSuuOwLrmd8YLuoRRao24gM
ggM9dn3dpADSezc7PhJYaq4/fIi83lvajXdKIlgrQOKUK594ReyYuMnxvzYSHiEiGlZSBvbbmfO6
PtyxXBx1KL9l/WE9bt17xzHVRjjcuwOyPWi2x+sH5EQ4a0U//v+MHF4j4ontsBirvUyPnHfsDY9n
5H8S+fFjebbAnQXG/2IflZqglqj+P3tBAax78rOm1cWTwsDj+gKU3piVOwldUpEGn3U8+3z6/ksw
KFY5sT7R5J8aQolHbpKYOCJDZgZcph/bK3eHKjquG1+CmV+Cseuf4eyAo45yg5hc99KO3fLHTqhZ
g5GSIojwS4YBwheWCXwJU8dOeubq9pK1MupvMbYhIIP7CuSXZsXTKsQFrfQ9adrRlmfh7alJqIG0
adzbAYfOSqX7bAdFwDsQhzDqH9q6ZmYUE7ZnWlesNzU6v9to/W2gr248Fq+83tKSYuGQan7Sv/0O
bwaE8+y8ms3Icnn/8CpXryvwriIvcpTFLlNgM+Bw94I/2eJjxlMHUsg+BKboMI3JNSgda4YZKn/W
v5eXnpSCiF6Ifsw9NQ9Nfr2Uq9114TAsbKlriS+paD+hGzXLCbbnzLflouB0zbboKjlIIFfWRJD7
R6gR04tb0v0g1RfCzvslFYDRAnXbGCxLw+Jenq29IsJrBSimutHet1L3ccZnq2vE3NzFFSxCwfP4
aWIKICkkepDwTanCZUmlvxGU1IfssEy6DFkFSMr/gj6lwwPqmnGNZWRerWUj5SojOlKbxb1dkd32
cdT0uJQ7Epigfmr+nsbrPzXD+89VjvZpDfQew6LBXn0qpFZo+3iHAqXs2u0/OMswEjXAv82hc/Hu
SxZsdE1hIJaQqSpm9QaGZPtqV2tMHUl4gDCjGoQ6IJasna87U2pt/n0uSF51P8IZBQPd3cneM0kH
qMYfqsLuYO9vNDo23/WTujAKns4DBYA6vfZ7BFJFqDhMy8bM4A7GeIRYwtFbLNFPyLpxlsae/j4+
NRSHwjRDI5968xdefodGg/Yzq4I9LaQ+UqfNe5EvB3a8Hsa0VPR0VFb+roROFrFTdL113W1H+3O7
7PHLdqdBxNEZOSQigcm/0jXls9K7MoSFocMsZrdtZz0I7BX36Wai10P0Iq3zbiSrfITCzFCgmSh+
WvD4/0xuAZcHjly1SWvTiyiyPX5F+1RaZmYQ5Z39oLVfEnUJ9PZ82N2VOegHvbjl2ruIr2tSGBnE
zrg3BQifGXe4ypOLPkzNJMjuf/7d9/Om8D4ARWMa0a/zlCMnz6YpHNfSqfA8rVz6MXij9PIH1ree
ty5f7+35Jm430s7DW1G6c91P7hn66BvVHgFSl8f/lqCS+joNOVN60eedNU9R8Eu9fTzlcNxyfRUR
gEsmKjH8ijVhAGVuqGXlKwuT5YZvhVBuXmZrFT4mYBxPzr2I9S4SJkr4LhjQiVGx69jZ0q8DA0Vm
470D7cVJ0Dg9UPhPW0UUdPKHW22ihsazJ3iTZGa3BGg9wyeUisi77ox9xMl43YlK8Zc+UMWnJUEX
QBaIMSQsFuIh98CCs+MJGtsjWQhQ93ngNVd+LiI1ZMsWH11AeQ7rZSwRSKMIl8YvceSmRg1ElQqe
GdaBjB4DhoUzkozL14xIOQhZgCHhaAli67O1e/49XAQzjjETjzX/eG5QvECYSyefuwfLhwlueRKF
2HV0M1J4J3yEhuFqnDTjpTj20uSpaydUJ4pvb16pHI9c5dA6aN6fJwuCbIIvgSd4bH3kLiSCbRfP
V4vZ2sqL+5u5vmidLjHN6XW6hxM1FzqtpqSfKKINgZ/EB96PTmjllWSpJkfMj9XS1cOZYynL+Y8O
ZuwicJYUOs8swDv8N+7HhcdKjCskxKWREQcx5qWTpJ3ONb3JgYUowcuRZ9RY+cNYZu4cbHQW4vAm
52NzCLf0a9v4Vc2AD6wTANLMmnsiBLgn6Pw0hXWT3Hgy6uWFGQqtEeADoBntJ+vML7VQWjy5Z//O
5pOf/Ys05k+rkNICzHrBJqX6SEIErhDpGRldLBNRxFICVtq22vHP4dnEuVU3+F1udmJ7/oYYTbDG
ulBKE1eaGgic4W5TQ0pxcw9OO/GX1zUn34eEuDSHF7nAGDJr7u54amFcy6ucrx1ini3SM5/gRnll
QGyz5sT70+QKpOPIz6KB3SoF5XcYO2sGZQjQW+W/zqiEH9kvzWlN9bP4a+8oIimq/rtf2uvfVeSR
fBIJ9dWaP2mPErBjkQsgvRwctMUiD0A7PPs2lpqPv/VuoniAjN1ZJGkunU4t+vlNTbfR1knOAnvq
dOyL+/Q0rxapYHubWv/Jm/wIEBK5H0LvSFSwcz2EUPHCXIzygB+Mtg+ZqhG528fsCTiTuDu2erHQ
chTCWAKxnYOYJPkJC67AnedV1CL58hrAOsn/2BOx8ycMaLs5MMLuEaTnT+ujTc4hpHXUgVGhvmet
sOSdyi5f2mmoPl5KCzuCI6L8f/6JEPmm+oAMkHjcfi/p6xjowwcUkUglPW+3yPpEOWSV6NfOaCE5
sC/efDThM0lGLWAGpEYbeYkxSfpO7A9ld7VF8yd0Fo5MRBp8GkJkAUhGJX+9hYzA1kJXJfUcW0fr
tMKOVyJUngBFdPyRa4NACM/jfBY392c39BFryGsXSQ6t8s8kkX5pPlWug5R5+FgE9DAfHoXg8Fq7
DvJpmE9AKt/SAStyqY1Za0rRJBE3WKQHEbdykBLvTHms/nCvHRM75lrUYxAm86EZR4O1yFfGg8T/
gQj6Wr/zWCE7Las0K4wavbsSMepBCGNJvX8LYsoviuPFLhDlgnvMtrirKGb5SI4Kp6XGo2FdQvh+
SqAGyzOz2GnAqhhoN7E9FRFsryyZn2LyPfVMrujsspHY2fE4tH9GUo8zD8SbQ7qQ1GUGl2OcTxKz
vlwNC+5NMYxBU3cpbAu5lcjGj7FgdsP4PyUxr6ap22QDDuEmVaFFuZWLHCf7QZ+wlyVZjVYQ24Ai
h96uU3vkrc5cnqYgA5jwftXOcXgwHjjqcazKZMvSCD9Nmgd6rFSmgOnF/+9bdoLtY23SVTGeIlP2
S/KvmsckZsWbx7vpNUHq0c8/3A4REnL8Pkqb/NCmFsxMnwqBrh1pe6K33uzpXae6NGFBW+wrE5W4
ceWu1//C2nNbzy8iEKhZoDYhqqQ30C6UOST6+E/EL91/FvF/PxXccTu0kPEzkNzPW5LCDuWIkPRJ
th0jvkIN2f+/hsje7RLF5wlOPJq1lIRcRb1ElNz5JHJu7pTYsWtWh/dgXD1swKqyWmuW/LrIDvba
izcpiW962VhPflKl8ln+IgIfzuWE1ZenJ3Wp5V6MWrPU1fXqukzm223LtYMP5p314TPwkz4sf8aA
qcdVHoIy8TUT2wtCI+hsnpBclD3wnglp9rL52tW8t3TGCW5Xx+EBiS6WJmQnLVj/XtTWRoVchHqn
77fJebldwdAWIYtVe4pmWJC01K7OaQjLhtbYzZBcF30mZvqI/TwxkXIMzRCY4E1O0fMNa/Yx2aXK
FEOpPWQxjAajmp/Qp8U89OPxUji/D0wJM/SNLG3mF5ky3uhvWTtKpQWuhFP/t0Shu7Ajd/P1P7yN
8h6ibYk5XUhMOBuijiN5u5jhR0TQ5G26X1qRNmo2z6h1VR7Ksb4g4WdpyPLV57cnNawF/IHP8HUK
nIDEbG6bzt5eANWsT+NF4ltKEfADPR58qhI+4a3y5RYC2EwFxo+tMK0XEfYPG66IDK2qN8FlJQJu
MSdd1h4l1PHwYkMAAxtred6rN3J7qlCdC0jWi7Qzr3v8xzoe1omUUL2rEwbZ+iryla1MUXiWeHNn
7j7puw5g3/D3CkXVK1J+ig2neAHkCfcDMY0LRpr9bUeVo5Hp7d9RW6AoNNZ0DebgVel55sfI2at6
MdliwJr+jCFiBLiu89396e2FaXj1PlTAkhS+/+toDgr4regG2LzWVIBdENom9w99bxzHJ8jwTyth
KlWW6mU1ubYYtFsC6HBEN3T0eCMzu28iVHi4IGEZkPo8xTWP2B2Ra+ns52EQ+c3VJerx81aRCVNb
24yKV2HoiSh5jtoVVxVH3BPHkUM9cBz77Q2t57YTOCUdwk2c2JVFLZhsAj1Ue17XqjgNGKTKGTOd
0w2w1vFrU1hksLc9Hnc40NewpiDzyq+TVwa41Nw4fXo1p7Uz4PAiYg5h5sKKQPdV2SYq5feou6lW
qkbhiO4yDVNSZExZYj0NcCkvB/vqNmrKM/0Mcf/tVzINIwEa7Lh+VGWdXffxAm2mzKTDvCQHUbeC
6QlZjP9lFToliTmqrwNPPlWbxD1BSmCAV3UYPATqadavg2Daic5Gg+MX/aw7reF3Qcsuh1jcWhJs
Z9fDyuw+v9ad9vspJA+TiwYPaLZ39QbHOsTWmHH1+AHX+Ss/qNBizSxFKhZb7JoM7aTHCe9YTOGL
25h4HhHTRemuGXuOzv8YYUE/PrHtOL3AOvUrhr+e1WG7IdhqzCV/OpFL5CZN5IerHpCduev/Qwpf
a/XVVZgRU/7Kc0gguuPeEWB2U1wcuJgAgUjiIZEd0gHeMb55YlKLy7F+7gl4WecCl5g3ozUiqv57
vqS77Xzfnrw8KZtuDBQVwKN1qOjhyQy36xW2KpBYp3XOvhVMB7teFd70AceFTzRIk8qHIbz++lbc
villcYqWzZwB0pBdy4sVP96nTTvZciW+dRvXxFShQCzhv4ULtRbxciFBAUtospDhQ4pOufPUQGWY
ytSJGVf+8lWi/Tyi9nGcBvsoP7bR4Gvri/pmnt0+htzfJ/IIuu+93bKxK67QgXHwPJwEg8P0llqg
LS6OpGz6tm3mbRWBDEdgludi6NqhwwD+WbRao826EjKYyFQaJ8aM3f9O9ScOz5SNzqOPUZssF7kT
ouqnCmSvrZhfB1liDmYSB/HpTR2dxIl9r3Cl/lAkdYVeQ+qtyT/NgvbWin3NlAN5JDrTjuop5kDn
9Sf4+eofsUYe2vVZHDYzI29bK161OZ0vYFk5hWPkgFu8Z9mlkDtfgZU0UCViMrlnJPiYDG6X6MpZ
DVZP+RqpQNYLD2nZHuGrsrmv9bFwq+3cupZk7x1sXB5uJ8ZMOpn7JpEfyPSu6uixXn0081uOjroy
Fx/DtS6VnGkR6cqXrg9D/1xhXXnOyvITbEu5fpA0bSQYDjtZ/pQHAZ674X9fY+jBeQ+LILVap9ed
SIm8eec+zgzdI+QtjB2cQZXdlbKihshwbkQwZpbZzAg9X4p03W6AsvrFv3BZIEZbd+t9+SFekmfR
th7pt23O5dtv/UzEkcZtRYKz9p1P1t4UGWis5OpgjOafBneXEyozMKtqn4UQW16HvrTjB4msO1mn
5wF/u+GfOV6IK+XgVYW5A2+bZYjj4ixoAmbyLF6aSWcxL9c1wAEUmPQSb5TZXT0BO3FSOUR9qU1Q
tLSwefayqMShTGBBJ7cZ0bd6DoBNBYAi3+4MdKDDLz/V0le8t2kSbKske/amEpSS/IWU2cmUsclo
q8a+rYydnmc7ZxtG8Y7fPWsQp9r5uJlaSSNeP8rgxcraylGoSj5YHtoauxlmUcsGlyCofaogAEw6
wGmi4nx6v4Lr+ehb5zN5LKnJL++dLYDsRDJeMXaWqbBEhdJTjrLUmWn70PaLSp7V78veiHVL+g1H
SJa1i8AkKIWvnnatXSRXJXPBGPi2lQabNvIrkzJWtkzSgqxsH1XWFM6LiJov8OfE7nQPMDWfFVbu
weAM8LXuMi2qLWjncp91uRkHTcQ84mgqbBK4W/r6b3jt8O6LMaspkYVk/HrHFgrJcshYGlUmUyHd
SdTp6y5FalpOUUiEznRmXo2QSBtCPhd+5bJ5pWlxLqYSrozI/gQ8MVyPiehA6tnjhPbmFHS/AK2Z
wGNGOruPgV6HfFfe3vyNScdlMClbpWaoNs//N6oDnEn5m64LqzUpvU4Zvrr/dnyqqibo14zGU0Z/
okW8nfo7to9ZuRiqn29XTUcc+CU/u++d7nMNnyXhJoA6DCRbzdSunb1I+Q9L/xmi1HrQmCfiZ7Wz
04Bp/tdUH2gDWMAcimCaouiDOqg2MJmr9Ifz+5qGmszn1YUyrq4UWTolluIrFc11Z3qly3yQjhw4
BRos13wT/UUVyDVPcqxcf4yBqEPGXlX96sbyNFTkQTxorQjLROLRvaHf2MUv3YMiZUCz/R9WuqyK
hlTDvu4BaD2HIpV3Gvk7Xun0/FlzEiKqrw5kA5qnC4ukPJbp0h4cS227mexmnDer/uZst1vs6GM1
SSn/cDOcRj68h0ISesr61Kkp22XPL4RhPjs2/TzmZnwUda0d5IfSXcUCXA9ksPQ6kHfRZ+SiccLe
md3s7yr8entTkesZWZ9crBQNtX9SauVOZQD2rO/bgtgxxByH/Dyu+QZPue/wRCjvYLPXKFF779Ms
eHyzLL3cWHW6d+LT0bLAmnz2bCdc9s9iU4hcmQ2y9MDfHaBj1I1N2WZGK7FWMLyx13NC3W4elhOJ
9g6aXPkfv7g3K8gCi74fQP0eZBX7H1mEJKGzwWDepdFZGzY6+VK+jcL/akszRjmFNlRFXaaTz3h5
7beWzNk0mBuC7oODwEYxWI4EHceL9mRtgGvzMoyBgEBM2a4j0kJXKlIBqqQnW9+4Ze+zj0NXD044
56XJJyuBmEeGDaJEAs1kW/7aRMczaL3Ksx4uCGvAIFIqHrtPRjom1F1tWalN7bXkwh0ZBBFyCQxA
9DweoJkOcZh39c7/vs+I3jEizOCfMvsVsOp/hIYCc0tTXwEh0vKldjWFnYLq7ii6PrlMKTCUvzhO
FTJ06yaHiV/9/F7xAsITZshxxIyc4vUIMm8dObwHtw==
`pragma protect end_protected
