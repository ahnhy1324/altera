// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:45 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oWfHMCniE7SPWlqd8QypUUSY3kXl7yuCRkioAouWmpSAGDIVCbu2GqPH9RJCY22H
IaKmbC7EBgHAdjaWynpdA72nhW75EAijWFQW4TJWLnJMwEZRGcKiyVf5wobjkpMD
3dOi8tsvydr9JdSUvRUu0oVcwAgkHrnyjbcTt0eKWPs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11280)
tt5k+ponz4LnxBDp9SwjArl0fJIK/9wVh89Y7yZnaBEuIJh1Q6jJYgEcbYSo2c1g
zAUztvpMwLa5ZLd3dFwOm8yck/cwt8SCCisyO85FyLEacm03cBWH4iJJ37KJz3sl
6THaHaOpDJSpqdNkiJSYHJX51WwsjPntcdZl/2wjKpMgIBsNmFoEPHBJYmv77eSi
nb/Qr49LpNZBSiLddBBnbPPBj3NtSq7Bg8M1ewg0mTTKUrnKySn5NkRY1JQI6XqA
TUS0l9kkCphOoKezO0WDah8SijO7pDFTtcmtznDz3r/DoboLGzgblVaN0roNKjS1
nrgOwkDBdTdT6z9mzbg4jEH8n+yxkKpazA/xTPZHy6+SjuLS8RdlRPL7Eq2uOeM2
5CR6Bdw9h89pw6fdfPQmUcm8HrbTwtQ1CXU1pakjL23HaGVW+GGncXtGcg6+/zu1
yUc+2/wrfIqSJ9/nwsgtS702a8jvt9KGEdOp/h3qK7/UrXfwGK8tR6k/+reO03MM
qz49OW7Mr066rCYMt06v1entKU9t3wJBhEd09qu7w22ZLrjEO8KqNDaVXEYfo3JV
WJQxgttsZmUFFbtSQeVEYYJVIUnwe3zJc6cQJL6c2gVWtpssNERbN9nerorNIeSE
jXu+z0P98gHqjrgldv3oZafe7J3l/bKsV8K5filUrzB2G3wfzCFubJzKh190rXK3
T+5G9ffZnUJXiP8h86VZVur4oYlh6vx8afFavUD6iiKKAU9WM9P59UgD+11TvHO2
Nys6aRX4DhVGmS/Z5z46bIq2U4PylbJW3hVbTG4EgsyL0/plo8vQLxRFmR/WgAv3
QEWj9+tzt5nG89I/kGFm4TVBsDEY+oKSSP/69LrSgwyBWMqW/zQaHW4kfcmb5WGU
ajIhUAcbCgECuE4WWKtCDfUpk3O54qs6GGyXNAxOe5efl8+tb79pfnSDHbfZCVYR
gRNovB7soXS8v8rsXYN/D0XqT++CtuVbDzro3VEUNKfAs0tQVFCivMXichneu+ZT
dcW+tfHvyW27r9jgv/4UmQZQEjwd82q4M2C6aLnYfGhPggPRNKCaDMtOL2J3dVcR
+PawCFYpGUW4Rwh/RFWMYIixNgVXi6zBBrESCP630oa4KknwadX/F/LpR5XBeE2N
biOpgwztGT3DlBkmUPKh/ZkNHsV7eCGJ8vBtreLYSOK/FP2diYTDiGsgmsqDam6c
Zbu3jsfYDdfdbgTP876b32P/+7nb5qevLwRXJZuUy/RzJHqCozqYxaZvoR0oTlg8
lR++qjIvu1rYOAc+qiNM0dD77y7xpTRLueyzKIJx/08PNB1A/SLEYWxQoCYItSHl
aRjyOeoMrqYbxoAjzPzdDUWgAmDylvd3VcZgdJ6NOWevGAtVv+gmbXRGLct47wvT
0sYPQEenq9/FDvAsGLr99W8rKSMkXcjgdYME9rJagEE2IACYhiiwzqWmVLjVLVe9
Ixb2Yrmg/QskMOTIhiw1RBxo+WZjBeDpCEDSmUE3q8zmgLiM7nbH+E8Vd28Mb0/z
B8le0QgtXEMfVCHE0zPyGFvDyuFcUnZ2EQuyd4AeACgaUY8xpq56BPqTIF3seApQ
A7HcOrFD1jkoBUO00Es+ZdSStWdx/oby7f/noi3mvarENGEFn9hob3wTZjMrdYV6
3K4qXkd2MGk6nI8ewCZE4nyDOB1V6x4CshfGXBhwJE1srEAVlTF3hvZ+Kujg1zeC
APjZ0wnFtvSerYpm5RbHlEsewrXCKImufnShj11J8Fm9KatcobqYH5omAtTGzNNL
QIR+ydkrxVXeQVJgdpR5bGHKIayw6wecD/qrFLbeYX5VX/doz+FxtJ9QeMMPcHGH
kvw4VZCAbc8JdZfcmPiGI5x59m7asmhAr01QmtJrfVCiy9UnVb0MtubzUSny2B6f
xtRz6tiHoUsPECS/Eu4sNTwpczXXQ1M7D0Cw9LNmEWyjs5dAZ2D4WVKB4GWu/qZP
KJJxeviXH9P7TlM/6Ue7cDqPwNwn1DvUSd7wNmUdy/gMcIRUp+Ihd2y9eewbZ9QS
Y9nHz2wrs7VBbH1gdkAL1SxDPuZldxoE3zN5f7jPk40Ks013TC5kSTYhLEYKcnUd
fZpUSOI8K5yRs9jzUXo5BOKZ26b5Lbw1ZVWoNvbsMDostzJH82R0j76Cg/Ty811i
7Hsbp4jts6pA/wzNS3fgH4vIlpjLb2Zxey7PzMTNMoepq+TT9spD06mdPFvbLPKZ
fNQkgBtpi3hxEYuEyU6yKb4oIEVDqbZ7GcofGZJT9ZgbGt0ccfEF0o2bq6IqCn97
S7tHklbd9yPJUib+64i8GjYT2havKnN9I2P/INDMskISubB/jR4VzbdMGVA8ew9Z
iI+GLU0yf27g9+FPj4gnLkq4wvRL0v4AuTS5MZoxRIcVfji6fCqD9xGkCyOqlNLq
5eEabcLVa2++xzDScuhd60JXwiLYCo3nd1Lg8ZpagJbw7uUdNLWtOFRc3FPwtFEB
S8oBaQ5wVEzz53o9Nj2Mzv1/fHZb8UZAWva2GrhRyFv1a0nQUfZLIOdnbMoXJuK7
+Xyzoc6h+uqEOndKkShqkuq+IBUJJrgjYC/CI5upMKVfWnNMbW0MtD0HCJNq5JJ2
4Du/tFXfZOMAzqkTzZ0x3tPx/MAURf1oqxg57j9U8HfnmbzPOPIG20s07syTUbIy
USjUdBau52bE1aPts/JHhD27e+3IsDIBIpouvt5B7RDclrwJKkUkRLynzb0+THSF
DcMjTg7ksF3p8+0RAyJ2xNJxITcLz2bu9mxQ8sqQgj73UFULv5Fxk9Sjhg2Ss8if
xpzofLuyMLSvst1zGvR0fz6k0kRsBWijZ4eJsWnzEJRIomKatuUEI2pqkurMCYCr
IA/OTuyzudJzPxJCiZhbEjy6OPyCJ5RnyOmMW7wTSsm/gYnnJAZh3/6cIZpU7heV
r+ssZD8HMqTQ5Yq7HL1oMs5HatP1cOfwL+S9vmI9TY/0munznFw+S4/VmjdS2XXE
A/wigJthc5UdA9D0c5MF/5eBk2DtxdqLOYANiLACTLKk04d7i5eaUivpDfq+WXMz
OV49hLhUa/aCtuO7sNNk2HOTp/0HNjP+MtiHcBEQApJwFz1e9mqcFsCjYbip9Fzs
O/hnN/lVuEkDMYxTUz9J9yISFX8FzyyFpoWVHqcUXEWClRLFRX1zw//ypppnpind
V0mKd1X3Mu6VvwiqmtnRBGXg8jRtNXh46k7FwZ8CWDp8n1Obn40cTnjcSaMvXJHZ
zrCXaZLMHJRW5++5t8Dq/Cg4Nl+PpxXrawNnDOwSKEISzADPi7FMu0KWiMesT/w4
SwG1VbzqXabuhDH/JVVnUsZMVYIv9TBPOCecX85Q87mtihlFq6Uz7TMvc2EZsTI+
USVBFQEBiKhn6UdHqEXx2y03R60IQWYUKJV6JhmiEiXJ9MLDrCG7+6XZyvhMl9Fh
eRUtVCR8Qb2ZLZzQaFm24xq+X4t9vRIZ7UZQgbuMIZKxuBITUEEU03UAtVyGKMMu
xAa5bEyoWos5nnCGeZvx3BvS+VpaRMjohsihM1F6RerRWL0WgxY5/qgrpwP6RHdv
ml79W/pJlUhwi2Vyw/TsLnb3b3O+GhVmG9cS/yQiBqK6xQpqudkIMHe7MusSBrV9
f4Oy79Po+bb01E7Xwmwz/Ypv4zRgeNBezsuIY0pml+uStUhpX6LKV6y25KwW7teE
JGGMBOG8vlYLPym+AzIshTY8X+1VPlQx8WwhW114Fv0M2yI49/lh4zxWQ7Srp51g
UouKILmlYihrAXkUEcWCgdPNrnoqKURvEutV2MuW9VnDqMSvA01dsfytwy6n4E61
nu2CYslv3EH83L+7K4AFGMJtTZiuJgWyTP0/keJa7GTYdF6km5l1lSwRenDGrFTY
bcoxOSEolNsiD7Aj4ExAWNbPbR/LFBlw69dP3bR9wmQ0njJmhxN9k5MsTBn+2cf/
lZOY0kNmX+v7O4eoN4chNCaOHjjNwlD1vQQiLgL1+1Ru/dZDMSvZqStlliK/JaWe
0XSWFODz60tI4O2IbBikOyRuMf269ep2ylzph7wNaF6b7OkgdHdMHASrcZsYNs4H
DJrkKYfnL4GWYYJMrH++gU+6ui23KXvpfU6IEh6e02Wc9g4KJlcg6znV1l7tlI00
KayioadAx9kHktwaOIeYmWlwW/Ekz0tio+0J/m1dtS70rWlvJ+Dtdsk/lGxCBRvW
ddriEU/4QJpBUnu7YfWxcp1B/52InV4G9SjztDZslK9YsXfMmciR0+6J5SZO9r5S
fWD5Nim7Vlx6EyWFOvjjPOi10xxXnSjF2JWcXDINdSgQifNmmqXyzh8cRmKNeqFa
1VxNLtFJy4Q1+ZmweqnjXI2tqcnCQkpiayixzZnP2cn5q3OnoU86Sdv1aPB7h23g
zyE0eOaOmyWo23LyGznEx6vuZIx6RIiJDA2J/MKgSUkFKqjJWOVT0VxBv1TXww7j
9yQWegIC5uxeqtDJsUQ6s/hEWLrhUjTKi/d9RKN+iW+eBt5Dv+DxIGUOMDorqQyt
0Zy4D8kEt3A5SkjiazH1bNBiIt2+6Q0yU0Faj4y1ddGgrUXk21seIozqJYATppku
2nCHJhPM08FN4OpBk5KN1pUooSaembpBRZ8jvTO8PceBXFftG1M4tz47KW3UqlJm
5JZkRLKC1qiWpky69M57qiW/08f6jcqxAUvzqu7z9PXiSfqJnDBx67EoH77J1svG
dg8VYySoxZ11NpNEDB1lGZsfRGz9027IGhwd5iIiSNRYs1KTiOW/hN+nPf91iT6n
ULN/Dp0jddfp31TuwroWaELgFESQf3AVOkb5uTGpsN64cc9GI0fUpkxX6R8eI2UY
zTwgpHP6IeDflIVIusqH7v8zIPhPegjqqbO40k96BBEvExT320vf3gLV5OUWlFaf
jRoicNCj9TEVOqkxe/GyVc9cmV9RV2EFalz4HNbBIhK+uPiKLJKo/cKCTYAgnmc9
yBVAh5LNaABfylnNPBRX+TXurUdpMijVCPHEdvC63WpCCU3LTAgyny/Gif82mGfc
WzWswhqq/NG2/T3+jgfa0n8VKOkJ+Qmx9H3LPv0OfbILfKNnRAlB2OI6Lw2Mf28I
Lj2j+eFLoMuHhvReyDuG+C7j/80qB/EQ2pWm/1my60cbtk9UGmZ1vBniwMD+bYQx
1CK0GirYse5b8fdeVVNL2MAMei/EI9o0nCfSqvPZEy9wHPtJyBMxv2RL4RZ8MkPI
uu5wggHMnlYlmW9Ig0O6M5OfGMaCiEG23Mojpf+ZmsMglB4HbBuMoc2Qn4AUvneu
mpV6ZonoenXhhzr711NGm2EyejKBhCkZ0VaNu+zqv2+n1WePTHiu2ZrO6ss7cqKY
xDnaCJNoceOQT52qKaoqa1IPRbQfqxfjIYp6lSUzNYJ1D8ApaztQ6CMEEz//C9rx
/mCAE/WMon02/RJhVfJxwaxrpQvJPg2E0YE88X37mM4C0xs1KvR4JzVk1Ycz/4qp
DxyNKqAGh4/4DAuoIfev41h2AHIA3jO2jUOKkJXpfWXebsuojXPLXWZZe+FwU1zV
oAeIm+cy9xokrYUZfUBJsGcu2n2YZrmqeXJrBEGS8Wc5b+pR7tlAx+PipL2kr4Cv
GpivHMfYOUtRQMhTZ9YwQ/yLIIwriqJGx5czx3XoQrGNUAm9yKR6S9zPQaY7v2c0
NKlOw0dXUUG76GnE4da3sgTOfLgyDWUDBwEZhHNJXd48o7saYXuUyVXGNs3GQIHG
xn6Qau/mlE59dPdm96TyDLdM9G2JwwkeWmYvHrGZl8rPiMEO63IfkFpNuMC76lw5
eD/Nw0sGEtaqD1uTA2hZVchgzuGalWELGV1JQ6t4GDz1pOIQE3aloRJjJitjGJV2
pA4uS4+1Sby/hIkwz04dlLKwZ6udLxWPpftp6k+iW2dIeKpgAnxfLzdDxtWrOn3S
DNt3vNxLQnDq9jiBvCBhYb+t/guo3xEF/U6taF8c1zJUcBOLp9Vydg+RHvcg12CM
AJjnW9DISVDuM+Gb8cVEFFCW93NXFfzJqkP0P8eyML94RtcWIxdESq+4O4Qv0BmS
KKZ+9ezS/BC/mguj97KvgNQ2o5fRrivu5iP/VZmqVmxqz/MLAxzmTEeskuqI711A
WX6YIwmHkuq19efZIrbkpswXMeTr0q1Yo9nSgx72MG5jZhrX3PiAXrkoIcuok77o
OxAmCzhlz9VsXqUb5422He1+SqVad1PVPi7rlJdwOH+U5/vXdGENRx6zcWoF5nJS
sUpusyLYW8FPsE4eInGKLes/kEuHupzspV7BH2Ff1nSXGnTSNilipAQtZ2e32Ssy
ksD7DKcJEj0t2N5aNzv9R3XH1g2VcebwxaM0f0bX6vNvRDaTubrMkkqtIz0TEPWI
8j0GqaAAu12hO84fN8li6MD2fbd2kwRsv46Sz0bRS5JQ2hT0fISYucbqkjHULUEx
O1LrrRhCgHzz7EMz+zBx3sN9yM0W1YrgkjRlSay0P+QICtcgvodom+kT2bJS2rrn
G4ba+2MBw9PM6Z8rO1wsuDXBO2a1W2IasoKL5412lsS4NICm9RLFPR6xhc4EvQTk
LgOWBhvUB//CiT8WLQGozQsnD60AIfGGo4XASoL6wBZsuYpZSQt/ekHzUbI2X7T5
kz6Fa6TpImABQybvIyCd9jdji7j4XLFCnXoLPaJH/hXyP/tz8/5tExcUZz8m4M5F
oeVcR4kXZre015wibZRy7j2MUH+5Q5BVOMzeWN34Vc87c+k5hostU7x0pEdF8Sbb
5kS2m7FGCD9/v/M+Kr33Oo0pi6SJobfsJ7gNyM9EAu5Us6zA3AXB2sU1xGJu55Z3
rQaYdaZ8MDEGkFqjFmVXlnIxToarBJLOlV23Ot6dh7s62PvegXjtoYhylOP883eC
ewuUke8LpT6gy3oN2wyMA9cTV0cFGVg4I2EvrmJhOYC8d3/tYwo+vj/CWaH8bn+y
Dsg65Rq1jsmq8YOqM/YBc1X5+MylWlW1bTIrmmlP9++l+ywwmjhzNwDzD/6uKe1p
cgWH3pN8Q6+6gmgQr+7kS8p0ayb0IdnKFKOLJq/X4QguxYAqxtxhf+cj8JcgCbZj
yfVwXxwkqYHNPCUEGtrMWYEhQWywPYFuS5Iv6GN2X2i/wdm2d4YmJYXahGIGEVvr
ves0F3jFVUfzVl6SK2iTN0PCDoPL0/0+Niw3hUzuilR7EsqX0+0ZPweEqu342DUO
8L0FmXgnSIIEdO1WBUSOQqIXw6cBZRAwQTfM1prgsUbEl/X2Lgkhip6DcKI1Cck3
mmFQ66CP1Xmdmx3WuUEU6EpiC+dAYxF/sybU43QIVVQVBGkB10T/L8Qy1fgl3SyT
aP7/Rigybr5iIxEh3fk4ioG1ygURtGAsVxCIPXg8i9gGs3MXiGC7glvNVovvqjU+
2iJSuE4/eHf6Y8fTN6Kn6gxY/jt8tNO0Zz5XSBNoPTGO4/irB9NGRnoFsCOpaVCN
KQtzlk5VpnDgEYpVWrit2zaRI4lPaMMNib9eABkMwOiDV33fBpqUuGkyG3RqvJc9
qv9TCEdHvMkygIHb4xuchrDH0JIsetSPAASoaCtsUXVv8jFQ2oZxVCq38pDwihYH
bWuiieOyTac4DQTYUNg1vIwCNmdepnoJNJ1+hJPCZWis2o4iGlKFDXesOTUkOGf/
wWujtZxY8abcZJo9ZHrdToUptgeIdBG14tlYfXDL7OCoBuZ8YCH11c2FCqc4nS5L
dwu3yV12JdDF+JUXob0WHaVHTpGSEwXjHoRr9/G4eHTLcrEA5MtGi970V46LwnoM
H44rTtw7EBZn/++C5UYbqABVTX36FpjqgxMmv7m8MTP4XmkZ689usdtXO1xaT8Bk
fL50qLC09bAUgQxBKXyEcCFew38/o9EtT6vbHZmxyFTb2pOV98znQdy75hGMUNCn
7d3HMOTekTDPZPkz/N3PYcX0LfgvSCL5iVpNVH5zAJIbYpoUyzVi6ZrKR6MwDooH
6kcHlfKNBItiW6tsTxsVRah8CCuL9sQPR1X1e67a+IxDJ9UbwpJraDVRbDgXNCZl
Vg75wzffuNrq3S48B8Iv7y8CTnYx3DEM/zuGw1ZAPlRwUAXQiDn71Ufj91v5XMs/
/0tI5MM8xThmU4gG8rnPzHCp458uydld4TATuJAJqQSaTUGFZj6j/GplrC6HOTCZ
/Z9o60YHMcdA8K00xoyBjMsECGkkstYS4T6wG/Lm/q8G1FhFRohp5dZ31+dyS35K
aOuU7n6/cL0/QcvT5IpD+xc6VVBZIFmS1F45NpbBC3Bep57HkT4R2nPFUdWDda00
yjCuFcqNv54cj0aZa1NqtF+id8npDSFe40KmdMChcKeSRmAKbCLxbuJGF2KHmO1K
oJHy1h7RixpcuUY4a56NnNkr7P/KUGy68f0Rf9xUFQbwHl8w7hMV9Hz6PU9LUvWn
Zqmn5JrWwdST0KOIrDH5s/4sCMUtCUxzbsx2ng8ikFGwAah0CsQbRHipgZvMB13d
K2S18WIg/LNgkPo5sL7CQDhuSicAcpFJvoiUfZGQvpHT0YVEek98hXFmKhpc3QDO
ZVUTjkRKf6LG7BgYSVs4i9tG2Eg1sHkQM22ejGIVGNHsVwz9mzOGn4b2ceTKXvoK
hsVIzKOjPcOiJIg+UxM0NdnQ5dmrC7QTiv2q+TJ2gfap62CRQmL4VmERN764BRrX
pnvtUEg6JwfTEksT4oZ9pgdCTB5OremGpNPPgrvsZcPvq9okGsY9wsZiaI0ox9Ze
4MC6coE5/IyLW8fDN5wqGQtrqKtq5/47FFIqveTdZkxeLArFo+e3h/cW0ImLSNmt
0aYpQZax1Yvh4teJ/xR4xDknGX5/WkqaWa0vi4qlSe9t7UsE6oUzEfia8isj0JZd
cLwslSLwiPpqBkcK+qyU1bfSQ6ynINzP1XARU3VPlhYEBhX1KwwbIenmj0iAONT6
TotDUbljDUkM8Rl59mDsrPD0TjUEcHeP4YNrQNIQI1QYcavSpxkJhJQt4syhu2lV
Trq90XvwwXfAxi7RFtR1anowiYrKlNsCP0hjFZ5mj1aIen91UpHk3IgwT5ZcAqRW
ZYBNGjRZpdEUblOz0oBc4DV9M6PJpT6mRaGKkHzreEFSXmOq+LVDbJYmEv8EL+Tk
SDe7jKscOctizsiot5bkI//YdFT9bCHdmrssaFSxsP8nNBBMCFq9G9dMdJr+9Z74
N3kdHeygPs0In0XF1/AYCzLcalF/z3fJyfEkWvqlER6JlDlqs6wJjuvk70FXJzEJ
bm21CZ/BPLFAgXDCKQRHXcLuTKsxHnF+NntUpMaGh64la7kEhuRTLTkn5QGyCRWP
UYmXENgwMh7QGT3VN5njBg96bW0sCnFrZLGgRPKYkPshzlAg62rMDN+XR3Qio1l7
Iz+ha/TYQiZyvy8QHyyMrn7OzZeo5b/gGBcKb+6LxnyyR5afpFeIZNNIFJpBuC/4
K2hw3zXmX0Qj5ORbRlUCInqMWaPaIDKpzS+iqjkq4mmuyLmG10IZhb4HBnqZYwCo
GkBBShtdAx8zkhJX6OFLY9vfuIfp36NnKM4zQEiG+B6LeE44k9r15hPVAe8j6EJg
bILWVSglP5NC9AcqqkjSZaLA72xeX+W71oiZvh8/xWYP3Xv6FJMZFuuLwkvGWLwb
qMfz4ZU5bR/sTQ4ZsihyPVBsGv9nX8ek3dKAmrIq1j6yQi6ZXy2cpF/MNtzsPwDi
HWAUj+rKxkajJGgjTPaoBka5i54knDg/VNZsVbChzRKvjq9ojWkTgSXDBW2Lx+XN
pembH2aEovgbHEb6woPbJz4LbP6d7GQ4jQ6AvCfMdbk6SnTe9JWmTwoS25qBIDJw
DM+L9eN1IG05dlFIyOpZhWxR1UEeLSAzROt47WDPccznM3u8hpkrGYiZERZvy7YR
fghko0rh2QHCDEuYe61PhWiRIt9y2a+C3YKCrYxbnu9U7FBg4/+VD5cKeNBqN4OY
AFeRVuw0XLx2iKoRiShqBf0mxno1/N41C8eDAX0rSeJ3dK91Bv2VYJHDVj68/ToR
s2LqE1/M5eu+54RS0xd5w4WAQf8PgY1O/0HMzxT1EZpjd64HQVB/56v50l0Exm9M
sp/5yoq8YuJPLzkdS2v/UousmfG5gDwUZegOVntM4MjoS1KfnyaILktzlmkMF39k
jip6QbjIRVy8UQraHyul6FBqGbZFb9n8MK0Msw9wKP2ykQLZhprtw922xCivWcsT
F8y7haUtHHT13kVPFyXXs9ODt/vdxn4QLis6LWje7iC5/Dorq60iMsQM7Vpr/MIv
Qa2eTcAYdPSV4XEsw7WNmRpgAUYHdZDCZMnzxbDCTXk8iBQZJBTc4eVS/moaZwmQ
KQWUJnEEvrTEUyTrukN5XG9hXrfcoBrHgNdnCvtBDmmVVyovx9k4JyfMbXTAOQp5
fbSAj4CUtLQCQA1l3m1Z61t3XtMoQhtGuD0txFo2QlvGJOTraWoTYA51xOygwCzD
gblkk263zbzcUcF7H7BlFXS9sN6v3E6TySW3TmqjMjTaHUI9Z00+EsZ8LNdDr8rZ
cQ+xrOKN4bk4vCZ/pVLwADPmPCYjwYqpNdVQ6o6iN8YbFpbOWpGdNTYGx4ktzxL4
GQNzAO1ssdvMMbURia/fdKkzB2J3NJYAJXCER+rI4QHYXP4QPMeUoeo3spSZJtRk
zc4trfXxfWveLlqdVvMor82dTB01iX/9C02FAmRMG0RXTxIu0iZelilDPeKaPb3G
v7jqU8oaVOEOogDqpSL6/2qpCeM0YOHdDXdWPBa6AVkS6sU4KPtwNYfu6KZc0JEG
edTRNY5jqr9O6a6bMCnS6KyX2yRou0lqCzXNr65D9Et+bHZyM3xrsTZ6KTbKs2QP
LhdlIexX0kWeTl3QAL00AQu5eNPxrxCZDs9qEQLMiwn6i+mV62N4fBa9bbYGp74T
mJpFYzWtdHfxUaSC/+6hQ/aDNvA52NQKadwtTWZcfnIA5zR4K94tE3P36HqhtrUs
wqpRm1isXVdHKR0YAxbA5Gk3UJ2OqQWamRII8W1C/cXsj+fIlHVarX4rCKeL2ZWV
eSzLCeQ6Mxc+Y6tzvWWnXhlonVaSV8U1Zz5sptlxs98akvpigZVvYAlkvX3oBsW4
dHqZ2Wg96nHJ7YAxZxzt8sfbdH9IVLkLafnfuUJ6GRZ+7chyO4ai/Wmfn2RZufFG
hTeBB55r57brrmcUFTPlukGZXuwBtH94bvp/xrEa3J00QfjR9H4nZPYwNG/8iI31
wHU/9ZjTjOux5Z8yhvp62mrbaxjryYUb9D0JOkZywPuE+GbFr4aWFuT9iAiJ3bd1
elKFX8RhvL4OJZuzEOwRsFabMrleBP0hWx4F4olpqzLOJCNeL9uBzPg5lJS46QiI
afNHVytOiNqlWzxYgyuWsJuRNZM63bnOFjBn9njkSDOZujrgmQSmxoKB/MTUn/0D
LqF570+569WcIb6Vh9fuTcI4Yi5DyJVHjMCYc71AsidpCV7mMRlyrpSRRCoFsM+X
IfzAMfTDdEPghesu47tfbWPjHAF2nESvHXvO0cfSQxNIGmKj7zz+yADm8RMG/Y2S
efQNO4ZrIPlJWnJiyNxHkib3J3rB3LPCdeHHdHywDuip5GKaNjDnxYuGQPgRi9Gi
eZOTyZWTsvmYOleqoKkf/DeAVmeNvrJhWdLWCrGUaKtgaQdvvNqzuF1RvTHShUhu
rZnvfPTyNNMjcy42Lt12OJCXeQeCtEj4SJhVIvGVVG5GoD/qkjsIFeJJpUX9+1Fg
kDFqR0WTDMhawnBzF5j8/kf6+7XcxIiMy47mPIVVZ5PnLap0FcV2dvOgeTFoLw3F
PnoLcp6sw3SASv2xeikr/foMP1Xln294mogjwl+tE/uCuyk0UQBBylR5MH85+XJr
out0f0VMYyxnH0nnqxgARXSZZh7o8/c713lVpmDnZJwDeo0NQlB4mY2ztgnfkris
yJB+cZC56VFmv8eDUe+178BWiwYun1hrxsvlRWKxHArjhQBI14BdNXDvS2aGdC1h
bsb14uvfLGAIGD2lOtBTYAaCyL1Gmc2ZGW6jCVxxO61JKRIeWucoU+Qb9M9gF07E
jKe5xZe4qtpZhMGgP0jCKU8RLDlAnQiNjQybuad8sXSp959tH1zufut9iVTlwrcF
UW1HHng8jHjVVnO4erlORB3W3NOZvRIyaEqVkkGrrRzCPnyrlCD9S3b0zmsbia9B
sQ06SQwNTFwCYU9DIfw0M9MFC5Lw2x4CT4kOZmQd4XIfdMb03DS+Hp+tEQcDSVB2
9QPUWOLJ5WzcWu5jMnxUfRDlOADHmKMkapZ0J7g5Foy0/n7bJl9PprPZIJ+ZKM60
DnHodqRHF1g30v7WtHlMQZldV1t7SEq7Xb7BjXIjjLinb7ZVTMxUXiD7YkbSkyD7
4hDOqFPcVXOAf1shp+2/YcUQjq6tvPJlO+dQsHFGTA/R+rKajLu0VBZME/D8Q218
BsMVdW/5H9MNpJYYMMDxYMqrSHVSDdhMU5WUw/CSpjpKAn+nXXTrbNoN3hWwzc+d
brrPdbSJbArtDTw0RpAs0mMRgHwlP65Vttc66aTUWur1wDAdn+9fbgxWRUtMK/fE
XWey2SHH8ok+VIG8f31ZUZ7FaGZ1qt+ZL0cJzr0WPmuCbSzov1Nj9/Qu49oL0NAD
+PCzPibqqypRUhCC8wuzqYzv60DjrYO4LZ+6Sym5EK8fZC6x5OrF0LudZIAykQwV
c5w8v4e6W4E/kUDPhwLgh4sMyEg2ZxF4LiG+0ztiNittfWa0dnLgDuzjv61k09zh
UZp57AiwvFpVB9wpPReeaJGY8m1jFdnPSytMYfzPb3A/fq8kqsRNHsDw2093VECB
Dg/TIOgSOT9XAJ0YhpJ+e0Umudo/FrZvfFXZnBm6FItmi1CO95gbd+Nmcc6Ze/Q/
tzcG+Dahjhb1PupADXqmVejidfUvw8okQ1PT2tuLjSBFvMimEAnMwNJXj7mIJd/1
gv6vvEzhHO/O+Wm9v68n0kjYCHA5XGZLKHfj83F9S/PpeyhKVO914seRc3xGlEyL
vlKIwZAm+SKqF+vLWETJ1c6jGGw8hGWGfXN41KZCcQhuwf2yU/5g8vfhOLOUdI3b
08bwKXqfFViR6yLmMYr8suHu+FZBanIwW//Nn5APmf8izH48pxWZ/nSi+7F+fZqd
XUEIg1oy/pPRVTGbcqZ/CHvA1yc70dxYaVzUFQmzq/QAvtdNI6MfecKiKqDiOir7
im3baxPLt479Zb6BVouAQym2i7pLvp3ED3ckCNK2vmi/PUtTPYhrS/KaJoXVvJsc
NnJ7GMVlvf1ZHR0xITxYd7m7MCo9QwC8jBdbvTbhzbPkv7uTcLb/QSREecR2w2j4
bVd7c/Tx2CzrwAmxfK9Kza9WVZzrr3h6smZ4K0Rc05P6IKLFZi7wO8Dmqar6c72D
dGgtmW9QD5LsTt/cW0Q+4m4YvRdlkBkpyxc5GdWrvreyX7GikzHh2qP/gYnjuYAQ
CfQd4KkqxQWsx1nEDtkL6y05NVMrfwmAa8Fu+vd2KWDbwAla3VQNqhNKKPGNP/Gh
bcE0O2Ww+bTWQtnkP2P3j8IRL6fjVcnhtqsJk7CpzYV/kDlPb+4DVATF68KeT8xx
AjMmJ6zvjzG5c5gtDbbifF+Rt3hzso40Wj6W4dEFZ0KkIs4tzVAHZfnbAzSmESxk
+0TX5GYk+J8FdsCCqzu27h5KaSaVmTVwrPUuXtv5Ru08T0qXkHIKL833tF09u7ey
P0Ye6IJhI5L3JPzFOWKmZ1F6LPNZYRvd0UBL5Fs+ACJJ4y1OaK5eKve+cU13B6O9
cditLFye0Qxyx4of1mpKo2Cz9MP5yaTUC6RQ+XTlIRBiE94uFKlyKBsEGgCmczQD
ffDgtGvU+ZvjDtMjjaaK9ArnXxSuODeLK0yLlEwhRfu1qIy9X/6bWzQI7UTyJiR7
0cyCH8RCFNwecrW3+UBYtA7Vys2+Lh+s2okh+2/7SkjurLbwEEZG5hBfOuxtr2KD
WFNo3JejR3EM+OFXQSKH/bpfOUMLK1DYatHl2lIfwYUkSWrhT/YZrWe6LFuXevAN
F8FaIG6DVUcXO5EJgdvjpnUEdnioexy8QR8ljgtHhFe3GAc60pbZeuMtUmciE2Jr
oHfF4AfOO8xDfS+g0ev8Jg4xgOi7HPrFfOoqAP5J3Zi9M08SroLjfWQ1G+60c7ym
Li+9ESJv+b+/K0w4VjLLymiKldqT1aXzB2P1vQgBrKSOyBCPAw3p2bWtWW70FQiK
YOpeZ/zy92UYP4d3Jajf8a0tmdxrIDDJp0/8pxmHIGA8YTKw1f1ivHDydD32heg9
rv3VYuF2SQg4gdyc6t1kmm5wXJ4bhKhehrbzEGh8xl/J9RGxsRobudfURoLj+u7b
z9E01xv60xMuv0O3HuRMvThslNzh1xh9mllKml8/4BIXc7hLI6u7+nkRI+dAubZH
yvd4S72JFL46laxZqgK3NccrHh738xGfJC26saOTT/Vmq/hd0BwXMls0eXo5V1wp
NOcZBvaL/C58/5W6lIDigdO+5dz5032Z6uRLCMuFxH05iOBHwPELyUiiBExDD1dg
mi/uzUg/T+X9P9yP0ICjsw9dxBwa65ezpRTYgrEntGI8ZKFUNc5HMRBtCEOZacJP
fG2CR9fompMC9SrtAe9kSIzlhWl9YeVmVl1bIXfo6dNw/K6DIoH0L855j/UpXG6Q
RF+nQiALabRAtqPsxRhuG9nmYl6tr6sjO8tquY1p6PM8satOWhsMHWEPLj6NUjH7
1e4mFJzaOPuM0I8XZeUSF7JD5XRPRxsaTvvXjbn768+8sxi2B51w3qMQiMakn1kX
smCXs6/CKPyosDjQc8brvFj8i0GWyO2G0sa5nyBmWo956gq9HOrsmZnRh6AHoGKH
F70TRzRmCA4wEsj6WJdXdTOFaemtx6LfB8psqwBwdTk+mA+39pnhZgJ7bvogdBeX
iOQY5qLnvYx9wMXlnI3sxNO1eiNOarQrpASoZDOG3xAvn1qsgp+UmG114ZEoB6GF
`pragma protect end_protected
