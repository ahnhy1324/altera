library verilog;
use verilog.vl_types.all;
entity mulmul_vlg_vec_tst is
end mulmul_vlg_vec_tst;
