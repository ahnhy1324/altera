// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oVZzt8XAApXah0Y7hK5IB+GOsp+xi1OIoJYHdCE6UkZbx6UqWStJ+nOyC5nYKbWv
D2vdbXwo1R2j/KKzJlsUiTnXJeDMAd+XC9CAqL9a+zeb4PnzcYei8bt1DCxjuRMA
HRmolPRI6w7sqApfLiKlfHZRB6SFpVFs4Th2Zu5bjNU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28320)
jPpGvGd/1WDfISlivqvXbf+SXhbAJnmpf/M3ZdJp/wq1QnkVx/33eOmNEkOa2+Y/
H0aSbAObVd72rVpCEQvY0MmNgg19yhmet1u5yUZkBkbRknYsoy/2FFFOkKdAMuYI
mIlRGWSHX+ZPzae1Us+rO7rXbSU1Os/qa+lZnDgXQ7PYiROHTfbX+yHrzQebMS5F
LAzYshf95dB2SY5mMTneWcHm82iuro2n+8DN5qcg3AgExBmvekSxBlU4ut7nvAgo
R4Gw1jnfA4CEpwhw6S5CWEbQPo/QZjBbrQDFKREiXyF3QJTk60Vef6d7M8x7/A2M
A+yWsVkcZQyWeYszSt4LWx7lUXPtaEacHK4NEsEFBtIuddxcTPzMACb1lrax/Esp
ot4mju63i0AfXaKcigY47KvOZdUg/YlbzHvxXb76CdmJ1XRMzD9bGcHTzNjrtVi3
i2McSrIsCa4oAor7H013qyKRwUcikVAOl0SGHlYZ/AjsnE75b/IlLYEHzhKxOPTy
9TdM+P2NDwHuoiv99UK/J9hqyrUDW2LbRirZ7X10ZQl03Q0isqCmxWKIJFD2DrUb
zjiBuztXYiYmr1dk2YwHuOrvKaBHDz3WGVFwj8NTQgwD9rf91zkKTkMuombPuVSg
rlV9RujuUc8XfHvA3pOMgP7OlDqpvzUFa1OwHk5BvZ2Gi4vlw+RV6FWnkBCq7f2d
hk1mbcCdREKoOMQBsARx0SwqIBYkHTdjc3rl6AcVYESTmqRJkVLnlUj+/47YnWAS
lJJX6dOLarZt+0sCzF2toumzomnj3bg+NQWkFqT50FpJr15wE1SAuN6/R+3HSiDI
0WU2la+0pxWMZmZ8iaQYut5CNH1Ak/DVt9cB/lNbkHIs1iE1Z23dAcx/eWprRA9L
LYyBrrFlapkh2qY2EXLGo96dER4TFVi7aNhcYlqLm5ne9yKPZh9/voKI/n6tOnvf
A+bg4ynNOwBAupAqQsJeEFsv8Djz1OANBlihz+kyupPadT4FoCMWFlltIUVLlNIf
vmi5MetrOJwh3syU6cnmMo4JTKAuwy3KjhRiFyYJ7eSpYXRGHO/3uHrXdohDducK
8/BY4riGNvz9K6zj+arXlmAjy6YH2xWnNCzUNAccjabE1aQrsMNBNEkmTNiDgsQx
XY67KOMoDpv0UWZsNsF7tbSqNIdItND4PTPnzv3BXftSrOC8MHpRyI3+NGPBW85V
zgkG/Gf4rBEC1fBd34JnlVIk25/2RwtGKeKrM+kIkYvsOfLdtdmmqo1+WlWThT/J
9dejpX0aJcMe1XKj4JuJwNKxbQE+c6fSmedMPPwl19dfu8w1aTzoswqich1WwL7c
BdftMdRP70PinPs3L7HRukM6JngwvuGkVmpfwoo/v83VpCZB5nO7XSOjZZg4eAYT
wz932iXBSNlQMbUjGNTe0kpbGWL0J/oHH0NfV9SrEW21fG+TTwTRJHIx0AN16aMI
sklte7l4/daHagRzSmjbRbVCyEYpv4rWfMNLQkm3WYJ0+/ZMEiZ1J/gWkloLYW1X
rXSoP9ZIAzjqHxQh6FDVnlEMA5FJWT3su1RlO3p7BsISMf3T1/MQzhWKKWV6WFcr
0EonaBmTBO8uTGiLXwEcPI0m6P3wnVRHPMWgVv1t48LqcYfxSzZkOVsFQXPbCGVn
TneTAwB/Or8UGVxdBPYNzXWS6sM/nV9aVNfQdZzk/maqu/t4on/CXA+ampD9jXXk
EjPImfRM/hruk7x5M+q3hy9+jIFvzo2uRDGCNoNVVTmooilZv4K/VrDfaKq1vhyO
fqPPYQu6GApeO0pweGTVD6tWy3co+iJJiE0AhKy0zJIrl0kLL6Bep2qgSWTMxRbl
uQwqmMRDNEnedEtIffJh50jJz8bkUJByS+Kqwd69U4ev+/qRoIcYhLqL++odhfxp
AnTNwhAJ9lOE5hqaa7JtpM83dpW0lrGLIkOeNQr6ljOjySLS1cXGNaIqNq624Y5f
lowJhhNYa/w4geEtwvahi8JsI1k6x7wgGqOdwSagZYHMyZxEbOxug5YkdJvEWe5F
YWRKM0ehHIKW+oD/kR6qez/4/z1Cr9FPa2ipvOZzwLbBrqXcw7Z6L0/Fq04srO43
m+fphYdvW3Uy+wWCHXpLM2j6TT92J1zzn/m+fpFcpR3bMbJJqGXjeQ9LDoOTxzAo
rMuCfeR7KCAbE6mws7idYpZnUANUnbqzmwlVpj+ts2t5B0DKs1qGG6P1xjhzUNkV
ljN95TaiQIL1xjl2qbVrgMFO9N3YUzqowiJheZC5iPSIjsTH7ji8Qk5BxKJTM4WS
p1chq3T3PO02qNf/5Et8LwAMrJnI0qNGqcy0idawJlOltMHrzfozNSzoMXRW4PNx
Nx1iMSg9QUzqWPqvRekO58ywAb4GIw9jJbX6WvpLumclu+4aEQ7yfW06VsvicP1w
GrKqufSbqiRff8NRjcsNU/Th/Thvc+gRJhWKDlaeRZFxF1BhLnlJG4TEcebg3KWl
khhuP9AgAnZdqPWKo+bkrpsIpSRukBYZNdXetfdJ1z/gnweftln2s0IZt+BSz54o
2DwV1tMzZZdnJubu7b/jvvVeeFDik55aaKoiNputfao8r56rdscXWv0CBLeFMfRt
DK/VLS5xDwbKNg7qL3I1n3FJ4yplwjQj1d/5D09bMpQaxgx+6ynE+VTWeK8IW3bM
wYCPK/LKWLvFkGqCjJWK3HFZ/Uzp011JEoztZHzQX0TiowJ1ciBRXJsd/rPi50/w
RXeZBWtOHsW2VkOAAUrn4WFcqtt9zFriuIb8IblJnziCbIdr+r/NKYCweW23fzj2
ggg02gsPUYeRjUjH/ATJDch4q8griYjwQZiaVEAHO5NKyLWTTU9GCt+RfKi63Oie
SU3LbweqdrI09NxkGB5lMUzuP0qZ6sQIrmEpnW3/q60uBn2uriDV+o6p/70nR4el
bHwDOaADIMtjB4hJYo90k2aIjVmG598Rn9LHtM05noRy8PahJGmTZnSvvSGc3uFm
uDrJAuto73YGsPRq6f1VShT04roTSAQWORtbb2NJlU5go9L9SKvPDwFIBPMnY5fr
biLhjy6N4zXFAk8V6GYIHxGhhI2ntuxWYYCieIM/oMxW4X8i+awFeXKNk/RyWoYt
SLi9+8FuXrUq/YUqZ1gVSnhxxGqCZJIaO7T49vCnKOSTH/6WIZqk/icURZmBODWQ
PiY04GgEIxDpct2J6wgoLk/6fFiHt9Tcfcn+k+n4BzpF90bzyBuziU/2X6fW/nAP
k3kVIydQsDCeOApXCQ51WVihElyaqpQwNlXo1V9k36I2VVEyOpRUUSGcSUVklxSs
TULiop9/IdPG+65SHSQTuGPy+QyAGroqrI2wgxQEuZcLHRH4wGADUxOavxiBG6td
W+7f7NLdVIZbsCtmG3DnkHgS79M1T5Z7K/zDKrHL4BMB5pAuckFOr8wBdKrPNzcE
VL5pK0TSbmgqtq8Q2wD/83ehxDOd3ZdwL++Oh9yleCvjL0OnGKu0S2kpJALwj005
bJHI0/linEOiZCizwi8CEHFv8+eImZz6x6jCoQ1zWVLFrU/OTf060r2POHqnNOiM
mNhUkkbjySEh0yGr/pXEz9slFqIJBL7qKetu1m4D/UpGMz5upnh9qh44T1wKF0Jj
87LKd/ynsNE5tDdY42v7rmMA7fhQ6o5UOJFwtLZJLB+hp3b562lJrcOkZ/vyHlXe
urJa7vHCeOBSf1csAN11r9tdYJnDmoIXltJVjFGuBoyNhxz9ypkkia48gK+FDmdB
ykl7bRdp5qGmy2Gw6qBinNCGkZNhVXqIgQSDbhESESFBvl8aS1NPsfCQ1HIYlQW6
K+pqEcuNxZBPWxrzvLRtD9oTaTzTShUkbVEJvs5MnC6bPumOL7+CUHofDXvLOuFl
lL7OYYgNaUw7rbGi7Ru7LObZubWPej/mRxjNYNe8aHUwl62UCUsxPKG+kuzlc003
Zp28zNikDJbZ8juIHJ4TpioUg/5OMPRPxEgPk1BKGulvhHf+QbhOsKZvV7R3fypl
d8ViBDfShDd7s8hIfxHxBhYvCfOtWhq8Qw0MFcc4mPK1qRcHr2YFD3/rk0BBieUv
M0HUgWdPjlQqmh0ohFrS0+2tO/SvllipLvZbBosnRNEG7N7NyFuGIPXrvXJpRM6C
0J9ZjARigcz3SfQgqE68cYm8XHGx6XPzqknWVlvQMZT5dc7tIsdcXCkEizcJtQD8
1G9Ey1xp/8Zsw4kjdCo3tmHPA5NbUSCHpgktCbUvNXysELvYfDwROHOFCYqLb971
iSW3p3JzfH3c3NIyrUafuLl3zQT0ui3hWQC5jUnJVbibpLyZ+7G7lfYH7YNrtdox
nakn3qIMxecqkUSpE4ACRMsSxo7MwtqE4LpNYhx3FNi4VNs76EznQldaMyC427Lz
q2DQV611kuY4ARxoMAx6kHegh92TJEDGpozIydour8DV2jiilg+bWpYsNyKYaC02
Ex4CXGQ5NwiVgj+T0BgNRS8Vuh/HTHT8j6RCvsXTkSNsNcSDrwz5/UzBhR7jDVRM
0kdtkSfPa3UweV8mfbXqJBLhYB62UtXo0X++n3BtPxavuNj3b7JSkwheWo3WHels
I2c9VwkSGvsw9pBR5MM0SJBDTUoijo0fVI5GhQ7HKiRqa1AvtBgLbn99N1bHBj72
n4cNaWo/+Tkk4B6Mzx4H5QTBFQIjnhBT05PN8AaEyaQFOKriNfiacJZHYA64yyEA
MFFKlIjxEZ7tjR0o6RNUyjGIW+i5mwxFsuqvurBUsQdJv1k4A+OKQ7tBQK0jVVgy
9pBHCb91Kr45GwAp7Tqrm2C9oKI9N0TqDrPtpIk3upVIQMi8mkgu0gL94M0HOCjH
eDmcFEdgi+y+0W8GspJ1sam9kKuF5JgOOwWTLjSQ47Qsq1+gfng4OA/aAIbJqb9X
3TEl1+Xbec2SEOeCrt1q16Ui+aznXx1oOMdGD2ezQFW64IoPAdAk1f3Q/HZHjGDi
VjQlAJpQAkMcF1aAdSDykXqjEAXrYOoq1GwYeIU//QYR0jwhtjdI4SqopSP4bdJm
/oSFdoUzisgkLaiKOWFV7xdAcTTPFkUCubPL1mODIEAsRgIMRJiwb1KYOxGjQL0p
qVlwyxnlKxjNnlAZwxa06iTkKDMGs21hhl6jVXUfuY4CdsEuBhIZvNHmaC0Dr3g3
9FlSx/VKVD4n0e/DhghKNXBvP7HOXFyGLqLeNtZupgOdQACicmSU/fdZE0Nw2Kk8
ePcFTkpL0Y9bB+0/hel48eZpnwqZrs3zdHUiT+OIoCxnHCAo0oXtnT8FxHrDUPx/
l6WLiDlVm905SnPHH3vdQwdT2g4lpzOvbp+Gxu81gG+a4FpaljW5K2Ib3Px2Hlaz
fVczfuZSlntP2dgEK/KjXvTGtwXCtlNDR00fyRPtl0bMq/iihrMJde6HL+YNxx20
o2eNfrgSzui2rNu4b6ywZbnjCXfr+xJM1JdV2kX2ty70F4xxnJHbLKoHyLUMlrTM
lanDqE+ZrMyFxF/mq6eZO7gc92DImz5fSVXZGM9HpAcDWfbsNzAbolAp1Om0yutQ
n/4You6h3q78g6tCzUPbHhKttMfeEowiFmcgUfwScTlTqRHwAEe/QBcuTWOdy7cE
aUSy3XXqgnJFqfA5Jex0l/Vmcedu72jdrbrfEy1uZA+OQ7alf/7dVNkryTFTmST+
6N97rRIqoWGzb5od22HemItnemSGN+Pvp7IffNoF6osvZ9Dtv0gV/DLxbOqiYRNj
mDtQi5M4BmHPW4Nxtj0JPq8XnBE/6mAi9pE0tQBbqBJhcQ+EhkPtC57cSPe742K/
snybpxDle0UZwUAJfVt7YV3mmRMvyMqnVVgTmO4L72a80PeQW0hKycc6fvrRxbJ6
qWdw6ahMVwTxd/YgLaY3GQ1cZQ/Ny/dO4U4FU0MheQszDpUoo5cjh6lXXoRULJMs
bmuSGrWgGhCNhOTIYCYWlCGE5QT96LZ6BKDrpT35brYzMWs4h7gnnbD1sXONdASL
HCaN0Spbg7/1J6SiPeZBHZAKeSclE/rQTH6foIHy01jCMTCvw4+xFkpMd7U832XB
QDMINvyxteeKDuThW1tJFoYrRceQDPwrDpGcZo2aUewiOI/bWLOaQ7j4n9zGWhfE
GCmYxDYU5d78nr6irBU7ZqG9zKy6+fhWrKXFSVFUkoKhEkgorulxcH6eatFL3w1A
tGHCBrptlyaLeJEen/zgsvzVDot/Du2fCAmBmCF3kZXFbIct8h3tBEcu/eNhYVOz
HWnHevEEjahreymSOCdCQIJoLATA51XQpN7KCrbiQDMJkGHq8mnzrY3o21Ttev3M
VHjXn62fa09Y12BAMvJm7ltf3eqpVWRQOQQwcUaDXTYomTUuJmWmU22+gzzeJAf5
MG9WmjIekaXejIvqMyWlEr80coUquzLFFpAMVLYV7yPkSwSklESRJ1NCrbG8lkEc
4RJeox8hN0HRr+w6UHnFm93maNTnSbSwfCv/DLCnR8SvkxGdcqME32JavXjvkjYo
LHvqHewfdUjExFOb6Z0dOcEONxgCCFFKpoxqSwiEbiybwdTXzGAZOEh8MRcvzaXK
J+pwlyTnzPy5ojEBSPCjW5OIIDfaSvCyvGyRIqGRWAbWXAZgQaJruuITPCh17tTP
lNoeKZkTfHuQHGLqPiGkvaPN3nlevqZQWmy5rJL6EpmhcYEWM1MiWBTjbTKP6OgP
ulk1LsvWumfviUAoVU1PaeJUT00rcARhkuy8Gg08qKde/KD63W7Vv9FaG6wu7geU
Y1juIue+uKqztNcG4wpS4e48Jtv72FS5Fc/u9t5TghUKUaR9epC0yULst5gGkS8D
Z5EIghYzbXGfweB9MNSni5q3xfaH1D2AayRuyaQhhguLhmyw5sB8bnIkJZr/gSkE
cc4c+lPSX0sZ/z3mHbAIdEw4yLzkaSwdGTFzeuQxJ7h2nZEjZkGV8GX+RTtvizqc
/kw0GtuX9fUY1JeYj+CH7lXn9uBYxoht4r8EY4vwn92BeL8CElsfro5Fezeu5HUh
qfImHYYrOH8JCsuF9JGLQQOu6zNhYTAiROlP/wYXw2LGp3hqdpKCZ2gSLy4diSTd
fKzBirSWqIgMe/fY/CMF3dSAD0Upd/jCyGQuzPwe4LwKONzm2pUzZocb7Q3YhzU2
tJVIUWxsI620XLYd5/Jz9funq/COSmAkMNif4HnuH5qxHO+9gDv8N/qDZbB6D7gK
cpw2RkLQ3wNMdFapMM887BmbU7Z5dOx+AJ+GZW63APfYUcpvOkS9iGdMHaNljCtq
i4D6czEx3+hP8el3f3rAqR8Mt7ovujz+vs2xBui1cPvamGYpWPI1rq+c7au7oehi
HjYtNbiYhz7J2T7zr1LTiG2BMkoglHcWkgFNOTIqiMKcVKkOMdQtROeUhzJkwiQj
iNB1O9xozA88i0BC82wXHBo01HWd8ZUDJs4Cw88A4lV2u+8PmJ4Td3UXcBPNaYPr
Cs4gIltgXROkZ00gCJkoCqHw4A64Zuh4dWOfgwSLh6Dr2LsPBLLPuCe8UrhZqa+l
dCz4SQPKA8YcTqgkWzxTPxS1PPZFNqde8aKyBYKTbpctMcKXw/iU1KPHRML2UTHX
ZzrFnP/uctWjUKO8/R5IM/lQmnQF5VDkwhQUa5ngAGGb6DGHFi++MWjYqAbYbl8D
h6/0QdT4PuHA8kMQr1+juCnTlNT6ZKPV8qnboqgMw4x6yhvwQnnj41r5Jsa69PN0
IPIVlQjE3cXJPWiAcpSRkPI4YhuTB5gVLKFgvYJ7tqweTLLsxUvSRpGgM3WSkyBB
cIqnxoqjEkyJ3HgyMQ2K9Alk3M+w2q5hF+M0Xzm2NVBfsqIyGFT36HK/1m4k0kLf
TlDpRT2DPS22rXuWwO88y/muOu2KrfxfTz1+06NrfbJAxP7LlosxKRn6RKoEUXXJ
ZVv+TyMGNAuhrdSAWFPuwHwUJFHLMeVTgeWGOd/tDPHPjB3xNWvdLnxCvCf2j6K2
pVjPR1iJ9PVhcTtdsSGRwOOW1SqUXw+1efoj04E9USxyFJggsQD3O27ENMPNVw0r
FfwIJj+rFGg1uPJ4NeThKPgOUNxUrxD/kYuz6pf7Aui3CoBqsp/eC1NPLRVfBXyl
KG6FWxW0/dhzJ/pRR0iDBqrDYd8VswW8sfEacrxzWvkCrTW9raiG11uvWLkWQGiR
pf+D/Rw9zG8njkgVuf2mWdpZkfknRC/Ke3x/my2aFSj1bEiJTfNwcLUtOJQKqxKh
J7N25FfjAGnS3Fql4mgNkNt0ouy/lG+yZfV0e/c/v0VDMMnUC9HdeUSBX+3c6l7O
S4jG7QXmL3fYp23D99+MhhZHwgDo78EeCdH9tQV+DCNOT0hQIXIjjh4T4cOCgYxL
IMe6+k+GtvI93536/9jyqc6nWTvduXE4FRt5z8f660/5X8FJuAygDh/1snGkxkI+
PGjJAGnogprVZ7IXtovikaI30mrQrJMWFWl21zZVLVuPs1i+hGu/gJpKe/gvKEw+
e8F/8wUGu5XwbJ2+Hen15rAS5fT2SwqXqJgSXAOY77F+x4gdRlxirq970EkVGliJ
96Ff91mrXqRJio76jCK7IuET0+8uP6WJxmFK/0Uz7ZvMz/1EE21FAexoSXBmc4b5
mvpC05wujHrUjaycgO3edvyHC27Kf8+3EEmzMk7A1UHYT/cvnzQwNi3Gs+TEpJ+b
LAz0ByusKnwGP6yn4fjsHCXsnCI/EJNRQaLSgrflMz+jWmy+VhVx81WBmIcmkBPD
de5otyt88/e6gFvhoSCe4AD8PiqL5qSDBkH8HkaFy6Zx7V3vHg6ZYcrTodOY2coX
plPZAAjTXYAacQeym3j89NaXYPMcQrD7UqihJlvSOWtvElyqf8DVUwdaDLbYdSHC
RmK6CUyqN1kt7SRytLOXjB2Leype3myMWUAAbh16VedfgNGygJ+IN9EMQhBVqXlq
i7ranEK9v30xWxYbfC+mU92EvGpIzjkxhkOsTNgQrwndAW0+sDU8o3zw8H9qUI6d
eJ9Jv4msVVmg6kD5gY9jqF8mmpsGnaPs0LVaAXw+/OyYrniAQgvvOGWNt9PT7dAp
LQv6Mr7wKFQABqjiflJAARGAH67c1JJmzqGbRUGRA9aXpio/smXehylJRrA2qGok
L/tad2e181yqFjO9e9kD0w4aB5LuGsZBKph6xmK7Hdz8Rd36EHvRmKwpiHUpTq37
EgM4gTJinekTzc1huIt08ZcRrEEMBpZ2lSJyEA4hChaJoE6D0WRr475Bm1zros+J
CQYkt5gn9kGEbK3etAovTIBM2+ZQ2MT6M9OC5P92FcGgyHGK6DE4rcZg977vUsff
MuMwcvped4+KX3NqeVnALqVB6ST/aMbOygOZIT6uXxPS2kNmcgJV0HX3Dkk+w14Y
+15RckD7dv3Wn+AfKm3jaYBgwNubI7wDk4WRiCS+PCGAuSzrwvjEvjR4NCAMhcIo
HvXgGcbKDFDnntwc0+krlKfsIaE/OArrlSBlK6zyIQn0TjsA7u1/gLftSppM1YIw
C+Gk9OnR+aOHjQW29YoO0ddGPW56TlEXv5uqxCKCeiirZRmjSjHsjsEh91ne2WPL
eQiNx0/QQkFFZ6E2pVaL7UDZjbaqObJwgSCPov/RX+n//cDrs05TwGCx4L0wP8fW
974TntqSbSV7w0v3eUGVrjZinFJnlXqgPysJgORvqe17trGAOLLbEMic8sO/mcCr
gwCpX2O4Zdcs3in2z1bDmsM45v2ZOIip/5mrEdPPBnCVm8VihybAu71oXNaLczh9
Vp67JPZCj2fHmRgS5atlv/GsND9Zv+hilH9+QwyFtXVXsIjBVJ3TZiXbfENWCt+a
RqcOqFpVWTLZh03X80kVIKlMe386epZQd0PQqh4WQNnxOo7Colojp458uicB2H/S
/zrUrhkqZX0SHZO9McmvKofpyqCz5TJ5qk5XWmtQl95uYcycveXPwds7AIfABXya
rPKidtf3knXfyBJUgLrqgDgi8uSFPSuQtgD7kIIciFo9QlrD6+jSseSy022/TsDV
tNOnsUz37VFpoGyS2u8leGl2hdyuqlYWNujVjL4GFbP5926zHax4BUmTa4hq/aWa
FNSQ0ZQQUgzAY1HNKbuZzL9CDwWPSUh9kRML/DNFhZrLcrGdZkR+rU7GQPnm6LXU
78fSVBP6XJT6e73gVot8t4CGYF0YL/2GMjnimvzVr8MH1CdKX9zsWNCJ2KrYsPmU
hBBDxyLI6L9oU3k3nq7KJ8zOjYcTR6mumi7NVUL5Ax93MBPrak5XTxDu7/hcEEAb
4coMSRYpmJKbwjxk6+tak3OUryDwl7OwJm+GoOrpFIEPRjXwVZ8fj6/71rCrqy0v
Um/qlQbDaQkC/lTiKy1dH+xKWj7BwCkAVAW8/mTB//S4lOtOOySF8+WZF4rooY65
zVfPGRevdA6TTEgHY7Yk8TpDYqU59cOnAfyukrDpjV0y1aFn1fvEYthWjmCGoX8D
2MVc740RxR3aUYiA3bME9RkXQ1Zlknv0ckRi/SwXWTtPMkCWibKeoysK5Q7gJeuZ
09M+Ux/9exLzAdUX77pMI1ziBKjY72nei38Lrv4rIKIjzDvH2ZoYXfvFEeL5OIU4
7Hjgk/UnZDmmVirGUpD+0tE7+hdfWdUdtWa5z+6mkoLkhRHts/6D+5fzbCcgCL81
sLr7dhBaKw+P4AQpzSXpv0tBLC39BUXEV8Qkihz5h9R8srMHGnu1elXkjhuhFtlZ
XcvH66qYi5fPqmdsRGOpM3J+rKTKaMlV3SxFt8PRGewnQh7I/+yc8Z6gmnXLyFut
Fitv9eTnTn32gZxWj3thGFYueVRyqZ9PUYtBSnTiOiQPdSd0FTHSMtFRSLLWaqqO
PO4+WrlTptbwLq9Lc+RSTU6168Mg7gRkTnt90DMOGHdZtSdnM69xI1kzmmSuxoEZ
kPETO9QxZGkMqDDpRyp2TL932TNftz602setam2nhmOB49z1oDhPpa6sA+qBDWNx
uRN0y5F79hBNi3F9Fs2Z2SjvNbqppBlgGLoMAPMsW9smllV8rt/8J/EgIIkorac2
pOd05cbt0V+9rZYlNwuwXNJky9QjsP7ycuTBYbP0hniwfohEtnRwY8nx/HboBM1m
gQyOz09rz0uRQidvDzKWSb9/77VMG8w0YYXLaJtlHMdYH+HZ7sYER25AzhwrZwhj
/m3E9tTMMWC9pKsiv3Oe0whs6yhNwuYS111kL4FdCTxMg6j1+mNIeV1CkgAvdXyr
Sm7+FZC0/9NpVUMzYPS0JaoY79KEM/kG/P8K2cRuoblo7RLOlwq/qF3lHBW4ww13
aj/eyaHdd7pwIwjEACJ8hRVqm7UHFC+z/YgMla9nf0sPkka1J0rI876ivTOwnB4d
+TJqNb7W9jNXRsmwaVbhUL9G70+ifJGlCNCK+Q8kOy8JCnmZEwFqf8I8MqVyxChC
q3ezdhv6a9rINW2J55R0z26MeXJoiFy7HRZscrg4lWOB+FgB2t6NS9kCStGhr/rD
92MJEfWwjLYWXKPgaCBezuZtgWl1aZvj8ytSh+JyuICNCOvcO+XcE2Hyg/h9M8zU
lCX/yFPXzkZ11rAApPk7Gttlx9eaej4cnwzo2eCcVbBMw9TXhHcmQ6t3LEp+o2Uu
5sWJkNciLCNDWf3t0lvZZJBAlxF1/WXXzGqhoHUr5bC6xWFw/dEFY/Eb+t5ti9K0
nVpbqzL1e5ucbDRANF17J360nLs5EOs/ZbacYMdPNL7UMYcr/68JHlSpvTlPCD4R
h/L667Pwg38yG81kRsf1phU9pFe8f2aCOyVZvHqAHD6JXBYlYmg15MPnfNmdLbjp
+akYwRQo2u/O6Nj9PV9Due+xMRHxEyALJCvRcgnl+fA+SHNPpICChKqLFLICqbhk
zU255MqXonrJajB/Tu5xAaPb9D5bthEwdFoarby0pc1WFKmoMZ6FRHsf1c/X3aN+
m1/q7idKrvCO2yFr/yaCBuprMzxLyUOi2cfdkhH8OBqsPffdF+SkiI7ua5EhRnzb
ph+CL8P9jAFvMNHu/Hhl2Y060Uq9oJ757K3CAgppzijcbKHm7pKlVPBe5MtCuMTz
/8B4i8lBzdQrk29WMTmDPBmcoDFZRHsVDhJbU46VXEqREWx+IBZIA4VRm4SRdnW+
6wfnsSXU+K43b0Nhf3K4/HibGMMi1hv5vUxNAILWtbXHCqjL4UpPPMgjbAWHNmEC
3OjBaZjvSjtkvDo9XwrsqppPGJpu/UzHCwXscWzJ32uqLp5VKrqQ5OUwl/s1DRw8
WNB/SfSP8+ZalZ+3lASN5Y7UylQj9O0W/IveQY+diIvWX/NopcP6Cb05xKot++SA
PSNaDvle1cW1lMpcmdNjvdTxehGLUl4WyXIik9Er1D0cz2amDTgf7xPDP5gCVxdC
E87fdj0/p1OHjFnE4aRgdsJA+/DqTyLrxutJYbh4gfTcoRX13dqbRHqom9l5qcZO
71K9qSGh6FxHGao0X3LY96LG9UrzumrDkSOAm77wcVRQjG29FwcFIfwTL8sQ5bfh
jgWHjbuaYTdLLLe4nwNFlGkRCcHEIHIM9kj34+jKjdbMa3D1ccRVsXoRAK/Hizt2
c5+vhGlYqkgvx7uhDcKdjNNQeWhL9Ryb1uOBBRl+Y5QbIUpyloULpYkn8P/ubKw/
v+zyEG9g4ZPQcnD+2M8hTD2ofancXbHmlSv45WudvvrCzyYkXGK7by/bgRJsOXip
B9ZnWk5ssA32z3C36KceuQ4BVUrOu+n3uO2SiaKtas9FzITKUW14W0mHkNKXwpOL
NOMEXRBXLXOpL1EpYk7EOS+Ty+dnJJykCCYx4Yrt6EgOCxylnvtPeZV9e8ocN3XJ
bY7QvhVs0aZ76WOTrpejZyF3byQeF5/6JutDW9kTQ+k/3K8IbYBpYiCVt46CJfF8
L4qlHmLV83WXpLaQ/mZMsPUo6SI1IdiQs2b+bCFZnUK8V68ISbL9WwU0Y6utHNWG
9m/BO4z2pCdcjQS29Q65OwxtOz0GwgS3z7H2+VqHvpevJxy2cCt+bIiOXoN328h5
KEXN1u3kJTNAwxNkjB2P4Q6P44bBwyk3r6DIOBm23UN8udM/OxpW0/d87JjKKYGa
VUKL7RzTjHuFB2QzZ+BCoEK7jD5fZjgZhPPG6iPpXO38syB72l9QjNsCDZBzNCfR
E0UTPvH/VBwSeDf0hN6FajOixNserxmuBZterSXiv9ytW4VY2aqZP2wDGiTXBlkU
nbwJTycQqDusDyR2k10lKAq6GdVTI2PClTM/HzEy+yxOwy1Lc/+5ToisYg1YYmuV
sxokXRBaZicJFl3ZLv2gTIM3aOfniJgxFNUXuWzT4CiNYP6opt5DL1Sf9HIlwa5M
qLWR9aO7+JOG5yoDjwNbwemPo5xEpN7ByJwQshCKic63QiAuvXULgeIQEhUquKmH
l47hI3j9PFGgFVYlxFEf+dhPowYhrB90Mlgcx5Fu8CLNlcivOCyrbHGot+lf6IEs
62y90yfzFzIP3G+43tRplOrf9MKL4iY48vS8yS94yGB0USY0RAGnXOWg2AKomPRz
33DoUKHrLRY2XhxywpDGYBu8Pys41nxlnI9MGbBU9NxRNKeu5au5PvErR9gWSqO6
WbNY/F7hV6mdCxpO+bxOfNLPItpCaQQO+nFiYX2kVMnX47P/qxI/8xIqJxagfWIL
IVBA28HbQjcex3q806M8ZzIyFTMIjzT8oeZvIX8GQ5odfmozhMbeaH9XnGVSvDPK
/zuGY0cQUMoQpKdx54e9EaAQcsyNlWFKXmucQeejtSWCEDUqtyMQFTBftrdYAiDQ
Uhw/ITIUOJ8uM1szk1GoY6hDpPhJUXCUtNBxaVKUXJeqMA6K9CteDVgkC1fSiAjx
7SDU+JHi9uv7igyhsE7KR8vF4RVHYd3ZBmhl0fMhe/FfbRbtiPZdSLfw7JjhCC7k
+zZrkjgGp+HpiPAQ5Qg13EGvc8KXjZJT4dLoJ/hZUjvpvphngs18ftT7J/M78pE3
yPGyTz0W+kZkUsWpImawEZtK6UnnXpkJFGv+zuFFHZEkGsgnNQPSvWRwlCmJnzmz
UnQ8X9+2imwfVFNO+4kRGDOcDapHDlsuxo170Om3Gh0gOFC2tKjLvuQgSDAuLA2o
95OriA6vhnPHHc8SXRF3BmxVaYv0tL7ouUvvZHUUug8enxXXjPG9vgmQWmIZK3je
e6jfVm5V05oj/BLjVKfQDpO+Xo3dVV0YW23+MeXa0wN3nLlvv3leekpkbtuqclxr
XuzpdHzpwD1ZUm6x1WcI7MJG2BThZtSaAhwvYWqPkpgoTGzwVGGuqeBO6PpvOKFj
ys3zyRPHhZWeL2qhtlp2+LR6HNE2ucBf+eb7s9E4Hji8C+bVEJDzdQHM90rqfWmd
NE2VRfVbYsCARsSWDpyJJdnZeCq8zaC6X3dFuDtJSuaYdybS1Y22baDduCRdcDdM
sFh2B8vZmnUMr6zkXXBf7O3eK+GYwrmfvt1bg4xuxjfnFvDGm9QyjCShUj3GPTaS
2/wPTJk3V3bvKWpjKKJkqLzP2a6beQPlgBjC6jmAWch+4i+GWARMdIkxRipDFb8x
/ZH2ptAs0iSSLRZsBaplvVRvzsqoW5e2Vl00xyPOmBjZrn9vTDemTUrxMAdiGotV
9vhCRAwVGejVTf/9rtwuS6Ylv461ckNTCaq06u551YAc4r3X7MnrLvLCfb3N6xxr
z8idvMawrMwA41PJ/ckEiZ/FY7MrrAI8hz3yFZnRqi+OdyG2lAyglbxe+2V1RnXG
I/17uf5Nrdq6bNNFNAr0PtjnfG0v22cz3lcF3H4iCD09kHSJGHw9N197xqMapInp
huZmGWrtailzQp9dF8ad3Izstb4ZYpiaROU3xqZ1E42ztVIG9/zEzcuz1Ziy3UOa
GE5/wpcrhJO0RbMmGYPqA8taOTDBjDRvkJWluXpF+++3iRUesbkFqwn9DSxikDGX
qBPn+0DBt+X+fddhVzlAoOLPde+x0ulKBgsjASiKwxP2iA5AgSWXBlfi9UgURgES
Dm/DHMkVYMEx6PiepupGVXilfsKIFlzVATtDhow3XW/e8LPwHvC+Xme6lVwssDm7
eFEqwvCr0NMQm/FPfsTjbpIbiYK69jNmy1mQJaH8lnY4iqOOzDbbYDlvhEmHs8aD
oBnfRAAIpoGUEWv7M4a357pIUxF/9r2Eb+8c8TWQsrT335t9Eb8P3S0Jzb2HQQlj
fQ7Q0Xe6flK3Nly5eR9Wrb4VplegZx5tdN52Dl/44kIGu2ea1Wpl6yY8V1Gv9esD
ip5GZjWASnJwYD/wr+Q7i6g/SCe1YPGvJ/1VgT1tbLdnuINu1hnRK9JDcqEdrTjR
taR+IijAEMjD7lDaS5yiiPJqPQw2w++rY+TDTOnOY0bQssTARJzC58qNdeWcbLVF
yEqJAtNAzuYEXoXBRu/S8rNUsJ7y9DDGFn+znbd8dUObpeC0/F1BQq9QxxePeLXX
mfcvb2CeHb6aaj/OycxlG00xx0MLoDaAB6BWRucXvw7n+G20BwIO9es1vbhbM4e2
yQwtOc89tu88wb2X8uA/wfoJEyST4vgQ0naCelfD7m3iJ1aAI3Wer20a4xAhgeMS
za8wSM4SdWaGyX1q2LmYdAbbQmSoMr23bN0ULYkNqUuREePXmdrkpxjhatG5Njz8
I5W3bcBN4NU8QOsNM2EmM8UlLbkMUO9Y30JreUtKtqf9mhujK6/WB8BGfVhh6KnO
lDN3Cg0b9lw25hv1zqp/yHQaRJiClXcCiNk/LGlgf2L3hqMWrek5yzM56mnUMSJZ
cMJKG2GAULYaa3tMrcUQIcU0iFZH8hAnwRaqubt28man7fuVWpjCV6wWQr+mM0ou
9tHMAu+rDAkFhbuh1KnWb0ZD5eObO6ySp8o9NMocuqmqHOPZapnFwemBSwAiqyhu
8jD1oy6YXrfvp8EvWsmgevH8qVn7P/XzRDz9g0qkY86IhpG4CncLB76XbLmQnKS5
6qbUsVrAGccLQ7T8VYhkUB4tGGa/lmhPiSAVAe01EIs5/M74sc8mnvaeQ4fxdAjf
vfpcHaWScaOW03mfHGeyIOB8iDHU5JV3bH0whRxGsxF/TTJZweB6IQRNO+mTNgMc
fytUvptPV7XyJu2+418YOPKQT1sXzJjtJ0t36tlgkIXaJIMRBgRnTTdKyUy64cQe
r5ckrnCON77TRdbYghxoMgae9uZY5hMtoPBHwt+BhyVj7+QmwALHEpTjZebAg3oZ
iQeAi68i09LM4phQyByKvS9oJ+5LSE6BwRG/vGIxQYOCm3Uk9VKemEKy0/VSCIVw
XKStV0btIJnKTTMmTyOWUOQRqf1NfB4VLeqMEJmpTfXGhu32xYm7VnuCejrfWGaF
m5yU7biOVwH5zMjjfmAIrGZ4ZOjaijnAKDVytNgUgswi/RIkk6SajsJrTPJK58Bj
lnYUvQhSpY1M434fzRsub0X0CD/bgYfO7TYTMUd/kw2Z7NGPXh7wlV3AwciOuZgG
QJYM9fkhDbnJSfQ+hrDvqNgOPIf2nrnhXa9La1KvPXv1xQRTI96JKw6V3Kfr0cx2
t84rF7CaO4sGmjT9J+2VI08kuFDSseaqwVDNHbinvGVzpeAHnA+2HMtYqayJr/AE
HlNo5vbL7RHoE4uZPa5GXsOvhHMCKwj0+/w+KnVCWyZXce4D0fSzQmIw3s0epd6H
OR0OdsB+SdpvyRX8NSa4f7wJEa9aQvDKtUqwxzQDcmYlAh/oA1XG308gKUh7U/iP
GpBwYeUdpr3ZFK6Sec6VTDxKMgR0LED4LW+/jhiHT+S519vRWxiDanbS3I74b1ha
KhUbvQR+L1hAEvbozSZdWhkx59QYuK9Rs6iMP5twaKoqevj1Pr7dSxmTRUGEYl3r
lhgFxas84SDotaqU/90x2szqsL0vJ5uCjcDv2GX7buUqOq8qlVgZES/Q2Ga9iJbQ
NBKQGH+wf6fBgl3RqPZHKstHi4REF0I1DBcJcnZUTEF1SeTFcBlEBNu1RD2JhY5i
g0nxLuqyZIQt7hcgKSNKYUkET2A2f3PziQHbUh2Dj0COPC+zb90A8m8l5V2iseZo
++7aivqKu2IhDozBSMnDWy4F97n7xSSmWBSeRtwemSadTPl+vINVVK+ugjoAXOQy
U4/LXx9L2PrLVo4rTWOSy9WyhjwicaxKxftfJPs/i3NZBHeZBLy+I8IPySNPXEvD
znCvpGykhG3Mb6puxh3zid9/4NaQ331+HgMRb8N0YtmHzb32uS8IbWVGSYFdmT8C
7m7JDeiEqR4wM0Uu3HYrDr09d5xGJSLsbaHoBr79vUDcsq0ubvL843J8ss8BgHqw
eXX/0NNnaQXxKvnp2RADCMOFxfS4lA3zgM67smy6eQVkoVgrq7PWw1jaFf+x3vRV
Tby0uV/25r3wmmeDyBZv1/HEwIa4MmUZ6lV/XXaR/sEQGvqKsicobhJ0WhQ1emrE
3iT4uO4VMrv8WyUwjbQr92+okLVsWR+p4nXgJ2YNx2cvTQsujf/QdvnTjTsd3ITS
JTl9/0ZlbqfahEXD+WbKV8OlyY1/Vbh62ViUoeZKVgDxFfgp4iIc8pPiK3eW6NPy
4ink+PQrm6Wuds9p4ppEdE0N/+do/m/oKN6yfSB/uOQHO+rTWAGUEAvzDdFd1E9Z
P17v1Ih2goG5ePRcmhv3IoBXXMqL4PYo4OfI0QmNxYQ33C/bXUfjBvj/rn/Nbwj7
fSW2XDw4x2eSi8L7RmI6Ym8MYqfF+oJ7iO6QotuHdNqHQYO4zAoW8MNXoQrpzOal
kS21fvxX29rXaM+/hEMM0rEqGYKieOlgsDvEvEEZJUmVzojV7ciRCISbtwVe+pH9
pQtZYK3p0aFtzo8Hoisl3/GigWaTPsKwBbkv1vFzWJd3xPBTS3Jg63LwlkWKt7II
nWfMZPHoyE7ApW6P2qOkVPe6mpwYcSQb28SaFsA8/fzH4iGVOj/iJmSKkHEtPDwH
9Y3d/EJDf41bM1KF0J3fEtL/8P8Af5Wrtctuef29ESQirff/bCW/ULuhX8ZLI4Jq
8vBjtnEHLjVhaEH2mdGOmXcX5x0o7XfJ2yg7OTomnoz36GlNYuIOiUaprnpVEklG
riaU8shVx0DHl0Ybl0OUSgF2J6sAOz5tcL5WVoM4RHSJ9PUWJVJgRyxANlwe+ENx
TlKR5ZGUPC+NSGd/vDsQFrgnRta3KFtKt+BUUZlSYabCg1n5xVFzLIiVxQpiZo4S
dNz3BJQuEV1cdSS70YAQ7BWvCiyua1uk56AW9sJRjvFBzsvXVPlnoWdfl4esd9Ae
Edxv8ZiyrUQmZEBTMrT0Zb1tB1PYFhfOTElo82c+5EGiF/rWngLrz1kFabw1gErG
8K9XbYlcRCOG7LD1Tq1AhGhSya4sf/Utr44dyiv62yW6JFdbAIqQMSfhImSTgo4q
DtxVjZuVkHBLrYrI65k/PCQYFjcalcajab2EMnLH/ujCxY3J22eZZJZ4v3sUsK5b
Bo8QCyPsoG7Lw8PAKB6eKHiXJs+k03SNzr3GT5EeOu4Gyyx6UoE9tTpLT8oHCbaq
3xQmCJfOrirEwNmYrQwLz7lxtPKeObawhK8UFxXPVf+n9vk1dTVmfvn2WOxdB1Qs
mvDN727SLy8VVpzmKAa/G0Wb/T2+urzVU0zyreztj4Omj0s4tMtPqtPMoayHdCBo
odTYcuVuOUKxELXRhDXtF6Z+snfoMwBH7ybptxGc8bfdKOiJPcWZmH/uKLJIZOsV
YDqpLB0DxUBS9AF/yIwKjAWRuz3l3KnjMWhowdVxOt8KYnP9nnzo/Tru5VdL4nt9
tD2y2YKC7mOONrQINMjeYEE3M/m398vA+22j4xRYWBb8LC8NEslB4TYzvnwiwgSE
OCI1aZdnXAyPIvpxN4qVfYpJRNkfDFRDK6YAFrFtbCChOMTVPqghGp3RV7fvm38u
jfQU31u+PoowWV0nx1YQbb7+xLXA7eXUoCKsrxZMPHm1Zx42ic38drlvq+W9e+wr
/bTZt8HY46Eu5laAPBxELyqtU9bHNwR6czdB5T3n4uwYZfS0LADOGeqmPNQ4Jq6V
aMkxFxQXdnTEKE1uZhs2llv/tRhsbecqQsOQIgpYORAnOjDmWhmUghVUkEtJsJ7N
15vfhJVc/0rANRrWnh5wesdgBJRr9YXZY9f3M3sMNBoybpZp26SHEKsUim1QJJk9
H2jbg1UhurR1Gy/LuHJK71cUMMwYkHJjxKJXVCbDc5wd1LGZ9ASsqZ7/7241cDwc
ySik29b7NFA5K6v2rlvhN2raFggTNrL98b52xLdSvABMD3MgS2zHtOjGvacUwwBs
bd0rmi0t6A7QyOLHqOVBFLjyJrJvWoaFZ2r+topE1JhJ3chiR5zJOIJAPjI42nDD
dzt8AGU8p00tc0fS03gT+z0gT4flyAV+e1y2C4Zmj4ZdKi0z3y9PZ6AY+dhOIojM
OPA3n+/2ezB3p/dQTsUah7V1o6B1NzWDblSfrPvK5TvKe+41qixUowHwt25fGOGY
4+8tWnmsO8Y65aUYQjARiqYHjaJ7gwCJZobzyiPl7aatAkCAe4HCegOjaizYcuM3
bD+HrDDC3M9Ijyp1IaxARWKZDQ+1ea/mEickRbwpxN5Fmxwqeo8QMKHWuYM2wrPM
vze+pdhEiQFnkH9vCcxsK0q4Aeqh7hrXLO7FAD3E+rjLu+px3bMfzxP4Y67NMQ5G
TYjowKU78NO56IdNvxs6h37RQKlxXUl4YruBHX3G6E1S9f7VvJ3q4UoAiT8RJWot
sGyyGI5cu9vsfIaAGq3gpHfnW7WX6EEQ7RQU4H9AEDWYdjuu3i2eaMlMhhXlY3SW
PON1NhQEbBrw2nL7z0zwhk3haDokr+BSQsJbo+K3TpFBkypGcpA9wJNI6ABLZzyR
qKNSjt5j6ScKRpgmmAdWg93j9tWvP6GlKlgIV2gHtLLOszVPokgJjfYUQAOjRMYP
XXQAnPka3DHtBYoXjpg8qi1t01SLjG+huq4qyViz4qNhNamv95X9XToTdz5DysjL
qRxt25IVjIE7hlriKYdOcUcECnu//vb4e0A6+s1wGHcI6o04cL3IwQEmpWkfWIxT
dkdX/t4+7NcugsPdLb+go4PspbAq759KPlQqhcvvx3dCGXESdori40FTWTwGrhdV
vRfeIbnJW8hMY+ZZ2PDn/NHs1iPkdGW8IhSCOzWWlX8+Y6QpRCV1OGgkEAx+71Qa
OlzwNiBPqsxzfA9eMoPIDdtGK7f/DCjF9mfSbHugmEigZUcyoOz0lw93fs4qldvH
0T+IfYDJgNdONlYvpQX9FTTe9lle1mZhnnGxtFnKbZt7gtNIzWtgZonQj5PbkTKf
UkJIpoWsT4uSFrYarUlSQOq39CZVS1nb5O2LtpanNpzLU2HFSMIqqZMJocTqsVAq
5H8fvV/En0j2NkrfnPn1Yrxr04aMUKzO3Y9EETqJhK/UiA1dwkbIpTeJyKrYWbmo
GqZTYYVmP6cscvJjTaY1WKz90KmN+xu+Un4QQ+p8YFHpUk+y5toLt51UF69elcSn
RtrUTJW9Rq2RajjCKJ3UP4a3vUoO5Iv1Kee2XVxfNuNpbLaf7aRvsAeULlFfZGbw
E/YYkkR1XA2DZO3GY5XIhp9NyZnLnPx1KZgXpNA/DTIRsmO6nLG4IED8bttwt8ie
/5EXDVeX1r7M9ZDf8nUOjm7rBTvfZA4mfj/0YJb3/KqVyEp8xqE0wx2bKJOZZk2I
BgjhOJgvK0AZGSTQhmgYbeWBzpVvfR1HzWy4SVfaQA0nhcxgMBzFiBzyke4Ci/ub
mTlnbGv0db94oJ+w56i7m4wzqMwq3joqtnxGbo0lEfmwjp7QCFsd/Z19xLnEJqHD
ur4paHlRCkL2VfDGvsGK6fHVqZkU6Xrdy2krU87JoapwRbrHcM+JYEyfzS8pZjnZ
ej+Xiwpi2EcKTdE80dmDAGdboAN317J3YVj7ufeMZ3gPr2AAw4SsS3rQpgfQ1grT
MKG2BlUAkmM5Q5EKg+XIrHKx3ZU98dzUDv6905P29uD8sTYBpWSod14+9O/jFDx3
oCQe0C8AQc14jMvJMGYA1gmU/6wv1mEFfcHbn70l2sII6TOAWLxfZq+dbrwN220W
swNnGVwfjwqic2XSOlpU5svfzq0dJ+65FsL1uuCeKpYW1Ewgwb6+Fixf4XyC1Umm
ljbLfA4knd/frvXMzOWCahE8gP+x+8nKc4KMFK7D+VgsPhqZ4eLtWiKFeo8NX2hp
Hhk+RGnPfXEwHXyiQGnADGTnmQjpww8deaOjm15DxwjURg3P3V+C4M0nhjiOhS+O
9gnS1ACi8fMIbLajMS5y+ipx+rmddB4weaRo+AGnRJshDWXEgdJxkBtsDIATPdKD
ZjEPK8M4rQ/cbtEoIPeP5swCMizv0fPjjNKQWU642Q3KGc5WVyhFhMedn5UgROEX
IwgEWq4mOvfO9ZnfIPpo5wpUip6q32xLausjQv8yQJjLgJ6LiAiIghI+RvKvIppy
FKc5cKyTIlx10B2U1YsvSWd4NVe2fgDm1sK++vLUbTdZq8mqY2e8CqQ1Il8I8bsm
+Zn6W5w5ZWMYQmPKVWlSaTSofIFGsGorju4Sy6VZgys6ejMiF1F1wGBNx3YGAl7D
OFD0TmJd1JhDTUPvAMoD08aZFRNvbfnsOVXqJL4VwmDvoroFsfJT+6GF2rR04fcF
6cy1HK5qQj4A9u0yt9zy/sBywF17r+0woWCPze9iKlHTp2l5SfeG5VY6t0eOPwfS
4h/06/gZgXjLdzZ4B5lZ6YV2cqaP3z45l/Eyo7l3n0AOioyu/2LO0vg+9N7f4m90
pxy5VvM8UBGJRUe3PUPwW36O1ek9NrVK7BMVme0ZVhD/2iFDV61JOUbgUqSZlWLy
8NCyaOaaP9n8HUjNPkeWhAFn83wNIQOZmC6DIEsIDoLSRhg0wVVFonJLg6jyZMqP
Co/S4YiB0ruthD2b3IbAYRLf3zHqwGqf1EOSjySf+RV9kZBOQYfJULiw0snkgELi
nrhi9CwCaN4Z01ml0xYQIRRlpCCI3PBoiIhM488sG+A3LmBOmbEMc7/WcS6qikzg
QL+RfgTPLnhYuvoocmXqf2AZOcTk5tuHgcgsLezY/7LB0GlZ8B9q4h0QWHQxgRaY
xqyg6Ktw82NWi5biTV5QboojZVl1nwHqJczh/TFRnZgKUkz39siHrZLtvR04NWAc
KzgSxGOUxxM33U5PpHrkj0bYus4P1/OSZM60oWEHD8XeG2Nn+YuMF9BcaFlLdOvG
Ay3YctoUQgRZ0FcAA3RV6CFK9PQ0PalnxWviKEvM1SkJ1OunqJeCBjRYovxT8rY4
lf20e05y1cIzBvyQ7ZNdnIHNdN23u8ky4e/s1aXdhUXfW5uwO/wLfp3NY4duZKgZ
RAhli8Bjhznfjy97mV5rCcr9pFvjuVszV1bXKnRdV3uMCVYSINTcSDGZ6pTzX8DZ
x5BVUO74/mXe65Iijq0rZ2IG80IY4euYUHI83voKbhy1mNlA92vCrRiYJ9dQhSWI
JbKSxZvF1mgMyr4Zi0kkmDolGfq325mvsah5Xk9hTKRU5DWJLJkxcI2IzYbTsaoq
pqZ/hDco8Ljq61NuoxR8ptSmxoVBZY37gMOwlAimz9u6sfs0KXZlz8f4Q19QnIUL
sBBL4Ge92Mu2zfXO+kAvSYwPKZdYVFUQIRJEXb8ir8MoL7A5TncJHtsDHE2eKSgp
0Hst8mtx/R3f0A2SxOcxhyEGKvQB87XDE9x5ZELp0RtbSfKWLD83itdOhcx4ubUq
9rfSUZr1++f0TMV9l9rX4C6gw0FuBNjhkpqmi8Hx747B7Kn5AvBwLXlGumMNdRnS
f7BTN1mnzM0AySdZmtEzXyCRJJ5wPqLLxsrV3SsolVfWvgr6Lz4I9dsSr5qomW7w
hNfzQ57/dvZzm1Rg89GVcIt3OKMkx2v+rP4AhJgaYxwpQPa89TXeKMMCy9dXith1
kNRsPWNo0zKBaQRw/8WiPJXFOFQ0sZ+RZcJioSEOH4dDeHq/tBcgrDYoqa5zjw+u
I+R4dbf/qybgGE2fDYGGQ7QZyFSUHoSNUbYL21dQi1LTp+V/ChPMjDIwubMes2ui
xnq23XM3u3aY/wg6mSWNZGX2Y/K75+4ehDyfP50SvFs4YSV9KhnKe2813nrTo6K4
qoyVTLXLVkjKlGrlwH0q5hTcHGMKibTyzQI6jMSRQyEtIgtCjm10LVznKXsTB+cy
+WO1MGQp58aGXjxjBjQK+yKgw5MX4GQWxEZRZ/joWHxrtancqvnGynOFEgly9Vsz
iuHs7o0dTpspbbIbTwz3WwtdUg6FfStInK2C7LUC6P4U3htG7ZBAwS+1B2kdrxTT
rW9aqOmtlx/pWXDAkZqJ6IJAf3ZLEC4BjHYov1tBJpVqgsHn9ZiI6Dv5VyoDJUZV
KqlkF2XuPf6EASjJ7QkpfluTtWznEE6TttmnGPJdRnFKg7n3fuz1kAKVcq+/ffDQ
x+Xh0Im9cr0ECdg7nRo5IeKfQ6O/y3Mzd+7AITRUELYiw7Zqx9j8sXkxnrfQ3/jD
XythjM0D2V8G1s4eIyat1np6bemiYFTyWpbTsbpXCHwPmQ375aqmR1qXCgOqeG+f
OW6tNuseq3/6uBnk0gtqpAJ0YwQ3xnAj9ZsC0GPnoa63f1brpZcYU967t17hEPlD
IAgQGk+85hZoS05HO/7IZJ6m9PJPIrqJ07wGWN/V7wTHdbLeKFM0146bKd/M2ORl
2FPBmrZ4H3RJB8FwdbLzwKCBrCk59mjAMP+Mg9WvQQVmO2QKcT51FTU+SEcQlr9G
+XyhmjeJ4MRN+UIJYoLywgI0aoDpAIdDQj3oBNJSdxjCT9ZL9oJiF65v1WvbZ3xe
x+tPCy6RTNcJLmGzI2O0rRcB45o6/JThbJ7OAnUx6mwlAHPGAiYlrbpKVC4izQk9
yMOWOZ3or5RZETtkgMYeG2WrHCWaVURS4DLP2kHlMINUxjUQpgptkAHISz+vYCjQ
auU2EbQtxk3spyqSbDgpDaV9FSM8yQOuqTp2IYkREwn2sTGV/WgV4HXu490yZXhM
g1yVZP/loP7Wt7ueg758L7YGmTaC8RpGr7qmR0EjVrrx/+RLLYjcigHkMlf4dVDB
xF0BLk5U0zxioN5BAVrJzcqXRYMuMv8Kw9vML7J064p/sKfEghZepm9G7iQcrMYY
7K2zVH2sbT50yWmAtwjggvAImykDL9JSu6FXCoOXrjBxLYInjXpDAtExbMA5pj71
0kZJ1rz8LnUaGx1CvvRqe89Tqz8XRDm6rkuDXGvhC02e81muIz6ZnNXaC2lD4oo+
ondCMq/ItLQI056SxBsXIJD1N2dlOC10dsBzTzpZ4P4AmaVookezr67b0lo/1leh
JjpOld7fEVr6b0YFppPXQCLZuijwnlK31jP6wdE9cES6q9UYrbn8xCf2AIyKoOTa
aLwzHS+KEofmTMctAc1uBqcudVVWjt++YvDVrpy/MvTXhETGuCX7dLglUb3U4PJB
RXYINpZP21KnAFyh/CefJ/3KRs51g+YWe2qXms9Z3Dbi+D+rX/mOQWaxHfl2RnQF
FKhg1Q6ytjm6Hoq7OOPXsi9yU4cHo8wl+oxlUFp3v1OVfIKoTzj90nlNALCl63Z4
BghCKbM9C0Mn2/4k36esQn97SXSYN4CuL/4GisD8I3eVPyGY7XAaNF/B1S4h/EQa
PgI/LY0/lLjWtsdF5CrJKprguMaSE1tpZougNcjzq9uXMLl8XyMqOFdzq1CjnzIW
hvmlBf2SLOZB+JSoyaXuQ9TlumBa2OwaLJ6JpMMU5drM6uw8cwGcWdnrlpHSJfIv
SZfrXseu0PcAWnuDsvKTbqf5MKh1UdWkK/6h2ekUSdQKP02IA/3fYJZjzAbUjq+Y
3SrKXFB0KyV9/8HQGUZlDDfYvhSdK9WfhvaBbauhFgcBIlKJ7+q6TECFjN77Bbuk
LhYN6ZBTJbBSNwvVWcXOam8NRvXRXbrrOflJNQqdmU5SnqsSZUYy5ySI4uYIzGoA
XQZGMunf2x45CXZ0lYgyikyVuBcK4V1havCqTpm/lhnJk3M2+zHbraBtwFPpbYO2
saWnblAF+XFAe5sw6GpuZLHypvsyciiza+CnGaa1Skd5kfx2/+/bcTHvAse7I9xq
AC00XC9JFtNm0PkQ73/ZXgYpck5UOuC0IRj1qeG1nEgvjU7pb+xSA6wmcJRIfKHR
Hj6QjMx7YlTMBMJ+FUi10I2ZRKJ94hiutxF+nZqNGeS48Taps7VBMw9EqdpVIqIw
JJwFAkf+K4wmhbVKAAn8n1QOhaJCAnMyuooUVr/32yJV1vGnUwiVeT5XTUCGi9Xi
Pyh2IPUwxVg1cot70zINWv3JA09YJm79h8exCNgpUytBsmmxjkk+0ZPdGMabqUbB
hVrY2pb+KHM+v/uNAUvIHpIkiVBmzauLRkMASyxkSyz45AK8yHXoMb2U+7HmuApQ
vGeP7MEcTs7VDNswIbaI5GeaDS5xrDH9bGnnHfDpEYFLPya5MTLvw+8paQ9ey8De
IJ0ND+SHrl6puA+shAbtuTLTNEgojH/CpUEajPnyjkIEZDqgttOBdD1A1POVlhdr
MQJQtta2jKpzdTvR/IesfcfSd1yP5gnkTx3zaXtPbGMU0D84sP6hER0rhLovt/PR
sMMq758+DIor4DVcijZrXgk4hCBiY0P5Iz2FcB6H97tUy+nFm7gpX38R1P1JaMzO
mSGy2mdoYQgabV3bEmyML7w4+prfRSa5WQ7TWXlghQTRp9APo7OtAsxlC+NF0TlD
uxVYrTJSSBeW6RoXqCf9qx1pLJHIz9LQ+JEwra/75GbIwy5yBOvoeh9PY46hSB+Y
lOcJK4t3Sc8K8wdUB/gkDY14PhMf9SOiY3FXILEoah17TxmIYcWmQt3jCYxNSus7
hy1q/AU28CC9n4YjDlAjuq2gDdJtr56Nh3MmKU9+NdmbeWWvEOyEdO/yPFW21+9v
1zapIzCddPEhbFCXs4kau4bsLdSd9AgPW3hsF1A7PYfBURB/O4D3hGcqBvJq6s+I
LhXMj42NdLnFw5+mnr1Uoe6gUC6nlXe0DJE+aMLiGeuOmCnjghNDQl3Yh7eKMXzH
Y1o3FwDjUH/kR54ws2lEtMsnTWenbMUHNYyYZkRfJLCij2sc+pRrVGrdBvxpRqDu
2uO7LmeiVE/w3zHMn4Kwr0sUUySnapWJnmvFSbxPsUvlsl69WJAo5l4fuYgsyLWM
BJ/VgPycbKe2ZPvbY7h8mfZD9NFBgH9qQbPNYdJcU03f6eVlh0YVMj4M7IPnxcY2
xjAfjJxyBMB3tSh3G1aoAcN/CPSGrkPEk30tH3i+Oe9IQw9D3LHQh8YHN+EmDg2V
+T+tfiBcaZDt4OOOAV8aCWia1znTBUoCxsaxQG1Vcv83a6TU8yckfH1INF51n5/t
9fCI7sEPiTj7Jexiv9Z0oieRdMDiqMrgNNykSqujvSXMQjGADdAXmLtH1S6N2W1E
quFtmEMonkaYVU69MCte+bY6l+yV6Q1bE2VWgN5GPMNWHXWuNvY2y2SJ2cXpRZiO
/1CgDZqG+FJ8wFpwlgBKsPvkAiZQDxESgD1wsPEuLz2XDu0VEs6IzOWRdNyiJIF1
uOjBBFef2h+tLv+xAMvXWDKQUKUNqD0X1P79XnVUb4Rem30QymPCOqy95tckMqsl
XgxxCVzOj1ypKlP4LCTclPVeBgaH+Fcy/5JFe4zdEt7nUQj9mVTS1i7Z4LpGkB2h
ezOkqy1P65P3OYTw48KCYjIkSjMeT5b8reCYjYcJVH+5Meb9CrymzeJm+YHfBWAG
PTHerAGi5lgPB1GKEfj4HRSHiayzONfl+1p5oAVwFNie4bfYrvoM0S/adScSfC9b
XBhVDAHyBXtmhdAFME1zxkOmJOssEO1ANsYIXdwv0zNeMRbjrwcHEKqdXJYAH2ZW
TjxEoMWh9IY/411+IF2bb/NWUU+DAhUSNSgyWV+cyWGWJKBPH/bcz2dOS13DKhZs
k008rAc8phfa0CTnn811c9VQlCIcqjtS7wVW2gkqTwQxxQx9x6pgK3QAO9/OGskJ
qPCbk375yD61Ani7PKfLSnE5fHXJNRGNpyY5/UCY+M/XGaRdzTmPf8UBcf3ZBU/W
RMvcDMKBmf4vUJLtUN3buiPwPuQj3WzfZh3QziVUTZfHD/kstRcOCU3zNjjRRtlw
/2FdaaF90a+y31OBpAtRKd8PxZScLminRS1igDFNHTg/1h0zTaP2cdnlJLpfXfV2
ZNfDmFI2CRhA3nrmPJNjQwhORJgHeSYGt9kBMiLtTd5FtBCo6VB9R+XJy0Wm0lix
CjQI8V+8M5Vio7E3rsY/FKnqRlcR7H2Ky4YnFYV7CyhnJFwb/AYxB7fKmEt2SnAS
KyY7e3uSAS5YgaMDNymZyZ4W4hxlSEy3rj11veVf/6usRcE4D/MxjPxqyxplVAuf
FToYBt5H6KcwRjRQExenB+BcBUHkzoJ/xAqxxC1HVEgI1ODsg52TJLswrbRkEAvZ
B1Cy10ZJ+/TiFKdk5rN+YZhgpZgj0GbzUnRK7p8EAc6sMAGb2tkg/D9I0jpuJPtD
aB6l8IXxKTV/hwHuAVi2vj+/nqQwHee/mk0TkA4MN1HmhSfMoeQ3zVJBDxILPaTG
GlVu5z91HWTHUTGBPk2j3rfvOeIVpVqCKF5cl4lbHMdw7BnijHnZXdLVfToXwuIR
DskOVl3SFcmPwrwP3nndHlARiOM86ltnvvL5wrgL38UKVxcPb1cDp2XMu4Mp+QEi
tE/NY3WuEOfnTqqE1nDviUGaXkA9Nf70fGxIA5Derm8o2yLLYsnZHjtGLDPU72LC
u2hukqUFYGa+6qIFQidnnmSN3/06qWp3eJCOEpaeoVsETJkOUQgoxThmadwd/mGU
+OsekcuEoOh85BeQbsti8h+M0nogH6DI8qsjEhW2qZCINEccGfQEpvL2CWtkyKr+
8dOf1MxagFF1zr084ULQFwl4BgGeQmjRFWOuGHgm6RIIyk5S4zfcpY/Ni9MiEV+b
tDYTzlC/Rs/79pb35pwvalUpy+dww5ohza1dB6DeDNO/bJBmkX2IOk4xs1PlDGUM
T99Tl8nEsElp646ptH9XvfQLwwIVfiGfuKaukuuY4/VwqzUVnUzINzvUJYA/f3MV
yvK4AnQ7Xi7SkZh46nA0ejQ3C1/s9AkkbumP3xxWcE1Ubd88XmDde9VQGOU4u7Mf
VoWPB1XbC4dmN4Ag/3+jncpSw5Vqy2LdISSczRicC7GcredYtRXZhiMP28Zm97S0
B74eHr+BzYSbMrrSxuXPmOAvw1v7qAnUW4IMcgZ93N8xWhxlSN3caUwcXBj1dLzS
sebfYs2sDDMPwJzP7//5ehCpNbpiETtQGh/+ZXZWSZfmIBIUnUkYyRlwZT1Is5Sk
1QoIX3ggydIr6lW/uiq7k/JvYdHb2wZEmFR3SSm0yVdfM5h45qnkrY1prESI1QxI
C60ZjFg+WHaLnHJavcz9ifkvXjrfFp/ity6PlWnX1f++DXabqxrMBtdN3MosM71I
KkelIndMe554mlnzrCPO0rZtzqF38/PFHj9W/NNbk0wGvvTyh4Xamtvqxb7wDYeA
CT0b1nO3nuu53GfdFoh6y1GSMviZFPkBMgiIfbrHmypUDQzFQCzhy4s2YZecNInV
ykROVaAd7edowOA3Z1USgsyOGX9DJST3VqheGBLiD1bd3bGmmp75lYCTpWpfN2Cq
VY8vMlICoE0jxqdYsB33M74ste/7TcoJcKxjh3bYsWsGu/8qEgHfioOV/pAzvzbB
d8At3iRRFy3DyEbvh1+r7Hz8wMhZCD4FXeoJMCfI1nRfgQBkq+JDi2axhh+Y6Pme
WLbOLRIbHde8hViBPZ/xozMtdeB+m2HijFyPEuY9izBBhMCZbByfxDwN9VLdilHD
RN9hYQWwYyvseCGPw/rLKzNxXJ3QnWxlAf8PWritZGbcTS6bt0NbSaXQUhctqZzr
UgmvNTI77xyToZ2TmbG6VFL2pmk5vqJcSgxkR43slNuscqBjUmwvCRIPToJRNYu9
/19nY9jeBr+TaDA6iaAYsBhO9I1SXM2f2Ct7dKd7UDZIppA4GCK/9CK6rHYLiWSm
AmS57ddAm3YvdM1jOi/8MIft2cf82atCQH9XqrVkgwEaF6AzlxbD03rIQ2cuc/2O
rUMOIVLGEdowWwRAmAKHiTdvssH8DlQn36k8UTSLuN/f3lmxptQrzyTK1vPyg8CN
3pHUxCzKwJAP0Q8bN0KHGL6b3BbOCm1b2dY6R7qRP0rGD1Dzi2N/SVfeKCuK5YGD
uH3K6M9Bda9ItwZrkmfQ0sEyL7Gkywty83JpEMF2J1mTmFyaJ0Zhy5tjWGnx/l9m
Hfyv/nAhvBpjuocwl0Eah0tD+IBxsJm2pV407fXE4X9b1u8r9XEbb31/Tx3I4saB
x1Dx2lkl6onzNpkdzIScC3mvDRoffwzIE0xgS4XklPCLBm/9qig8UiMviTiYRr91
K/GHTDhss5PDLTKQiC15dN7QFexeSCcbKwX/Mwdv1y8wDokAiPGiFOLsZm7RuOmX
2IFEOwP2tvnnBp2a4l+Khs3DCYAdJIC0IAZk8k8VZNfttGnxlSR2SKWeyEDIzQw9
/j3+asv4wkIftqF5YKkXPOSpeLhUfaxPKZCrCWkC09OL0IqxXp0xiQP+xJV+E2sL
cu4jRD/rDDqKX3mXsBqjhCRR4BzFTXdBc9G5mmztKhRUMTlu+55Fg2oTqyChjIVP
Xy3ZLDJfAWiXx9vYcW0g/FdNK6ivwpLQRXaCLtYElS168BuwBjy9i9mpCoSuSxeK
ZfTZaMVJEyn4GAG5zCF15dmqpYduy6UW1Ok8aKuhCb4Fkow5PXqQ6wKAMUGvxdQx
zqb/3zfhij1k7sYJQwjGcBfGQe6fULjJ71zT3D0cbj8fVI/5VmiY1wjsRks56zR2
aU/i98US/VP8jJiZTh1KrAoaoEb/QNyLIehFCMEvmXezDiyN8Cam8kc4uVnROgXL
UMl0IgNtqheKhBCNUU8Lf80cgBA+x5MSlaXRkUpea6wKb1Bsx12VPdl3BfCmo+8W
E3u+/5JWGhFOb/sy0/SSrcFdT0LzJoN9nod31RqSl9VzTsB6tCfa4sraKueLp1QB
1kQ6V2i3adeQXVi9YyCWVeZzw5QV9uh5AZCt2urZ9ogzAEnFIfP/55vhvgr+SDMg
KTKRx5b3q2V8xZpEZgbr2EemvrppoNbsshD+3obzSW0ursSFO7SlJ6yvrh6qjOb0
o9yuImYSPSOzumNrLcETZvaZVFfadTcIYodeSitVVfcRmRLuwLymFcDjCCsMBq9b
juIJ4aT/ZcYRHPCn4AXiwNn9S4iWCSr0k7T3aGNsW3QlmykIvcpXSvXNFgsVQ2OE
UnOUAUnQJKzyyEjcRAAPPNNMjngtEFAVTy0H62D2xvIhOFeoUoJ+2JIt7lyFT2ky
frx/QqoIeSb7/pZFx3sZZW+r1T5AfUtN3gZxf0zg9f+uDWayWSANF8Ho7vSMd8UG
RFHzSGKa4T/0A3jCbrR/7uVkXa9e8k/DMa9WOW6ohTOHaLKNLivFtxlAQUG7oE6h
ILfXTjWiE6bGd2cwsEsqUlwevRJsWFWXvFM4uthrkDJnk2wGK84h3CeZGQeW63no
sXbEg+a9FoeMRdMZ1X2Nzs/1pTccwyvmbTxlb+2UfmmhEZmNBebEBd2DZI8AfXrw
kRxbhNofLaqdLQNJ5fj0Ck8p6DZWhbGIJSJl+2c42a0yypN8H+8fuLXnPxY9aMqB
0208RGirvNqwP7i0buSyLHnRD9w8JfTlQIRNCKjWxhOUkMxjL6c0L9xA6WBhniiv
6sI8LctdPOi4DCbFhxQGtyza5Ur3mW7seCiB6Qwcq6RG7RPb313ZXRAMXZM1Z+D6
CXUgr/4043CfCwvmA3z0VF2L2tEw1gPokH/z3ar3zUVjeFSnc5J3QdemXc+90cQW
BKn/4RNHihafAqZ+p1pmVbMwvLiVtdQZsFmbU++n8sKuaHUe4RaTFBWKDMnlAui0
cqw2d+4PGQr9tQv/yLho/GpysvYCYh5q2+u/4oEATmBBx9uGN2I3MkA9e+n7jkWD
vmPhN3WHRS1704qG+wWIhO2cG6RSMwG61BCa/SP5Cx+oOhxdSRP7mqoa5qX2uQdG
Dj4kgYy4DbH+hoyAox+2zCQ9wnw4BSuiJ1Yp1/4H4sp6PxmRuxl6jFM2MW6qctAz
8KOzWvhM/ZtlNj/xdGVEhoeqjeFi1xX7LEfiA5sp5y0eCZpJiRHplF+XYij0vsoo
32YreaqFC+y21dfifULKF4S+UW3YgGiAjrzdCUHvz4hyD7Jk7SMAgu7xtCUaCuZS
LfAodmGAn0HduC+RpnpJyX1dltbqfiQGE63KfB+4+DoEIWfRPPzROoabcf5n3QvU
+5tJj6Um18SkhNolpacV4+r4e8HDY3fXtvF8JrIgA3/UCExSDyNyWZrA2BllgUbD
CyitT49KJp3sLLk3/wPA5kF+pQgUTlDSfIYJrUICrV45g8Oes9sR39UkMIcZYauv
gbMX2hev+a0W7opJlFXWfYSdrjgBaIfswaoeNFpLuTJuDz3BL19zvjDORiBT2pYm
2YzIG0u6VFYCsMSfqUKeoQJj93wlijzQxrbMBKs42aSoEQ1S5OcWiZekjpt/V5Wv
MbH+PaCXv/M37snTAjgaAs02xAygUHRa3DHwdDDtiNGJegp7uQCOyJI6b+D1UUYJ
8Wge7LeCXOI9I30LLXN8TRiQfv40w9Vwy40LQw10a6UevxX69/5LELbbx9xO5ipA
qnVFRJkWnkX2AUqYj/gxdYzTQLB5zjBEVWHnZq3/jjgdUlSljFi0zpnkkQazEUl5
l6iv1OAknq7G+LAzkD0jkdO8BVkTlSi2G1rWWcdsfcWuSEJMmbpkPeEXk+zz9RBJ
VyGIPiBeJcx/XPDotOKHBKc5gkYIQAT+VV3bc2PNibHo7C/mnV8pXExFoco6FATD
bGTQeYKlCcaJeSS8ae5yAyTu0khmtdJLqGBnLe1Qydu3/Z3IB+TXfcil0VBK/4f8
3v3J7BTG+xL6mbz/kV7shujR1q0hSin3gFJJOjABQK5v38ooI2EY5ih1jnDmHqT3
MiW9LAJzPSTrDgJXQrRo78lGJto1VehcoxN86iyb+T5Gxdj6W4+H4q4nDDUgN2Q1
vYvzDOM+V+dSxt6AD7RZ1ra1fDmutV83k3QsG7peOmrxKwMDS9cRtM3qGsnrv4lp
2uwZ9QGm7X/Kvy2R6e8JAQypFQ8R7ka644MB7XwRxTZcmdtdytoCQV+pdSivfuWJ
5STxY4SAde7bLGIdkJP6BE11GDdOXuCxrPF/FoVGGGl1ZViHDkV3XDfIiPCSbCqw
Snf+maoOdCTR066+DB/ygmdRT+Me8qaPB0Y52I3NYiFG3YUsh4Pd0lC3uN5/dCyK
4suG9k/pGWlR0shdmmt8uR9TqYK9UnRRF39kXjv7G7cT9i0tXyHw3G+PdVuupHoy
v4L7E9GFsF+SkjF/wgofUaz6dDDqDUXFyMNZWW/+MxOxTJeNlvB/kLVQikW4wIHq
5OMVYTq9P4cHs7oL1xlIZeEhtWKm19a6qn1VusyE61iU+KMtOAMHhzvHtzUiG8UQ
m5l9owvGDOvzE8m9z5gIfy8gBFI3OfWce3kfOQGrZ1IV3UJM5TfcjJKHeLFai08h
2YWlWFgieXWrdeu5HhIYdfQ5iJjQuVz7TWbsZSR8pmrcXrEveFW9yXWQAd+ySKPz
3xVz4QdPIn2I5Vwl9XqDmggbKSSAkfH/B9JvWjCBbQ6Elimt1G/9tECPGpktF8Yi
VjbfX5vuI37hNDtW+uZUfDpQdmBc0jmMUpcqNVgIf0NgmaNuddkhEFh4X7v6/SO1
/4SfENR+Y8w7iQ7anL7BElzzYfmWKu/s7+YN78vil+a/2hzbrcPwHZyhiEe2tSkG
dBWm66iZVva156VOUqxGpqJZq5LgPfmF2Kp7i41LiBhfW3iVGq5A2wGwjMFcPIFj
nphG+Mz9mnUENcNamaMMBeqsTKfHQMP2bYa+ZZY2lY7Ri4W6a/9OgPS8Cybl4lYF
b3M9VFVbJcrJGXdIO3NHC8rxzmaAdkz+QFTgkre056ip3ulPa0tF2DCrjusXL5eC
ezBRYVrvpSVJV+GKo0j+67zdy5F+1Jl23FSGO74yYxghlcVjiDnFcFI9xZCJg39Y
sS1odFmo0vpBol3LcC1goIV5rUCpov0oKnALi34BlokDvHTKD83INDfGYjAVFX+0
nU470gqt/+VNoACOU4RtMBgnV1U3CngQ/cPwQj1ZG0wv9Ra2IbJR860gvmzwGh9f
GEGfR5EsPChjfZV/fjL0I95Uk8USxDd7Bo6mYT+YjK5EOoN8LoyVuX4JRimO8B0Q
t73FFy+SywaCJLXtCJBIOTNih9VebYkDOiPBfT0LcnClj3d0BX9aRubANw53b5QW
t9YOVE+osxTTAsdMZ7f/aOpr+g6TeSMU21NK1JNgPQRQ/cM2i+IsHnkUpTQ1xdVX
ryqSj1K0qlHjiD3Zv9YiB9a3JZBkgeX/bZ1zD9QGyhCflveTVUlNJiUGc2Ty4En7
JC9PB8h3jPZgqLm+Rg3iGTJbBh0NJqMocsGBWV1tG1/FIrvYiTa3jJwmQAN6IPv0
xkQun+dIto56+rMCjPdC+j5WnYyHAII7kdZ2ZhizvJkDtgkaZR8OR9GInKlBeCGA
1ApLtv1jY3daSgCHBiLvH03E5H5BGvOPF77ztJcApkFoj/EaoeDKKBwGO8EZpPv6
lRglJBqnNmze2zo5v5ua27iRDwHUbhev7IUfbjg/6FOy9exHOO3iV9CnXxtubYZe
V0oJsb+xZ0+0VtEawo1geexDPkjGoBKe+M0JI+9CaTxXuPdjS54GnWGy+Pi++Ger
qaTj5dZJZ7DXHTCul4dRfrWwbb8aC8DzZVdSVEJtAw5SGpg3374tjVXhb+AZG9BK
UijC7NhQaCOZ31wfZeXFtnVCqTuEpD3XVPqclM9DG/oO0YqWpwSMoGcII89ObENG
h4yzxmoXlIxOHDULmV7X5zTtkDi2d90nQC+l6O3omtN5RdPvZ1cy+fXZDVxoQ3gX
RUdAPd5ZfnkwXE8sTLnpvAGfu1PDdKJrX7JnXQOfNVs0fjuQLQf66/NQ+reQXoD5
VmdyPWMKWslgBIm9vSH3g6bfS2/QZaDY2F9qoo9GZNIboWvn4nsrfayvXnE79Cxz
TVpiiVjH093aolZ98jONlG8IxL04w1QLIG2Us1IShJNOmkm5FqRUCqk6zdhDY+Xz
uPC6fzKrJLSbERTJmj+H/5wM9oUYM+6JLrGKcLbbhL6UQqt9GHGAnRCczdaWQSIB
tNzgL1SMlX+ibiW2JOwg2jtIrGrVxOB5ATf3AWv+vZGJVLkjDkHZmFjCtgbLYBC+
1cnrE6gKO5ND44IrIE47ZhJzWf5kgkh9pnNSCLqEbIkw3i1pbHWH1uOhkRt0J/Ya
10rxqBce3s59kTgilEcrlK1AkRRdqgIVC9lZTeMEdUCjp1PuIzdZrm/axkxedr3S
4I1ZPm4NhTdtatrPZG1WWr4O/eoRn+yP+1nl1nnerNkbVIUIxeshfv7n8o6Q1j/U
aOMHrqkcQvE6TPNJSuLmGNg6ShHln33l1DrIxtPMbi7jS61Ok9DvQGfYrHvcZtbb
0IqSx2qvfEJUVu198jH7mW9alSLZBuaRup6R8nMfHdEApNSOEEuyTX6+0CGMxswQ
5poTnn528TDzL7+jPWze0tP3RJubMp0wQJhpJgLnnb2xyHbT6qeWJhVeEhxk7UXJ
9/7e3ItLNHGbli+yqpQ8XLlWENwk3F7CH14zsG4jm6Gqx78hXgqDwPBt3OztPI5g
7A843kLNtDQiv5srL3ftEI6okapTpGIGW5ouifs6i42/0zDq/tFKdQKmNnbgThzl
jsK5p+HvHN5qq2x9GfVYv5haC21GwArgNQG5ozwPCpmWoVIlMGR0WOSijm2oPZUT
FkuI/ka0bzzMhI4HctsSslSp347LeCv997cZJM0D7H1uVauiVLqmhjwt4mP/lHgI
UONeiL4xc/qlkmb4UEenXweZI64/xdtSSt33d+voo9mjgRMjJCQ6JQpxxB/FVc7h
Qp7JYA81M/XQ4aEW3JNZ6LOsO49NVe4rEv/sifItcO5rtUcV7dbkv7BK4Lk5iHC6
IIytdE/YvLZGfl74Lq/Keo1gc33pMLTI7nXwYz4p94O/BxBnM81TrfRztlC8DKvG
wTj+LBbRpXILlTQ596AIiQ+yqFYQcZXYfNZ539WrVkSRX0LNek410xnLWY9oRirf
4WoV2rHtBmljuD/C+NSo7DcuroM+1kQz16ASoJoH9R3QGW9sVCxVpFnrN6S9qhFu
/Tj8javWhXCf+LrDDOioF5jYjgxgtYA+Pq8GVIhNM6D15D3AkHhU/1UvT4m3Qbte
TaAwBXazdDT1YWm7mlGd6JkyGLo4dzgF/6kvQWW7iXGjRDijr5eP/zvDwEuoDdtN
Tei4han7hjbH45LCfeob5DMhLmwhFqUMRtDr/jg7/cI5KH9JwN1hhwWI4CzzvrGq
9wxykCCgUUCFfHWqQPlE/7g14wBHJHGTzPCNgqDOWpNeKnEHUP5mp5p0xLOyCZkU
HQMnmQHVAufciiGl4IX3fv7AHsUmiAosBaKzPwpASDq3qEKhul1bijnbNsoAE3Vg
LNMkerMX0hJBhSv6DRbMM4qz4ewZ4DKyr6trihZn9/3uPvHVDx5u+bwfgv8Lfc80
IjtAOxgFK7Ke/fD99rceXVXNuQWXyq92+aRKHZm8y03ZHZZwKHtTIRjkqBThXKZ9
9ibU3QevU+6Mv42cWsHf2XFcWHkQP9uPB9JMT8GUeG4rirN+Xqf/142Y9OlsBnvA
T13KnC/5KAqJGUz6J2IfuuHxNSbZh5RRvaHS9R7qzfA8/lvtFq/AsXcsm34L3CYb
dUYojQHfLZZO3sVbPndrdKpA6xW8AAn4yxxMawiuSy0NTSG9bHoU1FWQFebVG74a
++37GCbjS8krtem+Qv3FSBnH6Bd1pZLA1RhJZmstkogzcoz4KRFCazbd5gIXurWO
OCJrISW7h5Nn2dKmBmL8tpfEYJjVy2h4mzBxmkszE/sh4A+xOb/XT2Dyz3yDGf1l
UFkmkoIEfiTPynw+GSUq4KnnRJzqEWJaxBmNy86aDqzL2SBo+ajkeQlrOHy4aYvE
sMBhOfrXx6wfJPEPM0J1HoKzvAHun4U7AXo/g5BRMzl7h9fCSUhzqriUu1PsBlKG
QUnbJzW1WU6Av0ykmGnZk0c9XdJ1IjZHlmtbLXs+UkAbKhJPCqXj3dYJCsXbb9cG
4yvjj81UPI+b56dCN9WZeb1LIOJQcXqZGLe3QT9wCYO3GnVhhm/rNI1PQ6nG/idq
9xJwjM0xK7pyrxD63hJTLp8V0n3zwGY6Lv+mcOe3pfg6u+SuUSdS4NB3iBUk6oXG
Pe2+6W5dnVUXGSegqKc/i0lYDDygXtVGYcKzR/OxfISgnIKizzx96NwvOrJMX3FC
p0jRZVqQIveM0O7bKXFxixbPpYvanKcVDT6s/ERVKs6MJeONo3PFmI8XNZ3FZpSb
cpfH1FGnhuFHZEuGAjcC/jTvrQlSmFAsbx+s0QMmjO345wqs1dQpG6vn/4aMVHlh
Dw2lqMH/HIF7AebPehpaAOz5OVXQoJ31+9h53Pbp0p5HKOEqyACOzI/BSE6DbPlW
D4MVQrm739WFqWQjWEkDnx4qUqgZUGEcbnM2ALtOagti8Ix3EC1Dq0SX4UKtrDtu
FKqvp+NbK4Merne6kWKFvu7J7CtOWaik2/uGFrVxg4oekH9qTfcDRiQGc9IziFbN
uOrOnSLVdwsxumgz5hxwpTvMdjmkgxewhrRO/Bw4D/AKfI8ikwDqbzoCUvGuNmlw
vPghQu5JW/PM61NlEtrwj7sBuQRp7r7JY/OIK/B1Y7wSWGAQdsQ/EDdpNqgJwF/K
xuyNSw0Oc+OCt/M5QznDvJJ3ftXtncEdx5iMTmNEIlDREr1qc0MEWrPwbLEFx7IE
xPzORnhv4B3qCSTFSZP9bLIASM/M1ycJ+NAMF7STWSeGTgA5g1fexUlc6hLxNFUD
Cb5fr0fvCS72/SLgaIvq2E/kfNUsuUD9XxATGYwvTqF8x9mfTHnS7GvCQ2n0jU3F
b2uN2jtOaJ5piW2fSw62ZcF7knsln3/AlC51D4yAq4abE4/pgEOn+8rcFMjJNkCk
ffFo6fetkYDGWoQM8oNP0O3rqnQUIuHIPxn4+U5cVHd/xEgOM3cGW1kwz2ZEtSkq
Cf0z1/wWu5od+jVpJ768SY44ZGnxJExAc5NTtEvjuaiJ7g9EcYXfsh5bjfuY8zFN
56MLE0MY7VaArdw8ged6e0Eoc2VKTOZBmfPYOMelqcih4ljCXJi12E88v1/1UCat
/h4xq917IJicZAcG60iiUyqFMAkRZYSPn/npdxz0ODM3WGjRxXI6Vjvl5svMUsC/
FDCpxSD/dLyf87BWQOHvVUtYyTaes+zLWiZ+s5Mr9SuounFKFkiwWUmXnCiZdig+
lNEybZyG4S0dRUMeKwca8pNGNgei+tieDgLIHVzVQB4zEKQZ5XjTCJelLAc0iHGv
2/4Ptl1v8nInB/J7i4EdZ3X+H5LyVJnRDhsvV4kpDseYgIjA62cW4Za1ugIf+JxT
PzG1wP8A/64IGks85/PVuTouQPFxnpx/F8F5xPHrAHTtfILra2U8g+Vk1hmiJcnZ
`pragma protect end_protected
