// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tmN31/bfjWlc9zgM1KF2C9pzMmC7bqlvpzdEQpHa3YI46owYWHTZLoGlx9IJ5+AG
hTVuHdSF0ktSCV8748O040ma452w+z6A+TnPfyehCSuam9USuwN64yIc149ZZZRF
rww3iffIaOF6FUUxmmN7Ey9Zullvylr/8xUp32k/W1Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6400)
KuFnQOV6+BYGfXC3fsvq2Eu4o/5XTkywxEqEM7FX40BCjh+i/BoxKzSa3iEK6E9p
lCcCRkZmZlY2BhU6SA9J1NVQUGnQz2sqVFtbwX43cDD8krRHEaBgRpqkr3ywo4Yn
0x2yz6TkCLMJViiYr82Pzc8sV+UvkbGiXhW9xkshJi/Ii+VKKYxRAxvCQ2oircIw
2tHiaP2XrL9itpvh3AQNNqA0CfwF4FOeQuPO0CBMHVSppe1SOnDxdq/HQi2d+9M/
C+3GjsXUMqE0akrfVKJMQxdGW4KkLWIzhUR8xQE0KbkIRj4u9/2CDkfEI0mJyYKa
0INSxogViqFtokM3tqfrXdGzzizuikyuQpURNuZtu2Q9NFWx1GWzl0MOVzFVqsYy
PhEXnNor3C+ip4lPUJ/ehSwyecsX6AhbgxcczzRJ6fxDrbfj1wDu2SmGobsWw9vW
z4qdOtN0yk+2SxnO2ifHGVVehlPmcAT2ub+EXHpoaIiXdwNc0B4nQQ1932kdsF4I
MN9zizM7Uv8nFznGXQs++r5Fshh53RTD+Iluox/04hGwQDYTOtWKlIsYvKWNWwaY
eaXGajDtoRGEJiLsj3WFjl4Doi+4+lhP7xRgMQlmIZaX3kgUSnf6jU4klwRSThXW
qSy97XFZeJar3AqPlq5oVZ9B1a5co/guI0zonEBPFEYdYTWQFXWCUepb81EPKEQM
HH9B/8M2PTAHNz5kAwAAM4oPIXcniSVmLLwQmCOCWK8HBTq+FhM0rPYL0dOu6reh
mti+VMZAmgN1KIfhXIikSnRZthEZWoyMbHALyXvmZFyexFzIAfWPNIeuxNdkd0Yd
NQ+2cMZw2KSkp7qKB/X3Q6W4tRy1VnbIvpufNMg9AlEGI12FLo3YgaJVPopnFQtj
qZSu83v2Wp0BcwG29yfRcA524EMJThTkQyeYsQAKhcShjVqIpmCaI8UqZ3AgbhnV
/NEBZtYWBLGuJFEfyyPjo8X4YHWu+6Gd+MT0Idh8uvju2YPDNd+K6KEFbpV4gX9X
lNi96ore3rbBz6KxcFm3iomVcGNj+veGJU3Su/j7ajdSYeti/pQAWlY6JEiNDDqY
3VAHHHkOZsva4Ms+h2Iu3osbLen8uEoBcImUIIQf5RhDvuF2yA9uykyr/TmRLR7N
B/eLfnGpdM+fKSOBvYUX9wI3NABMRmpFzObpkjG+kvg+4iixjRlewRn/5pZ/Uyl/
KLNM2pd9ua3BFOAdtv6guHg1Zp+FcmwQL7Q6+TO9LDZLFJ5AHgb2yEGcQBcm6fHu
NbrBoXfzw1iFcwY5K9XtUd41MuvxU6M0n+mlf5dGxFl3lbODIzE2VzS+FjyxCytA
8e8pKmzj/rcVNSXlzysHiJ45tuOcUvRxr6zx1+F/pv0xwLnex/So02ChUd5Rwx/c
T3ckxp7IOTQlQYw/w10QChiIGkPeviDITB1HjCCS+6cShTe+YeNh+eWzYE91kZ1t
QtOKJ87Y+rcZqCiBwC6D8lFqn2ivAejvyc3I2C090GfDdjwIgWv8EsgsxRp8OF0a
k/Tb489S74zH8TybB56SRmA6xLjifaPzCVL1xJcihIssy1+hG8D0oXxg0oJKXLKy
b1+hLpTTGbDmWG7bIHA3wBX78Pa1q6hMgUkWonJt3iCuSVL9xSv4fA1/v3H4oE+V
8Hm3RyMPlPAyXWKKz8VR/55kKY8qMK0hBgOeAqMQAvgmPPxg6OYwbGGTQKhWJg32
j3SULT46eGu0CEaBplv06Xxfxc0KJMq2FQgmOKXLpi9pedjiqOFPnWNkdFW5/1qy
IPQt2EBRnq18vkB3GpKZYV/QLMCQhPiMmUIc4yMgRqrUVugbry96XYLnGuoaHuIl
33MvdHWymfb2SMAVrTHU5uBpkZvhrkvdEU6Pwhy804jJTOLs+9mSVnG+ZleD3p9G
02RdvlCNEbRaT8dx105y8oxTnXvLj2Pb8su8oX5ZRlk4EvqH9o8ZJckAi03fGM1U
gimzpeQQTCfXrFH7A2sFdyU0NgJttAlpExa2T4Vo+KDzYaTGMFBFpAakQQXRPJIK
tDmksHuWk2VbvRgmmtsOQsmZF2uYMQwF46Ov81sa5m3weONYCiShoPB9ztSSzKn+
iKUDv0DRMRLvA+u1Vq75BCvZSr6HzeoqDxQprkFxqa4DZ/fNxbcGbwI4VPwwffd7
HrN5xFhXDey9/5TwgioFkytVyLR6ziZEWr4gqDyEYt24UZ1/t3dpIryoQJ8mf06i
hjK1kznkXeudDS/u8I6uZNhETcuPE1R290Fq7NhBlEG8YAhR/h+6zgbYhNdh3tYI
d6OpZWOEnFxkxixYZIhjw7gLcmRBDeTeaXeqEN5HfAj4HWTciGr+JxU//4CIO+FW
TfvPO9zQvDVx9IcxEcG5t27OTdVwTW71wWx1i1LgbwH1Mw94ggDntYLUuogbymti
xATig2PGNw1mIJl7+QzFgpqocSEuI60ia7gxI5zy5a0nqX6fbiHv/D+lvO4KLyMB
p4R95IIm6N3xWo7vfoX2uySRaAMcIuTQrW1yd+dPdlpMQwZzHEie6EcR358kmq04
mWYnhJJDfHeewA0orAU1+Sw0XZ0d6/ADWipgqjMttSlaR6JNI3Ld/Mvqjt1gwtJP
tpyhRJZJn24QkLgVZ8PJkWK/2eTaU36OTY2Lq6FcXrpMXx/G2pa68zghqZ6cQ2l1
4tpT1sRlO0/ggJM+iqPo5s28egxrsp/kHHMzdGeGEict3NExPqGSj8zq9Ocsgnv0
dHa5hqK2qhDGebNM72pXEK+UxGWjWYNXniYLKZf/tiwdywxuCIsPLXUsFsZBhWLn
rvLTXK3kolOBH/m8l7bHoeI2pZMSogCvxwwhGp0y1n7OoEVQLN4GoDWEVoj+VFNJ
HISYOicYasvafXYv6Eyxsdc2oA0dc1M5FsXEKbqdd4ittXmmO72k7JLWSlQ3aIIy
vNoAp7AkIJlm5spj5FDDfLVo92MLmARd+0SOsSSdDcGU+9BzJQY1Sl0JdAD9zQXT
FXAWH5cjFvsEWmnECUXE9cjLOSR8k61Mhcd6IjNR3S6oo2AHPsYcCt1Mn/5i6fy4
Z6+1U+h/032CHOGF33U+l9ivmgzK8KbItRbTS50A6Jqp/mVnvpDRc444aErsDR0b
R7cpPhJTmrW6moHsQ9NFGgw7v1zPf69x1SvzhBsjRoniRhyiIuUJXTupC8mP6nbo
+IyI1jEXW+pxd9MkCLkDBROmVzvcsUHJ/IK7dX4B5ni7cM5O6bu+gR351BI9TytD
Ieo8BcmnPvOBUKV+1hOW0g1xEk0fs45IbOEGlUiX1gYvNrgWaRvhJlhkj5XFt6RK
JAcXbSP+1109DAg3JsooLl7Kt9B5QFHLnndW8Rkcejle/wC4vTHbymJLlcEtp9Ur
a+sYYQ4ieYuXuVHvTC2kMOXAIiBnP3xEfjXmIYLZygc5rHQlsbuqeZHG65keBoMZ
DdpcEttoChBxzqtzuVo+H6l+wzjtd6P4iXq1LDTWMi4cuI7Yf9m5Y78nvq55+u9i
c4q3SlyiM8a2TxZvsZ86FoyrTbom2gm+XiqEjqg3Z9mwhIvgf/EPPwmoc6SeTgl0
b4y5gwLCJZp2UvyDHvt0COdnOOV/juB3XezV1wV//Fij4d2ZlFLrvLYkZkZMuiB8
L29crKyA9tz5CVqNoRzjxbDmgsC4TkE2O2eGY3rcClLD+WDfUzg5qa4Qus1yGqZQ
bKxM5tMxqxE50QIWUn7O1VRgqWv6pRrBMEpuUlLWQCaDL+hEsUw+PpHcnb36qhyC
UdDRjeljT5CX1IT8g2ERxMOF3GrLLvXfzKD2JbEgZhlXcQzOsCkTuIepN0P9p/64
cTUTunEemSrbyKxqc7f89rFF3T8bzass92EyQFqLdjSXlJVZQbGAPm8+50UxEUWi
zztMFP6C82dCkCPhd/o9B/VX7dhlf2aiPavUFCX6Xe/roG3HR/qdLpzA/6knKLoP
inuwiieekw2PAmm06xdWk03gPWnnKbZkiB1Rv+y89LiEEzuWE/Vs2G6pvnXQ8LX4
7eKO3ABex1lRniy0TnxAR3uoVgR3H9EI7DJzM8rzxzGu/bEizTFS28XI+gIarDI7
MhES+Z7qbK7tIQ+QD/jEeaDzdKjdXYQFDONOufYDwylMZ1HYyHyuQshOQxhnI5zS
QtdqeuAH+vDsE6C9AYekiPaVf90uLg8pPhVmB5wGXinBTsBMho0xm+XNmFJfNHyl
yHwSITTgqcmZzeg9IclXiyWtbyroI4w0rwc+mxLZfaW/ebz6hlVusBRAFg6oJ/4L
X/PobVERkjScT52eQcgPzrfozwHgnVKMQBqmmnl7jpglXSuGEGP0rmEJnc17YrDl
mTSBpqDTu7ajiGasSAuEmNgXtL31krQ2B10LAN/qN0u/M4S3nMeiviRDgsb5MzAj
9ilk3yCNp4/BMIbR5WxwOqJ3Oayv1ZiP9Kwxvdp5c19+B+54IH3yUBwfxX4X6GzU
ibsxGY0gzjTU+b1HOvnMgexdWIW152bQ23qaxMSEUxRQGepOtE8CEdBts5JIbOmA
f6v+Q80mvrzhJ3nhmH8kT1c23OOMpJ+uliKcXNlzSAD2TNstdvJbc3F2DjnlBZGh
Kv9s5+bEkKZ43Jm4FKPTdd5mnFSwqiM8DVgT360L2hVq4WUtfu+Ni2y6UAdxoDja
/awILQYDVL4Sp3mycDQROGlwcPmvrGqotxQCeuMpyKkX51+HxsQ+/7VhcoFz8Jsn
DRt8+zbN3YbXop0aJR024sJ+sFbt6X3Gm5IlO8k6yXFr3rYO2/9j/J8vSny/XvS8
QVfcTfLSGQGEFlWXGtyxICDfZcdttt/ectaes9RzFZu2ym5/g19cwmZti0p52p+a
Ls54YL8o6cJPmfNzbjC7NVdDx+TYN6Xc1I+6Ya20xF0MikY0skOhMysGx65kLTVL
NlG6ceNoPTn4VJyTQJSrjLTPeFkfbp4y89dTq2c182RyaaknrfnMP1lhLuE1UYYh
M4C9PzudCBR1R4MT2ZK5OCwhfK4/UEL7uunV/90UP0sEiEQC3E7lLfkKvSkLBrre
9OKk9A3u66uCUf4ZL0eKTNKbyaB07szT03ALX0z6x6pTvHVJH/xd781OjhQRMeMV
biMOx+9Tj7y95+cFmzqxbOW5gCAv55pQqB/wemn5HXevCMirkzz6StJ6fieYDkT6
h2WTgfufW1hiWnn95/kBR7Yrj0/xdfJ/z6aZ7pJYP1Grb3x+pSDyuNT3c5wU4rdm
gu1fQdMKZtgCLych+VJgvJdTJ7JlV4UtOFDaOTqFmkDOjlfEhs/h1jOcsYlHXFWU
gbnWOTwLUnSdAD8FIB9eSeccs6/cQksyQlYLYwjQkcg0c4p7IGM9M8DW6PWroLqz
xKi1+/WaFFjDJMSl+lYzbjgub7GxwMoyVQc/3ViBBkvSiwHovVH9mXWbibxZ6o6x
CTmJZ2qpygQNgLbrtzov7yxEEvI8uVdlbpH3KtDgxfKH0/CMp+xD3rUAZkKNMS1V
qb6g7LOUzxBhvTmjCiJylY2jN3dywMEJj59a7hL24sPu4QCHUgz7khAh/meg0Iw0
cCCT9P15F8dH0a4BpdvklAiixonVO/cAdRJZXZWjBDQi8fKf5HSbmqEj3yv+/Vcm
Sc7FfCyjJpdHt0gpGhyUXXuEZuS25+HSB0qAkGM7B44/rACMebE5FmCLgUPY21c7
tOId3H2tDqHfaFPyb6maICUOCFpaHVmn6Tba1ZtYBDvrwqyyWJxabUpj3quP9xQr
HXMqI3la08/2ssN7CxrDkdF2xf0Y9vwKxEncHXMYu4xxLMB1gZdu6emcpsVodRbA
Zdv3kSVDQMdTn0r4Mw6nm92QPowqbgm14EuFfGDObX+f4CEhfqaVf5sjwO+r5uwn
slYdGEZU89PSFNIutZm+bBLV3FKcB+giDoMCb3OsYkn3731JB3KCCzV7mDS62srH
lnoO0M1o6rH0ZKzE5vnAct9w3zImbMQ3SrHKc5z2v03Fuk/+hAX8W5HDkt4KL3Qm
fEe6FFAzUifTqtnGQMUdwUygEJs16HNFMJGLUF3DJ8Km3MU0KQCHLt4NlM4o208x
DTMi3ZvkAqfuhFvU+5tE0K4z0/RjbObTsnQ65qjMF5y1uJfL6/xyr2n0+wpERPcx
9YuievZypR9ocldmxg3yURZVr9j1fFSN2lWGlmrENXCWScTviYC0Pf02sSA/YmZ0
0pCPf34bPFsxD+MbHElci3PjHS4Cf7c+8N22ArzrOKnaf3QJSXlNCgdR+60Ut/Jj
/GZlrPW4GxU0sWqqIAcXJbt8rOdzVJydFTHiHDRHG2JcUfMIMQHiLreril5hn7+V
Ur7dzBKX4NtYxaN/YdAco09iiygdX8KCI0VMSFBlFNyTVgTHzBxf+7O7Bb1zWqZ8
cT5yZqcGWqUUMHG1lVKZR3bc50kMDJMf5oXxVBI1vYci9LqSwI7w9EYzY9GVtawS
dfW/XzvkYiyRcBTJ8xgnJRaLVR6hKQhfTN33Ipy9p4/ok3GzhchBkjl1oc82idMZ
74c3DCj2JSx3TC8d2vScQ7rvCmeDkJSI9/I1n41TD96ktU134x93LrGIIVw1OFkj
ZceC+iRZYnf0RzHFd2zNs3eVBx+DlB/6WohUxz+Z4w84ngsy6llu2x1LnjBmUymf
T6hIlDlgjOFx/uVNz06zmaVoLZNshxen/L3IXDQa7tdB8RO2/Ef4PZnELYjurr66
KWJ4utJjkOt2WkHB7iEKX+Snh8al7JzZ7JT87RHZtuABn9UbEQvIUs94EoG1e7L9
BlMKvmksV3VHmFuQkV2V1q3JTWiuPh7RxJV+XqlpzdjOLq2pDMhejlfAsdO/LHaj
8yDS1UFzFdXK8EucCZaqWJyDzLyd8cmjrjEjzLkBqG+SapFvGvdxKrl6wMQU1xdn
WsV2DXDdNU+oqhi20ehZ6U9PEHGzWHdp3EpR08O2/2eNLXqfYlYxJ9cGjAnML+0T
B/vNhiSfYO3kaFqqMpKjiqSDLXxxyyssfK7l94KO+CGMMLbSGAmG6U5C4tQ/BqpY
WfVaI5hEetpW4lDWGYM9j9pIuiyjdm6KcM5c8sAWEtGzfhRsxZDgHZ4HLdH4+KGm
uZQkdKZLoNn32wNZonksFR0cVt+23NkG2T+DmdXv/d67l/8J6IAFhc4hV9w9GZ8C
Yqxv5vxBQwjsEAbKaenfSoMKoyjjAQvN02GVLV8gsliEACZ7TRhw5tXhor1RAvHd
FoBF/p/+hWHL8PvSpbeQplh0SNhdCMLWfqUFhQ9fT1YyevvmUZ1Z0ttqur9zS25d
QgSxnxlLuc/nJ7lOsItUpfUtJQHbmOiM0fm/V/oQQ6He7eOvR9ybTlXSkn7wx5ST
MYxjGbJdwOrdshiPRA7CcPpuJg2WIgi/4fmIAeSLMP9Uw7tSxg0J9i6KoXBdmMNe
2Vu5ztZWSF+89Dwj/tfGBJPwOAkwdx11SdQWPGgrcISAWG1UMp/RgrkTXrwvUodG
yyxCVUGgIEp1tnA8NqeV6KnC86KHS56zLkS/TBbOKbDBq44mgy6rI0PX7sarPqlw
xLyaZTpk5c7MA9SZEVNB0wWJUq2zvD+ej7GEgcKEQ6GgO2HrC28rSK6PhJhor72T
txASrkit7TjUql42LdnWRT2dw+B7IXMt9nMtqIxQDz+4dLJ3X5iToUkWNhoh83Lo
nzGAybTk3OVgOXOVc8/PQ8pH8jlEZICclRRW/bzc8naSaBKQMd90TMDVXYPNAdj1
4Jo2G8IYeMyJxKj3oKW1KAqsX3N0PhW5RhIKfaiQNVqWUQy2xzf2qE/u1p7LLjaZ
zvBcqC2/hGnIDWSANFlGdxaTaql9gjPfkE3LQhvO8nOoMt4V9aQ9nqCTnRSW6pma
+jQ0A+7ZEyrbQqSO4HYTmSg+utUUTU0P1YjJkV+EnylvveRvxyKDvSchscphoQO/
c8xd5dKCmLsLjE90ouSlo2cxTrNEzm6fhTQ0aCgs/FGQj2s/m0zEnSlSJ7e5vUK8
QDutd0o7p1WmJD6U8ikkWkbNHvpxmGdLlF/7c8nYxfW6iO0K6894IOCGsr1rIq9w
3J7aXTBZJ/wE4+2R1nGCBNwZD27kMrZbc96HyG/zh5fRLl1Sh1f6uwsyfkmFHHbJ
RdoUw2nSGuz1unGun8rjh49kcdq9OdYBu2d3zWuLquIHvo96fBgBzRrnTX6zxOXy
l8TRL7T2dqVrSfpebOCf7lzG0CPiRrWZpQGuwkciJ4UdPHozxMGcfBOySyx0L27J
A9jHlidxVKpFCFkI0Km+sGhnAU5YuEimHut8CTnVFLV7hoH6FPO7d/VGoWi7AHep
nNyKCuLoRRBuYgwMxSVZOnFo39g5Nri80uvinx9q4uMlSgNkMUSYCLKqrGe/okhn
81KKYNcrh94SazjoEoLei5LUXpIw97sIDwLUxbJy5SF7gepouECA6p7D6YziT1JI
Rudw6n/iVrz+c8nTwt5h378tumTNXgUd/1oCJUfVYwa1hAp6ImSh1l8zzZq60LTq
9OMeQMJZJQO2CLLxQAQdrw==
`pragma protect end_protected
