// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
X6k3Cc9hU2IxsMvZeRQoQ2Nq323LhFfTKVKvem/V+22ofOX2n3mgyFlapiifThfx
BFnLvYhB6otXfYPNa+EwL7KVn17Z481wTZZ2uGZWFCK6O5zXHEPXWHw5kR6CW+qy
njRW7Xv5/46xuj7PJEYfPiKsGrS9GgqklkP0wYTtGpw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8048)
VniKG11+C80nmno1C6ysA9+PKwV94LLZj3NY7aQx4dIkcVqdUuffY/zwdNm5H/S/
1JQQW58wCnpBoqGeLSIOSsh+7vlL7DbB5gOGONhQ/D1cVoo55HSM37CiKGjtyaVc
btHM1t0b48oEHPPPBbI7n2YoLH+cztsxsHxdZ7lJN8Gcx5xBa9BR3+1dw72LvxXY
vQXDPt70bVJ3tnqwavoDG5cAfCUhpMkbLZDTrLauwAstrJ8tlOiaucvSn39La0t0
AYgZw/YqBIQEBDRe8AhnbyuwplmzTwMoiJfLXJg55N3Ah+W+Ngu/XTZcsRXGgFUI
P0VERCeR+zb1jiLPARGY5dm/3aQzgHc1AVRvTT81L08rJ0SpLEtax8fCA8v2CXQl
ycFEEhf6iHpWWCs6MqbgLgVt/dFTNO910HPccio8VUKFiphA9nHcU8GjhnLbc8dD
upApI8i7XiIkmYoWopgU9Pm3MCm3W7NNv++Hv9Ez0/tcQjJBgLaR4mUD1ctgQJy8
deNV+vA1Eo4dFtQGheva7eo5C5RJEQKw9TLHKYdVCPi+Z0O/GCqn70c33dp2MIA7
qz//OtaSBBNkL3udE/blJPUbvDMVwU5ohx1hdYiXmwo3UEcrnTEkDaAJYhTzHLtB
qEL5OY7zlTeS7VpgYIePcIkXR3go1oDXSnCiSKyLXaiWw5LODkGPrb8tO42EwXLB
Lm9gDfXv2MBE1TyULjefXJtk9htlw1wex7lo8xyWEsBH/RLlPnVQW/ElUseVH8YO
AkN4WVqhwKw0s1uIg5SPs5X1BPW+b3xPWnE9Tebk2ZhCrZh4v9zvwS9mRzzsrfyS
STGSD0is6i1q4LYm9NZE7h65m4fXeaB3AkXEMGJ6a4eoFphG3FYllZBNUf0M4vBr
bygNjxiceQk8sH9bgg9nvFhA58lcUvpKxljxiB668J03Zv4QHgn0spudmYnRNfba
ZowUz+jjeWgtbfnnJlFUTSFROKU5inr47xV7bhQIz2/oorNTKKyt+NGuUAjlAghq
AwbyUD024Ww/a+1cWhp1fKosOQ4OqrluVQ9DzutSfSW45Tjtmo5QZnQSiC02uV7k
LMjAN2nUWJuoYZeF60h9h8KKR9qjGg1AIfeaiyGSiZl+/gEKJDUhKB/KeK3G7Afo
b5NCQ9ncx0QWlrVs0RoSRciE5VlnpCJRu+K070lgdHvMVO3OHCrVYjIjgQyDuPAh
i1o1o200zgRi0MWKEcTUFJ/YMOFFGOrHOtyfP9WkcHrOECpYrnC1VanZMEo2Qt+L
gzQs4GUOifVNiWvauEGI/Jq99NVPUjs0FdGqAdGWbabSOX7175C0IX6a4G7rIjmb
Gg6K5h8Lphya0qVBOvFNJftWlsIpZ+OlYCF2/Gr3gKJdqjVk75MI8TAM/KktAz5j
LQollIYPu/g+3vZ4HSAwOYVycJiGqznpkc1WHBZFMAjeWLDN/M0VBUw0yeFqeGLZ
cQS6/l9iKCaghspJTcKN86UHCTLxNzGyiQ/0dwLhmBxLdDozSvD1ZzCFFwZxqtNC
cwlkpuHzY0eD9GM1woXohwOC89gngauJzILjTBLKFLx1JZsjDwR4KfYdDJnWbxwL
cB3R37Dr7HnfCL44b6ooj5b9YoDXt0YNEkZXBvzoz74pDzVQPSncYHHotcX7IYSS
MS0CrF8MAJXvjQWgFz0kyt3A9R0KI3oz0Vb8dhioahpubpRvSpwRPvWfMEEiQbho
bSN8h0f1akvqF4FH3O/4RpXkjRHcHSimgLimmqfqopaHprge4EAOHljKU7dpSMgi
aKQwSPoVheH+6+zvUkopN4a98Cc/HaL8vYfRJdp2z/hnS/BNtz4iV9RsFWST3N90
g3oaxuidCFTGHkE032SIYWam1LjvvixJn49O7DS9NbAJPZh5zA2hY/2nWpnC+CaU
N0UmSTSM2Sm2fL7UeLA7GjsB/ndEVdSawfkqb/qJGLtaXq7m5aU9Hnz6ZrCF9w95
SfDYkvgfjYLacV3eE2F8ygIh8+i7aaq3PrfP9ox0c2K184biNZ8N6SBJFYnQKIzb
27hqbcXpWfp7L2YNjxWDDUeMtoFtgDNQOuQ4CPoAtvXfwLWVnLmLgFst9Hg5npTj
Gzajky9FmjgPkwMc5lM1cyFtvJOReQZ8Y4wEaYh8fjkVXGyXlLsYeMTofU97dl3P
mE/+AnlDOmz8rSaP7rF4RDLAJtasjeK46el2vbJ0loDbtGbCKDeyyAp4zOILQ1L7
VZ0QrOsxFrgTIxyb2NgryqJTn/8o5m0oTM7QwMKP9desHQekW4t9CuRrHjfy5rtt
pcvPFzwabzBvUaSsX7aaxvPZBrYmVtjiNXdkA732DT5m5mACz9CiNh58RobhjnNk
ScNIIg4S1plcOylK9qHef50ZnW595s4vat4gIyEI2K5jT05+SLMjheQQYzsN5nn5
GmXehSO9QUiH6ENC4iYRtvE+VWTvKTjaVVRN1zW2wPskUxYJzkZhSSkWSxaP38il
aZc36ZeaJETwwQvgaKPQQzJxJHN/TQw+qP04Yv4lc5NC60Rmnp/peMdhlXt8++oy
4WlG5KwKlbEi5ndD6awayxBYEfqr7qWKLX/VvTQPM6GUPKHIkryni1VL3GxCT40I
YXJkFQmxlSd/VicTZfi6VEyRyfPKBp4OOhKrfNeJgeTr61sqhXKlSoUmT6o3VCu6
o+kReNNM/uYkeSujHqMmjSod2ti9a6R8W15yPraScXS54vT+vKcdF9uBEGYg3svm
iqthrpAtsiGN5IL0gRkza9GlJ72FPoOzrncCNxCdW3f9mLe/wqMQ9IhqBe85Qerx
fioaOEVikAF42kvHT/7blpGJJUIn36ikNRtbfmb3/PuHeSgheta3x0T8mJPxvufk
CJw1n6+zSEwU84nl/Zgxc4kXP4BYbA2uEcrVAdm/RWhixIulDU864JY1voYdHryP
wNVmzvq/9WaUDls5SOWOEFyStJxFwxa1kV/df9qZX6RtVtN2C7m77aETv+7ere52
4HVLETu6Q6sf1uA8CWTC5icnqsyjlejvIbYjSQBcZtQCVYIuwGGLRyAOG4GfcbET
Ki/yxPtPbC6sOXV4XL3tBye5d+OqWvZhVlCTXJ4R7+Y/oefLa0jBO47yJR+vP36k
iyGbEm3ua647JJuF6hV662ki12ZvbhPAuArMbNrR84rTRklO4g3HrXWbzB6nDKPd
6xV2QU+bmvAN2U4L95K+P1olsToYlXsPNom3BQfZ2y0x5yvAvOUETe5bvW8KqAaw
J38jZ3+r89Zc5RVUSFPg5fmqXMCNf/xfkO1JXv3SCGAf2z/RDbk2j7iO5tREYfby
orDQn7xDN9RsXlY+WPgIah/MGqMEcCuAM14kosmHVAZMj6q1G24TPfy/f1P5HiPs
MEnYIfEidgmlUFtR0JgY07DLpurYXoEUBGABbZaPsAzgMpBwqnQUUOkmKYnbocMx
1mSQoH8dMIk5JDh2f5LjIkrPH+pkQW+P30o0yhiKFDh41EhdULCZeGwKd66KKx/V
GSy8Iji/JdjhuvenuMueKZ8Tv6wVhJKt9ikzYfmhTOgeE71SaSM0x5OlQkMTjw5C
TKNij+qpbBub9b2Cyup47UC4y8s//8k6lXa3HYnlquzuJGk2tIX+pZq+yGgTqjm0
fO9BqDKjl0EbHU9wnf0XG1KAQsImA3yK3gS0DTiUZovm3wUBDQdgWJaQRdPZqL1H
i4jfPh+hwS3VD2IXyKhnSRSHnRVsr8NkLth7BDcoNt9cI5wGy3vzUwkIM2brQ4gW
r7W8Y4IBiJi0dB7K7xLlMuZ96RfsgJVeF1nocWwHruMiOQKfE1fEZzKsMW8+FvUU
XGAkJk5FV5YOdZmYxW/dqFrHQEg1EfUeLxJ/VM2Wc01aqhEqwAzJlDNTnBMPe/cE
VWkNCqUv4plnutxRxIka6v/hqDxDCxcWLSyAQ+upYXH0F2MMUAmYurMISyL8Tdlu
Y89UmQpaI1ZGscQ4lE2JF4vNvW3LWTzeCD+wLVCjs0XEdjfMX5uxoLaPM4QwIeeb
QYdySJD+xtmfSeUEu2Ewx8bVOSU3nfErM/klJzXJBh667DzRVgTnIztrrYwkjD1Z
DSMtioEfezlRwEqnxUWct/TexORBJel7nWVXsoAOuEya4Z2jQ5XwbRQcZsAAZ7FC
YedWrc7IShwJ5BgSotdVOsMP42MmVh3JOtIynCcQIo77EWusuxTyc9l9tYcnMp0w
kOsII9dP3L3W+6vjRUDSSm1AbAAGj2/nAdMLkLcIIJujwCBkO92Y+4WXrnbak09c
yZdEwyrhdaNMlpNxVbmW1VZYDi674PkhIt3uZOD1EOXZX797cqEO/3CrgD+Q/G3I
2cPDYwUvNKbCaHkDbU3++Hu4a1qEe0aPQQTVPz5B3F7u707QOgb6BfYD266u90sO
cy0ikoMaJSAqnT6w/V8l63fKjW4xHCgj6/zWvwYqytNZtsLS7L5wylp0HYK+1UA0
zErgWKxfAXSjWC7GUcbvpvIhsFz4EZpjomC+zNiPDUE74ipHfjEpNYuulTaLdiE2
kCWnA9/YilslR47S/op0zpeNIuuisoF11UYT8D/WsVDi+h4iXE/ZQ61rSicS8ipM
kflnxKdNZAdxTWiHr0prpgWLpjLxP7BRNVOEGgWBHGxqFRUht6Wdv1OGyCcJGKEu
Kpvg1xbFAW1/e3s50bU1GTEFARnhd8eA5iLmCk5xcYocS7Gr+vcF+Gq4sQKej3l5
WmRHgNLvC2AHB7b0N25FwVLZek8U0kFQnrSz2jtNsfZ79TOC4eELA4wFzLcKcT3G
mXZgtaeagWTayXu8/Z6Ns9PMavlb9i6F4/+UaE0CKudYNwwXELYQvrch/Qiz5WL6
lPPVkligupbuYFB0IHFHUJfgafACAbobTM3YTGgEmJJCmx4YkIi2CDJUQrbgKkxB
ET2bB0KfZt2gR7Mf4a0WsZR/Jy4MbQY+llHs7kUkJ8Hh5uLOpz0+smEWDdDNAqLH
e8RuZsoIFgc30l9FWqEgOhJYotmNyai4eRVIkNoffbHIaAhP9ME4FjHaxdsfaDQa
CJ8VlEKbDo7vMdmYCamA67atzJK23FHzkHqu1DHkd8eSmxh5t6YQ8Mw3Djosuvs0
EgyZuBQt7/2xthbmwX4h1DPEg7qUB1HysBaQtlTBCboTQi2xmZS7aw1r2TbgwDfe
JLXdjMD3J2VIdy/W472EZ12FvRXvx5i3hI1muO8zp2/RF7uZ3varLHLySp+j9O+x
9JUYmvKQp+l6fdI8mXPwuxPahki6OV0FQYVUrt6tpHAxBsFyvZ61KM/g9t8NpOfD
Ny4gvknyIhZcwtyUTec8z0d7o+UsG91y+xJsXkrdPHeDvtltNJ8QqkGj7bzz8lzu
YwP3yjBp+DbkpllA481zrf4W03OpZTIWRWOiMB7DjKEw5UsW64MrtkG+NiiU/D2x
VT8k4WPooSv00jBwo+sTJxCTRmmXkleN33MLltEDPs3fiJRQySWL+MheVJ/Det4y
22ICPEQy3uqblG9c38ay2bb31ckkO05lxqp+IgOQMFZhoK5J/RLRDK+BoLBrc+P5
orOcoTxaMLotIGi5DxMIZfCUDjJvD9x8uq+3YZNLGHGWZenR79uj3G1ZNpIBI+cx
0kTG54O5JoZelbx10EKg6cCcJBgwZZnWRjrko81kuvYIlcjyW6mzHoKxsILlsmyI
rFuyoED6HBE8Sf6V8EdUqFh6yjefCSOgbGNUmDQXpLIOQXml1qD/MzJr/ENX1oTl
EepoopKn/9Ti4uXXjtcZMcDj+CFhaa2EMKBzUMJZCkXgOgelq7T0Q7BPJxC0WTkU
TI9e+5DDyGbgdPhN+2/V2S51yyVwSARDck2Mb/yTaTQuyRamqgL9c2uQPIOtKYKc
zd4UiGnPsnAJ0Tvfj5YPWqWHfWAYS+m04f23C8MFil7p3zFvDgdqYZbGdZ6yKpjT
V14nYgUwO5Nr5vq9ZBaZVaWeU8h5NlTuvdZZvtd1KkQZ4ysjM4Kn/c79olKMdnhL
5J2hIfYPScSGuGMxIHC5BVVL7WYOtLdGeqf4RJimzYq5p07I1uC8USlG0/sQ0TVM
4DMuMD3mXqt0DbuZQ7qEDybRLDTNMW76lFC3OUzS7omf3OGBlWfdUlRLIMTpPBGD
DaFOrUlKY4bKVeJjk9nVkIIPHqKeJAMBCmTIfKrnxeSZFXPPu2wBVr+/lbVWXrSL
fnAl55WGdwlMpV2L8bo1xXRQF4l5E00t3wUGm3HOvHTq0c5RCKSVaOKICYmgtwj+
zznx2LZb/5AMglsqhWdnHpUQzxQizR4+4dHWjtbxQUI1YCWIH+RJ3xRZITcHmyy/
fXR5KLProVvYVf38OWK9ES1N4mWzC4mXmAC1OvqkySZSWC7bCQxk0+wEpQ8+4SCh
Mfdz3VRjih4fLAW7oDGsI4L4ECexenZ0zSWrmNsviSZE1mMgD6xe5+O0Jhv2hw/q
T2MDST39cTLG0dQ2mskt4l6/Gql/plADGWKG70LhR0kKz5qbfkQW/5ZjpxA+aNEE
Z9kZBOpF/oln/Hg6nWiU4bOoFY7UKmSb4LRWby91C0J5mMAiyrcS8n9AjDxNcT87
FOOqDf/OVxZXuoMhEOh41EN6+/6QXkhL7dA4WvrljZO0TAVQMZnAvOOLpfmoZDQ5
jrzaHlvxFgCIRMUKT/VGSWFihZaxfqqHkOHNB4hLmDqwjo2+5ZHncomAKlL/QbGe
N/NxWjdNMy7Ee26E7HwM6tWJ2G+PEriIt+fTyx5VGRK6kz8ASo2FV7V5TjAZp2tQ
SrWF9ExiuSLGM+ZFULezbEMrRwUT3JLrx3aokvQpkJOUcKbkkhR7KRgAsyJS+xwf
1taKSucidCEejOYeTPDxdGWcEpxkEY4jvV/kSHJP4K9wFjfZPk3aOOetYVHNKoDH
6z1KdxSR9d3WtvCB54u34z5ywKRLiQaUq3DAoiNG3avuiTdFf2kmR8zu3HpBjMuo
rC/2QJG7Kb2hbVxo26iWC7G+MJQW0Br/gpBjBWlu9RBGEUgYxffq002cqdDKfuZ5
t7dh8WpkJ6bXeTpsRLQ6ftvVDmJe8/+vfCSWHYzZz62yEg6iwFyQ3uRK+HhruDes
v1vA79HrP12BUMPCXs4RkwVsSwfNVqgfXtvo+fAd+n7bG1gjGp567C8qaiXKhdsi
3hD8+Ru3HyD5OSyISXVT8C5Wyk3VRlpT5aZx2xYIQ4W7K9zhoTh8qLQzvmcfgepp
N4B8Ja+ZRVd6hD3Bagk0hbMdUQhuokON6Jzr5Ypkw8+24bUva14afEu395vj3h1C
8NoOGfggfUj+Oc9cC68bwk35rUjU8Sqn9MftrsFRkPo+LMomBArtghvulRiIZSkJ
/rHhb4Wg2fmx2DFanayhFSyjvl/bYr8aTXCdtpby4Y22+bYGrrBaL2FA17yHo8hk
3yxFLlSQ9rQNhvZJIiJ/+pNkOGhMimH9C8Jvtf6b10nR048wfgQ44buuJkrEjHpQ
elcryzXQlkvZWMB9+mJ/gXfvzeMe+ghDwc4/dUUNWG+Nto68juW+xVUySvNok/ph
JaU2nxclJn6aR8pqAoRz2fCiHP0gmg3GgnbTrU9zxqG/yEkzzJAzOYqkY2BML+00
Y2CgaE6GEP/V41Hicqi3JfGllgB5Js5IQmklKSQ9OsijGasdA29ocF88HRCnmM6O
dJNUQYL5ghi7gDn/QXXvtAPirJScp4YZ7dF5KHbgbEnAe5E+o8DX5rTSDrRMqIPL
5UwdI8Ya3m/Nfa74A/yBs8go2+K06/u2o8zbruLat8UUXIVZZFzVzq/o2rbK7JjP
0UVr7u7Ba4n/3gagkZ7DIb/+mI3JYj7z30upP7aNKRHbcyob3zOFwSb6wpE8p+z6
pmKVwblU6MNx3Sx9hfL48h7d/7ztzxVFfH3MOnrO8IBjodjIJzNF+qHfBs+sSKAj
sZEEUpkJqgaidKOm6JqsuA1pcob/UDjOwSpLeZ5+9OYZpKJsiFtgY9XNsXVlj21G
PqpSJhGqznsoko7uAE8Me4Cf/yIZ/rrMvEwHheWAuFEvnQsbw97Pey+HPUldZeTq
Tb7R5ZSbVZQbiU0KN3yCg7MGRMme/iZfYXULSNryc2GlUxYNHOzuU3Ji2tRAEsMx
YZs8SnnlY/VFzjQaT6qF0HchJ9UodMD+8TvOj42uNh4rxNWUfb6dj2Pvzpif0xf2
lcaSYnuGu9IZkEbGGt/0xRVCs9BMprkQw65eq6F9KGZyWmthCw2ol8Te9pYul5Vq
kAthe0Hb1pfMnlxn4DTATfhZWi2CGRjlgF/pNEh37CQ32X0JDORoGdnPGiPHHGG7
7mflpg8WM2T4UAO/Aq3/ckU5kCmdUU819KOVNS7YjHdHE4bhw1JNTCBBb4tIAgmb
2gcteokqRxsQc3rFFDmvbiaUkmBhglrKaJL5c+Ly51MJ5vhWnd4umWH2JrskhOTm
srKalfLRlEW43j8K9rmlqdx6aabkxlqg7/MWYQS5OJ15spBsjb6cHtnbccqffjc7
WsCOqar+EgEmEaLqaYil2qYFkE4DPuvjtHZWrXxh5Rn4CPffklefidq4VAAAabT0
EmvPFa4NeAIVq3HX9dROhGuFuM8T0T7uNCavOMiyKdImEJIVYzhF1tMxw22FS+0l
KYGFjxFwOxJx+C/lU1Za7UsbT5QIAz7fcSxpS4AxFXLd9PG3tKT+gr/yGNJibno0
yd96JrP+sAb5rWs2ett7v6OfzstlgSDJ6lBt304acr6W0ZmADaIL1xUbMXovwIM2
Q3MtfY2cL2Wk0U3A1A+E/8K3kLZGiVgTm/gG8UJoJ6+QI97H1IhK8pQTImlB7wDv
cjHduCp+CzxOR13+kaj9Ns8+gcz92WVSnDWYQ8YXJ3InJ5UdVig7I/Y3e6Bj4VVz
UDvT3fjZ+E5Q8EkICgDolo4M0TAHcAr5kWk1avBfTBkDILFb8GU9kzV02TaLRfmD
KEzuKb0lm4U0YYKTUMD8J81azhqTMZz/WSz5dKW3mRn9TeSt3EHlxwX+IHqoKGyd
BilkpAyujG3fzvYXefTFs8zgfjeWXoh5nZ25mjT9rpZ7XWVKyPEeNl1UnteS+ARN
N5nTGO2/qz0MZ6jd7ZOwcm/sNo72KR82FpwKffheK4opKWaACL9EHZ7gvS0dhS9r
cN26rTV7CrdgemxXFbdAhlLyaLAvRErXt0iDJwzgIQ5mjQqOEqjgrckGGDfknrBO
mI5ZBG8587SEBjzPTD7hZ/qLSkFmX24QjzkftYV+OzPUDh7keq2IUXNdd0DmAbhl
pdi7+cQAJ5fWSC50Jd6C3IaMK/PRGhNqTNtJYGZQcjOJ2lFndEiOEwwkvbnoJHLa
YsU5/awkpa9IXzQQWMbJ7yC8NMoGicBF32X8C9LnvQ1l6GGHD8vTtlmJ5+f7Bzfs
Wh/CgY7ZBP3QF08wa5T2ZH60N2cY102Xqz/gJaGxaRvyOS41fqtib4ExCeefqw6K
HPUcFImJKkztOVZLYhrQYrXhdJBLqqSktFgu7YJUvZ6W4JXSEoUstcR+AaUtrft2
WxYsd5M8XAzgwTVesDhFJCjWBYFa3RDZkAPsjCCK2V8lBaWh//Yq1ymDpPjnHIQb
NrVwnL4GcUSds65P8DuQfVciYxKldEd2M6ts4cVAyTHF+FtAbtxi6SWoV4pAltr7
iI5CwCX+flXHsRRclWS2xuJKQnAc7V0ZiyRRqi6QuKmB32kFfkiGdVrEf1GxSHeO
HHFZ/ouwrrk837em4Hv0T/cIGwbs48v7Ic3yQZb7KaKWFS5B6s0Zam7m6wSBOW3G
vhjh25g8P4/dxUnrTaePsLkv0pMUl0ZAuhh/eDoMtM65jxwvZhNwzvqFSeDdGJ8i
xkiyNTfxCmhl/5vll4oO7R6PhaEYbQMz0wdIWOrxYIW/XRA5v/oedOxSpoYm3ocX
xpeLVI6TW8x+6buW6V9/aqyQ5U8Df+YhEml4GLV8gMk8PRv3S+37mRw9BtnWSvYu
5rtk9/pFT7nCrBT8QBUSiA7+QT7h6lOjxWdIyESBpRvuG3AG7RMsvNFuLXbwxVIY
MpnYCVcdBwjgCERIjPDEuXT77DZ9XcvTAIlsc9y4PXe9P87zDjgXzi1nxOgVfaI5
Y9GN/wG/2j26KzLDdAVqDR3r4IYNAGRTYlPyFjP124p1hje4WD9tkWYqSqaZsQBi
wOJRLF9E4F23sIxBas9a3oohlTiBGXGOab5gXl6d1XwtQ38o1C6jr65UHDQ2UgZ3
5Ml7MHfcF7wPEUhVKj8Sc529vjXGDBde91OH31WrjRc5mFKruo1HwU3Z4y64GVHF
s2rQWSVrQx7pT7U15ERTqivbxL0DTlZvHMweb092eksv5B9aKgOaMnSlprYZ5tYP
Wpzzjf/Mc/mCqAnNs+CkMcb7wEvY4X4j0UbaIzkAh/X6sQLlS6fAHN5NrI07p+qI
f4hE62e+6lBJN1lvxSjBCFY2ZMIQcJI9/VlYfjOcNnrpMJ0qpZ8yrUoeqRJ2ki2r
cV8id0/deqORN6lljxq2mMwq9BmCWI2+QXHvonEHM2EPgPgo+496drqHgPceYdhC
ReN8uym+Z7lmvKWb1m/Iq6l3X9fvR7eN+Wu0EDQVlgUp6YefloxdtbYt1IwB91p4
Sf++3w7oSAGRbeBCG8esdSd3DwIfSVW4DrYnAU0G32H4Af+Q59RPqj0XcS3hRWNs
XpYD5+lHDHVrTcEf+1sgd8uEaxJgen6HyzJ6J2fl8RA=
`pragma protect end_protected
