library verilog;
use verilog.vl_types.all;
entity unsign_vlg_vec_tst is
end unsign_vlg_vec_tst;
