// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:52 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EmGdKbLvZg1XPcOK/Cv8AIaeIrUoYv68Pj9lRESsQJxLR2Xb8bu54Eq7S5wYfQ9D
cwndjR3HiEVwRmcXhRja0tGLOQ2VAVx/wGhirkINelnzn/uAd/hTWYSfp4K1Sh0U
DFEv5gDg6leyaZauMJw/V2O1a7S8W8RJBH5lHVpXs5o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8720)
pHN8/9H0jgXjQGpCjvrKcHeX+mj7cjxFyDyEjF0X2sgfHYjJTzpD+q7Vt/3yvA9O
JvTKzWZ2lHqPd+FiFNFr4rpd5N5Ju1z2BESPfseIFh4XL689AtNqxcT9DM6Mpzn6
QguobnvPNg8bn9eUfYqxIYYie//eO3JnYY7VA01CNntPiz726QS2J3NfcMmFgrer
OuMmA0C38ZTwjHE6Kar7x/uAKxYPK6LRjFWB3qASdIuNa/ewR5lRTdkpfTkGSCzT
Ebv6xjr0C9k2PHDrNJ/nL78Oo0GPldqY9zpL/uwK9J6cVP9NfH9dDBJwChbIyYj4
3VMh0ZniM0TLOaEVAvDuaeW8Zqy0D40Ezj6WdRa6m4SZKjn9RstJRtEwaTg1wrwh
2c0kot2palNDO2pbLyqhichXQbT6l5bquBBoEUdPtK/n7GFYiYdHKPByx0Ca5pBW
UIVtxQUrVxgz/do2X05gn6tAhcGutShjgTgRhuYTS+w0PbPBJ86eD2mY2365x2eE
qOZlRtoQDO+MWUuhgLTX5J6qLA3cCRlO5GFca+m4WwlBUbNhMgSPlJ7IFMTxFjEk
f96kgO1YNhpbCqdZI/JmHrjvgJFOqBYqcI2JbOoM+5o4Kt1Wf2UMensdn7/Hnak4
DvApj45Laa6VRhjb5nUiOoEJR2FOa7IlP1UHlTK7FACoZco9k5yN1kgBXtox/XgI
8Cr5vmFgYxjPXNRFCZZxMdY2cJ+jze3YUSd1Xe8DAi6bXcUFKtPNOMu3WzQYL7Lo
5ZQJ+g/hXAO8YgMXFhWlLNEmeiNqbESPbu4T1hFRZ6GEAtLxWzNOQxdJvyYa3SmD
eFQDHPk+Ir+TolFTW32Ii0eo3G9exeOc9/9iseE+GUZB4OewVhvJHDz4+VP9AuLD
kYyrmt37TUc3t/6CvYB1Ony8AKJVfn4cLyHrMp/PS2fkUevL/NPHhnMPc64LmnUs
xfdCVw9Ir/vONC9eFbAmX2U/k6elEFesHl2IXBydnNdmc/EItcqot0bnAE7I4RhK
BlqMZMRPSFQlMMbMMiPnOUUkg6Yv11zPfsTjm7615W1620s0fNctg/MhI+G12jp1
11OeNvDz2XrXWdEGyjI9LJrExbHo9Si3RV5kYVNS5UerjPgj/uuY/AMSjykOrkuh
HV4QbVgw+GqpOuKJjAO0LktcipMrT0HDCbHzYKG2eubQChW/mdA23gXVbDmvwN4S
oH+VCQG0vGyGb6y9UwSYk/lvlrwrRmzjqV8KjpkpeeVAVes6EfP6cbxyKpo3qg5F
1Gjvxlr1ZXH4Qmx5kBpUQoJDS9ZxaogdO1YzlDAp+QsN7bTzBXuiylnLRh7Nb5x6
Tporm7v1O7DlNuV3w3hLGJLEUeA1Y/oWir63Dp7/isnd7ASTFknuKlgRidMmVL8r
+eTK8tQRREy86Sv+2g2gsw7Rxo9Ylmu2nNMPxrP8vakvTqCHD3Ph8EYEjc0/LTNT
uJioXISfr6q7spXhuqw1jE5jQKXhyOclIfqkotOGJXNHbfAtWLh1pd1q6KjA7bWo
ypvpib8jul75ZsnK2GVhfFhEfIFij+WYLTwkhHMwsGDXegnsWCyCq/4HCCd3qrxL
mrX44tKLXUuwlKCoD6NqfcnnCANdYP+X2zGoDKekxaaUm8kIoWD/A/rrtczbvGqb
1ZLZl5AF7kffwMRNk3NMkJWZWfjmPtXcTcGEA1+m26m6OwNU+MB52UTS/kotp7qX
A9+2jpoHdLKPu2uESbdxYW7Juuq1P15tVhXjH6OiMEfE4g/XcyfLhWSevIlhH+qU
wA4xNJCUCJH2Ozj5422cxpmxQJ/HjxVVZ+WnFyHaJ+n0EPfx8MY5tYzu0+7kfkMi
U3eJ35+0sJy0D4g/gCmASWS8g4+9jSFfSZ+kVRRB4UIcASdnbH8igtYQJtJ6tZA0
fzK/9Y6fKbmWXrUE1vlSV+H0KLM0ICERiwn1n3skfIVO4OOW2naXaYPa8B7Ug/eA
FWW4ODx5Jit10Q8NHv4JIvvnI9ssImeibfas+w/rHtOwqLpR688ikRQ46yQJlF3N
JdnPLTZ6asw+/YPrsbZavZ6fCp1KDbZf9F2FQkd5yuerqVClpoEjK3Q4Hm3SLXlR
XDA9vmEdS6DMl/W8rXLsPOH66VPv1y69jgyUPBllh+FyehKW6fcjjzNXfy6I0Zgw
9sAD9CnwoSCafv5JycB3sUrsGZb7C6VrHgGQQ/EM/DDyZzVA4l0PL7gjDo19MbSk
jKS34HzMhYUAoWNVFMcqAPMLmA8Pqulo5KeOiT/Hk/cKobGfATKoCaydqBus9Qaw
1rz7OcETS3mLwnM/67outmDWJYr1LYfXq+lhZ0ViyIeeFy+HcoHbYFZAGyIHYFfD
5k4DOaRB/kRtsnHAhF3w3gkj9j3YVdGl+BSoVCfnjtlEKBJgnRWGBNC0MdytZxPr
VgqHU1ifDIGHSF5IF+k3IpDN74ehdWkUjUplT4bTgW/1z+EJHUQdT+votoGJBR2v
LBoCFoDChUdGIaTpTh7/sdkD2zpcLzmZT3ehCjsYob/hv1kRE1I3/xMAo+5hZwOG
S9ibGEk15FwLgJYGwumdWTMaqzpdbvOVy7kkhNSJaxrk1vkMQfzDc76tVsyCw+sx
hKTJ9dysDrgoKtZ1WI7BdFdCwS6kdzFsGycH2HisLhiqV8tjIyn758hBaqgqOTrQ
GboVigWvnTS2yBkAuCJ0TLDy+NaLtuB2+qq23JjHk8FVG9e14e10LCB1Gg9YZv3L
oGP5lMkXGp9Gz2AgoxKanCZHZyChRSvn4PQMhQFBF9IHM3f9GuJTXB2gFmxRArDA
B3u7yJOjOpgXkOZztfzkO4NtQGXySB6+TZYqGkthJnb7Rjbflv3KuWEYNTKjLad0
zIJ8uxNPYKiP75Q2x6jE3fqkXP3FmAef3YImEsYYoFEt/yN6QSTIL/xj17BG6MVK
O4U9OL65OmhdB7E2ebLpV0hPrstN/vmm6rK+toaBjz0LWjXQ2jKV22dzHrOWk8WB
jBMxoAlJCJKRvIaPANhJ9TgrL3Lh3Xa2JWZyajWrd6S4EcX/28v+32NhGHf429jc
u810F0i60mIVfRYGEw3J4dMPIoSJ4/EgGaei4k6UnA7LKeE1O+yvDqcuSvr8IoK+
2IpahlpaRSNyRAg+MBSSBqyDRbtITOGk4Tb4me/9RhEjGn8TGK/7+WtHoIzwDPFF
FZxByFUFqVBy+tI8NWr9enozJmJdYAqiL0tJUPZs4+66RuRTIslO+Gkg5DHTML0m
ZHf7wHHv2FIyPcpycsTLsXOfXmfCMB2sIURzNVgAM1xk/EqzuRipY3c/8La4Mpau
xDhVYQgxpNIY9I9e1yuEzxIFwxjdx+6kgYokpXxItxRUfKPgZ2ScHBBZ3cX/qsik
pOZ9Suybu75IGGq+imkjCSGFL3FGQLYSiNCrmCTuxmKwJd4pgNRfnRVGVGHbry87
YF1CFGDIaMG2GO1Ohk6+R98xdAg97buamwOadJ5jbFosJlqXZdyaD6jd94ySYc2+
399883tlkOnB6LqecQ80+mwowkesve5Q2FbUCnepp42/Z/3fZx0D8oi/hZ8K2dDj
+7a8GWLMQCkqBfCZbLE7i9ZFclPmz8qFVeP61U8Pt7yMQSo29tVq59hHU6u8FA3Q
3kCPBrhoQt06R0Z7xiv3cMxp1Xb+JBS0k4nqYXOwCAX8gfBqoA2QtJrjr1r4rrBi
n5K/lrFeUECb6N8TFcyOVuovd5zdKnbbtRV7hpB13JEO4xGDBxdCwNiWl3hxV3mZ
lsqztjcoyZVGUgCKYDPGBy6UCc60zxppg3VjI2DMocY0At32VACvA09q5RfUzMEJ
25dzDT6gQ4/EJFeUuK36KiFcGu7whtJc6nPqpgpUxoKdrTQuZbZ9qCKIVuzElyV5
06ZweakPpza5/ZihRr7Jfdw18AZA/bieQ+3iAAvtCWaZWebOA/Dw/Zb+SBKUgZd2
EprF2hz/55bWvOqRfbsPNO7VKdADjRKEl9bbkTGZyo1qnZ/AR9xt6r2VhBYHifK9
h2SN4TiNrt3o7QWuBiflzeWJ4LI19eB1pnXnShiw7BjrPT4mX+WWNe5vqr7Kx7TG
5AteizgxFeKxYbhqqy5A1Saz7OZetycAQofq0wMZjE7Tyh8rxZHQ10n6Hh2tKtaK
Q/QvQkaKwiIFdbJMayhnY0XheJFFOj7JFJkEm7bZQA5tRbdjpMxBnSAWAOEBhlNz
7H/yx9Lfh02yxzvNYOArFI6EG0jWLq02OD/u9aGZTxWWiPhhH+LQk5kf90se8MS2
HrzWT2MrD/AgeAZIZYsg6TVOUp6tPEaYw8ACzySNC/C5nddlZUi7hif2bd2oJOgP
mHTOo+PV39r7LQb4JddT+iZlbRXrG8/RMDa3fz+isew14XeEFvHUgKDaMIxh91DT
RebB1KAnbS63NyeNILySB8ncMfhnwfVLpdgZmjjkV9Sx2DvpOjLlx4mrjHjhyEt7
LMRJqxSyerWpjA2/wjEUZCn66N8xuZSyJuGcARP2P5iM+UO11kA8Nda9luXfm/0S
A0YrcsvzI2BonQ1VnFV5T4qdbWdlemojVpSuib1VCgf9CEp2JM+kYkKeXYsWYO/+
QRfV4XbRnm5rFNLyqfFjqFFd6J+HKAP4SEms95Wt1aGFnwDT72JJQP77hYdb0CMk
Z1EjkHvnSp2BLgMQmrfkzfxVX8NTT6I2mqLRE66KEOZm5KCjIJL2r3g+gW9Hf8jv
3DV8nvEGwG18tLZ7NxX5UXihnnoh1SYPkgyKtQBw7nju/4cfd7i9VgpNi24VpBKx
yXo4RXu4SxAavOUbSX/bCmKsX5ohQQvp2XyLuOrYmSxUbLtMdBUb4DboPIX+T2Or
cv9PD3wJEiAjzPmq8Hs0lmhWnOjYQRmXMCNynWG5XOtHEznOYqBGhlaAOT4IEqQJ
udQavabiRXOpyLCWRRxinGot7wFr1IiO+QJ8xwnrkgG04Z7ZOMK+xdummXmi3Aeb
v5X66uDH6NhM4gtrUJ+iIm3qwdm6x1FwTPC96+mWmlLPOTtB7apmUiB/IvsuYPlv
+Yb5t1KoOUWLbGI56CDyfpXysVCluSULNgFEMlFBX2/Ve6M7YKNzSkp3yOUmuXNL
3gkNjVROOHowdGUBz/u5+UPkhtmKyPkgGxw4NMpyK18QYeiVG73EkGzRIUzbUnYp
TyXJsFW6+6N65yS31HPp2L5pC5A+Hos8gBGgalj7x2wqE3KHXyKSNQtzpJKKgMK5
oHtl9lbX08gSXxnWF5oUlMaIthKfJT4u58/oaVjUXlq17aENO36c5gMZtiP89Fy8
owHAaz0xGlSZXFQHXV1caK9hdWiIy5SQDrqLlO4IYcIPgTOmZF5usuqHPk5Zr/7U
KxB+m5zVFFnEU68sTPKFZbjTPbVO58S1M6Bke8ONV8OCRG4mx6w7oCFN/1Cq0trx
2LT0mH1gSwOVAlLXO6XKHPeTugTcz3QkWT5alo3z70iIjHbF3xn63zOK2EFnTQ11
iFifLBeEzZfXwh8XXfTR1NnG8qWFdp9RW3QHXmmYr0m08mp9BlyComy0MyAKUzjP
F8XfgA7Ke/Dik6Un/n6U6gJJt59VtkC61LC1oovHHImx8+XV+J3K8qDQUFEmttYy
Ngld5305OD5NHmb90Wh4FuI/BINy3lUOf54QNKfke6bCTkbJb3IxJJw9r6q/7ZKV
6eWKyL9qEhhlzDci2wMoY7n9TXTV7AsLHENbcQSmLqCfo71WlwI8eMCE5IArcYaK
eqiRyqP1glPLopJelBL3jVNSkzr5DhJ4eLINvg/Ztppo/5ONW/6GhFbzsJj6/Qeu
PW0eSltus0E3ryV5APsrbRx9leuURprfG1gk7bEfSkvqOkDkvKTYnh4x5cHxsUum
uOk6/sa70LU0NRgxwy0ukN981hk3OXvZmOWxgeymx/DFiVSON9lPQLAEPVcaq7HX
Le4JHYR15ces9N4W9TDIF+NlJh6dIbWcyKqoy8P/pbmmXn69U20VQtVzDye8JW4C
dyLgZAMwp3h7DedlULrE5O0T8kU7ZBUjrRlLG7jwKt7paN0V7o4kWdfpoWy8hRdK
gPnc/KuReDC7TYr/l3EL213YswQzmL1k7sz2aMpG3H1Qf0utUZVLgDz/PrEgkCp2
tnD4iTnNXic7n6APMWDFk/gmQJUMnPOihYImHLTnIMkv/oqG63OwZnFBf0aYooZ7
V3+GQnvnkQtwamUcGp0HhU29KbHUSO7Qg7p1Yx1c04W5JX5tmseDgadkGQxRIs9j
gQyXjje8nVxNTLpRur8m9Ng/cw7tHaKd8lmG9kJJRxricNZgU7eSQ6HXqq1cG6y8
DI1cdzbHVpkI8blL9YnB9BfHmn11NG2AR236a3d1lBivXTEai9nKNDjkloiHqyzC
rqz3ZTH9snR5phhfEyHknHKcd2o2PI00uykmoo0Uzvvl3PQxLPQbj9p4w07G0MS9
l2S2uSwmzSHegdboqYJrtwzm/vWUyiV8D5O73KxhI4bQOH0zWwUJ/xJJy3nsHT01
5UtEUQVpEWxFpOUXV2Je0kYXELIaJ/KqP4uW4EJrlaSNhQ0N491cI8ow7v2gNIbj
0XEpD3sip6HtAsMmRIJ7j1ptSZGIU4TGuYUCSonAH97cSeKClaPvCcqVeGVnKL6J
myavPou/FifjbiTjVo75Fst6goVLaY02w7Z0pcz5PecXVKzcb6a9frjeinfmJtHt
9uC9/XqbgGkglgxD6uW4uZxCF4cTJNWwLeVykMAXw4T0Xo0eyoAwa/AZ1cTTn7Yo
ATwIlVc48VHTCZzNFKdJGJykArqPwtedav6WdSph3afpGyuWq/mkh6I4K14kDVwu
w0q3nWhVqfGjXKQ6dSvBzruoIW76G0Z/NSJ0lAQQ4DODOhD3DGLOREI1OZSFX/OX
utBt40HYPR6M+6+0lDaGqgPUx4mi1X4lqxeDFbDVaJlOtQNxOo3Vyq2Zh/pjONNC
hyzmtNeO/S3tAYBU/5idn2wBdxkg3O89YvD+AJdEIN6QThye6kEz94FRTXJD+B1p
EKXzpgNDniuacxVRTUJZjBAPf4t08J/0Bn7vgzhd6J5JeJL5g24JpLvBQCLsi+jE
ZQjHTK+ik2qCJsQT32VdkHRcOOQSnuiN5wq1VSLG8TzQkcQg2XjD4w7Ha7Xf3l6p
r4xmPInpfkqM+TbbNWNgOnCcAxdLewMCiCJeI/0/Cgohre3WKfUV3haNAYTfQzZX
3rQUgFoNbld9irfB8l3aceWCj97a3FurdlrEWccqGmi5xAkN0K326NxRp0nzHzRA
wlKrXrT97+KzGWmzQSBv2WkJRehI7eeb/mAXxIUy2HM1mCZoO7CBvv51poR9/3qh
hZEkUttpo6HzjfesvjKGtt01WpvhgeVavktktMbxy27jSavRx/YkloafFF/6Oofk
SMo175d+G+H0l7awkY2OW+Yrkssil6yn1cyBMBKRws4yjj8oEKUl7za+x4WG2p+g
NGumFE0NkzWc6JYEwNKGd1yB4OO2fq7gbGNTvmwgGKHLvpk/vDP3krd6vZzQd7Eb
KYr9G3ngwIr8o+cVM8s63MjXU0H4d0pa3vM1RedMMm5uk92TXSb+Dn6GI1YMgCiG
Qd7SOdI8TbGWFL8oaQtO1RmsEC4BMtRQTtU32E6U5XhQxlqwpc2Vo36Httn+yCbC
Kvh7GYUXbx83WgFedQE29FGdkf3VMTDkH0nHfi4IUNv4ZCvLCtc06sF5LN4NWVoB
E2un8kYt94HpR+mj0hN4WCHUQd/E98Ohz2dQFnlJAGwr2o2iOqR+ekdqYz/eA0kI
sRQvjZx7LezF4DAw7yvslMsqPvfDfLET0i+UBkwxogvGemc7bg7Jx+2F7PddujCq
7eYEsiPNnkhIcw+A+fvj4IYFeHSSJ8+eKBHcG6oUTAn7ff+VT+K2Z34pFPBtsJoe
+vmE+hJsrnimfgmUHWbau9KU2leXZUE/etAsuvqXj7us9/iY506Pta0QaZTiSl1A
Q9f9ETc3AQP7lc4lvh/YXkVoWvqiKoJVl3ftwlWFDDiv7oZ3GYqeN2sQBsy19un7
hgPUHNDhLO5yE8e7Lb/HLNukujbGyhLdkkaHBJot7qgAHNkqwhMHmIbb8bvzg6OZ
XbK99zcbXpc8kcXMa/RlGDXZnTyCskwx6gfA9teyHWlEC0lV1lJaxNGce4JQChTw
R/f90Q2Nz3+z/mkrywtWDiCBSnrA+xJWJ+CRJk5sKQzZ2fqoMdfEXs9awDRP4elB
1hqhrvqmHE38orz0zINk6ElREhy2FcJcmr/DCEOIV62k37JkHx6FDPj9fkoHnx3S
WkrSKdtWc1oLxbGOlOLH+ytNQiMgJpklgeUXNmrPogG/NGTPTceHuEPUBHMNCNfc
wrarzB7fyWuTBnSCbB3dHykwl6G7Hpqk59gZ11BuQW1EnB6WK4DQgeVRGDd0vyAu
S/4aTcKbi7Sudmsxbe2vjhZIs8Fv+Q4oFgCmWwnbo4JZKwu6OTMv47lDWbGFg0Gr
L1TaCk3i4gZfAGpoUezNS5pljGxWolgcbgoPy+j+QaW8EzUZhcU2h607kXPGYoFq
WchusVN1oHkyt+9LuozIgyu587Mj1MSned5UOkTweJwLovaldZrMrsruS2OaEBen
+O299zosYwCInXTm8Y+ugRBYgsDlL8eXfH1zXBMzw1AAlCJGKYlSwvWNCasB5ERQ
x5U4FGZr7G0nit26T0YjEF6kJHXTA1mEDyxty2einZjqngMUIQvTg7s24TrKn0iv
GrVlygbwFoZoFfiojGFW3dXLuOGcOWBRHP2RUMY5rd0Hn6UHl4RAp8c4dyiV80OC
K9F+sAxchbqnklPQgKhIE40ITOcRSEMk0oPochulLp5g+2uIbvzUNA8WFxj3hBRn
EWvkNnKYnyWElF6/pvave1EGdgE70w9UzMarcNe99LGNigXs2TSLkB5Y2Qe97W0s
LLE5ZgItssIgeX/6g0yE3Ij/3xOICX/6fCJU+YnwcgkGA/sJRogy8+iBSyoq6TRQ
dzc7M8I/lCDKxDwO0geiXT0J9r7sZ0jRjNNjEofKWJbHpH2Pq8M2YIKSDm9DYxd+
A+X+mgaeePjRDmQFUseK4E5Q/0aE/MVdEPJjE22f+zfncQFZlQ+ltom650+Bn7oR
EyNjDprJaFrm9x0myQ8wREq9SYI2Wsur8MrQ0qFDuOmJjO/h0bzi7NMokLJJT9gp
iOfe9Ub1Kd+u5LAgLHXCBAfTumg7C1b0xmTgVNuuTw5HC9ul/6/XemgNyqib+A9v
k6bdvcuY/Ja+d3CyxNMy4DHmdpJkmvq3gbWK4ge9p4hiONd97WQ8RKWzwlJzjUsW
CebF2WV6wlvyhIsO+Z7HMReCwmJjFhoEW4Mbm4+nyc00sBGChRlE5UEO4AbEsjuQ
uKuOCCrJsenBn8SKs0HlZSnj/2o9+07Ww00txC3B0UBp2rEaEiMsza/dwqV5NIcJ
sFJPJ+XaJPgMhGcCwOwEpLvHso/bG3kizGaHZlXElK7jiJXWv3SwiFWkwCzMg669
9TyVSaQpt9NCvKRK6RRe8phFXZ61vKUsly9eAZTCNkR7GbRZTVq8PQ4Ybt4UcUlg
dZvDG8zlZa6hnbiEykPtMlHWtScFKJ1TXSWBs8nlMrWD1FCn69+g23pCIPuH8zVt
uk7sYcHUKPO49skeguVivx7X60+AoSKkD+b0vzdDIJC/1m0l0Zu/qZN9xQvPACJN
OBJ13G0X/KW+BXn0XBIwBSNbhjTZOg9nNkQHhj3P0VbBBBDDYag7TjJR0rnUcmjW
B2rFD3/pSTc50gTGn7viLeOgDn0IEXG5SEqyJuCXdxO4PzAk5ub8E3h0z+jUSxq4
20GflqgOGjAQjo6evoc1cIc70pa7fPxktbdMHcAXYtQyw3ZpwYKRSMc4c5iAmXCR
y2ux3FzBH5patYxPSrtjEoHc/ZQoVPNrsHWty5xJTxjmjvWDfMdSFfmQYgS2HlvB
8dJhLrU4c3FgYasf41FAh4WYd7WvJOAiFm4rCnYk3bNsBGPO64wvnLN6Q+vJRA6X
xrhazzFCG7ZESF+NjrNHwtfSgKOV9hDhM6ChKGhjYgJMQaKWiHg2NTs+Brar3mBc
5wI59A2YNoKs5dxCKqY5k/TC3kHQeEouqjJLciDPHadgB2OeGXo+QiX5nkpd48Ct
J9orqRisKZ/Mv9NpKpZyVM6gsshP+aHtBscn71wTsUM5z1fsPLZXAvV/61kO0KyV
EsJTH8JA1vKnVakRzVOhrfZxtXsOc/AZqnaWVtwsDLYhUwLA8b3vWTVmQ1ZMAbhL
9EfHAuykPKFkzt2RrkSbbHdXBM3ZtKk07gg1dm7L87W44q7sZq3t0P5cJ5Dk7WY6
i6Z2n3KLga27nRwAf83QUGOp50pqOnxjXHU3rXePa8yoU090L8MCIj9k4hqa6LnR
nzAbsQohqEhq7WG1kuVOwrcMeti/jA+xVlrTp7c3TVwCPVtY7IQ8LdrbX79GNjXg
zDZNxtgtgXjFISUlLJblMorHKQMaTlnH3hUXxghbKs1oOTzHAEE2FOvi4iC/2ldp
4OjhvkZrZvujVrlR+4tbhhzw6bue0oh/CV8bVU618YgE2YKh60rg5E8Al3i3SSsT
sefjrtM0ohRWbXq97cGXADvmqxrmHCz2UvTIp190qZhHRAtbfYPqjuFLrsUpjKa6
GlOhEUwEFwVNJaipDT9vSL3Kr2J4vzY6QSC/A0wG7nokxgc9rOB87VabQvg+Crjo
uaFszMXIvp2+XP3sj3KxqnbBuLd8sg2c1k3zQOUW58tpqN2fMDVm04C6SN/UGEDq
ft5y/S254sMMTLyIksD96YlhXuYBy8RYgKHTD3xFtpajldVZjiE9nfnmBq5PIle2
JOToX8nk53Ulr/T1+ZrFt96+gA4YPaN93z3g2LLThQ82KEGcqoL1rRr8MYrt747y
Q/IBrcCAwfI4N/hNj45HMQK3uwdamlqe66IIOz2YoU1IDc2j3DJGmgVUxj4hXKJV
pULYDV3awpRbojGGlIfeUFbQkNlqHTDwIbad/jPhfuQUE5UZLsWOTtyFQOYjMp9p
yHbOUuTrjiZ2HFMXNhVYxFYM5LVjRzSHuUSAtNFZVtZ77rpHPe3yNpM3cicguT0F
k5C+whsUVmrU+C/KD46oivo9C8YEslD3tnSOiIsFHY1u6t0sjqNBMpXA9cXWL8O/
9/MuneWM+CR6wI8I+t4ZIcGDToXBJG9UTFomKnseL3jSBrHK11uBl/mNFjrk2FOD
PDg81zDnTA3QQZl3j6ubmrjikOz33MA7Rmeey91tzPEIbyJkZuwoMDSPqHTeV2dC
91KE5iPVu3c5zfNWWxljdbmuFQODCbwwuuHZUNbxde/U7rXadJIses70orP4GDeE
5V2aYnQlN3gF3XFgET2WEjFEfFoNZVjql95hzAV5Qzl5Y6hmGu1QVqQM3Dd35STj
rdQsa1F58rSXAD4c3GBvanDVk6u1QBP7M4GnNSZE1iV20PH3zlnIGUQqB4E/kiq5
2Yp66wwby9WaxTTuXW6Vh9ZYmpzpSG9MnBaztn83vPrg3GwAq5ZM9bulHBqIXyZI
NmF2Ji6q4W8xgTTAXvnVfsFn0k0Qn8NaOps3ldr5Gig=
`pragma protect end_protected
