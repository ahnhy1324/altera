// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WddGt/BqYqGeHi7jAmphNDQ84uXWqQ09BYYB6a/YLnir1/m6vBqyX9GaUhvjDVen
GLLgdB8QR6vd1nhzctsIsOyrj+GRn5fqGdCaZcJs4sC+cls3NhDtpjaMMAW6yTKB
8HE6S6qHB66ugqxAwyzjZpgq+zYhCI/3iL9t+WZ0mFU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 61344)
g25Y9WaUPlrEJDAc4DlKdISYylAH2OnyTCqHXQuBHgK88FFyU/8W93Q2G4iPeELX
rehJY/smzGv07+cKPxfM6z2FKDWfyu4uKzarpJkk2j4RdrTvF0Sh+8uyLSwZkbsX
9FMwWbK0dBGl/MEwyAkOoEJLQ1prVk/Wf3yG20E7fFvqc9z9ptzRVsIlLUOS5OvB
UGV55ELdVWToX+HCpZfhsh9QyFPezLx4b6a8s99oneSsL90DPj9TNVEgZ6i0UXbL
ctCMYQlL1sKZbdmeKUDQyt5KKUuy30cfFEA743Qcjh4HClCId27wmh7zv9Z3IGFC
XrNewNFEkZ3DTA01dqf3X86ewUq8ksWFpjCpE78C+Y/NmqPC8U63LjkS2a6q4+rM
wmwRRdUuNbd4YQf9n/Q/7fL4BL06whboF18rH4j7uh6HghpTU3BlyGWkl7vnZzjE
zTpJHZ/vXCb3aTFuvkZMsiwItYf4AeixQKXlWEppz6EKLrEZW2YoZJ3h3xtI7i05
gS+XgknppJG8mWmD+9/xNi4X0Ie6XAgjiXiXImVsyRmEcPQB7H83+gQxagT1YCRA
3dAU5kJo2RapVbUtwpH8XrlYO9PC5RNK2gQpCsInfTndNCcac3vSCLACwiZahZWr
hl+LQAd+rNHQRvK8kxv+v2EAKTBT8IvAUMPC7uCsSSOHtxE+Q4sJ9gjG0ispfnQM
MhiPkD2r0fhoWVjonT8mxA9q7+e5W/Llt/PuoK0unvKfpdiYgMe2k8REqH4bf89X
NYK7yowWQVRQgw1ltj2dSZvJrsKUAJw57HAy4jq882akkfST9BiZeFKp/lQWhFzx
GftVmrsXsj5W1Up8IgAHZ7yYhQKFJmNiuhs7/aymbL/epqb3Pl8ljx22B2teQ4rH
EVV+WB9p0Ta7YHEd9mKUapo6sutsktojjMo400nSDbOJukujwl3znp473CUnfzgi
YCywyeqUBl6UWTwpjBqbEnODsLVNOgHQvfIslwJODpWlgftURUCJOrnK0TyRpSUS
0YFbAkaMVN7Pn//+FGMOjwnYMPYvEDb5wexh/bmHuss6Mm0nfjn9SFAsngfvcupD
3DLLtEtfQOM3HwJE69pbe3OHLSwCCmEsTLSIDo0fKuh7GiBp2ovtORZILzJr5I6L
fhfJSyqP6/tp/U0al0z0lMPzFldTryfg8E04gAoF9wOTpxs6UUfp6RWbTL8KIM8r
jgIgqgUESxT1NHIjAJjMHDm+oJQGvi/FNh0DxwI040dn2EAkfLG2Z46Cv535AZ0V
Dcj0bsRpCb5WaYauJ2+GesiWyalAvmjyAK7FaYvvfeSPQultYnxXKsq/8VlhkAGG
mQNFlii29i+tLpZI/lIWcMke3nmXpECQk0cOp5MbRCVUwmNIfStAUTQqnIe8ZviP
E65RH2qcPZKzX8fV1xT3YwakcPBxD/fbZz9YXirzJUGcjow0crpWzXqPVWZBGy89
iYYhPWvONOxEOXE6ZLHeMNOOKMAppERj13mnoxw20NxxIUGl6tC+v2DvsWOKVmZQ
ThIWFR9rHFR+jsmRJE1sDUxEuw9nPoxnCP+yxbNjdVy5MpOhqBcKqB3ZWE+Er5qB
bNYnMPnIFThE8Cl18ox/R+rw8f+NgAWWliOPKG0vEaolYZ3xtZLp+P26KU1VGKZL
XB3QsgYPl71JIOWuwUbfnMRDyfU2j19YEhPC2P/Hw2Kh6PVORhV8s25sEZRwWvZi
bp+330BJnx+0x9LS+/3cFrAC4Z0TYgp9NOwRfBnmz0v4blu8XXVKDFFahbh5wJzU
4hr08G0NqTLNoRteRUR8W0JF29xfYsd4/Vkn0MVRT/NA2BDCo8J1RtXquIbvv/kb
/z7MIEyClhxE9KfeZTjzSn+6QxlKUjSmmb0shQpmE3H0Gvlg5qzNUpMF3KRQbodc
JoV9g16OlBvJtDB7DIeo/ptFEin8sigx1WllCMYOLR+SmCpGzt6jVhPZaA4qVZ/v
NRhoKsHV7pwEoml22PiBQ91V+1f2oiAybVI51//eO1znQE0RFb9dN6mRsOiba73d
u0GItv1lVCiKD6qi4cJRxws2FIiQW6dokQzce1j5uRnCO2HP8cGjjGwKuA5b9hR/
v9FAUg9W1u3luJc4Gll2Yc1sVrya8qi5StN4e/FvUm8g6ikOIff10xPPVBfrLzmw
1jRAIqk7oDvXSx5J8JySakpFYdYqpXT5+F64irbYdFp6mg2BfP5ck5ByUX1sbkNC
KYzLCQ4JCROTC6f+cjQNJHhmHPh8t8K+0ytLVBGrD1PATByxGWdXwq2wTuUjXcUb
qIa7qqRigpummYhJDZwsh7kN9zmCdYME5YLcw/i2VGme68d0RrGFDhvctfjye/8N
mMpf7nWJTDez2Qlf4aa+MJaiju9Y5jfKtj0thUgxV0pNJr98xlP4aFkhBq/UggCS
2ZAQ50pvZalDj4GWVsOaksyISW7lTtlTxHpPPUOjJBY2mwqMByNcOLNzw0TivVvG
q3URXgmDI0bznkHuFA8Y/y204Fj7L3ZYopVhKUn+Rk6IvxBYQP4CM4cXiNupOVvI
qTjIKQazKPMv3Hk1NFTASapOtubCvjXRU5cvyVmAnB8kYQOyKZSk2tII6yUsisoT
H3eJ2BesAZ65Fv64R4pOGxAegMTg4BXjj53V/3NDBWzsN5ml2cyllqT49UcIUG64
J5OhBClMWENiQMcMJnoYmdZdq4yOFB7ygRF1BxBqGckkMErA3OUzp27K22MVdBdw
uqzqKfu+n1XeVBWKKLZz9DRAwapHb4aCMsl4pBNzuPQuS4Cuj3U1JDAF3W0LFC6T
1Jylly2gzr4wUFcFl/uDk8qOdt00y3vw4MAcbxMOOgx4FtP4Pz9xRDJEfCM+DlCn
ylV8TGxuoeN8PMpsegxPHUP6WM+aroKbMyM3wwyQFHasTuzZyeLvECdnzErLamni
unDvD6cO+MRJXYZ7RA2RINY5eWG+MTSvu+hpM5rL76vT6nPSJ3AxSLWzoyDNDbiX
9Vt9OSnfmHFm2tOkIeey8upTsNN91NgR4lNUT1o01fyzQHYic5LckNEUTqhJClAj
yD8xdqzutWOe+lUsSGkTFBjuwr5mOYUrAAf+YxgLkhUyV/+u1r0nSkVA8XGmh+er
Jk7WH+3DCHQlBlaumiqZ2b2K0O8yZBKchznj9yK4ZsowwalnlOiy7fYFzIJuP3HS
AdP9tyoxWu1K6LimMjeypFHaQmZIfAwdSK+0t1R462g8qfi3mbY94W1d8z727GSa
AMsFaLIieLXSIrcsqCDG9PTfEuHUbwxURAMrwkCdzKS1NoMIsJM3fTO3GGZ+5DOO
5pgbDF07+tiK55GrRfXzOyDnat87YMJ4vFCrrjnjlXUbzPi7NMWoo/C/NjnHLC6b
+uMrDe+5zPnNAxr+Fvho1ysikLRLDdBLTkBBAKfq5I8L8q7Mwnn+yvWktkho6ONk
N3EOb5ONboWSLoELwhymCjrl0J0S29rTAHtgv3JBKYCiU2h9vrLAVgYUdyV8OT/Z
CZVMQaJVRLRoRzSX457jwWdfv5gsvyQvNvCts1dkIt+0zvDlvTd827DpHIyffB/z
iOprdT0cQyDDvP8Ajt5O6oBRMFenQ4qnxXPa0/XmQPsx9UvivJXPvWaxEPoovDTZ
SOkAnpM9r9wT/TQqPUzqzJms1Rouf+rFEV7qQXO27VxmdgnAtibkfocDz6anI23w
1bi3vNMmcDMesAq12e4hRC08E935ir5102cJPefTlyzIM8Q1iunw82e3K15T1LA9
wLbgEAHHw9QwkZckgOvsEym5gOfWeep7s56fJrVuQZyCoDfV1V/WKecNthTNfdnE
x29Ctg/TyCiEQwHI0mFx3abENITlHSYhOJRTuohfCH/SEDIQBj+C+o32G+9nIQbs
20NHd/CYau0H+S6UDrL1YPkBPQS+WtaNf4CaveRzRlS58vNRl5ftfYYOlJs5azNs
yYkPyVrKd6awgI5gnjVAO31QcCtXFLlijZTmiwgk/DVBXRB6m22YSwn7tTetGHlS
SRALceiUOfQKbutEwjcu7qyOStuaR124Q7r6g6MAD0Dpt6hsHcuVcK/YcL6Tm9VP
F1EXhWe0qGPtJl9Z9+OcuSbCWYbF0XRstDawkZd2TpzJe9MRLXiwoAF5ZHJCIN8U
xdrvbz1YcXTOK1/d5fpQ3VWIrFy20vXvcFYjVVIqSY4s0rcKlpBCxYntIK8tmoT7
yPi/MScony+oDBNJJTByJ4yqBZyPhuRInBveKBcSVuwjCibhlRCYcGtmQIBncE6k
xPMs0LF3elp9YYYDI6sIMok5mY+xHC8y4f+NeemPYcnSXIVnehX3EfNKfIyogMay
7DT6HwGHLbs+gJMwbhbmgp2ph4dFDGJAUHCW87TDUXR2CbGurXGRA3MvK2mtAETZ
f2ttGNW5JgOctPFcTLukGC2Eu2f+Te4ao/qBVStmkm6p41f0FQA3so0M07GHlVVQ
+BDAToDIgyC9nDss4B9cTO27I7keZb0zUD099VAcSZUwN4b2nNRDL4N9gqS8wE/d
1wBdfdLvORMT/ecaf8pPeSMnr3aDkNLwPLjh0WZupM2QeZe277K6Ol/iA7Jq3xFR
Ic5JTuGSFgEfZtVXN/PfzQq6HFbQlMFNi+0ZhukLvzvHOL0SOgmC5vHxH73bcC9e
EngN2xo1+KGGJ3uW9m1EiVw4oQXjXrle24uXC/cYNzAFMaA5HL++cTwF6ilk4jTC
WoAfLefUHc4a4dl0gmguQwHx2u7yOklIrCy/SOpwY3TnCaq/Hc3z/ftlP4RgJyNI
hm9/wJOVjgyYeXRh1bMC+R5Qi5j/6r7EzgrIgUQh2yYPphNmt36FabQ8WFaLvnTR
gFwLLaXCZxbOZtrDotkI3WnZ48GIZliosKagheJpiiFAMN3jqJrE86F1ODawid8m
bAWAyOv4bQvCBtf/zRYkhjXdrP6yBlsbh2Ii/sYpu7TXB4ODiebf4IU8LwUKX7vQ
dzdFaArUxvGtD+3FuE9814Xt0lYfbLjlOLPUBQMYPPbNvsxk5/wmMe+9hpnH98fY
9kCP/SshNgT0tlz+/7xCmywhS2D4VKmOsPfFUZuh+0tSm0Pm2TaD8kbpROqks97I
Gioe3kNWHgdzDDdvNcdSj3OvV67MottHUklqpkBrTx1Mts0105/r/G6occf2Lbun
Z13uPVbFHtvSRRmpqhsLrJjJOmIBpJ7o8hp2WOYS/MTYBvjztpWxGBJvH6e+bly3
zNc16PsRW72Py0QageEe3sO6YK8xm0w+WPm2YO7QwLarBA/MCn6znbKXlnCripME
7e0LqoF6fj8kMiEDjQ/tJNPoZ/MaENLV2ZmihutBHrIte2YYHDhOHIyxUCIveaog
4pw1c673BkUdjzOeibWrJ5VqN/kGw9iLH/MnAJfejM14mJUIWYfsgWDywVQ30PLF
6pd1B/7KWtCr+WK5O+DptQENzexFDwOcNYcAqU2oN9fjHBGJReX08BND+LpxKM6i
vHlazBnMPBIhpKjQ4fjQZsSRdGsfMqJIvAydSKt88V39rxdYRCHIK9ra1vYU/KmN
tXlbUpB/8BJnrQ0DHMM9oYhgp5YM5FIAZILdtJS52zFM+DIebobtM3qymclsyuKz
KMTziKd0afI/PliZfhFMPTY7vRz3oIsSQaagNW3PYkPEbkx6q6CDiNu+o7Jx9Uw4
ONLfuexnmM4l7AdVw22LUo5rRNQCVGHPcXPGsA6U2TXWoMD94xEEWBpogHE9yg7P
Rg3FW3BXsNBm+lNd7jcWJ7W3FlqUzQwFG36vczoBdIK3aEcfEEqCBiDwHSs5FsPL
dzTtmDcWTaRfMy0gnLnWdSAKy4V1GibTvXZ5q7HKbDv5f76ztAJ2m4vMPPQwCqTg
zGlrbyIJIf44BrolxPS0rgVf6f7HjefV4oinSpa7lR+Ze2K+ku8oX/pnwmOpCai6
e6BgU6AyBMsdxI5ojGUiLFY7//VA+JqzgTOSB3sV3wHhaABN4qy1Fked+fjcLXUN
xeDKDlnp+LHZSoCUdHY5TIiHaGaTnXaJf4/w443HN01PGF4XlwG6IP5q4eXnCYI0
YE9qLmWhRe9TrOkA6tdBS1lErlfdJ8JqLfV7R38Yb1fD3Kh96B4T5Bd2W69yRxoj
lUmARh+AGYuFvSaLKYAdBc80har8goCeQmxgnNLWP0BZE9ZiJImYnlemLQgem4BH
TzZK/X2qLIXurkBRibkvlkK6wAPTIzVCvYgUYPn5ZQwQma36stI4am8kB2BmQemg
ZujAPCWboyKvAursHQ9YxA0trwXjwzRbDnYFGYnP+0AzXT8mhhQBCOTfkjMj1tYE
JJTemJSacIrwTKPeWS06O0UWwp5sj/eaiWn3KUVwUDwmdSq4RFmobl+bQYq13U2c
mRSNrijZjC4EdR7kIES9ErIQNPcVwODibUKidUox4l5o79YpbjWQ4WE6ZTc6yo7U
a8D50xbnuEMWM9nIBJGC4NablnQH0CDVfC5deGEcs+SH2kKL8tOldm5F3/d5CR1B
/xP9PBkSJ3o4Usmqq9WceoisMYFnLm8IVN7a+I/yGnZH2KIWSb1QA8+vVcxI5U4w
tj6/xKNI8WiEiQzESkwUTkveOvApYEamiDioHuJKzFwoHwDdfooaeNqH0I+0N1uV
8uhsgMM31VqGCjpweqwme9sNqOKLE84yaDj5aimlDe14IWTcmiUPrvmKED2xPBL6
M4j/M1BvaLgpeb/KZuU8rcNUpWvaJ0aOLBXy0x9Y/SHDAxiHQ4RO9jqhKk42azi7
sPfpNZeYU+6QeDF5x8zkOMlUU8GsSatJil3ohf0mng+ucBpis3qB2amkdTDKBQz7
t6qvo3tAbg/7VDWMsNVWP/7HGlUUCRrHBzCwRQ1dkzxuv6d/fB4iK7uL03l1aGH1
3oG0giYPvoWK5/zDLufFlC8EIK9DVRBCib0noQClxEmXbFGf6A3oTxqqSzMZT0eS
xKCFwW12gVHG1qDbgL1J4Rf108V+LOaBCz2V6hQV+eAs+lVgrEn67GxzDSDGtS1O
ERCeSX6TFdfiOWQjAm/faep4ZMysmuNFQA8pJ9bikKGABhb2evTC4H18xn8i8GNN
2TGJnKGoCP0inqbT8/e3Cj4qf68mZllM3+e/gNL81Lqidj3vsviZNdPCCs7m37L3
8Ar9S3I5s4OFXVANiQ/7aR0XfNkUleLthnhXWJ/uag038SoIacnb0+dZDAITiiQC
uCTgVy00WTf0RVam2aHqHqpm3GJon724UTZWRHrT3pXfFUHoHlcTn51bDuycMSRi
1pgh4mPrKpXEqyUaQQwxz1m2iYsp9nmTw0gNUIy0wFaEaLSN0gxh6127ZZhuUqbs
FO8yD/ULLea9fSjfSVjtqS7toD8yxkxOq4qcv5/aXTZ1QuYGl8GigH9MHQMSB7ZL
2hX6G0clm8s5sg8h/Olj0VgLUTLA0qgrDGEldSvNPzIeSFpWLG/2bnin50Z4WbHt
VJ+w5ZZh9yOE7uF+F0+5RGOLxXEx1StT8786YQFcwcH9d0FynvbQo/n78pXdsQ08
NUxQMDT7oUHpEukyXVed3qdB7DGvXjRihDVPXCpxLlKummG/iPjIF7c9pcqQHvUK
853ZKuUsWKwme5ttv0gyJeXaWdzUVUvcs4qk+gOHeOHcYfA0At/rVkdAxCwwpMi8
H/Cznw4wCQBPgXQHj/RI6qnspYSzr0r5GkiDznDddUi0y8CX4JSY4ACAT9jR/lHn
xz8z2uswzbt9M7eI8kX1VHpI0GNSSdJ2K2ndl3/xLHLhzWgAaUe+mK1VqkkeP0wA
OV8shlrtwowe6Ns5XOGNZd8ChRc/lfwod6XX75HPR/Y3AJqm/9qHEBB0Z83wzF79
RQh3QVAcNnPmmL1XIs7QfjynO6P7Ku9vpHqal/3SC44q8TwY4/RNzi8sm2p3D7Ba
8MEeNs9DYxIX1itQ57yfI6YBLCb1wPl+JYJ8crTkyW1P4Wryi42D1QYZJDvfOhgb
c2ZoXRoEnsZgQA5Pf3ogtolwYzto1TLo2TgsJFVth2z0iDpUcJDfFIZadm+Wk2s8
1W4anc1CpBB2UOGZ+6UZ/ww0XxaW6p8lb5Z8OOYkoINTlX9ZCiniH0l1ebb/XQps
ni0/YXi42vAYZbQRM7V0yBNybCjsXsEY69IA0u3asXYO646q1vQeRHpmUPCrqc3y
IcY2jTySxhqM68t5zciXeWX88k/APhKWYLOV8RNYlf4CqNI8HDFYEkRIcaoKSsQS
HxlbV7UDcRFyftEtzlOwhFKYHByG2SyDqz5pTnKWAMTaIO+V5qi90tAqxN+aLVTH
a8/mABPpdjjMiFY14IEqMwfqn8vmy2jk5GK6g3koQsBWfNVp9PrjG9biS8qbfVnI
U4/y9ZSzD6XVaIJztxcT1KZiDDFSmoSiTss1a4K2Bst53J2iZ0+Hbs1LyWaukDn6
mv1jgcQ9CCXCeubKzMEZS5SMnAHufNSaN+4YUKjfR4hc/UWOKDBIOooh4s2BLVPs
W51Kbwy9KNWpet42TKqDDtt4A5V5OUuke9rhO6lN8S1bW1RsXR8sMHFbaoPkr7Yz
EmgPUM/OsaZ3EkV3JNQoowkZzCx2Q6TBy2dVqVqYIS6mgziqNcQwZ++r4Cq9FoT6
IT7uFnpafkhMhBtkqJA0rDrJMzlV0tHZ0los8xaunZeHrF+6X2Eo8O2wS9Ny/2+Y
QC9dG89jyi/BdsltTTr8YWWT9k2A6UQ8YMzcf/8b+gjNwhSxyz1Tg7T7AfUiN4AD
P0+t5OS/2ezSSS+QPc6mJztyR5nVKics44xs1jC2MBBDAWy8KsjIykDux7odkhBL
iAu9Ye5B8oBWEgNzYjyFZrohC2e5wmIcQnS/brGK4jcqMpzRCsFsxAK+8yJhia5f
+2CYqRl/aSmjmtRqHh1wGImNc8UWt/IFhqE46QwatJK0qiGqgm506oSWQH0XcRTd
e5JTmxggGzNMggyfJNPDIvy04P/QEzzQmg/JkA6/O3I+Y59SLpYPYb2/7bc62j56
YfOhPPyBTe1WR5+TaB9Kba6Jw11peEjCX9pzdj+7Yh59hwcivJAXWk8GJcVSZSSx
PaeaTFY0W7KGlivXHUfdmMknXPJGjqTXO+wyUaEDcu5ngCJNCrxeEZX1tVST5m31
HoYjIjGbO6blqdfgTLi/2BLN1DH9J7Nl3L1adBh6CU9ZakPaw1DOd5LHo3GM3mC2
MJV2JJ0JBI9LHLQfRoxDraoZT6xB1mwSqDCmg8OuKCOl3bxi8HBJBPrysExvwOMC
wisNEbaNBYgHEij2EPOQRh2gSNJ4pTOtRLnY5VSszG2VUYqk+vbGK1fkwX37qSUQ
AX5/WLe1gfK3L5Ynv5cySbIW7ww2ISitZjPjr+q76xiJf3bhh0WeBbgDb1naBl0K
hQ/W6s9minka09jeBrenXI46MgcMXBloz4Lp9PA87lQTxTN+a6LXbb3t+TE8oD5o
TCBx7IY29c+Ni6O5glZq/fZ1xugyrBpVs07tXQzvu+sAyhLE0qF2tFiiCk7Nd711
8TRcqODP5JQwfEJc7IdtpXwv49nO5byE/90xQxwahkq+mFG9He6mUBDZmZqSe8TP
EpkhQeQYS/U53m1uS5nZxCE8za+C5zGoX+q4cxbJpeuJ5Yupg5grNUI5RqZBmUZv
uCpSUU7uIePkeL8WxYGEs6c8nS326N85+Qo7ndYvHpWl1BoGr+a4l4zjGrfLt68u
tDR3DPyB5Hx9bEwl0Irp3S0p4QSFrnqC056MFEfGDo9Tvo8RbWodPSHnePIO1mLV
/Ky+neFqloBbKRzEP/TwBHpDoEyOUvwnoepNlMfoj1Eh+t9vPi8ComGf5WJkzLx/
vYyAdPJvtO+Timl7jnDsKK2BDINz+UVWyGA+c4M9oJZV1OU/6WMWnU5G86BjD8aC
DyJqkn2nGpwHGOQO5MD8S13i04eES5br3tj2uAfSfXabNQVFt9MzhKg/9w5pSEZO
SV9/ALTsVpFIqm7o7ouZJjR2z9MVDrjYI3aUt9hJ8KwxOkzduRlnEJu6Wa6t6Xd2
af2kFpfJHYiXvSeyzRKjKDuhh8VmIaq60N+zgHl/mBTk4m2bByGG8j6imU68Z2wB
/j8Dr56MZAxGG550NBG4myO5+jj8bEHH1eXSdnxzEzKnZ7DzGwtuXyDa/iw4nUbw
RDfH39RtVVLYMbo9GEmCotGzrXrCT4P77x0OJzM4noOcAjjCbDznNP+8XsXo9lMA
mH7BXorJGE6h75kyrQDiio0sE2DorkUO76HSrC9VRTz9LhXLYKwQ+ceAioEwVK/D
f+nWVaOdfMvMleNEfX27eCP0kkEVqs4pKQ6ZTQ3zybwEGQWlBIY+UCSb3GMGp0fc
oyJS5BMeMPrVoP3AZXHus/wQ576hwq5itzjJm6ktVioOaj1CSblrxNg0+idmfZyo
HfGG8VhtB1LgdOeqUBpdQAT6n2phxpiUBtKByCR7FlycUKXQUzpfpTNJnOkcXM7y
i7RhIwjtEqegLOhvpEdUI2pIzcD/cxZRTFCOJHjSySFatTg+iAR0iOv6j6x5fe+7
a5Ig37pZOEATAKZG7d9CINqVYbQFfHDaysjlW2mGU64QNyxBhHzy8BLMOMWlvSfn
XxcyvLHYdgYfOyyRNIEqncGwmR1lZb2BeG92yopBeEXuMgfU5uLCHpNOeVFWWLHN
gwYuOmBn7PWX4ZP8a3HtDBD7Z303oFg5OtK0yvEZobBwrxPjKc1aJgi8+NZDIVJc
5zxapQegbA03v+3F6kJeQVJy6xpUmG4h4vuBaH5NmuUqzlPG8cYDJAjjCUG64GLn
DCoo9xZ9mCNEB7X+c5NQPGzBns6hLjdKT0pSUxFuTVsOkXqFHfjZfAig8hnGXFrQ
YfpF4vZa25gqKaL2UPfEX+Lnf6h46YeYJCHnr3WSyPh+hUbZIoSjC6veaAa71DAn
3N21+bRuRbZvl4CZ5jIJ1SxUatOUYTSYg78AFxUgUfr+kWPaSUmmBwdWAIgc9YIT
DMFSceMfqc7Jv61+q3ZSgggq1DHuvtsll9GCKS8d4v+hY6zVKEvyY29MVQDmuarb
eotyEM5oUwmLXZkSt8HtkARfv0RBaIIcn0DtWhPLMJrFKBy//1ZpRObPUuTu8yow
OcMbn8qmpp4B9UGQWuJpDg3njklxlHoUKPfs4+Qa+pzVLLEryvB1JaJ3gm71xdKA
E9hmSseor8UYJKc2ufvgh61mBswKG0q3m2HVfPSNJzSvJw083uAzOlaXqOPaNfvb
CYTgVw5kuPbTvLRgs4izNNH5JZA5C6k4yjIrEcNC3Itzith8uK8Rp9YFKny0QqQb
+/+jWWh1ewPIBcmfrqrQCvUDZP00gfi8wA4PLHxELR17w2BDdY21g9haVXRivuDQ
RudLQkMDrUWO14G26JrNgf0M5oi4UpEY7fM3czbr0F2fQXtm21C3Lvee1if5qD1K
VB/lhErbX8KzF0POO8WwKtL1MdoisZrYJBPZ0mg9C1tY/ygbEpSuufwXMxirZ67o
cn4EvVC4731JMdPscP1pgMc6/jDsMkIbCgIPv9MvaBf8s5kRIACZ4H0EahLKQOEW
bFea9tB+5iO94SRx6ZWr3SS8iEfBuPw7v9DtMqI4KRA5QzpPmgp8yaKSxlX4aTf6
+fDTn8pyxqqhbtHYYw6u7jwe4e9W7Mr7n/fhZPOhpc+m//r4vHBln4plT9H/FrKp
FnJ+0CO2mqYVAX1pTPHnUKGu6A9ytzykdLILUODjDdOAxKZPf7WSXjRzISBUJIb7
GPlVRODHYIeUsJp3K8nC+lhiNLhzzhdJz9pszkQtExuBvltgyKyHbmwJl0fo6Zgn
JGDsP9eAX7rDgx1LNASAMc3b0t5FaNc9TrmZUMxHtcWBYJFGhqVnBuB/CTwbwYgr
0BK3WhM0Yi8hvWjMHZo8jRU7YsCHu0KCZcZWW/FiqocQe3sqCz4EWTtas4IqTfHV
mXA/W8p/3XcFGUaUgqL8wFllHdxbZGtuLEDfesamPQ8uC0/nJYlrX/NflMTNIzsD
ixB62VsjFIhYHxVB8mJ0Pz15HpHrjKMFXmWXkStlI0/7fkV/vdrLNF9mBwkjRGOR
JMdxwDH/FCbugs387F380dxBEWg/rcBw01TpiIeRJlapUWQFMY5g/3qNJgDpfLNP
DXMMX0zAK0VWPaFwabRSSdwR1l7MAdCSvYKdtgwEbmjxwlzyYap8W5Z/CtYSWzXF
cPwHNcmFoCIZb1xu+KNgI6JJtGONCHUCI+FFAA33UtZQoME2TUe5nUyacPRRGJ+P
K+vHjsYN6qmWxPIE+bpiB5qRZmff2w79a36sj+7vZmFbsno4XG3+AvPMVNOktdyv
PVEb03Oq3A8eMW1E4+Hz8zfFEGas7VvW4zZ3ZeLpZWCO+zxJseEK79jg/QTKKprI
wcA7PBcms3W71qNaO7wjWkT05c+yriAA61coIaOB51a/TQMXJ94sUS87wiUX9OL/
+qWkuTorF5SqT5zvHONwAQb92yp1qnV9KCYtC8QPcEX8nvbD3dQMm1JZNT6M5M5i
PO3qV/sPhhi7maVqS8fhAils1jKP7+r/WVwM9DODS2oiCvXOWUofL7KmLdg4FExb
4VnZns3I1kPRVsUFiJ43sIHw+LfYh9G3L7/S3DI2Cm64ufBWPko4PXcX6T4WM2GZ
Cno6T6Uq0aLSUPAVdwZgnX10nkSFNlR3Ee1HoUIGfMhsV/FEcADPC4YU7Znqhliq
zsZZYxUTdBDibAQHzDLs8Fb4wd+lIhGhRoyQJWFSIlpX4mzGrjwAcDaLW92c58ra
YwqlOghR2bse+qDtAQ0BpQxECVRExkLJQkTcoYtoBYtEOwN3BUJ879FgzjI0fmeg
apkQAU9674SGQygdzbc9V02kz/DPHOXkFyMQOlRrl+84/O+FtqxWgVX3G0szNA/d
RLskvKvnnT5JLwHH9A5iXzvfUOB1i3E542191HVX17rAKqx5iq047a+XRG5KzUDo
KocGBf/ruJ4s3olwkMn0DzSCZ0jb8ovZO3xbDi4HUxURD1KsuLx7zADu7DZTuwAU
tL2xg7YYLvCtM+IShb9OOMJsK6udw1Qcod8FwBTCTAho41NCMWgiSjS2g1Cby1d8
vpoNPd6wzBb+ASZMqWWXMjnpYS52VTK61mZvCIVDiaAxfbOt8efWT/xQGxW5BovZ
zjCP+0zGAhHlEUp2uQWvypobrC0whzAfj7Jw0p3AQgrMXo/MKxDdVZXNLJL1eTY2
ZrEbN2SV7vC2AAjC3NL5LnsZ8FH+88DxLX/1LyqmVVBThVnE2D1b46ao1T0UEmwo
fu1o2r+cotK3WL896HYnrIK59iplEF46CkvoodjqIfWcOasjf7q9HoUPET1ZAv1E
F9ZzN/g+0Tv1xkpa30STf7KINNcFUcrs6RI6wPkDifFuwV038YknnuWyLA29yOYy
8N5vphzklW6IhG2AiZ7qk4EsH7aF05CWitcNBIcwGr7MvWMz1TzyDN1Iucq49jYB
8mu21mIEI0wM3D6AFyiAJ7snVvPdh5Xuk9X9yh9FyNWYfSgDXfXwrAUfvhDzTYKD
dxWofryXbhXARb3jOR3rvwj4Z1V1UvqIMGH6w6r8ir3liE3/m9wnOb9tTyyD7fe7
FqIagd3kLWGf9+eg33cZl8MnZnVz/XF//jkSsyM6G9vTJgjBbluwjvQaWPCDmtY+
ely4tvhHJNrfxsORtW1fP69rA9uK3ohdR1a4c59eT9hYks6MjlLxM29TjqSTJtx8
Ygl0hflfViaQEXRGg8vVleqYzKoUsnovlb7qINSVVOHFBEN1ZPF/dR5vK/V7cH9M
X/Lyt1EpN5s6+Y5cUHcfOrnjYtYBURSknCrOu9pG6i4Cfw5gB8GIpirJf02wvs7P
HnfPZo5Rjc7qvklWBhFm8lxaxHPWHROrtbujCbBbqiuvvtUnVQFu9SUEcGcI72JB
Ofi9gPl28CKhy3e5IgSzHZ4wT/euJXs/uxyjxE2Cfn0wS+1MynF2qaWrnG0ViLVG
rIKJbBNLW6c2Qd8DzqCvKT//ljGMJhBSnBBS4R1p9872kjLuX3Ar5bxAFs5aDwtH
NzhicI/g7doO6Q1DDQ0+sQp8tjBb3hU+0iccJYso2Zh5byyUcUqt0UIk2EsOgSHw
nV6ukU3oUT7TGxH/0vaoELc0PlX8jFFVVyb3SFUJJTo4OiWAunLcr/TGv5m1Wlbv
D3JrUzVAzeJlSfnnHvPj8GIKfmNPyDUoA67FHHzrdYSCC19+SDjBf1e67NNNYTLO
jT2gOinlYw1I7/uLlSobnmFRJp1+8dqUVKQ+eRpcgru6tP3pCgJ+uE4mfOR0OxTi
7y117fGmU/3xf4qmL3wYFN6VY9US/c6PvXOCtplSu8+RcYjOob/eMoshaEZ2UV1G
cNKvNZ96clli7Zo9eMWs+8nhVsZTdg70tJfNlzUH7OdUHW/WkCzQjRDevggDkww5
iUP6rnB88F/MkVXklQNd7TeaafM8Yo9EJeSAd+8EMx8O/u986A2rvakHVKI7kaDm
emjbyF3ScO7EJlMFuUUhD4vmjrNXT1fPRlx6pmnwWgfUuduM//7caSvpM8Y5PnP2
KaMiQ6Vun78SUAUJVOtHLGQV6vNOA7Uee3IAKHmVcoM+k7Y5pn8ZrWndI1UkAAr6
GStv09/sxWqIxuzU7LifkxtWEmZYeprOYZsdgVOOlr0FAGn9TKV57dB083EqJXPl
TxkHqD0IWJH4cEOhM8fNTspW0uQlmKA3CNkrqYTB/TNmOM4vPUo1czXiKmuxGrNx
45+G1aY1YLwTH//4i4CLnVWBZZ8WXWykBoJLczGcVOCAwRXRqkjDdDZOkz6lMY8o
htsGzv9XIvUxmLUzzdsoMjMV/KXNSxxKDBDXnsI8OQq4+BUqhrRleyUAoxOg3+v4
9drXZIxCQ5En9u4t8C+p8jN/h+9+JjjiA5kBBTdtgfA6nfg4h9Qw6Y2QBf4t5AoK
PSfyBNQMgohc2qGpJlImZcgPT/NnzeE8CbsLiV4H09T8t4xgBTurqavxy17iYLWw
q7izr1HLlZ0Oh+PXLpqKzbQoqPYNQc72SagjK4WpMIM1FpgxrAovZaRavpH5LgYB
0UFufFZhAfygWgwI/5pLAjwyuMQLvh92KjOgZ/KkkZkYbT9uKSGcivMxOGRzI/Jb
WxPimjFc30gTxJhs/C9DUrvFg4nfCSUrvtOummpjZU5obKmz4nR17FOafWMx1g4n
h9kN+f0GJhkN08w5pqCmWps26J7wW9hFPG0D7vcTb/p31Km/pZKt3s72/ZS091Xq
RK1w+MqjcMSiNvOgnE26D/elt4XFRqrh+na9Ghva7o8GWBKt2IGLBCaHoaT2uqB7
v6f8/6VarxiGx6jD/Aqbyx8bmyxSOwoRDfuarfGzzAe7u7G7RqQkfGYJPCh6/bl5
GB5rJMZTnkHqQq+ENEgtzBGjvI23ajV92ioVaGzZsyM7C92TlT6cT9lNgUFajr03
PDu+09IQ9tSx0uHthSXagq/wARhm6iJDOvm/KV4DyL7U6qXgS8W9/lKthPClVf13
HzkIknDZdMpW/slL9GDi1n/nJW0qa+Femcw3j+98jogbKCjLZlLR6wuDrwNN/X49
hOn1JckUGFS+n0xRhbJf+FBZ2kki4VSdqFiCZV5QXItLuuIlF70mH4qw7DMF9bEm
54YkGChCbqALCXPnQ/NT9OlugztYvP/kExTGNFr1xUAOk+EPTUau6rKTNjpLVP7z
5/0w5m25O/YRzLsMt3DetxR0cHkuL+s7c5NQx8FGDBIDWANW+Hd/ZTBE0Ur2JVp4
UkoXLOV1XayBl5pgvULe/ER2CSZHe9Y8OZrsSyTrLSF+plvGmZDzKMBZWNOg9t+m
HWU+1nBZ8TDgwnXAsJLmw6qfD9v38mz75IRKsOo4drDhO8XiLnj4AhLsnuNI7HPw
VFGzJqAw+818X22NccViTIs6Z0aZXLwKTbSUrFCltP/T13+lN28cqTditmd+ZSdF
uVcrzdIzBEaMq+UqNu/YOVOYoTr3wfsJvn/EJUXu6VsR8wH922Zz5NQPJpC1fIQh
RH6yLrOqG9KQ3n86NkW9QB0Pj4v2lAkwLFimt1asa9Y6FjpBn9MDLPTlBHRf/c43
E2yDq2MuXRV4GGf+mPUiVcmdRNC5CBnmWkdCrqT5qBk1rdbJZDV4j0VVAs4RFop6
hDjzGw4i8ZUzHkgAYgbavwb67cFLfIYZyA3UtiIa5RqTRlIY3QsZmu4dzDtdsvCW
Bm/Sh6f3iSATRkAxnbSgp8KzuSykogtJpA07t9lCo4QtPcYWjWFw9ZdamY2GXabX
4YYs96S1cdV/WzTRj6fzccofjt5oYtoV4J3L5zhZGPXiEhl5WYaO2R8KAS6HdYng
BExivZsMucGfv+mUAD/BLzUGRJZLPHQUnGiQd7580pOaLBmDFP7eTwu27K3x4QOo
TTPF12TKwIzQLe0M69ey5WedXC5YnPBDM3eg9PEqG7pumaOdYY/cyMpBufxjQ7vn
vBNVvC2lfvXGLImtYu3kOMxqmABRRkRg9UWbpuZ+jXcvfpyhaEAH3JUc2m1/oPcl
J7dSIS/iatdtwXM27GHmaAAVnb/hc/Ady0VGmB9oXIjqejBNVrFOJdbbFceknTnt
omCnS0WSb9vmNjTlKC/v+/nTf6/TqvWKW9M/69BzbxKD0GgmCfgIpCUMDX3X4E/R
mV2Kou7jYXEFZ5WqjZ6ddlbhbXNMZxl3P4uC3GTERzsVbRtG72GxMXg1Ow8ckJgP
4z3sIJMV7orqUOBmgNf1gs2jWY1Ek4KwxnBK+30cVS6LNfCqI9cv/qoY4/nPKtz+
Dxt1ClT+CiMZIHdGOZHQE0oL7pcBLzbIQcI9UyFZ1PsW40gwSHlsOVpo9kXGxWUb
QIvP/6yI5QMJ/dkFDeohyuJTfDLupJzY40SgCV6hlvpqDdL6+3wFjz/nDKuWgPTj
ALk47+5xf3PBMVpF61H4jC8Vt2cLHdFPzUnT1eNVxnIUASccMZUR88p4maE5uK6Z
ASKHCjAePWXjNS+PSEm1+0SZNhHzOGr31roFTP/KKPVQ8QBubGJJLonn/KEl2KVC
J42EFuoahnaVkS9HwiT9HpdI09pYOHkHH8UZ3aOpukJzxuofmKewyql9vJX/dJCu
8wWac7UtPjVS8Osv4Aw1bujWrjS6KD17RBBEG6FfTPfUEjkS1TRkZd5OLX6sOgy2
EdcbMw686h5PJmscdNKo4pm+zJctT6CugRtxbZqsArMJj97atFBbZzCVKYdjE/yh
0keEYyYT54CBc7rBboaXMNfaswTrO9X951+3mdHfgGJQRQXPqByYqmS8oEVCUbLo
l8+NYCqK6TS36wG1pkY+dDCz94hzjExxOpLlw0rfiuovsVQo0rTKC+L5fjeu6DP0
ZUHvJ8oWhbjVweLSSlM7dCP64unYsCGsQ1dxsWdnjq+xd7lPm3ovCVSxbKKZLQMI
TZvL878ZgC17GQ9oHwy8D15odDVbKnKMwwjp3p727Zs29ph0gcIA1LeYd0WW8USn
SoWkC8SNzy9HMw0plDGkX2TanFnAuJHZzeMpLutm0RwAzxB9/Bk02eRGX0tZJRoH
iX19NpCmUO6tx2VS0aMeLScroTQTlX2pzyilKwlYNc3QO9Rj/7jmhychg5d38pSh
Kboc4rWuoRui38b34lkGudK/BLPmKnxpI/8fVKY4oBcQ8EgIIkB2UQyWvJNrat+8
YQoayq9yiisLP6PT2428Kei1NQmRwH9dH64ATIla6lWrwAfo6e+qR0te+KibUrMN
n5TdQk0eTPGktuWVGWTZpt2v09b06TSreP3k+w003G5AEzIA5tMfKDmLEZiQ5MPg
35+94i0hbiLMLYlCXVePqV/kqIjW8xuXg8fRh3ZgKuhIKask9gBApL7Iu3JH6Fnx
0u9CJGmGjQSC06GA4j6iDhc2AFL0ZlLb7rwWJmMKZ2CqE+0GpqFHKPjtdKWYNBiH
w6K6gIWiT/OQaQxIfm04I/Tc60OCzHZPSy/sfPGqv5GiBqO8hgBEFk74w9Pgpf28
K6DMgODRFxz6wbWuJuZPUPMlPxEGuB8aJa2VuIYuP7cdyg/+gnBT32EVwt/zq4Ym
tbFuW0X0mSHwe2suMF6PawRIA9peeDcTp/j6Zp9jSyqnTIuVmHS7tw9ttD7adnFC
tmBXLB+uqxk11AHASHWPCoEVK4oqFEG0VzrA3L+vD4TinCnsQ57yeg5F97To3PZm
FELLfkNd/0+nH6X4uzSz1tom2AltQRTte7yFDaBquxML1vpM7rcXdJBAwRswKoWz
6QUZXwKYULhAUsmJ4hJaO5a5vIdQ/d6TRfc4lLbMPJdE5DaAu0nFkxCT9FRWgjhJ
j0H1/rUwwyK5eUNakXICq/OCz0Q2Llffv3kRGF92liA8QkpSGPQGb24u5NqrkS/a
LrZBdrpuU7vgjpVbF7Ya/DRSoMGoXHyeg28aWTkNsbGdKsIRVZ9Ks1bxZsOfsuNY
eVNNQ4QJ4pDEqSih+IALwKqk6qnMuua65HA3PBdWPWhVqvxKpCtOwjnk97WyDzup
LEZxKmGUS+phJiU+CyMWei42KfsclKJSZdDOx/SlGg4A3Id4FxD7l3tW44/5cwHI
k8lAIRf9KpEmk37gbtc8Q856D/QBrZC+IRY9CqHDAhVEV1idwtVwCuD/i/aT6Cys
bfTmhrW1RGGgmOJKw6bcgqA/p82itgA7nz4UUlQ5QOoqNOnwuv0RmAds8Qc7QNP1
8GbwmKwPQgu8jxwWNVgqBaTbufZh7e+PYzgJO/EQl4jTgWqF/S6XH36R7pVFlys1
cnT8cOcmSBcIY5I5ohkKs5k4ZKk/+NUBO2ZiXKZbyg4T+CJgvhjDyYflUVShJ6K7
OO+5jzX37PVJ3BIrI7Of4NKfsMxuXuMoVnBufojykiKnGVJOOZFl7U+FcAKU8AXR
J8XVcv1k9WohtqcSvD9IzL8LjSoGHqgIGDmxmClyXYIegjFtdl8swY7TdN/UR7GF
7K1nEIuryCEMMqIFMOWpo/vcUFX93Z0CndoToVSWeddpeGFLBDnFXdzvUT9VgWzu
oxkhdAC8XyBoYTydz1Wxy+2l6YIG77XWH5r0DHhKXPonDYWMjwNPq6K8D6Zm4Ouf
V6xVeA4msIhY3/SmdEk7jTjuHQu33TxTJtIG1u84KPDVCPBVE/NTIWiYvi+oxiVT
hJyhlhcAn4qnfgDdD6LeKhyNWsEwtsKKKWspPta7QQ6MNLV+hyPHN+z5hE+pBGM8
jDhhsiBlSOPnOaspcYcHhbhsspWs51/YhnaorPRr0+B8ZeWqxZZNas2FyMyG/eAn
zue+T5hbcQOwd2MCxP7klHKJRiA30/MGD5+07lr/4BJzsZ+O6gK+vrWNqWGy2zCT
iMfPcswHHUKeHulOx3qtgvMRtcZYf+NJZHNmpW8zr4DBgK70h819gHgZC34fzVg+
BYqN1K2J5PkNbesjg3gfMLX573G4Mji6jYQ73vdDa0a193FHykpvjFQxDWZF83al
WcuKPzWfxexykh3gakSbPO+i/Ley8LkYwQL09uYpRrXLPZhi+62w+t5o6Qy8IOX/
Ue/8QcK2EiEqMb+QhwwH7eiWmx6H+o0GQj72HLqXrmqK5fJpH9zm0DHAO1lJ2vPD
YfbTr+1SUTYRXZr/dUH6J2mLgnv5x0/HnG4r8wxphf0leeV3QpcZebWyrXnjKnRe
px33VYR4XnbFvuX2t4YKTRzenhNCa+ZK5v9Qa4eCAu/JuIWoLc8G8QKLk2Gy+kOE
011wZ/x6Ykdm95KjCvScp677pCFkRZd6e4vy77HMZ2DXjkOpWx6nK5BjguI/5hII
yrMMNzcSXQtan58liiiWVROJqE8Qp0Fpx2DkdlCAvIMqF4u5oDzeaALUJB4R31/e
Y0BBIQsvnOBSkbyGJT544X7tY3I5IosaveVCQGDa+GMov5A8D4s6QRwmdRhqvDe4
63KnnqJz/76bhfdUJZcP87EppgP4yPmZLCT02ikaKa3vAQU9w2tRooTklRy/JVgL
IYeuoqVQ0A5L6f/31tHYt+xH8gOAAD916qiR4LsmcIj85yZjzt7XJc1XomsDGxEb
o5HkK1AaEWY8wrH1/u1k0tqRoLvgIrFStFee9Afs7MKmvH5vbsL60h0A4O1cXqJv
zTSte3wKLA+2dEHZ+lqC8NNIMs4CNIipz9V5FLPSWV5fLyAFiDsE3/kp6n1BWxVZ
FJ9AqJq/yj9FefjJBaqg4KvweYPemBY0cpX/D6HLvLcSw10dZjQiFJPpx8UIvN5o
UcCRMJsUaafSdvk1lD/SSoAN6wI51Bpxg455aLwC7WGNYbqZwE6f1X7GR33FOEPr
P0A5Z/m/gXS/9oy9x3xpYky6rBTaTjJ1PPD+3V4vToPWnluBPvZH5rVuatVK0RNt
XjDM0AtvEsIqUdWOJfpSV3um8ez5BJJcOGoUWXszTdBL5Ylw6JsPJZqwuoZwDkrd
N9W4FxX0wqYyUt7EgxnfShOjfU3Xz7PYT7vVs9B7mFWmPk88z7UmBQA6LHrugssq
llucnIJUmM2VXxiQYKxuiDIBw5MWJnZHdBGsZ56dh5HosNP8zhu0qvwLB3a9aEq/
PAS0LUoyUfboB/WOf5xtuuTOsYJle8muksIdRTv2XPWNDO4Ln8oqz/8ZjY6y+pVb
561Qv+ofaLHU92XKXYSSYHeFWcIHm1G4oC1914Bi/UnIvjKkBXaNJ/s9ZuXeoX8Z
IHIytJdSEoHCEaP8e57qhArE93pw2LoEG80eIlpmuayDqAnCJf9sgUjSSLftpbqg
4PCOEwjNOg6E/9Aex8F65mDTJl4I8hbPVyqngP9n7wMlJ5hGuuZ81pHXLmjcnb9r
cpksVcqOtznFBgFWzal3rlukS/iP8WlZVzazkK2A4A0+8oqrrkEfSZp482xWHc3B
77uuotl0TvELPfWlpBEttO1mtbe+uVMZRhgXpFCon+Rg7q+CN3HVH9xGwQ0B+wpr
WXPiDRHt4TJc4ytJbrJUv4Y8EDYkKBWtpULZJ8Br6wFUymKLXomlQK5GwHg7ke9m
hjAYeKiXLrrSaKVdOtTnbGH9xRmtVIaKff/QLVlF3ROcrpNNNjoDdSFno6YxO3PX
rxdKjGkG/hYU/03e4oTRoM7o7hVkEYKoEUwfT7kWIkR8sDVUncQlwKHlLz4bZ9Fb
sgEFUkfLL2sFRFkS26XPlqdbSma2yZBtLRgnO3qWeId3acPiGl3yRE5fVjqiy9WP
lryBsa+7UHHdWmnhOafyMFjP2n7+J15qzr815QU2C5w06dPguuJWLdhrWTr+X8vM
lpcBfz+no73bKUDrwQuLVxkFRVSBsJOCQvudCPNxOTqt53uRXfp9BL2xQmBdcZ7w
xqQBlgw0BWL5hf8YetlcfCALvcvjf0nhCZeT8BsEiaP7r08BwD83YG2iIc5h+3Jn
rNEgzSnzv6HhwuBnMNZROzhvJhuwU8qQpLkPIvET+oqT7QZ39zG1uHInsIl0TrhM
YHfSnvYTWo+np8yFke1DaolwYOMgRfTmBdxXoHhq715JGEjCjr4QA2YcxUfBMwvf
v/IHFP3+ga9PNJ6K/kIE7eTfsv+Abh9JFYtcHCqzVaOcP9OHx+7wTlnp/oBQcsFY
jY2CQYIYiGNiwtB133uhhIjoOEKnzn/eXfEo/xTFb5bbKV2LJP56CEEx1/9We/gc
tbfA1Z8VWBFENXw5xqlAqfYlGxeMxHo4PICQILFKKypC9NiA/DZ76NI6dyqLYNql
TqGEXeUpR/VENJYlNpuLl6wUS/4rhLiiwwrl+HftHNB/gPjIFEYb2zoIXAtLinpE
PiUg+dx4SKtGGnm5Pyx2D7IJtO/1MJBFxnZcykUqudeAhWMTW4/u0o63OvEmWriT
N42NLtZCEdatqGnp7RVMBlQtiKucfGk36E1SQI6KLW7g2nHPcQvaQ4spWiR7DUtu
kX8uR8WDsoxyvecTKueBoFjqIWV3hl88EPYwA4eeZkXALJMg8ByBzyKRCw23hwon
izxaWuJkmb45C/Fh46eIQNg7awwV/khRqzveAEXckWEZgPM4ads8J/UKyYEgjKn1
+hw73Cr5eSQdKZ+qCvT03tS1x9yubmQDkd7GECpcy+LnYA8pYlQ9eStY/woUUmTa
SRxzPRMtO5YuzyHMbYgsEn67suM3tlgs7uS9bLFWUiAoc2VeWJuDRvL5GR37DAzT
PMO3ol4pYV2JH0dL4WDK0FTtJ6nAW0PkYtgCYV+Vt2YxBGRyQXK9ijc8PUuyVZqf
ZiBV5H9UsDP47RwWdqx3+QIqVFycr5UJo+zvYMiG4/H0y6MnT6pM3RwCzRYDhVoR
RPdcHLTfSJqzCMEM82Q9eo1zch4+IT71PQcuaBAyi7PO3FiO/+Vm1MInIx/fYH08
eoMrXbQzF2UTy+/U0tahVuPRM18353TBsZKaSc+Joe0bGgvEQVjk8olmff/bkL90
6QPMmIsMbKvXk3AKVd8loUqKwlXEExjQPIYaZmIB2Z7u7tKt/3Ah7YVW4syq9HRY
LrirbDoq/BD5q7FFzxjAH1w/6h7ntZah0njlm9FrjH3yD1WirnTsFgmnM1kHaYSQ
zPAPZzAzt8MlYqusiNlQDZfH1DFjQqUcpxUjFYFwqpTPU4FvaMYdSdBlpl37FdQE
Su570FHb3AmWqJu4ds+7lqBvIDWE5t6Ssr5jhPok3pvx892O6nJDBupa8NvBgGPO
lsz3PsHrLnBMQ6AG1qfQgvMz2mQBnW/uT8n2kor4KNMRok9PJgDYgB+z8YAJThYq
WU8D8V4Skp6qttecOaJi/8PL0cjcviSXc82t2HIv3rpcJS7a7c88qks5y3Wq5cRT
hqNffVKcucM/NWT6fjpQzZqR6F5l1t/5vey/JdMvBkMUroJNQUBYvJqTM6xTho0U
5ufNZoSYOiFB5t2nmgqsNA6zZq8Q7448njrlQ1N/966C7yS20Z4Of64zYs3UuzXm
RkYXqvTrb93IDXZVY9N46O7LMulU6BzDeklk3TrzUEnLcC1yWrxtXSaUgNcG5IGj
YqumtklHPv5AQMjGy0qEID+kblh/xsB3UwkhP89WjMIVu/fKor2T7YLMe0qhQvNp
OVe5pJ1BseMYxyBfMSdLhKZETrZ/IELvJ0GEh02CFHqQ5UFhezZy4mr8nx8E9f8l
Iam9ztiSzJxFO84N2uCZANYT1sNYHXFFoWJDaHNgwcdB7LX7bo+bQhCTr19rWINu
JDpkkuGWO+bmT9fvVaGkKr3JwMSP5/I2Ps0fySZGTHj+eLoL1D18kABcfTYc/eAo
7uVVspiuse8Iu3ytaAlHn1ZUxqp/U/HErvX2OUDvszLHST5Zb8TsjlHeaZkJhZLy
DkGcRPXgbqzdI6t7JaJRhfoDkzepwiO3potDKOkn6Uyi5RTanf9AUfl6zCiJ8SHJ
dppCJHaZdOAUqgR3OqeEvWeUsKxD6uNhCCrQb4UIFXI4Jmt1XM65sjVz/S8C+j7a
v6FB18+AhaWtpyFa9FU8nQAPk4jIjTPKphZzsAmWrOGj+I1iwAZsd4k5+iLrCmv1
2keTl6yJVUziGTRQcXRmG08JifGbMA0wjP4mZttSo8ge7XhTcGI9Od98WgHmYxwH
npl27Zb4T0KKQww8JMaGTXQxZRL9BmYKx9BsvRvAd+vKDERYbspKVpgXaum9Xgmc
dxie35HlM0jWg5ILdIFcXnz4NLmkhnpJu2KtcrE10klg5jTMqzrFpwfrHOOCbnz7
jijO8ZA8nSs3Xs8RnVYI0/2g7nNpl10QQA46Q0hLcRDOPx2obaNHUedWa0YfQYZZ
B9Lj2Gp6FKgpOYtRrXLs8Go8xtrkn2Gn7/a/hnGbqCwbXR72dyvxP1P9lJ1v/fBC
5qnLsUoscW/hMw6VDdYhG4imqen3djB5MzgkeHYt8cuoQ1itIUmw41Z8pi12B7Gb
36TUHixG53FDoXWTuarj3Jk+dzqmQv4Xav4aC0o/KXmzwD2erYGLiT32wBbN+Cpd
tb3/cHlPvEM6J1CHsAEyr5+t7MwlkySflsPioN4l7Xz3EEv9r0uxbFdJUGPrPwL8
f3v8ShWNcq2TizavJzlVFbI6IAeboR7bkzEVF6vC/4GPI1eerz4yYza5JivUEAUw
bH7e2k1DmavKk7xi/Liw6FAJaPPgT71Cc5ZMU7FsSI8vy/Si6X+GZvPLYjnkI/ED
6M+9VL4BUEff8uSvEFzd92m9rAtNxBSizWXlxAMXrXjMVbO0Y/A/vq5/57hwjOpE
1Po9H+hbUW1Urt5AUsOPecBvpg1VJYVq9xX3VvKZ2jq/WjIp9xbbXPGQK3JacEZ5
Rmfl4ouqpjVNGHecr9PwaPbGu6WUXFKgHLqepWK+x0YNZ+jrXvvqJiRhPiZuYyYA
nvZLG76uklshVxBgEMUrdwCFJpEMRt4g6R09q+WvdB51BRMFd7BGH1PNFezUB3U6
ifAt2NDEPGsB3PxVx3ounpEXOjETfxuCDhBQhYEiIXPRkEqUKRq2C5X45eR5YkkS
VmurqzvnOjjwx31A+ID9D7HLwLA7B3wgv2C4NJxJsYhbsUPZTC3/SmLfPXmOQcN+
urlsVLMpeDZs/QM9zGRWk2u8dpvOTI9813mvS6fhBu4zzciGAX6+GZBydSgv7Nls
IpvynVWIWBtxJAp/qLIItF87/e9qRTRhzmluscLLUhks9+Vp4maCGiVEq4WwPvW5
xcdV+Erpu6ADtYBvI6ridRBVJZPT+k/wPAeTFTrPjYb1ls2BmcS0moORKXM6PD6Y
WobMY6sZsgo0FtXhdxSIjYpdglzXqrPLksRES3OF9j51j/CiLXOzHfDleMSnk5uN
wPdbgRA6na04IGFVeBgqgV4zG3fFF3jbJZD3/21uPS4liPcnPMKDz+Shk0xXSs9G
E7qGes0g8eOOwJKXFHyH2zgZzdh5CSTiGpMJl5tXEWEi9QUCSzVCl2JHTmBaeKGX
qh1oRQXkQoBVBnX45sgDLhWi6uSQaQ7msl2kUx1N1kwVy8/Xvj+4Tg4PLLQO2uCw
F6pJi2lM94CPbXa3mkHPpGbe8J8+XksNBtlqZ+74vKstC7QRS5XGdFajL9DRTW2W
DCml/zTgoQOhWnPqebkwP+r41mLyXHAaTWSu8xGCV4lo1aBtc9b2F58ZGfvKgem1
zdOE3EhjBGq0hWBWKgbxlJ01mZbqraLao8ttUeHmBs25gvdrmvnXXVf1l+iiNw5G
f0JudEUkra5pifvAD3KwuDjdBoxl5tfG6S6BxvG2W8Jp0YAMRwBVXnLeY28KMpaa
EIIeAPhZBqZeVsUXmKSWQgS0SaaStEUrgi+XGIzO+XCjF/AiHIhMy9QChbN7AMbK
Cwh4rjy6AeiCyfouwr94OjaL1CTikOPd3rIJbI4yJl2OPrr0uBKPRIb3jXb2fX7J
q3G5+ygK744M6iz979de2PKgy2T7tmfQ4K5xM1C2mrsKsBQBvCB1ayN+A+dBTBHf
o2dtvYmSBeYzMVyS9LdVsF3SjCI0CoNUK7e53kOWdRd++KUygWaqLjbvRmkATu5u
G9xnPu3MSugwP58uFYCsmjmiK4xJF4RO7Nu6nuVEIOIxd2jalP78IwY0I6gXKX6h
0zC9fWIS2eGanUhGboTz6B0Akq8TwRv1aC8Hat4/E8tLWjAhaowt4Ym0onxybHxS
is5zuu3uHLh614YIhaIKdAr54QFv87NI9nCWnuqKUv2NeADy7a7VkHEFadVCQVZl
JB3Hc4LPniOYFubtfH9SzJmD0+Q4HZ7WweeFxx4NkX807x3PCOhSJxKZr2BE9szT
5DDttO9oaS5FT+LNBlkxLjMtBi9hgx0xciTeIWVRRPmbV7ql6NeMOa0nTfeSoQqK
r1f+QlozQK9hZ++BrNTw5K7DJ6Llw/r4D0nJQunnXs+kNsYalvsefWO94qsTonrw
C/Bj9ZxwDxOBOQ4Piab5sUlrE/QvpylOhxt8L9wZ3QL81Y9hx2HB0HN+/FEDpq8P
Tr94Mjilsz09NWxiWc0wk6F1t2dTfHbDTs8fMNFLNjJi17yYE26nm9+iv9HrIn6D
A8KJ9k7/uLUqHSaIb9rFnDoAKf7mHJJONfi5sQgnQZBc9qvavpjGj5ZWqUvdMtxr
9PFlX+lqSgWL94soBW3XGR3JHiic/Zq1t082kConDvf/dqcFPGmijeowrDRbdhOb
sDO3cwRRkpGBIXR/ynYk963Fyb+7htlEW2e8EyEcHNxetMkS3yIpciBpSuxM4BwJ
6DzoLWDhnOPilLBiEubIB7gCsfMoIHvsHcUopyNRiSjvB+5B3x9lz9GVxqvFcIqT
KdyQ5sDn9hj8RkUxANLH5LeK4t1dqfcIMIAfBfiz24or+KvH+JPZ3kttDEWPcA9M
t5/SZc/YENVMT6L1asGmKosNEsIkq6DW7IAOaCAWoQA39jTX1CJuE0BSdy/IO9NQ
s0irR2Pii1UKhomoVXXcRWRMJttBWvi6sdAb8kjm5mC/9OWb5PSw6ZBV5ujFMvmH
8FuITXOxTphOoGcsYLOtwTfo4DVswxYhM14se26U18uRtVl/GWML33Pq/1BCnLFE
NzlB2fXIq4BIUnxiD21aVFo0MTu2m1U26mkkrlS6GvfLbmA1/ss12QAaIidyIPLB
SIfWATl50anarZEMgQLWznrf5B9b68VvuYURaExVhaVvRgVhv4ihyLd7UYNHI59e
FhzDLQxJIrVwrNjTW6YqMT3EK7z6ObS4/6bNLVxYbckNEDBIsObscHKwMMue6F+H
A/8HLv2mAfh7LKT07uCzBupkbUqTKcSkZduRvTe5cgM5nQdAjFgIvKTDYnDhdA5F
qT/MRHmRKbF20r599yYO56TDwv1N4Bv5Umz79wyU+VM+ZDuZOfoqqIvE+pwJNWVh
kXq7biMclJua/i+Y5K61vQoQCL00mxfVDJAnoD36kHTogpJWz8NgCKtuFE0grW7a
/eEvkWf0+nACnn+T2ZAshAvfReILWdspJIg9TW87SXpjAtJd/n7JbUAk8gblyW5b
W9hz69RzcySiRDJuYKgrlhUFwedKcO1YACuEHzuKENOfZtYWq/fGvKAoMw/DIdGR
IH70UTdaIkShrinFHaczfuF8vxZbLdi1xHqG263uzk0ayROoLx0TpfbE6idi7hfw
Kon/I4Q4ics2UzS0Ras4N4KEcwqd5RB/CYAj7s1ALP7dg17M7TOle7khK4zDAgBz
zx8D9Ajfpn6zVp/UxeHXqLlbz7s6zMAi6jKVW/OBY04laT1PNucD6TOAWhq5RrPd
BujAE7LkXqp3iNgj1m3uYm3fPB4V9/7rgaPWhXLlTGm9EIzv+BSjInWkYQ3SP/FV
nBtBjx+VNeEbOm/AXe6UOY9uQDKEAMF3I4/CMv2nX9B1KRwDtEMQ/T/rcEil/dt8
Ah79bPnFhDdT8SsvPfHdCAv+t4YIONGwKY/UddyKSIBaVaP5j+tjOgLT5+Fma/z6
dCqC/iD4/gGI0/9fd5wn7EuPizuNM32RLEO58Vn+VMID4mljqLU7peVHSWI8Yhto
Wi2ZclfnnZf+sjrSWCeG0cOThQfKnxuvFYOnDBU66Oz4C4Ne88imlLgGc/H51ij4
auEjKmUJa8lJYCo5IerLPINUI4YzPDdsUrSwg07hcUbJHtNwIC1qUns0DocvBYus
nq2YPPqzMDqgWNF6XOSAOre7H98k3s9ikBy+dEm3PlnStyQiHV2UzAJsUruVOM9P
2jOLye5iR0otEpKf+I7LGNRvwSSDrdF3eEfEHU/8MCdSHuGSUXcEQLVfaDyKotRG
1wu25rQPFUAx2VlYmEMB28H4jRiK+6/7Q3swyh55HvPipMAciCg4PyIP1jeq6cRA
RyBvyaU4p6TklgyWdgOAJjf0kpbzFuZ85vXgFkIJAdFL6AETrE0n91I1rXzCDuq5
YvU+NFjfJmBUl39S+IZRhl31+suiwP9VHeLqwnyApwILJ/g6ZZs+2t4rj+9/8L55
Jf7dZ68pWQL9xz8wyQG5kUPQck+EcbE7oK71ysC02AhFa0XVk82Kal1lY/xOtChe
tn5U1neWHUvknXhbRuX/0hr/8BOFXtMcOfHTkoEBqq8uIL2ypSlCbbIfwoi7QcLO
j4WI6it8BPheBC5ma31Zv48QUUCJANd1Qfo1SWgzyCK7hGNHYao9BoKqjFlI+dXf
wGAPRMnuw9xTBB/1ctpCz2DX1y/aRBUt25pep4JnPUEK772KHNEzgUi2INUNM0t9
wUswVqiJ7AHsKfQodUPk2d411I8U9YKW2b9AOs1QLlblI3GFLUFWDT2wZtdeMct7
vR9emxkbLfsyZHart4/beG+ET/RFubiH2DONJt/bWo80+EY9dupiGppsLm3yAfNg
3GJMbF7I1/00hOgc/bxfwhG38DzPJqsM1mvfihbFVRvZOXmuaxlHITY497onIoSN
Ozv3/l6LPZFaOh/nTpGP6y4Bjn36gLefqIZNamsRf362i0z1mO194JPVii9ugVTJ
ZlgpF10ohCFxACK6gwlS0XLs1p4GCjvQdqQiQk6Jq/NF24ZoC82QVkRkahe//3ap
/WBYIVwD3cUyrxrDoqDCThHjzCSiGcpe7RUmtpvFCiJIYsHeB6b1nm1pBITppvEx
zNWT875F6Z96FaO9eSjSVIjEmiOaIbsLyeCkH+rYVdXNFJrv+F2mANvBXCwOcdvE
BOPZdqPaDX8uLnVWlf4yMgAeCyB+LLwuYWs6v+AtqDxVOQN209BLN3Lw8lA31tqC
C80l8QB/RZb3t3jdg5poVOhK9kilutxaSvP6UPqzgvzYOiEhDDaYUv3fzGovSC2O
zFjeTr6rn4hRE5AUmfooEkRKGLdbC3PCcEKahSsNRJugpKwW/eeFOjRUOCTyHyyK
wLYBnPe2MQZ5N6+IfOdmx2EL5tDBUIRnJGciQmmZzN5ninFAcT5ZJeD4hffBfQZi
QQUgaHgWCNNBSVZYKY2V7BR6eB4CG/H+7atm9SpDt8q5nqW/iDH9sKAguXvyx9/r
HnxQljbmEqMgfVA3I3h3DY+xX+kJHkANeM82nTNz3XP1dVkdS7vumh4sXy4qBcu4
u9/yJX/bi7r23qdOtsAKuAqktnSWlQO25hz+jytwlaam6lkRDPOQSMD+qMUDHd+n
P5HFnRhJqIClPKo2+yNkUGQWFeo5F8RkKOs99fqxEf9ZKhDLKMYMn/Db+WWJLhpe
/0cZNqQHZ1OSwAA2PrclTcsM0pvclgdInhqifWgdxCgaK+o58nD14Gmn751cG7Qj
HwWA3Lw72SGKmRC58GIAYvvBJYvB9ldCE1sMcRUFIndcdZJEXydWwFC71XfS+k/R
WK9tO/CI21hBHJVVe5+CSzdWYVsKNrK8wQpU1CZuuB9zjs+vXWw2VZbG3e2LlVKr
enyA9Y06vU4+8nk4E9Wd0HCg+QT3SBYZrj3rg/+rqcMYo2+8ACiXqo4NnZMs+nxB
QDAV+/Ez2nHhjvbErpyJtc8uSQK55MHjEhIsNYo+n1Er8sWhp4JTtN7+jM9PuVG9
ba58EmId7UVGB4QwRrdh0rGA+o1O9sOzltxGZJlO/qUkU8Pa5oe6e9h+CWE4xXI8
DiNj+Z/3zf5jZj/X5BQ0GaBtwYhfcfg81CnyAmYNdqjyrzl9+QXhkSv9bdErc/t6
SkUBDEIRqIvFF+8btIxPNrSyRMeAeGmneVhnUVVLuWGSr2IrkCNvXTBa4e5HKkzW
XZTJZ5D0IkqQWj8J1sANaMWN8BqrVdcfQwnyO4ipv1I1SkIrmgL32/j7Mt4Lkpdi
FBnwVWbBVaClYbZ1BIRL9oy/0Bj9hwBRICWXeBNNkLbC5p5659VZgcZC5XqJTrW7
ywYIyhkMcYos75MLtmm3STJX6S2EuBB9gUjdEtTWdX913PVNNe6WyLxlHkJRfTK8
pQVY0QJsT8rTM3W7dfHVl5edMGbIqpgvTc8XCHmn/rwf1UnPdD0EWHzYe6BkxvT4
SIksXCCBI0plgU9nPa7eGwL6zE8p5UnPvkw25hdWEBF5d5oUjDDZf501KaPIry5J
Y0mfUaqbC6BDV/nNP803Hs7tl33wM7t3yLdvDFQC+ppECXmxaUtN58IJc6oD2z0B
gO2Erx3AxSkr7k9JYdsEIMwvvC6hQn17Cz9KUUnlDOlw4fWYoz4gX09zGL/viQh6
LScMfSllCIzr9vke7OrxOouICq4t6U/pKaaaVJZkGnBaSFTS6GB8yGbvpaFUPvCt
O260Cf9FXOFf2+h9ijkTLSxOVrmm79cuF+JRdWPUzDdcEuwFVlNtRgz32PVlf0uB
A61OkMxQj6gGZPhOXKk5DjuNVSBfYhfmPqO1RPH8igDIfvEKqFmuHWerTaqgHKwk
nd0ZHAteJIkP5aBvX3ng1oc3n9Lt/IsDv+Xy2Y/LjApavEddBb8D9WaGr959Ki9a
F1dvN4ptabEGwOcjwPuJ0Yt1/H/dpPn5aKQaUVdY9fX4UajpKsjEl3GUK4FETV4z
XYPhf/FusrfvlTk5WHWXVJbX0hkJ7GD20FIbw/t0hZpT5Vwd/nlqcnPhy6b9lxB9
4JgQHaBIhPzwcMr/zq902//kCvMNZAGX3+FmgDzHDn1ci/gnu6U8yqDUD5mWnuOq
O4Gi+j+AmYOd7pgOT1xVHxuWKYMlgDnRxg52JfuP9iVaY3dwxInvkwPWD7IhVATN
Dgh9LjB/9J/F0WH1N4W8D5WyVrU3OvKfg3hTBgLIz4yOH84tVEyO8QKHBygbXNHs
GUb8y4omIiQdy/9XC7lpStSHXEwNJ9vLKep5HS4NrhULFJriAWydJVcQe3RFM+GF
jHu1UwbQpsm/x9F3aj9n4JVB9XKDMXoJTlnaJRD5sFyuXOc1sJkXG8K7f1YPMgud
kBrIZ60MnN3Sp7Xbp5gfP5sG15/xAFSMMn2SI24jfnd/JjyOzjKI3nzNn8W5T6IX
ucQz1hvvZMXuz6sJvLEmQXra8OrXnJD8CP2d2uhJbRdtNVdeShQ+7h7fTZUS5XOv
XrzSJS6fyvONiWDbiiVuvmXvH/eGXexf5DWvuTTNyJ8zfJggoGvv/sfUAqBu7VUK
zPG0titFmE5RCRlZMKF319R6aH6D5BkvRX0qF+dvz1emM5WwAR5aJMTtNFFllZEM
uNS6UhIU7x7E7dCC3RyHpCBBlyDYM7CB4BKpTHToWyPZ6yO/c61dMlZvnQWl6/Ck
m2yLh+HjMynAn4VkHGQbhFK/FBP90XhJQl1mU8W+sWPakWhjyusFGVafD1katpyx
oY2ZMIRbxcf9LoXiIqb5eTQ72mfSpr2sAwRFmoXhxKAggCnEpNmgymJrwE1ATQ4t
0ERqwn2kShQB33yaJ6xWc0Y7fS+1TP21vk9oIhxDmLANbDqasSoArlcTMoOyL6ng
Oiga++avLIichqDVoWWeOToljDstt8WmOEAYu/dmb8jD0kyq3X9e4gYaSal+fcxu
VauC/swf6770AtHNFtpzpz4mxm948Pj8a6ZvaI8uwbQPsgxvy0iFC0jk1BnNcUKN
xakHqnDnIRGbnM7hWM9ZV9FRLPOeQ0xOtBVl477y+ETrG9mziKzuOvRn/xOJUktJ
uaFUSHwLsKxutVqoNyUFhDZDqVLXeC8VGBE0fdrtqmsFEY+C7EV6M/kRFkFYt/zZ
TZmcABDUr7mdjw0nBs84ht6xwd0MA0k8pcOA27YLWrVUiwDQjJoke9DJTX6LanvK
W3pHrVuMKuAbYqfpA8tE8QcKeEKbVrqNEZ1LjVXni0kplNdC+lnhvHzARNtyXG3H
6xNG4Muzl4LDarcs20Ah5mm+/nRMWdhp8Wpjw9NIlRByiytshmLZQA4MNB+WUrSu
gZ+RxCwkuDHdf3ff3RWH1a1j+9zyYbkydjE6DKK3F5y6VG/B+lm3uLMx1G9o17n3
g3u7J3SslCSJlQ7U3MuCZuu1uiFBimcMoxFf88qJT0KqlCV108OnDk8n6KFfXekk
5fsbS9QvbSTyX40+mLNgXs69Y/h0JQOWygdjfRxvTms1X8hIRZuOy0mVbsIbMec9
1nzKhLqcGPA3q/GVYwvI+g/A037KlOcD//WPAA2BsITbGexCgWn1wP6ap/KRE8vV
JxMyfSPVoBezOsjFMWEJm8GAcaeOPP6KnYdbzu5/FTQsX5gWE00lNUgZACVo0VwC
5TET68pKVh7+GHoD1Lv/YEh/tdtK1MEz05QORUsAKO2MxPyOSlinlwSh62KJOCKQ
G3vmvMww48HbfjkdpuRXqEoV3x0g6XmrT9gUQ+WtyPuyM4SErKKN0BGSQt78yBHY
DQmFWHCLBzMoqdZleXfZ0ZglSarYmU7Vz6s2z6kMKfGUYizKd4BuUdGuIz80/c83
LAivv27m5Q+6NZ5X6ZjHqJx1mABJKObrc3CMX51PtvzcvKhbpbh3r2Y00zGRes95
c70NHtPjCUlcgFh58MRfv4CjskvVzWK+98HxWmTYjJOjwW88B3uvrEVfwy5RzuSY
gFMxibrdLV/nB0EQj/vNfl+M+MH/gpELWMBDyE9ur01WKLpzjNAbV0Ll8w2l0pZC
/nKAU0uAzkQ0iyvwN5gQGNSJv9WOamtOgZODjqPacAGkrWjsO2Hk/otavvUOE9/R
2LMSvbozfv2WeLgJ/l2h6+2ukRCEenzX/mEtoKenMRegQDdVJSfOQ814wz4x6I01
85NzpIh9apKrpm3f16qW/v1F2DYM73FjR9ZnEfZFRSt2H+IAU5HIe/15v5226rCa
3E2Ha6mJQwpB8VqJzRuRwjl3sWRHojp15YMP1qdKgZavMBnBIA1f7AdhMQ8d1tBN
LmAyCPxYFgL/lyj7Go5wCknwu7cpxoJ8ASrQDbSv+6fwC/1yUObx1eD1iZuZ+M1f
OTq6hp3S6+PDjyFbBR1UrksB1YeO5ovV3yuhBkxjYqp6fNZHkFVZV6/HTlhNOV4Y
iNL1ax2Nn+9LuRyI5lHTzjFY5QOH2OcdaETz8Hjk5yLBztjLDHgVPUPwXr5BvCt2
30b52CRv7LlPZvfEnIwbYA7TVNAp7aKX+KuqUHZnw8JBdg9okIwX+yZNQaU6TGqV
YDgLNlUMLXaE3Y9UJ4K0PnP/e2HNngjxOZ7PJ47Z21/mUcyKBgJY5HWYGzCZtj9w
XQVzbYZGdQHnUbWgFxlU7JXZjUdjgxqzdbq88O1qPDiMNJDoPXQRvCPOotzCbkxg
Vo/0doSvSv9ua2UoZz8ULarY6Eq60wyyfeTa9Irneqq63obicM9vGibpcM8IiUCc
0cFiBI/CMV13+kONxy4TpyS5/Uj6AXjCnBQBpi+kJkttjaUl+UPlrXYph+F4vvqq
jvmXFMNIuWVbCiNtqXD8+B1OqTu3xQl9P1DU1rGziwRzQL1zwD6K+nRrRBQyzgb6
2vtdMzedHdZDfxlwMD0rSQNLmxC/AQUBe0DLQ9nCzEB/Y9Vmr5KjJmyY4zzIQt+z
wDtvXf7xZWOQFyd2WDCYhM5liVtRkBy7fY8L202Nc/UPyGpl8LEN1mDZtxTiWZ7i
AIT7P7N3Z358vBwU2DiO45BDXKVcWjGO69yMsIs1ci3B0KW5XNy7lUCMSqo7sBwH
52yXKrMwxbYygZgCkN2Ckh4tYnQvGmLe0Qwwdo6WjPa3QTcUnzxkqYlrlG+zhlW7
ComlCdPg97ibFVO1LwZrT/JOq9ELv+4GPTuypVaqAMYVvOedV8IqOdup8pHMZzG+
JlXM7wnIyEiuKG0HqoYzM51hRp+VcmU38poMqZyoQ3I6n+UtxD78X4gl1g9TvQKW
/4C33FQhM20PKVhSzDtD1u6G5Uq2cAPL4qxTr6rMjFQydWBFl2RpukkYD/GiXbaz
J4N6b8a1g3fchgxTCVb/yliMhC7V+GHbGSw6WCwdkBuV/H/ubASROy7Hv40VGWRR
Eq6t1NlWZRr9N+4qyW2DcjCPeCncuPtyHEPDtZUXPoyCE+3ZMYu9saN7R2wCZuX3
QrYz0CXiBewJCefjzaIe9ytj40U95mx/CJFHxgB5XGz4aw7/1c75g8BrudQWVwr8
UTf1QL9Rfd6MiANK8BQGiZBe809/VeKK5b7fwt0sHmLO0spOAtb+R7TxYjalxjpf
pAcTXjG77JE7jFOHUr2HRg/c6MTbUgJPGkdx/mTyVkH3yuCIgLeEFJh9cCNOehSJ
AxkvQ53/Xmh/Ch+gtzh5gGjhyOu6hNdg/DlWENHz7dTBkPWs5jMMCmaidJxZvY7S
bqQe0AMZDvQoNFdQ5uoGl/6PirpMEWXLf6OEjvFZEeqGmCC/OFgfkoNQLitfjb6b
B9eqoiUpuw0urx9qTPJ4KvqznBo6IQ3iyyd/g+/zCBfB6Lv2MXCxVLLch2arXdPl
tDwphM7dI7zjdnm9OZzfFdXUhWDIclPNzltB0+brjim5OlXp5Avozs5QWirRrJk1
X0qmz1/ipjXFGdPSnymL2dPUxaSck0yKYaSfm6j60Qs84SaxTvP11grDDan11fHk
ECnQzi4Fs7GU98RCN3vOsJbNW2kT/OtPAnSZeGwMsEVNA55HhS+24CwIvbFmR3sd
p21dwBA9TGab8MWKsPO7gSDBC1WQpVntVljV26b3//F0HingvtfHM/NPg9pYGr+v
W/RVbU32tJGMukeOA++wEhqJWeChckchksctzpGllUZKwMaMP34Xm1Ya5/A5Zlra
rqU3HwDuQ806pQlpzKUssCs/PkUrNNYW10ip21b4LetzhfujVdgH6+2OKlwGT4Tq
lOpnSM3RQqvFR5i+s55UW0aobj2xsJWMNn/9pK0nPfu7eOJjBVvk6u+ko6Zcfzid
wFNgz+ubRueznG2i8V9fDZJbMNzQKk09pGLqOOHHHwfsJ6mecu9mK8VKXfcBpLRm
Z/fYNRx7i4VTLJI4SMHQTyPrW/jgz00ZSooIt6ooJhjiXv9E5aDCP88X082vD4zw
pmRpooPWc3Bbe9q+Co8dco4vnKEsuAzpOIbmh7O5LgfnuRF5VfTfKXf+BtKIv/hM
v+5N+vE9AY/Uu3+rbvf2XxhRCt/VxxD5ZNhwZBGsHXm3kG2LQTEtlLD/TQgRqfuO
rZOVFrBWHuA9cbmpz/gNE6cYxB0kk1Qw+fCojF+xWt88d46Np3P7Z4K+BZCUi5Ua
RNxYkvaESfHUTT1Xbio5FfoKaHqbHh7Z1DZkqAb5Yl0vsPr/ChbrxHOdpoWTBStP
cRIFLv3KH00LE/YQ+XtJ+CF51P8McBlpiF8FuOPJX8b3XI0PDvbV5uSKjXMowSte
1hKCih1AgHHPmGxeSxtXDgXqARRjFuk2mjj1Y08Y2XABkHs7Q8IKWdlUsvl0LhSo
XNhbp2xChQvOKLr+ER7Ud+u/oS9w3XxDbifVSl5Eq5WiorBiPyg8oCxYn1z74r92
wCJOg4b2fAYj0YeCxwnO54EFBlKzp+H0+vVVrt1ko6KDByzJcZBAc67JcjWbXOX6
/vqXVv4bLWvKEGujBws8XUtdFrQP4JOcih94ou6iwPklwS2DzG7LOYiJUeoJHE75
HdWaktqOqixtIaXAWkdlp2Bz7XX8sKB3HRLxUx5WL0ZJEDghW435ctzon3GlVHwE
+lJYblZBL52pFsm4yftHdKMJb3FjJGA4jIw5p/f9pb2OlmbZnsNp9jwuHP/y6O+f
btLYmD23lLW8+mBVbZtJcvRB/0G7V1F67GRR0QNhm2rzaJYzElqF2Lko7WEbKHCE
i9rdp83qrSdSJy8bMKaoJUOvYDHTz34aXNsU+7JB333PNwiGaSeSEGQTMc/+5Ejw
Qp2NJtJkaBXgPwIFeMCCxf2/PjKQzjNtwgEOrU8xXSiv2cF8oNxg+eUbxCDsDkP9
AMRdk9G4fsKUX+ciOiUz6xH5QGOhKawrmsVFUp2u5XQyJ2U9qOjJmrCz244d+Wvf
NexVwFOY1jOylJIqHC+wZv5VDEzDmUToNYMYQIXZKmzK7TSVJzezH5HiBM+uP4gw
hYY5QwgoJbgPEpQkniVW9mLqdKcSRYjhp36dkCye4vx98usrutCY71ikAYYxJxTc
PQgrtY48yazoyZr7DgFsLP5djax4wNkkFzTm9se5rARDCbYz66ey0C0GNyTY23Ef
JZlCSFihV0JC1ZQf0Dv/ZxsrBT4wLSMOYdk4FKBVBgLLnb72B3uhTIsb16w3skCG
7Xva1qoInGVPNaayW9jGWilEu0J/Jt4zTNs2K52P1/+pvlyZoqtlG+EBPhEKJpOf
wHYD62liednlnplkrFGpHT/9T1cXgi+pZ+AlQOJqhnNSklDGNre28eKuiEdbN0NL
YZNjwQdg765gGGbUDXqOovqmHnhqgR6JutyP3j3lRf7vM59yq+DadANpmhAsAz1U
Z549msCCijADZHzoQdysPeGnFYrTYz5ru266S/HPcJXYak+H6tsuLlNVuPVUxn1+
rSqqVPvdtY8uaszUTch9Iw+X89Ab6v6oVOM0VITdX7ywULJxjubGHxDwnu4INm2+
EnWH6qDTaos15xWNv8xgghv/WeuacCf/+OlaBFzBIlrgquytS5GP8n1G3vwVZUq4
5iu9mntJYEoGJa6ypHXOv79FiAogn9q24xOuH0uCa4Yt7ByR9e560AUKauMR/ggN
cmkta9On5+247aUjhjwMVrVNux+nXswmqe9CGBWOnobnuVIlxf8o//QLXvcBzdIn
LqSmf0m5uV5poDm+y4by4OChZfB5zhee2Dah9m4VK5YyiAVdV6Uva84SFb2yS76d
tV0T8tg8zIhYgrj6hzA9M7JWwDkUnH/INmXv/X+9ehwvqdgW6LK4KhTmR8h9/Hph
K95huCw0yIjxujclhSofy+AgXAo0Uj8tkf9eto7F+D+5k7KLonCg+t/Q9Xfv9wg3
xrGhPmAr8xLdnSvS4xxOHor61fJFDTcq/4Uhhnvb+mLO5/+rX6/SQUzHYyPt3BGP
EgLf/CBdNLgaeiJs01Fx7MzAxd29Hnl/d+sbAi27Qo3QwlFsVOxMnCMdwHMof1oS
3hkYZnJTnwoPxlMzc/3cPTl2xM2TzjxBNP78V0OwzPv5/hJE6lV+hLhuZ0laONM+
jVGu+YXgGX91wQqlDqRr8nq8pLIOoFnJDGOKt1PHw284X5LRd7oFghraPLmr5qBg
bZ2+dMEQ7QIwu9mtr8xALHYF3Ym7G9Exx3yAQxfF5OIwf7FHzs7w6K/MZ0jma970
49xlcNBHK64a1QWShbAtB0toc6Oe+cIk/FWecoxK9nYvyr3YbFgTy0j5xLGKzOMD
rEUACmMuKn5Mw2cTSqUkXZ9exsEd4VwyoZAFY6eADLp+zWYw9V6c6AGkWe8np61K
qu+0b2dsq0iW//eUF8uhr0liUBEIwXClDY0IvVzFcNWLZo/VKe2V4giUnSvLszxV
x/2lGBRcbo8ZQwkjAgEnWXOTT+Kt8srCTRPqbFCc6l4sJKyHVk0vDvjUb29w8KG3
H7oGIqca86mzJJkAMycYpLAEH51ZrNQ55DUFQwD+yN2bjDIwX0nCMOWonV10jrJB
ttfyaRrMgMUheLxpcF1NNAPtW5YZc3yWSMH/BKY+yzmMfkp7qCETUw14WYXw4ta3
8g6gS4qSJMyUakloLmDgAgYoI/BsX32Xp8FXwBhAuEybswAvg3LenLcFslsguzMd
lTLA1zeE+Zzf9XB8+06VCtt9DJv9NSyN+JLU5noAzmeYKykgAmMe3Ds3va22htha
V7GW/ho9B8ZZS/XcuTnoHz54OPcBPwnW9kmfHjUtn3Hvl2VZbp96UeRz4/CQRf0+
msiSl+PfGDuxD4wMyj+xPINuHfuHoi4v3O+6g2uq48ssWJORRBhPebqpsBw0+srS
xVIFJOZr0lnExdiJZojFZ4mIE6S4H+HFWTLqHIzBj88q/BSQsFl274S3OBC6yjg+
tUsHnORvGuPPMklvjdF4BhIDyo6cdeWQUkRpTiOnjqMOdWc/beUe44pOBur60u3c
lwXtbZC4P2trcJtFxrH9FYldWmHYmez6pyfj7NooqyytfelYhuSdynZkUjbPCMU7
z58LSi76BLhiWrg7JOSfKDZhaZD/lgsfVrTZdsw6zV3hcNK3dJF21zX69yj1b5BW
lnUQs2pPJmui7z9k0AxiPo3+y50bHWK4bexksm91cA06+hUEBauNmFrdzfrQ/2jE
6I1ZBLVk3ME2QErTSGr/PnKmLOQK1dGRs76jasxDGGKO/yEzkgVwnOOWrLOSzwth
4EZH3+BiAFyOKS4PNMjf6/i3xRvqrsEErl7+eP+mB2LU77hZHjnK2eHRnUO/VRnc
tF4ceJpe2AREZMShAho6aiiDsR+MQ4HKXEexD3sJDhujyF4+ociEaCLZ+HpFLF+V
iMhynGED/U6wUTh/5mFQgJkYxBeFkupavXR2wPxt4IEgRNnLNAr6Wig5zFIArY04
QU4DVN2SyqE3Ya/N9EeFOeTYtpUbg1RrzMeExmmVL/6zY3gcY/rZ2zYf4+61zxQJ
WG4GCq49EK64P76DgH3lL2/73E3mSj60I5XPJ93Y7dDDrkOTklSgxMCERkRJr0y8
eBfYaqtxyGAvY018HVyO8TOpec/4PCEZ7SJfBrQkcMhgvj9EsKj2aRIPDDUhylA0
0c5iAYYwk9JWmGfUgmIj+0M3CJCPUlqg69X+QXQXo8YtTpTKuzani60K1BX+A85S
hlDiiSd33SxTZsW9dmNLk1OIw+x2BZvgqGXgZso3y4yRwFt8Ub6dm0CIDFa3uQRf
aQ2ci8YG4BQqEW5zq+4sOYPXsTD+jRHxxwNPwSfow6szcxCYGv5IGJHP4O6BXPlj
mvfzwEPCTewSjcg0EfRHKTNLpwWxLZJTncC1PVJ2KNlMgSMmMfBQLLt/W9yrFrJQ
u9jVwyssUUUCzlQlkQ4CQ5ePoE1RQaVdHvpLP/3qDPqdzLzRnk2cZgYcCvvjh83P
duTGpAJYb9E8HR5oEXYtj0YfyVcDcd4/qiWN2QoCSw30AzoIN5sVcGjTxS2K6D/g
uHK7DPFl0Cc5vgertpWmvlRWeRXnYSaucTKKdKsojZvks0gCO8/0VgKRqX82Jbxr
u0Vey1mUnsZkj5r9a+IdFQ5EzXsR+LA5WEv28VunufaLtSpB93yKDRfeJECfHtqR
ABZT2gxoZ2cVQTqxYy8xW+54ng6ffbVDPf2UVIAjC0Q+v23i8Tfwd61Ikal2ElX9
qaEWJoF12kXdKDJs9sSuq99/T5WeYCWRJ3nz9/ihTFlHn5cbADuWYvcggsxlnzIY
WBZgni7mJLxEG8jhnztaAZIleDe99AESp9lwjU7w+SzE7sliRuIlGzBONHrmTxVt
VogNThADy2zh6waDdL+hroGjIhSGzmbuB1JmLIX452/AosCEZxDgTlNqpOUIL+Hk
vICVpfus3Al06Jswm2kUry2y+Tq5s5WdK26FeVh+zSI92YRCoOshkwE6PTsVSPg6
eqOQK8b70hbeTSvwvKv8rXwF6PRvURHXJ0uezWbxxMj+xsfWHqcpWDMxG8Tf0k3m
aJ8vrrUtbGKTW+P8Gpmi8uRq32XkkVwVbfjtH9x887V/10J7KXUP8wI3P7WTzprX
itgjZ3l8HLVMhK8iyuhdsMpq94wts4CfEBRRUSlwyGYP0VHQyOWi6EVYsURLC4xm
lsfkl/rY4DWKTMf3VxwRJL4HQko7t0xmPQT9We3iD7Yf2uobXqeOqJRRna/iumGW
sKTwumltHXDOoI7nR1pq9tBFXgtmNAWp+Rja7LdSQ12xRBn2yMoS2kw8HWmDj88h
4WhZyzt6Dy9zKpcC5xoqRxB74eeSTfVxHoBogxkQU2tjsAC61NTnz2a6GqDBB1tY
hIRNd0kbAztgromiiyIjecPAWVh74dVgKRCntTN+8kEvgATIAmrY2ADeHBIUjlWn
uR/YyLFHtbPfLXJDhr4l17xXPza07iiiB4vUU5WccTdULKC/aePAmr7pBR7HA0T7
YOC0etm9qtYPQKGNUTlM5saqrhLb9aCcqSmdEzh4TVcwMVAxWnwo1A6sRbQT1BM6
NhETlDFaW9q7tjRfsqLOkTZA8tkw4wdtY8eC+ieI37Kl3pRA/PCR+rtmuorGcUWw
seNn6ph6rpRc1BfjtgBFdPKOR6Ee0zN9MwgSWUsmqbKv7szZ/VmqYkEn0MjZk9Q2
fmp23uVO1pogDw/J/ZkYUcXn5yUQNt/tj6WwPdxs/4i/Ag/PyLaJ6AshArJCnUdv
apoz115nlwc5Fbbqzvr070Erh453q1BaI5kwxDJlHE2gx0cA+rzkDWZaDq51Q1DX
h2Jm7n2XTK5SpuZpZwmDwIUIwzhTHmbWo1eGg7e6zWsVz+P3hdKmW3Ykdd4VwQ3C
t5Mlqn/te/PqHedBExE2ZwZVPlZqdujtbaUbx31WwIiZIma0YtuEr0RhDGwGlIbD
zO6myzsKSKsf9RpGH/wi+NB1VgPUwbNBQd5vO8lOQY6Q5RXHCdvOy2moF7mHkESz
ZFDSrIIioUJlUhtqOvifsQM+fwA3mrUlGQcdR6skwp5QfzDfLlse54mM3kZXGzCb
kEisbjm60OpuSWb1Cl35SdkGvtkGBhSMee/264DE0KhNrWrdnCkYAXS/jhURlAbZ
DTvXRTJ/G496ZGohgORx4pefLFR14juaDIv1aISldIXrzxAsNzY4v0vwfCFSTfMF
UzjXjQn0lhu9QCpriCGQivq6C2BEAFxvlabUHI/6tQBBCyDkz3uXGMb0EKV1jgg1
SQ8NqxH41elqLRH45SuLtWUpduLIdwma/wTklT+lNcaw/8ahBLNYVzNZXUgrU4VD
DRjXhahDW2o9WrvStI++hLYEqr85SpZMyNwyy1lu4WPtefE73sEfz4B8V2AKJmvg
fqWxs/EyGj6IPltDPoAqMw7tElQFnnKj8AO0M9lM6KLeeItsEu6ysCprDKIBOQER
wgHl/OuWfYCC/VnDMv+KOKIXBWmR3O7h2xJ+3qgazSG0uQraO+hd6dP8ZSzspY/2
dJGNoUOWSDiayeJL6PUU1Yk0RBgw5Q8KJ0HBSuPzhwE7OWDDhG14eqdkrEejwhwr
QzOkHsGD51Xspyo83Al/pEjd1Segkc5Xm9Ou+lOsSc8QlBlgawPvPYoJjudZ5xW2
ZmRfQ4l9mYn2OWaFRwFEk958C+RWBzUOg++jpJmBYQQtq2L3WVJ5DBd8OX+rEcdS
Z1zZLwmawfFO1oeF4go1zwxnJQEs5o6cackNKQM34SVvaX3ISi9uIomCw5RT70U0
gmaub8MN1Tj1bbR6gXgPEdeKUECqWOOhnvkm2xcdmPV7wxKpo0SWcv5CIfjjq+VH
BQmXNA6FCx+59iXq31DhO+SB5ySlW/gIeEwJCUdsEVaHX2+O8riDu//A2Y3gbUd9
wbzfEQkfOt1DRl4b1/caZhWi/qgDsmCDuQgvngOMWXJDPbFTYZuVVHmltjNWm34j
W4hBA0LaHURxlRWP9LUXPhRF2Xs6eWYJxdlgyBkfG7IPzKX3LE9MCgdHkPzfCQoU
G0vIJesST2/Mz+FPx/S7CPHvf6gMZiMZHvGscQqXZblq2pk3rGOD+q/qdbVNUvDQ
rVMUhKQ6Cj6FF/K9ddsYhPqSf/13c40VXyONCmAIZsm7eWdM7VFM46iQCDDv6/Z+
ObeXMVP6qzLHhEyQpvn+4Fe0t7WsZpWgEFAjYhuNtsW3e7fnu00re+8CGWb3kg+F
JSkv+Da7NVk8PJp33uUR3Q78lMszCp1lebCQ4jqEAYbcHB7H1ZJAacKKzvohdtlk
zvjJLPFtVxlIHZdG98ny64mVZJ49kzjzdaAwV8ccUtaXafPARoGXXtNRW+7h3pYn
AWpmDkGEJg463uDODkx1xM7QfVhi4RvrmUkWZ9/6I+STvOnFThUGmOqYcGN83bJM
H0zhagWrHENNiEgpdLAJCB7YtY7Q/5E1n8rG/kenG0tqoBWPrrjBp7+fLhmF0XUw
8G9Q/YzgUfL+h1xim9Y3/Jf8CbA/IC2sRIfrs3ZoWYl10f8feU0pnrXrv4vkO8w5
4FZqqSzaWrc2JLj6C4AvOo2U54Za30pt5A1AARJ9QMzpzanYlCTvKdiMyHBKXTA7
nqDBS7v6+KjSM2V1/b9FQzB+GkPdOjmvC3BKMxEadyK5/cWAcgHJG/CBblAR13tO
w6cGNvOwGGpi3IBZgBruIeZbgXqFlu9DOJXKo+r0YyXwme8LBE8KBr8yNNAofh1s
qvcX8HTwblvQH9CDTt+4O/83K9hndlYouRLsLaRdgrQzCzGyQSzF4IhFrZzj2laL
ATnuumXGgbX/0mYXfJho9W1P5iplHJuuKnXpE3Bbrld4V3vsGlKduM8TsSqB4UIS
dHkK4Vjt6OwfXWBzmGC1V49qXPagCejgxqKfkDu+KEXQE0CcwD1astsVvPFnoGOu
FvhbSiDpahZyXpBzmctLvsgA4yrW3oFNhS1mhJhB6TNrzV5kVfu1JwTLF4NeZiCg
XrbXZP+ya8ZUIg3YMjesQy3BjxJGVEYU01YwchOlhv94QDsDFXqKg3aQJrMZRGZj
TFGL5Cru3DzdlW5TKAnA42LZnelS/gfHX2AHP2yEEQ02m3lBkkMJjhEzscM6Fe9h
45WppXasq7oXeKPZlL7wK5RdezoJbnfSD57HRUa1awISUoMTogwiR3Vv34O6Y7Jq
5OotrbLMg9oJB+qda6XrVY2E3m/OhUah1GXDHYEjb1aZPRGa6u5qbEmKBhOgDugS
+0KYu9srfqmAv0OUB0Uvg2ZP6RD2U2CQxZAXI8MUN2FUCKvjrBZGCJ9Ume7rxDZF
aA2g5F8n+RfsbCprUmfAPJyPNHew0hb17O14FS+NvX69mpmzE8F7DaTHfr/0NEoH
1fYjvfIIlsW+8msYPAhEPdzenle5+g07Zp5wgLJ5QvknV4uZhu8KoQo6v8PEd1Kf
hippmw/T86gGAHHytrm53UlOGSrhvaBS4DgI5x0irzk0YAn7wocR2Q/SUl5Fl7pv
/nijTwwRiI4U034YXBcvAWIEcKOCJwkar2hw4BKXwW3dKzVpc+uLcTM0Q3iUseqF
yuJ8CJsEZHMNL0egXCTuBfeSRgE8qoA2lDWqvTQ0Bm7ot9PC889ukgnq3MGDRobG
myMCStn7/W1TN0p0ILQu8+pz4EJuhK99PH/Cdua6BS9EWJMQNRVKGJBb3422GoQ7
b9JV7UuFuj6QJ3xfDVlMG2wJLMrg4dUJ0LXS/ZlZELGbev/xvXP4NRKeUMFEg/47
QNcb2U3Ldg7XjEUQ6uFYlApvb+m3HD8Kyv+Ltl4mOWO2nx6bq0Y3EC12t4MZlE/f
SR4xjc6TxYVYzRXjOwgvJxr6/lvSP68P+5W2ZWkQ3nyRDCr1uE3w5TE2tRApz/fz
v3Syr0yFWEmK/HoUXA1/9Rk6UcKwvDkRYgV6iKAE2PE1JEUra/euq313+LGXPtPG
+XLiUSMEvVPw2NSJsvlcXz9Q4aUJF9mMSX5sfrGJbgG5EkzFJgjdrJBO8Zel0Hjb
gr0tgdHXdXnZQyzR4rSK1aR88ky60TXtvd9sE2sYfjuHfC+DVK9f34giJ6k+Ptv7
4zCVgwr7qGlX9N8YUUZy/bWtv+cScwn6qnu1xk4maioH+lQYyD1k3Y8nMkq1KoDF
qsZYNiL6aDnfvhgPkIuJQQOr5iG3fKAqn+H/eID5n+G1OGJLIdS1pNdQ4+ZT+W6w
ULePBFx2GRLV+ILxTrt+zGq8KgdU4pO+rThb0kCYsE93DAUfDrIrNJPoMmd5y1qU
Am00saaG7RKZF6occ4HJiJnJJCf8IQv3PdelEcxg98XDtbRbWxL70A64cirDpssE
7AWp+ncTJnTPzlthDn3xnFiu3bTm/Vhe8VSDaanM+epg1fLLIyfxofl6Hj7soRIh
C8nNDth4qqY8BHUVR1xoh79MQqy5wdlK0yl9t8wSwEl88HvDxrqvY6qkVrQ7kfIH
1jh27znyWfauTBTrIJG1FpyXFYX+rdOR3w7DBDm2/hwJLwzVriAsVxUFEItNmupx
4DZFPmCuwJHOlXQxBrkU5XbFB3WABuLKY+zTLhIU+cVoGuHSt5wrr2j3jxKIZbAp
fmVd1fa+xABkNmD3kRkl15aoRw+q1XmWpc9Z7UweurKZnD2wWw/e+Q5X+dqx9YQh
gXacKtbcUpVIitjYEkV8ShktNNy1+FxTlQjO5aVWH6Ia1K7szeepdrZneXlmUya9
mjD+RojcpxPIUJnt1oeCNXeTez/q7sxmN8E75NvKuYlxVb5gWxwME6Lsq9w28iYw
BiagxuAKbLDbhgOSSZilpt++UAMxq7vuTXdTOvOFwKaZSQcw1MQ+PNyAohjF8KFq
opd3E6+8ybEEJJnMGl3LGBRqCp6ms6ujJD3JCEKIwhKpdXU5osl1hgHGbJoQOXyI
fHOvhn27ToisInLzMsi9MgRpTefTfVZwCRHgULn/CMDNHH/UgHE1tMpOUcnbIbfl
uz1TKeKhd05Kkd+WkOpyyp8GfBT3qWscaJ1UfQjKpLVcBQZ0KFEO3I+8N78GgKLw
JpJLVYYfQqtTYGYHfpeuRYpjvdkspU/c9+y0W3cG6ulIARZxyXB+uP8z007B9JjP
AWaz6+VAMIhfWrRndu0OUme5vtl++72lkp3x3hP/PY2frhd5kDXF3o9xxmZ0zJTe
fsHsRfWDdSj4AVH4hshfEk37gCapCl8ATb3Pc+qrWHPIeB6geeN7WgQHjeRbJUbW
v8dTooZ4OQJq/cBPFzq048ewBaGsAGksJ1urmz/8aRGsO5PiplbmVq300JfZH56a
sqCjzjCRZGk8/r88FvUSisvcNmL1MoNcH9dwZ1kxniBxoRogtosBB83PptFWm0QA
HwqPZXWRKVPYcG/cth4uY+qt7X6iRhs1eQ90mogbHzxJ8QT17XJhFf3HPQVaIjWr
FjNKC83C18o17pA7Qgs38UnWJdHKSRbo1X46zFtDhBv8u6Ihk4FcOhE5tucYrMtF
w/FdO8sKIiGjLRIPYGgJ+MK/gHkkLggg8Cd8HrdvkFl3xkauSx/Ee8HO8sJ6Vsxy
bOpnNNZvCtTJ/HdPbda6rmIFAhWoxmqbTKw2zOfo7zdzeMlFzHRAK3FrLsKJhBwq
0DHutgkQSE4sg1wkQ70gvb2fiXrW95frQdrEAsffXQiXX8l/rTF3Gj8OwvN4CiCd
KLQugBB3+XOQUvjcN8lLRp14ovJ51bSzyZoL5h6GwffyOJrPBwDTXtvETuD4zHiV
w3MHQ2QLoV3TpJgqHuFP+mDShdonH7osVaYxSTYBXJqKlAQgvLFEIQXSdQ2BEhD7
4NOhqQTlZKzZxtNOe9oqfGMrQpvBa7WfupyFxyGNmpzQLueNattGSKQi3ZE8K3RZ
e97cpgdIaDi52x+2cGrve783DgW1CuZNAi0tb+hrpphcGZAV1hmw0W1bgdc+wYNH
TSM7jh6cmNalHLk3s24gWnGrVLzcO0VmrvcL6NJmODreTuK5NOg2UXXHNEL4vvTq
RJVmsqLlVHwyW0CiOSXxqZRaDpI+4atO+J3FDK2dN8xpyxmKOoBhUtXKYr3fEoC+
AwdWWqHDp/1+xWvVPLg1qwh8a4jUOZ7NLB8GpAJEv4NgzXD+OvHGSnWggFBVZVv7
/ACLpLNJFUjmRNiGABWlgpEwRmPUnwp+StKTePcOi+GghjHJww5OLRj/VkBqZqFx
cp7J5n4NljAgyEuPhSuKVcThGNVepxyVI+5Ua9ZsiRTjPqTNvFCNE/bqqSvD7WVE
Kc+wTEGFh+y7JUtKbJ0R3nId6eZoFnDlpvc8GSyD0+7BVE/1prLXy6hogAycROU5
SqjTtgXuk57MHR2pwFbs6wBuOtSQpULyZXvFJBHlrSRVb91/U7ergWol1dvgrWQB
hWR4zDRWTNXuDf8K0RBPcpKNWzdmhSNnAHwlBvsYKoeirP2FcZhR458VYLEqaIvY
glhw2OjCmP3Sc7oIFndX3UmdA3ldukw5pa2TX1bTkiWJmUmC+0bJCIuS3cXUuF1i
fFwgIu7+tfRJVC1tCE4LGjmNUXA73TwgTZREL9XOktGlQG1osuBH8nuDecGq5p2a
/JbQAy4rSF2B5t7nsoAvy2Q601BU4WP4+t+igJc8z8U+5GbukpRZCKZ5LPWlT8jz
DTxzxMYKxz2JTZ+I+8XtQiKRCHWtsuiKxaAjaPPFUOY9I9C7rHe3H6byzV4J2zhX
Wfit+AWF5e7Ixts7dfPyo81sLmFBjKUhX3E3A55Xsn0NvAoHGh2Xa76S50ofdOiB
fC3StIGxsZYyt+5xMoi7VPsZFNhZqZa/hCRMEtGvDP0qPJXLVJOWJ/1WnEhmSW2C
2OJAQcN7aB8c8Amz4zvuh2Y3tzkQ+ftqW9nfgYuNNCEqc9BoBGjqP1Rx5/bC+ukq
JIAbGPVnTW+YWSYvmBtdGAp8rzOnLZrQmfHthH2kDmghOrWpW41HWZRyUXHwYy6e
n6v3VWBckq8xQxGJX+VdJrdG8VA/s5DgDPi83739lNUWpVICAa9yvBAcD1GXreLS
sIy1rc7LJGz9CohXGkUMEsAmpBQ0EGJ5qY34c1DciRx0pKjyuAQRZ6gfx/TyDS2G
WOiq3KmpgSdzN4vkPQ/jpRleEgHCHXzy1rImyXRWsXLuYDLXoenhDb4i2kk6aI5R
4NHOqILtA0X76GnSGcm1BNlBRHEGyhYz+pSLOmkYa3f7ziVa1lmgTFTXDC2C2Vet
SI10CtkdyxcU56PM8b3CG+BZBzbURCiDlFYy8dY97rgs1b3oyMHhWpMgGbBMDzzx
4fu7RdP5z5S7F7af0RN0nXy4fTaaz5EHcTl+8eeAxrluDWsnPhXbx52aUePZCccN
jevpryUgTFm0NK0WfGyg/gayuUkN5XSXKflgIh/WFz6JNPZluIcXVtK3Eil6ROej
WVbRbUjRA7hWP0vW2rGSgIMDSFaK+dk0MVs/2IoRlenmVqDrgBGJH3jJSjUl2YHx
Aqff0nNvX79CvZxhoeyhr9A/Y2Lctz9asew2RfjX1SKu185m7kW30K6LMK9if91e
LhMAfSKZoglWnYUDiIFYaPG+6Ah7tehrSBUmHiV3XPkzxUxPxqPe3Ruh/QXEZ7QB
2n5XHtyqg9rZsD267KItcwmhLf/pNP8hH2xxGCEwNeVEUuGoVkYLkUTFcLtIMJFW
Hrtxzwperx5GkPLivCIWMKu8Fbj4hjJTzQZwb6IA5m5HFO0onm6MTX5o8oOHoHw4
vZuVKwOFBY7rhcbXtyBPbhdSVIVxgAthnpzABeoyDklJLu5IfnlUTkmzlJ3kJUY3
0RH4VxWVSjbvbtnMC3RYkFMhJGioWoo3VWLHNCzKFmWLNTC5sPrKJMHtF0yf7mfN
o/qQJy9/H8zFDrTcOh4Qv9Zx9OlR9UmQFYcN5z9Q+OK6lWu66WmhdUyn4tziBhsD
k8+4j1NUAqyzTt5Wr05My66kUzw0EcKCZoYoBc9qx8TXH6tbWMYvRcbTLIZ/Uf5S
+7XmlYpKtX+/eY6n0NjRD5m82O04bmLfVnk5r6YeMkWlOetjEaymIVNtlwH5/6Fv
d1H1YD2U4HdUTuKF5ZrrTHf2D1hqF2hKVv42w0Q60hmr/J/f0zdUGCDKnKKXrFJQ
4V2aNiq4w4jN2pDjE0f6ArePPcGzbP4KSpdOEsSRtik1WUbYLNHkTVOs3S2VctY6
NZMsmdNj08cIJaJzMzNQm/XKjjZthrm8uKqSUxx1Y0TQwH7EVWyngZlFo4G5HAN5
k2fBj79ad0KSs3tu0L3vL1X5sEqR6Hei9LU5EGXnkXZD9xC8tJ97In7QpiYKcVpG
EOgsrNsaruQ9QQ9+t5NxauGUPo3YYKz1phuud2QE9Ao0bTvh0hyXIDHRy8uw4USS
ZmI3QAR9PkwxJu6ONZ+w3DxZ8c+ZalFRhrLYBFm22KsFaI6JQ4E8wdK4evvhvEpg
LKQhgcCX8oqkNYfMKpjWfkK5KAION84RZTCNKE5tkn4uvZZyVjp36OtB+jNhOcMI
Cx6zdbVAyxI7pIjf1Zuua+lWt1+foeSaLabZ4PDQL20tXwtigOp6Kg7TVzvaTBC3
OLeD2H1HhkZHrWlcJNetStzNKaonVfLUy16WOeJzdpXsIdCjT/nk4Z7Rp3TqWXjC
XjjMIws2QymxJVM4NxiLAhkrA7hIGyZTeyxUe5IHqVWKZ04JF8tLGvDaNuhOoK9o
DR9hRAbYLE6Ap+SWsCrM8h8Pi405aeqMK1ryriP2GsAK+bXRD/vi/rixj6MmUTmT
kqan43/Zdkgnze5JJHACq5g7oRJL/KLT1HEe3vjkRshACfSBrA9fwSdtqXuhEEjE
IMKr0zE7BRXKuQM23YU5Gz29fLYK3A1uRNa9TC7d+zA4RZfaQdFJE8ya3aTY52ZQ
2TfyCbrE2aisUgcawU3u8zRgVssxzaM+0wcUz5Uvnm1q6g/q9bK+EP1y7O20tDU0
qC16Yi4hMmQ/PUXhtzZktMbXgTdUD9tbNB+l+2R1YJN0+mbtUCVHXlgu2ip4UDHl
LOjsItUqjjJU4HiD0bKcS4BuR4X3dsuYuYVsq5pyw8L/p+Nv82tCT3DYCzxwnUpU
v+ajbJlewYZY6y3TQfNlECS+gKg3NJ2ykm9lnAxCuNVuvTGssM77ESBoHmhQ5Rvb
7YjTSnRrgbUx3v7jMFB8uRcB7TNuZYH9iAAWUwV0XZ1ajbTdOLQmPj0OPSvvKVWk
N0x8WQ6I1ATBjkfact/X7TVtxpA7j+UTLNEXSUftUD4M9AAfmNs7PE0TXyrSJ+Sp
+2LuKqv0tpksIeHjsvF2+bARVDWOREz5UnWpchiGAE7oYzr1V5SgFj4ZT8+a/51f
/GQzViU4J4aHBBI3ZCYiqnttgenMcWq9pGOwY6emYbw1kZ9WtwEl/Kzm3cKrsDmU
pGgiRd7qgl801HsO+3sXfbPKxDdCnJeAZx6TDxQ3GPI9/7pxDcf0tAaeIJfT1wug
yyzJsJy4GG4ioyVY44nEnX4kaBOXAxGZ4SL2h72FVcdUjSxG+eD0+Xo+ouB9Tfmv
1H13Fbxk8d0QSoLCCKY/IE7KU+3gEheweUsrT73EdFhkIzmUERGbqBehr9DFhGTg
1iAaXHrXjPwXdo3XaJ35ys5y7Q8MfaaOZ9M72/nIzaCGvZz6ntRNpmk/GyURI6bt
k/xdR5rIbtMLIAQpqBZWk7MzyEWt8A23ZaQZleOhNjJn3j8GZhrbqZeJxHwyQ83g
JArphE3ynLkxAFS35BY5kBPaVrTGfN7ZDniIQr54XR90A63aHw6IasfMl+M5qif+
8PekAqebD6lJ3pPrMl2uMunD6zVbY/H29Mubt1c4wwbO/89uP+FpRLY1PMvTe/EK
0kSP34sZmaTkvliLyVK1OylzBYQxy9pLTjT/fGC86e1bgkNJh2Ln/axOvSqVPV7d
vYRY1KOzC6FJe77jVufWZ51FNtCx8TjChDpb6/F+O0H46HMSFVfCyVM6h/LcJmGB
OuYsLJhPs8w15FfuTC2RAU5Ht+gaIaKfiJgszsIq8u4v5IgwH8g7GIRlJeIIED2X
70r+3nKUwEYSy49bbGltXKSMMWcKjwa2SopfxvJrHW8kJ+A1r/8Dv5R2MOS4gkh+
ELZB2AGBsEQivEZwXl+PSg6LYAYYNb9w1PquGQajKDECb2aOfEcLdYOJDejNbU2B
7QbtVL+uQv2umPlQTqzMRtkbTvX4koIA4ak2Km+65R6r5NE4OAMURfQxxQJUW5Rc
2pRplQ40opk+Hr9+IYAyiobkDg4yJUrIL9AD/oTV8bWQo41olZf0sgUVjaboDjT3
TscpcqNLaMjyHA48FNilIhP5Ql7ufTnwTJRbBzhkhH3cgU2UX/zUrmTpHtzTdlo5
AZ2A1OTu9WkOb+FZUWsX4hwOSiffbpM0lpti5Pm9GtrnjukBE22koIAaaluSGjOh
hAVe0V2zk+RPR9nBeH64PWCIaSStRWW/fiIrYZC1sybEoNxxz01ZJ/mzt5/thtYk
tBYdn4aDFCWUmhH53Hhp1LkhuY+oDB3bJnjG7hM9mu2aSDkGOCkPA+YDzpPriZ9G
lQ9I2BG5BxMCTZ2yDOcalczRt/xrj+tPfZ/L3EjrAHuA4S71TWmKG26TT1bWhsEh
LjJ1hg4v/BUNtttaU2OKR3YoGPWbGlzTkF3JY4KOEoMg+Byk1mZUf+IFIVH1P/hA
eJY7FZEWmoqUsIr2LlGjllyqfcpQ9pWAhVUXu6AYMYKN2y3mIboYGU4IUYrNmsl4
j9Zw691iWRUCFGzuQlKuQtALVqj5MQSXrE0q8UGD1g6xurHNb/eU9SMeaDjL7fcV
2hCjUE9GkjxcmdqQxDnhjJ8XCxJh45o7m7ouequwXoVMvaT31AxLGPzX59Q6JCaU
cWe1rPbpM03SaN3ufCx8wsH/5RJOAZuNpXyrIuRLDsdAF+KobO0KuKVyc5JYnaGG
fX7LzS45FsAQU74IzR5zs/j3xwrhVbtHUEg0TpYS+UIxPTw6Q8mlpBxBBJ4kfNsb
G2iYbZzl0OOe2r9uDOCJOtKGXHFumxDro6VO1/zPxVOLXjdkMkxHeCs0XiQSgDIr
LMWt4Iqu6TKyNd7Fc1xO+BejBZiXgYXrTi/zGvSi8cZeW0JStXapVm3ItxUWhFCC
ci2kjT7HR7f3e6zlInaHEdEywRF5Kr9gCC0wN2DWEtW3j+Zrom/CeXbZAOx4SF6o
Q7aPseAxEalavUnCLIBqjZFtQe/KzAOgzUgNLNQ+VePx0G91t5brBbRzc4jupxVy
MSpyMjqwHAclFU2Zzymg+tE9NuDGgjqCwpXb7bz2sA8muhqmNvjhgHvCBwVi/MBS
UkQQacdEvWQh7CFXJS3bcMcwtIB7tgzAB7wJQ+ZgryU46r65mOFQy888su1X5dAe
bd5tQ01DjG84iYdLhQRYuzH+lolcE4Jdmp4NFVU2EDg+qsyFAzn2+VV36T4F/VML
g4ADm0WPmLHk3VaS6ZwinEV8oCJce38VYx32TvjZPdeUxOrth+HW2mlIM52Ooz/6
x1swYQorxagbJkDDtKxl4f2HQ4/hpXeg2JUMnDn4IwVClu94T3CUp2Vu9saxdbKV
y+FPHHiWPCc2zpY/UZ5iUrzKiJSMK0N3pNkvsbQbVrDl3HutTwNTjAQMzdb05/0q
VSArmlLsZovcblSKx5AXlvnSRrt3p1uQcFHfZiqRdl7ZzQOp/BLpCkZJuUXb+7ZN
/dJJFNw5/xTXLHVfkM1DudVPvz89ZETSsZkkYJucI07ToStDABhuDX2MPrXW3J+g
TCKf/8aFhU5py5RbZ7o1UUOElsKLWFn8+YQlglrpGUsaqcS7jse/9ewnn7aDa1fY
uD14bcCTraHKTKm2ENjNUJzVnCS25/X3VpoIFcSN7+KF6GNSFrs8dyIenUvKzgeo
yEe9UecePuvBZ6Wvnm2XvQx8k++0n5o13vpIIHxnOPt8hknvJb4RFR1MbWnh7E6j
f3wMI6rilUcGpIKoXPkNmSXmN4qoktImYttyE/jCv85SDlgGPPbDMdw+mb9a4wMq
immi/6ERI4BAp8IomKDh1NCc2BSOCh4abQnQWd9HQtkL3Qb9DmdEGn3fJlo59KPA
uFjLcUKE0tAZMPekCeEDjGrERPMDLFxXBKAojZetWDXqv1U3RHYooXWcItbTW4dV
0ArYDdv3ALg0TqFLV38ZUJAnBkZQHLwJsekkzwP8Pj5pfmcG73IVE2/zYfjJEm74
KYeQ/CQcYuEddx3IZyXoDx2rwrrhM2eVfzXSrORzD8W7BAZ7OKuuejHjz5CT5v0K
NNcsLO/5gpnPQPqAMmy4aQzZ23geuOhQ0iNQ4hpAD9XHONK0ZsboczHZhVdXmuJD
dtaPGfHp43Tl1WkzsgixTHkKbSdJlIk8JsSQz7dmpUMLQku+rj15+3x0WmSPd2bR
nrs0DJ83Ihk3I2w2JlaNogSiQdULlI5nYs8WUOYkv5J0X7dBuPUts+wDAQJUwzgZ
OYxoe6gUKaDMa4RiI+LGLUcxT7yUNlNce/6cNYmgDzJM8mx+PuDwtE7OuFNuBJ4Q
j1JBsM5hmq9fiG8EGIYj3E8b+w1/W6ZREDGj55u0fUpbsBLnFxbdibuA/OdtzIc9
xKYvsFmpfgMHy3Sxf4pFtV5IbpetxSk50/gD9h5ie7aTu06uVz6KlrUl3bHVv3X2
upp04qh+LVAYhZ6UdAr5It2uneL54g8gE31yx5uiSyZa04qgU1O5lHW7snZPDGUR
SFo5ml18HmQxyRuvoBVBXt2pVAoBhzuVaC4qcBmGKw4JyvJ77BxdwehGQV9CS/+z
01g9M7/ts+yvn1k/fkwIGMG+3wfT9KIeKlio0vXt00Wy0UUAiJfeyMyI9Bq8I+Wa
+mH1vYCh9FTkke3vr2W55TJuVo/7FtrnpLYaKGWpanqMw5oBld82Vut4j9TgqD44
McJsLtLTuwHGjRn7UKzMXQhdxk6oYUaEEj9YBMwaIhGGEbF2Eu3074sqXg3TMbZb
zHSwr9HhE7amqlmHJqq+pQzOh6SQc153EgfVScZbm7dUV6wXVIWlWmFIRAY4IHFn
Yl9mQDIiehd1vDg+P1GZBx6zOv+mBP289llDxb3XBXP34YcEbNinzSG5kKSRPz0S
6zFm5WholY8As6D3msJoTkA2VOI4VCiAT3xLaCd+Tc5NmvEq+s+25dAsOjfzucPD
VronxyhhHERIXe20nARPBp9WoCjNtzux2PMtvgn+H/229rUz5LE8OZTUTjmsSLd/
JlOjw5XL/KIKFb4RH77cFSsnl+AWFLgI/V/ni+yaMg5QX18vbIW6vnogQNaoGY7I
Wg1B6qX6D4tmxxtPOXYQYjH293st6fYqMittPPQDqlDiEZgbYscL8oQOOT21yRwj
hzh86WUoRNMGbGT/BeZxiSNtAXobYwOuWzFGfgn74YXFtXfsSDSOzlFv8FnjXWfc
0jUt2KmeIx/E+kDp23Wums7cl1Nz9o0xK3XtxIyp4bjPuJQgMcs6msV0TGwVnX6E
yP8JNIaOgJzx+wFkw4vRCXVZTRPhU1wga7sKXiOvngbIALZkvklnKUzB99pKiVM1
z/VQwD6Bu5ldJu3A+FY/BvHkM51jUNIcva/0WBuFaRNQ3sd+47GAfcU4yFZ6/Zfb
uCG9xnpKJaL/0OUKks/vWbDEorfLrrMnYtEDEpewwOoos5lbjlmH5MqlFjxv9+MM
dXR7KtpqQv3e9IYXLjaOodgP7FITPlBu6NtmKzWhhyEp22R0mNUq/c+CrBZfKN3D
0z3n7+P02pS8t+ZgODZZBS3gc/iCm7uLktRQ5/lZM7M2WjY4nkzdWMcJM015igEd
u4Rdz63LyVCwvWpe0eyINUYb10oR7Gyu2cvzTjRqID+wX9ZJK1kMvHfBvzraHS85
ZsK6045duVey2/i7ph6mUXToW8EAgi/IJDMXdxLYRcj66/FK2jBIC14xpPDF4eal
PvTFj/53oUxnewEsRzHxyj9JeevLFM0fK9TDSmze50B9w/8F9nl5yqgFsizYvKT5
gaBK9m80id65WE6RlP7HJEd5K4GoTvhbgsiDzHiPp723r+ZZe9LW6b3GKC9FFhaU
5qzqO/7eHsKQa6rAMDNbEM3CJv6VYpz29kDiBpUQNGPyFTft7S8bMlHPqQ0eiJ3p
q9S2q8snUE6E7yDUFwjh3FalfOU+jqinSPrbgKX3/ufMo9qztp383XJ4fqA6b1v+
UCNdSEnZEu7A6wcbyat0h0ZIKiM97VPdDr9xe6VhcmlpPrVDpVATB7aVFvvt9uSy
IwYWmRxZ7X3/Gzt9TuRQP7hLUfQpjlqbgdlkbALDuWknIqIr7U1HgfWJTlPccXTj
fGAvIpPLkriWOLzsTPxnhGJMEIM5Q+yXZoP2qpsDtiYqoDc035vfXMsXqpYz2GHe
gbnpHJCRSLF9GfUc4/tx4aIBGbpqa9x+5pqE5tWdSj57CTgnqA/GypuS0BOjlLIy
rLj0RK83EH255miqMt6M/VIH7a8PkUfxMHkpkrXmB7g4Bu+3XxKrDLjJ834NCwMz
XoweT2J8xXFt3Wpl6DIbZ9g1WKw3IGKafTqred0iNpbN10wvB3grNIvF9UthlS1B
Al4X5XRxrZLZFSkeqpCgYgEYHOwcx4v8+3Prf8f4+4BIV9ediTnHtm3qRo26ToO3
ZpU3RmW3xFDa7XhPF9N9+6TQErYra+QAXLHOAdOT/Bb4fwxvkNqkno8j2pr3cb6J
+B+TYC8Nv7QG8m9CyklcCqMWis0gpeAOG7L1uxFeYyIzgEaDxrhFO/ir6SDm51AS
KCPp4CbHZH7rIVroCP7AAEBxbuCd2IgfJ3e2cBvgsUYPXMPENMz40Z6U8VzkhjVn
EwtEVvlNkbyeMdz4RZ3sKanYMC4WvrKPA67ne4cYY9Al/mDLG/Ss/DTpKqMyliSa
wElaU3LgZgB/XKhxc41QacEYZcVO1uvG4qj59NLNR84O2YVI9dyS2bjWGUja/5yv
uWESQ7IgQ402tdfUC1lUuzn/GW7jMK/0B//Z+Wg6X6vmgeNg27s/mkLLI8dAM3Vf
Bo66fOf4r3f1XKvI3xGRvMkyw9kjVyGqT6c/N51rl+wbhA85ZsVgptdIwLAsRZiG
zf1EdTRNzbELXgRPHFc5JGwoQTp1t/HbWNmhdXZBbmUStUJPRADyYJmtQJOJP791
YNuQtx9RR4gqYTl8baVCn8Ag7wDEYlCOZvtGGHjYlMCmvxOCjSYdSM563OK4Aqag
2XzPZfs9APQKyb0inxqauhuD1zILlyRcAt8tKnU/6PjzeSj5Yt+WNw4Q/ZalqkOk
gfiHFkV4moA8wmvovjRGDHk2p5S8jqxzAjA1uCLssoDHwVL8yNepgJgDPZgMJ+OF
Liuu3SgTh0be/3cP8rYzCzuliE476jtc+hvpAm7MVNDxtBXGD5l78owb69DKDn3e
oBHH44bv0waV7MANlER7oQe1PsoHEE8z/hdMxAaza0VTScNpBShh/EmBrf//fKNs
4PGVOLLn4ctXreDblLTXm00cILkaN0lErb2gXOMozfE3ZHtVJgtdyxbOwEMD2OLz
JxX9V7IAaBKrOyGZsY2QrjB+IkesItvTIguHvGL/4xXGLiWDSlkPfdT5R+M5C7PG
sxhqFSIBMo1FO8MmeTL/bnIV8thw4lnTOSSjHFK16QcK6S9t24Q1j2eI1snpFdgA
vMLkco0HHIiEP8PiSyCX/2g6iruAq8un7kl5gd86B3pcZ0Jm+xTZIrdh8TIiujjb
qC1sgCUxVIvNFsO+w8V/YpADkDy8dAq6qMQWVQpXq7TIDZHJRc9pNTMmDt1Y721Y
/hzXLyLQ3dCXZDgQjBnwMM3cTIU2P0410gfpmorwL9tDyk2n79kQCDHe95/ClYX5
tcXZ6RCD+PKms1a4xHbWlnYC6USAwcrGbpEMAnUBTvJLSJQZI19bb/KNcThDGzFP
t0MpPtMJL/MMhl27bNSoWUcGL5cM+z5wVIvOVQ0jx8tK+VhosWsOw1Am84JUw/0W
a3KoI7w/9vCVU3jKJLto4BISfdIm00kyYGR9Yjwnpto8ky0bzYX2ZucT/B23dzvS
vkkSihEF1Mgvz+qRRSJ8trFc4Xek5GduCZ8aqFUSBsWlQgdBAQCwVpoM9a+8dfaZ
vW0KWgF14Vv3AFN/nb4rmqlffMmW5aBlBXM0qs98XqqKBS24NbXwNJ+g7d5vHSvk
KUOfK672BNTg4Aqh7qHrVx2SidXZzGAiIEwG8tcTtFR4MTpCF98TB5HqL0SgNSwN
3k8i+yPNw9DUlcM9m9UKTuaZp291hIpEZc3Z4pwIZuE0eur6jzcALY4FnZ3tsydM
xY/Q1jdYoxxPHf9khxJ5gCrnTDy2J779bGcYPz4mSnpjbTZzEUdrClCcpG4DslPM
OTp09XCUgvWYAl1yHcnlaVjPfw6pPNLwYfFgld66KRqcxaXOtICgkH/dAjTfxE3e
HtYXlRQSpPTQIoxZNMHd3TQ4VUMcBe+1r0PgWgdtKsx3FZ/JG38ohac9KHFrsCzf
en1vVOMX2PCaywBhoC/GqzSYyIE5QrVeNM3uyOcXQr4ChR3MDyJPETb1mFk7l5u4
Uqj89y/+78eQbf6A8UKkWmcdyuNnEHIvXF5zT5IwQ1O9Li0JFZ53BpgI5oxrSPxD
BAWBF2nbParS+4wnKMc0Jxmt3YTxBMYX/kCKiLdyr+EWT5wVCau6U3/9Gi2oE1YM
iIV0S8Kr9uo/L5tW4BcROpop1j675d9ape54W/5znF1Y1CNi5XnGGd+k3V7H6BxP
mJBGD5w2H4MZRXu6muv5Jb8Ho8r39Lz49oT8LZiGhmzL7UDWkluErxkrXR1y4kqX
bsBmCxuCHA+6RYERx2tNFpPd8T/Bj+BPowYhjI+5AKzTFK8ZbYj70aEJSK9rGh4g
2RF9JJQkkBbbSFAeQ756x+gdfj9RWVHxzZpLL9D6Jwn/Hj46W7ZEIj17jy8/xXPk
gglercyH5Zo5O9l+Gff6o5Dx/Snjy659tR80jvakuBltpHebaRUb8ftspGm+0yQp
rKhq+gtkrqsvZC6VUrjqDRVaSipXeA3GFvy3MgfaLH5ANFWxw/jFcIJDfrcRfGcR
O9SI1lIbxDDFChe6+ahGNM3XeBhnjechOM4r0iHRtAHdCKFkfPqZXz2/H7jzIlah
+5+Bb/AmbtBojHbntnCO+gHqtSZCgsBYWz2+iMFUGSLoTyIR9d89Jeiqe1SZeEcZ
r/MPWSRwAjJs8HmJMRSRID7ikLYfEWxTl+lyvZ8a5Fl1UXuS4B0jCDvAD/txeXcP
wZbGCs5NURIcu+p8E0O4zll2yC/goSi+KWzYAnjCR0tFxBt+xos5dwpbu6n1j6PV
PXkCGZ21dN6MRWM1+4nmUoJI+p9l7WKwTfsI8fZSi78SCrNt7sGwLk2aepUAOU8g
6Ers/Kzds3G3moFailb4jo2vqc3YeCZUAZVgArVJ4/JKT5F7/tgAuBy/N0SjX2/1
AM2BiI8Miaps7Kq/at7azm2LlboBExJL7i6RBmlNIPvYapP7dRXITlJwK0Y4TXO2
81N5dPcHe3CxPeYqJ0kUV7IAn4IoKEGedn/JDR4YWz7W7QEHQ7QdQ7zqahkcKAiq
GhckLuXG/xGfoC99Xo53RV61SOYp8r8KfIgVKF6eZf1iYfZPEUSXkT8pAjL4FmJm
4G4pHItDxLKavEhA5sdYB3bBKIBleH6NlIB/shTBSMVNGXvafCCkQoEIrycgYR5r
s5q1a8F7b4dyUbK45fn6zVyUmETx4K81bYd4sq+bvFn2eWUEPnS2n77CSHOzYpVL
sQDBiqmPirez+mFJZ3Ic5tdyYbwkKu+YPhP2LOm/SnxqLfOrwmFLHYyH4YIwZkSQ
ygqqlk/TSqtAv47HBovxNBxpljFwLDL9lMzkB3qpsGvlC3boeAZmP2pnbBYmUB6o
XhRBX1KuLTL29m13kt+G8KU87i5vlC4ac78ZIBqHAOictyALAJ3ocVeZdM/cOVWw
c6N/eSnV/2wdUuM+jALzzKoEYjp8SeP50xHmyMPzkjDJZnNe/Dyv2lIEoI3T4mGc
SQ9nVxrduPhVpDhVYujpcubuxwoP4mKH91WUj/vAKB/vqdc/0faUqSjVHzPV9QA/
Rl+wbRazq5bBAW0JopoOCi7gOB89K6iMGf+kv5TVTpz6YQLSVkgcJMwnVzGcgpK8
Ns7Sqar61YhyMrUe/0BMiiSp2UZQZuf/60Wlvrek2/715/8sMV8NmTPJmYFZsdty
JLCH/BbWtzJ8qAVhr1uGyFumB55gWaKUG/2MgrSKM+E5P5oJPtZtAVBm3IqGJ/Jy
MkDd79ro5mgTi5tpT7Vl9kH3N9zVZfpbiMVZd26A57RYRRKxGTacpZrnF0ijlkgf
Ck9wGlny+62gcvNf64CP6hBkoMwG64TT/oOCTwTp1lJH9mMNJhpnP4lGKfmFMAHP
7K21wpYNR58lFMe2cLs6fdqFsEyYq9M4Ih2a0PWBZ5xx3sX8d+hbw0i48d55F3kh
VHFwW0CnpMmVJG/MV5QRLdhAKw1qDPeSJP5mzpn63plwSXYrvGH4E7q6d33IR1OI
+QgpDdbVq4MZlLWJAV1sHVELiNGViN9oy3T4CwqxyuBsF+81vWrf/gK/sFZa94QT
JsVs2GVsaWLqT5VgFSRDAt1ycvYvntQJbcYqors630FTMymG2Yb2SoB3gTGAPRRw
nykpD7DYO5RAooNBPspj/d3rBQR8pE/xwuF+XVYjEJvwsKyGY3CoRtwM2QZGrK8f
+eNrTjlyxbJJilppWCCFTG/awGJKY89mW9fUldNAiG3T9i3xJRY4HXQn3lwezrAH
uj7fKsa2kL4SMdGBJYPsscBCx+VgJwyHNIyvUiWLNomtFmQI1Pdw7e1Jsvy2E22L
1NrU4AjEZNATqnyt5vVSAO759Hm3W94CEJVn7t9IIwEld/NK2WLqRyeDOMl33Iil
FwkyBfCEPNPUenPTlzzrOqB0f9RxV2OkEN0gXxc8tZTy3PKvCpXW0nXEGkZ4XnVN
k2YW8cLdVLWBKclkp2DoFtNzvryBn1b9ZL8tEU71LYrQHMTJdedK7g6nx5qNFGJK
UD2Yowg/ALaToW8oaW27LMRElPtjynv3d7jEcxIGRr4kraV73e68a2038JaEm0D3
/ymdkRn+IBkzc/KMGGXU5rbfgSxpuXHqvfgrqcTPA25wYtPs6ydIsN9GSeM7kJoB
a6d3a9rPuOJEH1gghurFLrVKpVg6UQeobFGxdFWjtPuWpJRc/DB2E/pgK3wztxH/
8HcnC3/Le7UbMSFmxSugfYDOPyz4Zj/avFvrjI9tWsws639cYq9T2Xw+B/C41UvK
5jl0otr1MKAPxR13FwFzYfe890ZutE7wbk0vuhwNiwKH4BmyA7e4p1L5vkt2UhkD
GK9nZ8f9j7xpsxnklwv8/p1BJwBldmhfyRNefYSbTU2YfwoAVy+meJ3k/4QnEhg4
TLIpJu1I2h65JsZnDXNXIvpjHxdg9ZJ8ESBr4W6RnA2kOPmSZ6n8dZ+Nn4Uyjwj+
NYjnu1qvGwzJ9OnMTE6M/INjgDMainF6msnMP+lX+KZFNC8hkXqGrckBXrCwCJVn
sUk265f6rgMnPGfbC/8ExApR3pJMTRdEreS+l1d8euL4p2Dcbl2kUgJty4qtuP3o
geIEw42qC3rlyUIfg0I4sXDF0IYyYjBFzn9fN53YxlmnFY2aMqLT5gM520si7wW5
4q6PqGRvD89erd9cK9pMkt4tiQjUQvGuv+WiMTXq4PLi2EvmGBqmb3AFV8mIljOE
+2/qnKcHyW2Oco0QshP/a4KyS8KmVRnVmenM9PTXN+qpbR+ztswr6jNk5z79cet2
M17P28GGNTv6JQz+BX6EKe60Lp1KUUIka9nK09jahBZ9hcJh+LgniJxCXAhqkZIQ
pLvEnbUyg+T7OFtkjvKQwnd7lTz3fz2PhV4ixgt/7xPMZN0yTokXMGT9nWqfFGQ2
CCtt2X/V0MkkuiU8rhd856u1h7lRfjNh/DyrZTcmrhkYC45+rdY31R9HQe85DBPb
vyhLYHbncq9w6Ons9Z0QpOFKPf368GgyrUWdOb33wQ8iYmO+zMGZ7Zt7xTl2Xdn7
cHymFDdLCnidgCw/FR+UpabvkoTEuDkm7ckik8/XnVtGFRTe3hPQtylU4AmR+x5d
Ug/LEKcKS12luYtZ12QGeXkRPR7ON8l9K0hDepZ3kDSFuFDQnm5HwEC3AgUQKnXD
ls/sXLkb4OSRIguAAO1vXA1kcDcHszAIKEkaGgdL4c0aGTeOYbeMBIGFjm1trjyk
VhZMW6IuUfxds8Y1pHzjlmdQ9VYzMQIgGgUYwr13GKE3GEqo+q/4SNPNHjER9kkv
3WdJrOR5/DAGx1EXGDm1oLI/dHrK2UCxk8F7pMKULgO3URln5bRGAQBosi/Xair1
ry7bhfH/Cy9TSctANu59tem9/hytEckN0Z64oRmmvNVoyeKE6HQQBEUOB6ZgbtWN
KfmPYoIEDZh68+ya8SThCkZ/plAhb1NCVBXh4OYrqgl8fxxZoKPVZWIlCMfrnhfE
2OaLqFtaujLt2bRMT1SOwMhOoZcImVW5xZCnedwRpKa5ZCdDAwBK+jOBPct0Socg
H709HBKunjQ08Q4KXXuQcS0dAudxj6biR9nlCEiwgzSTB3FpnYh2YeCzmQRn6T/H
L7mIUG6BNoK8ZvrYr7JYp3cuX0RneA01R59/Lv1xkh/PCizt6S/TUqAx2GVxl6+b
ODiulLYy23ZIArdqVMJg9jQsE7+U9QLBB5wVpP6kPKUM950GyJxV/ybPRBmmRFiW
ppbWM9+OxACJXjn17ZfG9vaYZY7pDUtoQmbviQPJQx9KD4yRUHzEVmBtSx+V03/3
mz5Z7D1T0eagirrJbA4jizPxlCVmMIj+C+V6SkQsZP3X0Pm0ae5CwOBwkV3TFs3T
4Oap7Tueo8sjj8TOUVwvs8O6u3rJD+ug3XzK3/ivmzuqqiR/AhdEk3tO3nGu/UjE
SxNhgs+LW8EwFny2Ez1e7YLyYwuK+w6hI9rthr6EbVf44LiyyqJHZfQ7sp6RFXNz
j2W06p3HM7YIELcz2tJYjTD6dpCroHyuCQaSacwbTCeMYRSrzZ5kAUeal1sAPLEl
fhdoU/JLTW1q2kHcqRrs8nAcewKD8rUGIb4Emqex0r/B2hvUSgTUZpFe9hRuFb7p
jLoi4/McyZKvpji40Y2DrZVIJ1QFcKoWiXaxXjJjX2Kf+ZF6o3hBQvltymU3E7sH
dXoxfXC06ceVtLFZpgwR0hTMHPp8KlyPMsjc59YfdARLOcVFC8WxEwmj34Aa+FLE
vZhbjq4HmSiey6Uo/kwCd5JnudaMAqx8rdF+lgCYRYOrC98eCAQpHm3+M1twGwvW
UUApwKKAgQlYXD84h6PaFqsJGjUzP5HSfyix74vsCfcEDpYI6awkPpMwOntSN5Zw
U5sEIEmAQ/oVk1HtfQDNrpIgNhMcPnJg+LRec9HuRFOaYPiJ6OImQfkuJO3Xktvx
WMOzeG1+PpRJp5dGxL9LW4Q2JzHblgckPzDK01JEZpgpIi6s7MtTpz68D5r6eLQT
rhuaiVTH4DVp9tRi8iNG6Ex4redc2hf2L4d84SHMHeyrdSiNTlW0PgSlOYm8tncT
19mEjCwf/QYIvnMFxrxJc2MVE8KhGujZq+7ptet23NDZ2Al57hLN4gYNImD5UbWe
dA0ViWpcOKHCnTWXQwl+DbU22ddptTarTWMmE+1wgNpJDWxZRLR4P9i/syOOU+VQ
VdNT1uY9iij+1OPipJg87MIseyUKBRGi51n8HOFlxLi5wwmry5J0NXiK967ukJkt
/rcarmG4qEztvBcFaZQDCuU56+TkhTg0Oyu+0iV0mDrfi8z/mti19/xjg0sV/rzu
wlUsMjCe7RYPaDfmVSjgd4ZMV8s9FStNp2N5P/Fb+MUgyu6uFAm1WSkN2pKwYKqK
ywpzidbF1D5F1OKwPQRv4IyvMG7pyWDqj7bR7R1O/8RWx8p8vqcRdk27zpk81kaR
gD/tBb6WH0K53TKz10Dz3VPCMyRVfmREJ/ry2Nlt1p76zh9arl3ZT7baiGb0KDRs
aiUS5gsUoVo/FhIFmnhvXLwv0I/BQvexfLk3CfcxtvEMOS+KE/uLZeIVt+zEuoCT
KmvKkNNU5LmDNEmsjQUu+WEwp95y0AMbx7vo0Lwa+eUmt8ZrXSl91Sv4Hk6RLEMu
rSQCOseSGUsC7qWjRSoFQHo5g4lOwTBw1ud8zl/TNH0mnphirEoGARRgV2NrjzOe
E0F8Os0JLXts6u+QhlbW+3mrK/A7+wz2es3en81A+PEcykneA6kFWZAC9Jr0hkUS
Ib2R3+/TSJ7JrATgGUiBjR0zNfqX5wuvLaXwhurwkdjaP+5DV5e80J83BVE6SN2w
APwQGCyNfkcUg/2HlcEU+VV7aiqPZoj8rIe/PnMtc8wBb9bB0frCiwfpZkwcoBra
fqVkYqv2XQhbNaGhC+uJpc3sUwQhEtwpPHc8YlRY1Aov7ULo5dNrqmTTCrb4KrE1
naNDKMiMWuJKWcjTnsRax9lMbWUdeJsu2hNTEJfTR452Rmxm/vaLWA+mfJCFAjtN
f5uFZiMitHsB5EDBPauViTBdNeYJOK/50HMEolNwfGUZunJEizAQxo2O7pWZuM/l
PwNPTKbZUJBxEemO7h1YqbQHCDf5sqMHPzDn8yARifNRgrsTO5n6hFTRWCeTqUTJ
dk+S1PSrjh3MFnMm//U4PH3efL6WJ3sFHLYuxAYA3KufMvnMm4O7ChOXLq84Kszv
mj7Z1n54ho5KIjJc0BGNf2x2DTCF4PtDFKP2U0xduPWK1c2EjYnRJh8JcRAVVnUi
Kr/kdD0iKiL1RzWoLTs6S8XBtg7B87sHMTb/2s99O+LlXT9+muhiejlf2gLwJ11r
2PmFfwMX5zH45hWEN84NFvy3mo3wn0RLfwZ61VGMDhjnSEeBXKrm4VHJ8AiwEyNJ
bq4tvZOiz3GoX8ZccAvq7z17nNj8v1NiIrD+VVVuh0QkEdz3OjdGyDw2p1Og/U1r
+B3mkjZSATCnHQ605oyBBqrwN7tV6cFA2EFb8Ep9KN/Xn+4JVQCdRs4XuB98eLNN
JtPaPrYVqOy43hZ6RDcZKNygkFNedBJSrCHB0WqFszHOOLn40YMEhv/2yMTAImeB
MGj2ct8MFDfrtandGhCobnGjCSFbfyKsQ56VzFb4zTK+TPe40o0i9Pmz4Vkhdcha
m02+rdrHXRvi5KYcvbdcRc6/4CuJ/otBJ7cqrSiYa1J9HzAefZXROnUwYZuGmk03
fWYe345cTGwpxzYnG7GPmJFejE/M+r9jmPQBYJ76n0Z46fPfcg1+FQ5ofqTIhnXy
ziiwD9C/nf3ig4Juyq6gvm/uC/E8uk9NiOK3FsVMoMsK5rvIaFL6Yc7QLRxi5ydg
A4Zr2brS6Dql/wNtPMKEOo9IEEAqHm7J85MARriGM207gn9beD7dnOtyWsg9mCwk
mFulT3D69qiUwGkWT6mTnUROpGlTrGUvwJlQ7Z2YYQZ+pmVcJztiKgI7pYML0ZWf
c7va57kLaq1zPOU7XvTgK/uSRhQv4jMp/mw0G0G0LxZsjlUwEO0aIfyFWjEZSOVA
ph0Eoimwtx4l+RAJIPBPsOdbNUFN8WRfE42CNNqiMxGlapAUaDyCqrsjXn+rKU0e
UCeR5afh8FmbyS47cNJIdEOZJiFqgfPSBzcFUFiMJpjCrLJ1GRG/QP/QAf7ej66B
ijW6/0PZ2sugSuiUc4bt4ck+iRmzhVn2uAQF5nvgdRBEM+DoG6snwJEW66/M1cbR
6Fgw3L2F3swfY7QBrYL9HeyTFlpJ1oeB+kBRVD/YtoBxGOyunh8LK51tISVxSqwy
7TuIUMc7nQuX4dwL+KGsJGDeNTAjQefqZBywcsfUmw7jZrFJDsWzfyZTdUTYXnLt
SckqFvyQ7KfYHGMipxtT3SyomO/6/xZUPBNbGZSL/2dT3uZ7mQLxQkXITS7T+5oK
Tp2/aldsgiMWXHu2vLI0CAYra9rRNPBP/zsWH7ea65TtckvAfKY1ILsOttX3ez1u
P5eIdovC95F5jS96AmNQvXOEROuM9tQgjpZ186xb/XUKmJFFqzXTLeyz1EhwVJt5
lRbPGmYyHm4GIT/0QMjsZluEJVaUfyDKqGM7ZWnEhlORar5Oa5c2KCmhteFuybdM
cbQWtNuGZU6U5BI8e0KS9mJPRUgfh4okQes++9hMIoG+VABmGm/qws7tpoFgO35g
+U0hJXYRW7jJ9aeWbkfw0Xa3OQhhCinv/ewTwduGUrXfUjddvzMtoprN0H08jTBf
0goVWqPaO4EkUlNsXHEUi29d8g0grUz3V4Zx0fqi94c5GiyUS0zJ0badcpxiM0cU
PKItwP24JHSZeJjkNmL/T+xdWa8wpuh+jyyBGmQ6KFroP7h3HbgnzIf9wM0S6ShL
Oy/d1aJgetm/g81leM3PGmOJZGVKVe7to1AeRW/fhiw9wcsct9VVt4dbVK/uvYv+
8LADytyUh42IiC6s8f+p90fFtdkVjYZKliHvVUeuRD2m+48Y5ZXxqa4k4Jv4mJUr
If7JWDEsrY5oq9gIHwxtJuDvh+2/LQeTk21PBOD/ZwLDqwQf1/UWl3t7JkU5Q4nb
qcX5VR44jfZhxXnmpq8stE6pJSYFHQNqXP+ZToIcbIMONyLbjhQj4AEi6zHjaqS+
9nd3p58SdbAd2Y6xVu38NwaCNaYXEmgbDyjPnmQmjelLcrMppZkyauzzuPJXMG69
rrGGgbrxyPHCBQk7+mS5eO/AUoKmJubx7ni/3PPaeXbs9vrokIMZPY/POgx5NkOU
Jxz1N3eXOrV6dlXfqONN5RIjsjaWkXUwuHtdB5+R5j8lid02ERvaJq3qRNbUrAFn
49ldVdD5C4RYA9wBASZ33qxNPS2Z7Ef8P20WQxxPE7bELbos0bmaw9gwI2OcrQ/0
zqO5cQNUBw66N3BmMNz4jiZUy7cL8bE9aS0IRCbKlgbuy1V11BNCU6IHjF8Cc4PD
oicJgY3lr6CJC7TvjVLZLaxhYJTVnbkUL63NxLmVYRA5gVv7FDPQ1PBrirezuYEb
Y2G6OW0i6MyYlEEZD50qE4I4q5TTdSXllbLxs86Ty07E1XxhLTr7bSTO4v2Or1fH
L2kTxab+kaNH6U08EU4u506/lg15QP7ElqSvVHSXkce9j1uldXZN1cWYrIZwzHim
01AONCji4FZM9mdGI0ia417gMx5EuoCJjzARDzsNmejtHo0sk8iTtT6b20KutQpO
Cff1Qq5MVuUsSbXLvWwHIgzPpI03gZOpEPa1n6D3C8L4ZIUdLJZlom1lYtamQxsa
rdOZVEiTqS4ZZYYltpwccAyspFCavjefKeXg1xHHNDtVSwEYgROvfaTi+0msSXN1
xsCupes5hGwn0bqn4v/UehiYtffh7+GIXEmvWSjB/bFLenawEGFMAKn7y0mPGyMn
qrTlfg4Ayyl7wpC3/2D9kKzcaMQjVVaZYfR0X7Cl+1RzlLFrG5GSEeVSHPFV/VK3
1BOWHlGvQTgmF7LPjbmoZw/8r+7KeqQZ8I6Ge/QaYEs5qDKaSfy5HivI05Hs6lfV
yyGuhVY/m1nEB5THjVwyuO0waHtXOHXVRBN+D+jQxkgI8HqzhixcFvyQJD2MmBDp
hvCoN160EsxcbTNnJD949k7pHz0mCgcTPyJpxfuNYnuy4rgikM6Bl6ByinPc15IJ
Jg4RhNzTrMTqj0VMhw5eeolysedG5/H6lAWa25czgiDEUnI94dfNOsV3ux/otQBZ
IIxk3B4oAjusTOX4zA3zLc+7hNSewtSjSH4Svlld67KIpVbAxzBtDQHkdSprykh0
+qYrALx4rrCUelYwDHiZDFTLAmZn72MyD/GRgtdTUWo6c0Ol10+U8zWCliN3DJhh
J95OHjMdTQ9WNNH57X2u3codIkRm4OvhNtlqWsI+jNFLLLb3TgrMq2x0y43c51h1
CdmPZY5G+cpu25NlM1iq1UapuC3d0unC8Sa6wLUjuFG8nFt26Y20Q9vhM6ztZuMP
JzWWaaqHG48v/FoVfixdrvXBEh/WDZ4uGajtrnHNCbiYymXuMG4GBpBfAzPfXbhi
mkeZwSTkQ9tNvhhwdtSApiCafh3p2SV73n0FhwcZ96olDcQxEfWqx/uyag4jAXiE
9UBVFBdkbpdZXavt43g4Zz/NDedNEWQTJF7fHpEgefBbQS+m3P/9OMThGJDqoDax
ZT9j8fwTYBdjEmvK1PaAjSKixWk2rSHPNhBVfFbiFEDoVuXNp/YG21s2xv+hk/g4
LkkeOUIyqxVq0Ynn0bW0BA0twJzIF5ccRmVxilpvHxWAgQrENLmVFpmGJwHweyn7
OpVI53yhW7C524E2MNgKSSLvWzYMHNdnQy0khfUcdvbggiylemW+lAfxNbeQopwz
zKWcr6HnwSWI9zEpumuqxYofWZDbgZcMGi5YE/x5Jtvs3hBaASuMieqXbuD9IvcU
gEgKvilS5xqugkk58eAGY07q//Z0jFQoJHVEtLAArA9EaTlm4iu5r/dklK9/9pF2
2EaUC7G8vzWVcKfZma26JESzX3dddvuCfVU2PNnAIY0fudpeXzy62GHRRAzsz046
KrCIf9VL7WhOgQOnjYl43qiU20uvs35IeCssXOPIUZ8WW8imbQL1DNkqicjUe14R
At+3zKNLGl9hyYJiZ5gAXV15B79S7DMMSKcx3hG66PK4k8+VUr1+V0sBu2ZVpZ+B
dhRYGd5AOsZr3YBn0PUFFCVF+7JqoGUAKLuX+O3s0BtURS0YgEsRxyV/9joslySd
vWyR6Iz6aHXvwN6v9xar7JvKw9sYSN57I5VrMDULcKHWnonikM3nuW41JZLWyODg
X7HAzcjfXYWucq29AjO5x3JR1vZGkEIt5/LcuLkSluiHGw6oUxjQw8XCuzrqeza/
xJnckSO3RnFqT9HJ2/aySxVj3djvPekFXAqd1YnpyDGvDRgjtf27+XyefHOUq67B
IysHwj9+4hNQB/AE8hFCFNdgYTrKp6OxaBEcuV3lESFSKRmHnsTrPc/anal9jORa
eGNCRw345sYaRTDB8AOhjZ2ynYK5MkDPsf6dZ6VbBb2x4T+mg+GItfxkRgDzhxAj
W03/LI/ddPCiFTWvPXsCIMtb73TKV3ywkUOP9+Mxz/2jq0HnmKW88rXvrYDry3xP
RS2yZWQNwA6mdn2tywRhcCcZkUIbD4h7c3s06OGDuwaR+wi9xhZ7fodCz7mGbSzr
fBI//87KcU91vh+I1f7xLPqH8tU0oI55PF5W9Oys3gowlsrDdJ6JuF7HPd4OJr+S
K5/Ln+TS/b9KU7+H+ngayiYH3uLCYSzl8JMlb+dpeCQFy318DDPtHC9WRdcE5cf9
IuckfxD0SotfCXR1t+QliOqRnrrcv9XRR7Jt4pyepV73quZ7EHRCSBAGO83uBxag
IpKxL/uu36DONTX06L7Vx6malOyPB5tLJgG0oeO43Avm8OQpsSP4mnegJBjX/LGJ
m81KX5uTMkIYZi/s5WjtLScEbzWHMwhVHzIEAoIDipAIjiBXy+OI571Rh0LaKvwm
vO5IU205x6pEtUH6JaLUEwhXEpG5nEZH2sz9LNQSY2JnXPkGH8XrbHj1zcoCh6zp
/0jRJHl92sGcuUD7+Ho8/2uzSPjlIr6vHl0lhDjmDWyGlg3GFKxGyKq0DGfGbO7G
zr25KglFPsXTm/qN905ReXliLAdRb53jdgbtaaROnRxesDr+rHYNqgsj5k4WmZ2j
d9+/hALNF6kM/xZTtwwv3y3QWzAymeunpSOfkYvUh+Ggyhw2pWw3MRypyl1BfKa+
wanOndmlE2EM1k9iEBSV8LSX4BkoS3y8YdC3f9ACppKUYI+UN6rkP5P2jXuJ/Xyv
M8OBeFGYAwcmSZiapFi5oZlL2XrCevufyOpJwpr0sTbCzEHPmW9ROsewbgzfm+6J
KfrkRdBgMhyHOLEk3P/LyDLzd3OBotWWqn39FXYsCPt6iID5lxWLVTEa1nc97gW0
9flyOpVntKCCbhJyCsp8JCFObgE9UxJaWzcZjwHuyLTb+Zj5Sx6RZzvftCvt/cWs
4FIrE49iC5R1y/UMbQu26GcULYk03eS5B+wmWsQdbofex01GA/E6bBlJq253PVbA
LizEHadx8xlO9gM+Hadlt0QHUUCpKkgUhxtOebCN1LCLyQ33AgQOO2l975iQZ9rQ
51s0gvhjnPyUQfkZWYEunt/AjN/YQzTtyWrPUaps2sbk79dTeOCJK96SlXuYv2th
DU+xld3zO7cmPhXzJwFt+w/uOSKC1w+/O9yhBsoJZIorkvCLiXHpAHAJvG6Jrmq3
1SY8hdAOh9efs1q4hN0bAyLK8AkzMXWQyhLMU9XO6CZyZ9vus7C1Ijcw81L92g7O
ex7pS+kF2S3zYD7+wiEwtppDzU7NA1e5+qRsKK7jB0VNQF7cIMp7FOmEynoiCvEI
PSrrUK9u/6pnA/jCiKlSJ1AVuN6DZMOJmVdu6xJaOL4FZyRkJQbaL2cF0OYMOYDM
UuhhJgcM7JP5s7SkYPNbdcZVZiEhxJYFAYSb0DG+JO4shh9oe9IqD4o1QJfD1wgv
pTOjKFGijdmsvzWE6P2RGgmqAaECyWkGpve1p0MvPa8JEfDBLN4VE23gsazETQZh
4HBswYmTD2iKHqPdtinUQ6PVLjljU+YxRaUSlkB8TGf9SMd94SR7mo+EBbY963sK
BE21wQtzVkFJIS59+JH+ORjSJC6+iRiKMxWj626y2Wm892kO9NNfoEDBQ+e0J4He
K7/vdQldlGAkFjNnHdjpTAZrubeuJWdzUBTCpagQ2miiCZKtk2Yf91eeaF5JZq3r
II+E6FXy5vDjYK92YbWq2DkXqVr1xCUoGJVTrDnTc94g6lb/7vw0kePcD+hOv9Yf
LonJoBnY9NfejmNnOu+HdYmO3Gd/T+5Pfyit8XXPxlUR6N9YoLkF2ZktaGAuQAid
VtQ4O5kRYbEk/sZduja1/Ra9r+uTCeSNeCkIxFuAJOaQvfCit5NW1QyAPM6ml82a
I9TDh6dEsb6YDsrxnMT06YO5h7QXQCmdbMcmyakQ25Waqfvfo/MBaWooK+pPBw9l
PksvxLxc67g4yrYgNjQQKnoM6NR+fY2ZuXku4gRZe+oM73mcza0lIbSUtJsgI/1u
gps5CiJKTuPvHNzMJpeM4dw7LHEYj2ePn4EDQCAxZXpZ8v6E+GVEEIavhvPF/TCa
V05UH5l4WtXatd26T+S3nmEXRuaPQiw5lIK/7OY8tLWJ4gLdjg+id6kmkfcEgV80
qk84QoNl6WIYUbYEwyyjZiXzFqOxZxKKsreaqtpgpOgyPlYMnPW/eBQGMUh2qWCT
JMs81DW8ROACRbTvjbebd/HGVJFoXCY/k0t6vwnPo9M6HCdv3TTmbnJGVlaHJ2vl
mJaQAO/prkzNJRZQe/pHpo0hcZhBOU5cD51RI6/jJWF8H28TyzLbpxncJ4AN8QYc
jgmGTSszrpgqdXOoMP1PhoaNmGLye5JGcB9O5yhsv7zoBNILu4rgXP9bnwNseiDB
YbvAr6QS0/8+Hysv81Uy2+MFMMaA4/7adhPTpJsq+DuF4YO/jtx/k43lHfa0uydi
YXpXg/jVLJJod6zCwIud74seWVvfVDI9aPSaDco19oq89RI+V4BWUTowlHDkJLmK
BZ6XEweMtAddHi19CUpkJVmR+49kxF/w8ZuylOvfxWTdua7jofx7C96q30JwK677
QvhuR1VA4MrtPXkbR8Pm3rqwpMVZ0gei8vPLy0JvH9iGxXhRZGjpeibzy0v2LkWV
F8gB26McU+GlQzvEzE+0D5UohmGEbIFz8Xv0T3U9Xqptq+JX+MB38qj0PsR0IsFu
UVgkMBqngfe+m72xhvpFWmnb6VSvFezTuJKCeI9TgLSUrSwQ7Cp9cJuAOH4R70bg
pyxfNOjasSCzs/pxtA4+uyy5Hcjv+OM9XYKfQofgs3AHfeUnQMUSLaCIiccGfGpG
RkSt2JgJnfOR6W02Y64Q0uF+INCdHD2I8ptdOcRUjVe7+o6dqdIzYaWJ1vKqRuMG
cTtabk9AWunEj7LpfVxk57UoRJB2M9rpKuOukF96pNoI7cnUWnTXKXvueXbsIMvv
1c/moK04/16ylKWx+AN+LIayzChrlnVS6ghaVjQf/fVuCXj+k7rubjnrISQKFW/f
ywTX2MgzQ+4UAaCTPkT59fDMplbeyS5hvw9g3wnxxVZHl0+JA285ojLsKg4kyBxh
fbgmnRD1SkvzIOgjxLupKhtfkBycUzRBTU5P3m8g+W2e+88DlnY8XQ9TwbNnVTfU
jyPxw4CCQ+mRzkhWPZ4Ll+mmPLcfm46C/l4Odn/tHyO5U7uGlH1XCG6fT9N1AkJz
e5sk/K/LCHOOpXUr6sP1j+UR4qa3IP+2CdkfjbG6UiBLroidgwlGThp99lwWC8lX
JWItH/HRlqD6CEXLtgtaiGuFWQ6frKI6fw/QKG9QWqwj1qQyqN0+ZYyTuMG0SmNk
rptT11IdT1ribuzN/5L0yXmNq2UNrC8u4aVxibRmRYZi1gMwyuD30YvyXOV+m/fH
xPIkuS/tZs+O2vBTIjqzH3Cy1DiHYKyp3vjsJJo/RZ053iAsZTTFgNg6rdVQaa0a
vzBggIDUg1VliVqI879kJy0FE8riXO0w2MXouoADox+gZwatB/IWw1qQCJ5tNE6b
GPwMVZrYfHQ7aznPcAC9VRAlNUlGynuy7+uLv5rbt2Vd4xaT2NsClGL8vFSxBOQH
OfCg8zb0RXp6rWqBbotOpFxiYCpkXVxhKrR4mWxZcnokuVOavvepppbXWMZcKK+j
YtTxR3LGeBd1er8vkn9jeBVbCgN2xF3aj26qJlCYl41DSjgC83r1tn78GAa06D8I
HsKfU6Eh/j4J/NoOUY+u5cmzhA5AqHDffgzw++/XpSPGnW7vvHjyf5D7u5JC5ABz
4AwguyX9S2lDE6+aCg2HCI7w4aZA8D4kxAkDr77pS3KN4L0IfW4m91F8oktVmH7r
svYqd9T3203jbPvGv1fJpuGK1uJAhYUZbw6Dp/8thgoYIa4mzFnlL5fxUVnhimch
UaMj7aj0ovtHd4vxoQ0Je2lJBZphx2PxBKABdW1MaQF/2iBwNwNX0xDdikfjj9LW
4unX2LdutXBS7/23XTTrSZdBHVToxt1enmLgD+2OFikQDsZ0N6pLG0RjcVEKCxGP
iQXS2i13MW2InFcluKTWowW3crvEraSeheGk+V4TUdtSaeIgAI3UDo3IIdyQaIfy
dMHeclkVbOeoUERK2EoKcxPUMYgHADE7AMvi8EhdSvpFOVXRlvHzYqLow+vgSbUD
8yS8n1IDjmVD5EnOgQiWy2qsdDUv+9NIrgSEgxkzBuEC8dSfG+SYcVBTSq2FrIly
MbAbqXhiKck96v0Am8+rdDfb6fdJIf7mKEtHWGzkxOoMaV4RvveiEBcS3qcA0gYd
JPFefh2l1/Vtzk1jlLwL/fVqvfaSqEq587NXAkvW3oTRAae9y+D+eWDqclZoyUPl
lMbPspiDv02PEZrjo9zotS5dHOWYmwZDj/NmeInSyTXzEhlOdHyV1qJOaA2lnh33
UrhoVCdg76LNe7801esvOTZVq7+Tva1HswJwBC4dnCJytGRfEnRCIXDHYEm3HOVN
CKn2MqKwZldJhqRtsPSLLuQAP0qOIVyeFfvvPSfzAx510o53niXzIreAt5P27Lrn
1zQFRYiR1Fajd7bUUBA49t5uHYxlK+TeQEH8NnCz6EQ0ZszdEJTO9kaGXYGIHd5m
bYQ+Wc4FHz6MRzpujJeWZP2aBqXjj9RAvAJ+h7hLoY97honTSBbg+xrMPa4ZNcim
3P++vOrG5KifFbP88stodpX2gzq0CZUhVg1B0w1SB12+F1Ir+EG38InelwkWNV8y
HPEREW45s53tGfEahK81fYCB3CzpRpIxd0Go31zDwy/hPKd2p+E3VPnyp4z2t6VA
1iHkHtmy89kxklbHKjBBv/hxXpMNbrvos+qsPGKhiPxCwMOJeoMcSqtCcpnrN78B
8yj4mZNaVNma/fSoBl03WPz9cCDHlJhlKL2WEI4ihYepYnDC9t8Siavim6EMn+xm
sVB9zbfqcGe9e1hDtMQOOihwXesBQk5wphv3tgZzeYLoQ9ybWoGhv+v9zw0DGxM0
imO8II5Wl6g8uOlP7BMiQuZ2TzDBwxBNX4bIBc1tgJbD6fToD5PoDpzwB9Ynjo0d
AlBh2bsUFoa4+Vc0Ch07pTncTUXPmf2yT+ncvuYBEp9yi63tssF86g09aaJFp0Gu
lhoDEYTg5K9+H1y1OtzBOOE3+bmCuOLA8pa2Vus9HNk8IH7TbrdEEWvffS95jbeT
K7qqN/0R8Cefj8AmqedwvNhLz1EAgF/cJqTAk8hRIEchiFwvkLpdTJRgxlan6RUR
B9GOtqW4N3KENcUyrv4E7EMV0qAsHAwe1bFeZXE/n38Pu7HWzwC/fgTBWZpKTsMt
csUhBeJX4d18pl2Bebs4tNSY/JGIe2eLsUtZo7AtHJgUoJJhKVUQiDjQdh8Lfknu
kL8I0AVqomITmfdolcmlR3u9Ggd0A/WobI9eUIXtXqxsOSMylxa/Ef5gID0ZCrVP
ePdOF2c4nnMXj8Zk7cVgPacpai26JqCNjjRbCzhZyIAO9jMNCSB1e81o1jgXKyoU
vHnieu21BD4s+CQdc2NwWDeWBmf499JFHGi7YfzeU/psbZUOzVJ3IAfajoodRloT
xSuIHxg2ehdn7QaRPHn/1Iu0VKuJ11hIMqrvt+/SPSppnf2i7jA9dBeOhV8f59zE
0EBYWQhjGoaI3nNdFiX7nBAdPRxBBH9z/SNmCvCcVpVPNzLtSpcWoSAz+B1K9aao
p4JG/cEyYTQ2O0QKCj4i/WUf+cSDU1eR05L2rTysDEX7magTlGfAkAd9h/OvPnOE
FmGKMK/dRuV8wJDz9Se3/0ytkWW6foQ4wZHimsGxuFS64I6OYdSJWBmc4XAhSze5
ylL+OD2TxWcl67oykYp9rBySBpKfsJcLwMhRKVXmHWGeVI63er7bNnscb6cMhNw/
4+Uu2VI6uId23YCyJZh+QWHSzhkjeaX5rXSRXAl/F7Yid5YLm4Tc0gXeK2IkBOeY
ReVu5tM21Wq6n2VxRgafdOknXgsacLCueRuH01383V1Z8TlHP/99hZSFwXEVpzrX
jWqFTEdWEWL+5j9rjWg9H60zAUeWIsD9P9ecgzDUDmmrOq2R/c1pG7HHQp6kFHjk
F+UBlXE73H7vMOcolyfIzpEXQHHhEG4PW6VjD9/7O7NG/o3orQIQ91UR2JDHL+vM
GMJpbQk03bk9RSFI67JVA0AjwLNyc7fd70CA+2/gtWYdKjMGVQcoAi+kCWMxBf54
V3d7vhNTSW6lDTogyd7oTtJjn+sf7+pVZR768iekG/VRG0n7zhaG2FOmy0d2r0cg
rbxOcMA72ZJ3se/eHS7gldKb6Uz0Y2Jzx/rUbVLpdNZAPeEj5O5HmYu+rn6ZC97n
75LZoNc5R3m+DMgcRWHhCYY5h62Zsz26narN0xBaK89fCCnNNXDMMvtg5+HrvUnY
dnqZRYF4h7jeFt0NAcFiKe7hWzI+9cH4xpm2S7nmaGxVkDGNk2yU/NO+Igx/sO48
YHJiATZkwhQh03WMXWJbz1iiXocOBNK2dNt4BaB7NO5R5HkCOVIeOKha7qodPIgw
X0ZRmUrrkCyU+N2G3a4ARDX30Uvo1o5U948WSm9S/QwTksrC0gdyN9ITuWyoRKnc
NcdHtVRu8e7xywXohWej0wkpTFcs02XYahQGfJOVx7A3cz0ScOuyPyQptr8K90DY
yUdKS5bRCNR5xH30JUi/AvMi8hMj8eiC0x3fk3AR1L2Fb2rnFlCYsJ7NWWwWci4e
moGP7d+sT8eeZBGQC26b2ByOyl1yzgBhY66BYDbSKj2Et7Le4p7KqfC8+yequYGC
HSNDsy1plF3qrXbJhk9cebtn/GKvgiRNd4TyinthhzGRRJ8o4hhz1jksgvgVqzn5
mRZBdkqfuWZbGI107MHjGVNYlDGKVzTgQ2nGs7xZBK+jrIK0urzlt04c1fKMRbNN
XOG3R2qhFLNSIu/hHRyM0NtwPzOrwH4rk9RrOzsJ4sqVfU9895kVoIL8GtoOXq9p
flouXtp1Thb+NGkFupA9xYRHsFS/c7W+KM4b+G9zcDnJEF4VyNJxrOivQdDutOfv
g6xULZg2v31W/1PbQE2nphC7ltvIDt61TNbkTwdJgft5SchujUR7UzLaU2TxTPvg
4rv+lMj7JeRm0tE6xCsoccbTZkfb8FiHqJ9KqVW1aoeMlwPAcuUp/rJ3vo/slDEj
AYNXPDtYrlAp/71wbBlfcJqLF7OpCxWuqWAR1ekTLb4X8sAhezpDlB3WR18wIRIo
IZ78Z1KXaB8xabsvPXg7Wzw2uIXGaM0MIqv5DK+v/AvF+wA3qNB+Rgojcgr7UOYH
yV/pMTIWBAvrbA88ObHGe6zbQ08QN/N7Alv76kh/nVlTEjXYpVFgwlzs/pbhXag+
iPh7BfKMz3m0luClfh7cK6niF70+tRu0Ril2TivhdemEoLimGz1lipe0de21lb22
K3fDMuaSZIRrnOo2oQipQ4nAxbfz7Ghl9m8l7gjE4CX7VewKUB8+D8Ub1/YNCDqV
gOvSOndBAY/eKdLZnIaRxtQrVHTMJS4I5eEaJ9MTY20E3nCCtJhZV3fxogJ5b3va
tIrWJusVNozbyZOPpu8I6NzW4Qqb/17mydAfpLi/RSz6FQMEOAces2axe+H4/Mhw
BTkW4Ar6pS7CjAU03osb6F0IL1SPXLCEtxqBLv7ow/dxXEKRoBkdZeyRg5UeXY65
AtEpN9YF3pZTpm0R9P1GES85koNDbWx9EQQhwEo2tbAYcx5wtnbNTEFgFEtVBrx2
rpyTex8gND2j0MH6RyAet++r3PBrjJJ7LfG3Nq5LcuiBF3oLBxNHOTqlU4TgptCh
4LmvrpWBT8qPsXZA9x6ip3ZjvqtR1wfzgAsxiCNasVi6cxmUPQt/2+zDhF15k4on
/OU0IDu9dsx4mQ7diJF/hRNHROk9pe5bpM4Ot6zUspj6ZfjRRqXisU7jfdN5q8h2
1f2iCBpJ0meaza0drYQ9hYIvsg2jvWulwvJC+HdNpEf8I4kbZotzVlzOUmHKJYfB
A0nMwFK748ZVLQcqLwp8KgFsPqJ2JhQBqSRS7zpNdQTOhoz+NOZ5YFZRBVN6RgXR
f8PAdXegPhC5YUh1Ty+98It8UmxspPI18mrsiaE9nIKkkeRydw/4GdYgFmMb3uRn
/hrcgNF5yRqEREdqZ9ztWqEKXDz6b4BHYL0Zw5upVtahnM+eOywqi96uMtlHtOG+
oxUpFe7ft4Wu+LuOEM1YkGR99Y7yV4+7DZl4C4Moks6IAJFYXzXQdqsOfw7CFHlP
9X3Hu4v2usFzr46wD1p1eff/g3dtrFnXQY0+6CF5ZZLw8yq/7nXVhzbjHNnq8zRe
X8h75v7w3/vCFXc+x8uFFpb/R1eJX7zEjtWIrCi6MuTJnnDr8ElqY8NNuzBceUrg
a/A61Q3ToPVMIL7qGmdDT1Q6G8urZxYuNuU3Q/a436qwmUUBDxMU4TNFqKgqk5p7
c9gKuMt8fPfmPAhqRrx0evn1eohe1R+nLg5sam8sEk7Xr8It6XmDZzo6BboOD++l
yYRs9A6vrZ9y59eZ9vC8H2DPyrC03hB0gLRJbDsp4Vi4m0g0s70lFkxALGmAIig0
6q/c8rEDfS0vy0pIvhi/MTiFv5ec6O+QXNT+vKYTjXeTUyvdSGTYyHJaSo8VNEs3
XrDFYKyAtLh8sOEfy0ObLEAN3qNCqvvP6dVPqCL2BRiuUlaLsySwO5O1bF3xADYl
WHU+4BrwYCDSrSSY6nGbE72um32VNevQm8pqxOdzXt81bxWjeFXQygn/7v6G/jtm
rwMlG/lYpOC0E8U5KOH1Ixy708HKyUuIT1/5C15IvO+O2wlHR4znBXYzCEO9xLa+
ZjSWMuVSupMpRxZ22SxzZN7Gw/dPrLwG5cQNv4671CVBFs7yYRCWmSB1hzGh59YO
GD6Y5IBFPgQroMoM8+LdGRobXOZ8gcGaHYRMKenbFGN0mtTK8wlH2Actq+GI5rHn
nNGBB7txEb1cmgxC/1rAyiZ51/4vh24Sv6rpwzuf4i+VUvgTzzDDGVr9f5Ke5rq+
qbsnO8a/TfJTGgRxr3cLuPb3cRzCZU0GYsXMNPQD2czE6PCTfsFAvefOC4Q4865g
BOGZhCsW0aQacxdKjOyfABuDemxo1SKf1zEdE3UYozQULpKH48JhrinYRr+lrNr3
MBACoEcJ2kSMcLEZ94BM1KHwJyKukdCL59kyHikP9rxkwyvEpA8ZhYNW7rmuXUyR
54EqUqfLebXZ7OHplrm86Hzm2jJu9ZAuEdJE6Suzq+NXGPJGJW72yzdbaN5Rr4CI
cnUaJjVvZXwsUc22wGjlIUS1xQnf/v+c0V9gvdxrOZvKLbUp+JlgHPnb2YrsIXN4
NOREYbCoejwZfuyAfafNdcPzlY7vqIUJ1+R+dtSOlOqwJx6SZG5ev7K4138eJqP6
/gD2PdatbrR/BGykCw864cRPJkFfnxr5TglMgaMGs1wF8mfNZNko4ugNqtXsQa3l
T3VFSaS2GY86JNnkCIDJo7v4ji6BfWJYcgW77srgM4LQQQitiuimCjGWn29m+7XD
mQDio+2sbnUMpkpT4xookbOW4OeMkpSBypn54KNEcu3nWvUCJr4OAfe3vQg8kxv2
qKVjmgSsXyiRsaUFQAGT6un1nAhZZ38XCcP1Dm/JFUGXHCRlklKjZeHDuaX/I3te
sZ4vTFuNmmjKAFbLAa1Dm4VCSlbdE3+1G9ZiSG4y/E+3DzyywQvxURvdG/MRS/nC
cGKcN5S2pbksbJziCQP5fjFt7NNLtNwrE0zLKx5q/sYcgbYpt1db6EZypEcQBQ8R
AwjY2b6v+YNzEq1yyYSMtslY6W5pI8LCakFRY7k5j1ky7ZhoE68SbS60Or7qWIAU
TAZz4gO9lokIFP64yXvSz1IcMz0B4YBwssAAHt/ppa4xrSrVrp0B1JZQB37mRO7J
ooZagSZWCUUOdhfeiksppzc1wDVwnbXUtBRyIe5rUcWkWLPwf/TjQRmjt56YfAJw
QgENNIHlpP00GdbMTqj4+RUfCsCvBlQO2Ea5rbInBHJ7wnKaWxGUYLiZwpnCmAC7
a0/uK+emZAs6AcX4NPZxKxn2GsY3+YCkttWaA0BoysL7rxsnBWP72Q//yPStedYT
Ee81rm+coCWl/00j+Ah4iiAXuDayc0xHunPkHHkQo90oTlCPMgMaYa0FqYdMk7ED
syYYMHijVXJGYTxNs1bDaSKWDwfh9cQ3U5QsbyV+uNVIBefNwyjFiP+kpvQqvy+i
ZwLNjnKs2P1EfRWmB5K+mJFLo8JQ4DmMnpt/yyx3B12G0Z0m/wuUmEL+CmLA0rbr
gv52Ap0dafuhCrKv7Ww+JucMJ2NHUEfrjFHV3asORoSgFW/8O6gRfoWqDaLo9DEA
b5jPd9hmGlii8VTqFtJ6cur8Uu82U0pvS50h9thNlVv1zfCyHeaz8e6vXZH/xxe7
8Nx7EHzC0mU8fTsPUr0qC0nIYEH9OE2nab3u6RJIAMuUvs0w+DLvm7waWnPcWPFr
LZUUUOjkl1uYJR8+TZytkR8aT8YcJmzrPMYUftFB++XmZ1Ndah+ge/MduRa5sshz
wQMWVYLczJNDkeJEb0CHikS2Pzb7iBQQzLL81FNeuYEb7eQfoiK5VNxLPEl6eOEr
TXEU1drUgIEmNvCpu2W33xoz8bGrbv1TzZMvk7yHXTaqO37kEgsCE0te53tgkcsR
jJ/2Ko+8st+T87ALstirFksbrqoznKXAEjaH5l+PRgGUW1H1FVqtW1TqJJ5HLX8j
1iniPFzedqa1hI+3JGP+4p6Xkuk88KF3N5KsTdE1uBIKUe3upqNDNY4wk8PyQphm
Up9hahnW1e/69eWPKQw8dSy5N146GaVQsFg00ebXe7vTrCaRUN1wqlNE12+5y7pr
gM8ddSUSwspUZEDr9BXUtTr2ff7lqC3Dt2I3rggzG57K49Vt1ZH6HglB3CEuQvM8
RFiht91X1gTjZqIj4QiFN2YXB3D52WKBzPTg2UGGDq9/3qhTtZVt5YtCYUjXZwAe
a6jFUFC2gWVrPkDv3Fp8lfWyoxw+JKzzOnRN0oGmktoHIhMs0DL+nyemhJNCcfWm
GC6kRwny98jWKaZVkLYg+aOT2EfDnVYXerWUMJiFVRUWtiw7q+QZMAp1AczZybb2
cqc/93GeMn9u4C5kqyuLK3b19djJJ9SnopkifSZcZXcN2sTkPhPgLVLuCgzu51tb
nViZRWDXhzp3NmhKoV16QQ6cxrdUPW8ZfERONger67mTWnWEUz7gZ/R/KozOTfoQ
4BqD+1v3pDujmdq+m0D4BRtEXgpS2+1mZ8gDlR0n51+HojIgHdnUW422gkOB/WbY
/r4Ghasuh0mTisSqXG8yEMOIFOW2RnIvjdkxLHCEB7ugrX+djTLtQifluD6UfVbZ
Tk0ctYWWA/aN6lYrDtJmxb0XROVPUhQs901xkRBFFeujR/pFoCEKOIVpw5lzkMxH
3eUBN1UspxgwfNNEEVgi2WQsOOQrjwZ96P44kTh0te3cPtec8ZxdxRpNVk/abgf3
GGkLhzPM55ewvBIrxSTnCb6q237scwDBo+nhc29qMN74nLpTaULXPdr97MUNylI7
yXw2xP6g2R4k9i5sa19tzuD16vx5leiETP0u74D+karVnnapjBGcQGaID/H4GDw/
vMfVjR4L4cyV5m5rcmjHxCHK87pA6fTMEhEiYIPeNfinilGMs0ZODH8ZqpFyKsGG
J3zYszcBDey8hXXhxJpPQ84Pf0I1qQIXUPRNJvO9p8l9ivFYy8vQ3Cxe4oZy7roQ
ljH+RiHfDUup5LB5d0Bm2vp6K69IY3k8SOOs3iTee0pjRNqLSc+0aHTo6IpW2Kny
5/4X8KmLU5lnz25bAwy9tMOwKg6yzmVBMkn2RPtzjHiaNMS8PUpibTKTwW5vBljP
OT4MyjLUR8rH7yAZp+DJRroizTvaiGZ8dEedZx4A8sBdKVTM8Vme0BB+qZTO7dpC
0AUnn9GIZ215QC7zM0sL7O7kEGw2bB9BIlKlRWnXlLMEjkqqOZzvnrGpzo0xzfBc
RNh8bJBlq+mYUI5i+bGbc+VeOAGPUmYH4jtuu+Bl4SI4l8UaXskg+Nw2L5rmYqUc
SUYwwrVvyO+P3QupHEUQ+YztDusLyMEkCO2HGpM4/VTwArE+Y8XXQbpOBbSEfbFa
pEpvOr0EWxaUzgW4GtiXYSEKmbEREZribeS3LTr9kD9KXqDcKgms6JbTt1RQwBBi
I93+tjRBuvMG7Hp3rWZwWaQ4YmEbea27zzgRq6SvCiXb0QTjTMuKrLS0L9+op2TN
LWkA6ZgsIOPmqX1k1Wxui0QF26LVxh0fuLkS7io2SxpKJOurOd3pg1fafrwvXVDo
6UzEtPCHZzB6l28hP6mOX0/5TVdgtrmabIpJF8ZhcfyfLzJD4DR//jBueBawMOV1
6Hqh1XsGlkA712hUGLgzyvJHoTO96EISOEsLeFIR8Zx4SMhCWo2r6VnsdlatBbjF
nw7LUskt6nsPKFZz5Oy6/Lf6jCUKU9KU6U5Rt9iupFxBGKOTelezPHkNSjmKqZ4Z
kR5DGQnBWwvg+j5MAvLah1d1EmcK9ZIqsSBYPcd+h7OpIajMfPw+CNQPrNorUVBc
w2+mG92c7IjW2i+bopz3bndYYNxTsNYPQrWP5JoV52cSMA4SBX7i5LBYfdRtVYfz
j+0IeDtXmaDh58kz28BytdsluiQsxpAyfmbMfCdRmaPzGiUL9HJtBHMA7YXZlzPq
Vcj0FlPGEDzMbuUDaL2EwtbKdfvl67cyw+QS9+5K7SkF7yc8SNXSA615k8dze7SZ
4DHO9b0strHWBCUFXQJMbSvI9JrtAEeuQcGEWdJXu7VjsFNJugjuDjvWFFJbYZPl
+ibXTA333zwHHwXF7tkfOFk81/EKojPnd3t9hRvy548aDRibbqbZFrrUhNwCrKms
j+fq5BZKA2aqWvZx1qnYo7Z3YSkytsgnyBm+Kvm0fbBy1HXHoX1Q7lKZLHVvVnN+
H1nHSSEylhlNcZWprgdtfx9deMhGV5lOeQNoLukPrt8OdXq7SEUXxbk4MOspO2+R
NBbpdbPgGfGGgWplBevPupK8QXPhr3E5eBTSNzcba9G+7lFgkFiCfwzONzaonM8p
kvKqHao6Q4QngxE4RW4sQ2IBt+zU50M4D1zPGqzh9QDT4grtnBxAPY7mwqBy+ijD
4lhbE0YJqqrK9oseib8paWoN6/B4avLmWaq62tUUpnIWLvCk8+df9ll2lgR0hFSU
ib8ePzBS8aEN6o1VWb03gkVSLAKju0wOdPfeGonccgFuWvQLTzZrPQutB3+/FXfo
MTMTNgeDTr0cFXDx6C7VFCQksL6dnMaJzTjrBXG08PhuOYL8zefGfEJSLLgiQF7d
LTyp16EK/txapIHzE/bkI5SRS79zi5DXiaiXY8UoIF7FqvKHYO/TyaL+qq4xR6IS
w2AqsTnpqS+nBqwZ+CyZPdt+oqN/g00CNbXl6Ys5z1DCnpG0l7MRx2sYttGXbxeA
DHtFuwl3/qp3Agd6bMRnY5I587D/1Km3aqVWSMIDeHSXbKsU3t5nr9ACUTFvtQTK
XHSdsI1AlgUSB7cm7xZ8o9hh4OjbUNyxm/DuxGvQnkSlyQVo0Ghqlhz38ObUC55k
EDEk+cISec36JvkvTui8Y+bt7wi0CvyRROSX3X8v7fomSH/WMa43zMIbsQ4qEvt0
0dnZcWOWfhuc1GrlpMVQdJMBuulvcJ57WpjwI9lGzgvnPM1mK10yslrVqY1A3iHL
GMaCAI7EyglHoZ7Q7vPbSbaNc7bDBEJWQ26AABzGcLkUjhGlqH2Q5Vyzcn79WiLq
bFhwi5lQtAm3vC6Wb8LKY7/f+LL7OGTLu3PPcMEcG1GqAVwb4iw6t7+8rqmkLL2U
VNdcq24XN6crq5jG5NeG4Agj2gac7JDcM1FHt3x8L4syGssNwbHR79Y3Fgad6FYv
rcWS92Pnv/fqa/KEd2bAc0dpiJyyVTWWrdrhpOfUMRp039++Hhre6UpNH8lxbFTb
uFzt+jcxApE5l+GhsGP/LiXqJvdHuiFpLVeSYxBeabJjqqkBtcGOHng1KVHDBgZ4
QaqE/VN+Lwh+tA3fkftPW/IviKFQNryAq4HDZNgUHXJtASFtDsrXwhJesjzmSSsz
Gmw7VKs8LqQYZh27xg4YMGJAYwqu4kn9U6gX4w23Z38EzanzuLNstvkBI4nJ9qud
hc9bS5PpSLgbDkkV8mAGUswE0QWTHb1oZebcH92dC/22ybrpBq6Fgyz4DKW38CV6
VU5ltz5TcsNtLSyN2X7kFq/I4zKOVukzhAe7YCmMVjr0AJ0R/xHBbR1zaloGyQ6r
sMVlTd5U1skX5ORqIOlkQbnMmx7YU6iPjrCdQTVuvLA9IBV5080eBTDDP2kQl1mA
rvXfVkn+BDNcGaFG08UlT7OwXG5PrRRSTUrbhsOC6ZMHpKs+EJQx7EQkCjanArnG
9EEfXsH2t2hyyq/WtpwBoH49hURi5IfYhYlxvd0r+AKofRE0G+GyvYqTmOBX52zj
6t3nyvLktaTUa6d8SbhxC5aIe2eKDzEmf+/EeFrKsPaXYYy1xewl0YhdGN2fR0JQ
elOya9zF3u3thvOzAMhuh4RcYxXBHNWedziFsoiPeqHH9UrlwH1pDqngkBOUO0CF
RdzpPP24z/prK3yQcyfiDcAk8dg83+vh1dl4I7HhliZBhsnksZOFIyvdzGbgYt/3
89O4sSsJ07jIVyLOkxkT6UbsfwPHaW3rMjZmGEuJFlEpq6TbU9SplVJMhM5BMllx
rlYXd9yFBrHD2Vf6HRcQIjCJpw0r0p4k0r96YaFpC1dMRkzjRBtRdkm5vi7d55PS
Bu/aWQ2cFLOCERW4g/4zzK4tQCsb5OKlnnrxkFUlpRnkQ/YAlL6q5etSSN1szsPK
REfZZVNrNkZqW5A7GcEDn9MQZQH8OB4QRW71kbqZkbTOJUgFHaWTDjSNx41Jvg5S
wFhKzSLCHbeb0qIFZel6yOpKB4zLmDHHGGFKMawYdZTa+eVYQmpKtp3UXTe5IMJn
ozlYmKevUeCgd+QTid6Ux+JfKGHTCeYt09ib1YJD+3WKDEkuRmHu5xIhuEjFRZ71
y2mdFjCv6D7S3YFTiq7U1h0rk4pGvQMofJLnLd+GLs7fgjcJulgUlMi1lH5aI/Ft
WuEJFdtAXiXbXDbpRp8hfgkKdVCeIsfeq4qnwRcT9gSJCj5dNKDrmHcE3aUjwKC4
`pragma protect end_protected
