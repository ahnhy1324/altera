// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nyesLVbTxNXEJJSBCYOrxaoQ4WksNfUMhmGGnmupxEcxpeI8j22rh8FFwDzCRGNh
m+g3DMHpb8QicNNYuzARsmOXZJaALYpSLtw02Cqn9KkyZsWUM5JJFM/RrAovzt0E
u+WGi+5eG5nJ93KIgphG+Zd+OoLMQm9mmFSY5bvxTNc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9168)
f28eXWOCdJEzPD1AGL/CCUjag7hf8mTNDqqS9CqNn/J5ZOgcI34aBPVwY1bMDsAI
x21m2KTIGQvCQW3FWGQBVmMejawyQLUyCSKsueQgELFR7K7f+a+TvuKMJ38UaCv0
FwX7D2yFwjIwE9khdyk2Rk/r+8Y/Jl2F+v+TgeZ/aBjvPLn93gb/nMJCVak3OkMc
HRqlPCRaLDQrAKAPagMF2XEyxaRWncpkRY2si7p+719DHoRsh+Hh9WxcJBDSBR+i
+mM6lWp9cNv4cnrB16SQRTzQAqgZiQ4hW3cHeo0/Uhg15ojELSN1f+iddkz+krln
CacVzuDnpqJmifGZy1UXep2gT5cMENsVLFyrgUGPbuidOnSPhy/47K1U8yjAZvlB
hzG6Xzuzu/JfHyIB7KtPQTWExPClhsXZXJPeyWZoEvdWUrOGdfeTrOZQpZQWRs2F
kKoS0NoI2OqMZmrZP+cvLQ0tOVDbKI4VWmkIDB+g+sVRsm4MneW39Yzq8JfTZlHA
lcRcRUioRtFaaWP+Q1dyf1HdERjZZmRIL5BvaKffIkwN2y04NBn1M3XAjm9+lr0F
Ik41Ipnoq+KQf8okUlVrkdqFv9rJps63Ls8Q9Cvau51PbIC1QH2n2kc+Han+y4Fv
LC+fqQoq8Maquu6ueM/vYYq+mHIZO9HoniMUHovGdOKVltdOUCTg8ojGbkfGCVPW
Zp4xr78n/DkM1MLzIwUuMPclsu774T5eeN4UTS2WT9QBnMwe85U/uzv/xh2jJM4D
Tx/lP7V6BIcZV1TJn6MN+2b6VP/1foh9mv6KeZih3Y9mXPTLsc0i0GYALsxydCO4
dFqq6dplSKsT9aLaX0kfzzQFS+ISVcoQ3aHnMq3yo8uq3ZwrLuXAcZrvJEUmcp81
0MWIvo7srpILAbovc+aKv1iXoE1xwuC0A2t36hvPDn+cXoK53kVL1xR+1SIBuNvD
xmJ/gt94boGZIV31jSvjSKgT+tiCRtFe9KAs9u+SeLt8tCLAZt3TKfW61/vjfVt0
z0DeJPByJoMoUIrCD+6i/WwK2Jw7ub7bBy+bVW5w5x710btFwYy5Oa+rBBjqHYVv
4vUy2IoV3Yp8I8zuqezsX2nhhOkZzospeFzZh6gqk6IwzSiwpNdvwMTz24XVXxzw
UxaX+EMe94+x41QJO92S5q3ivHuWW0Sh8rtIq9bFu6ChyxWn5wxpla/LaVsMKrcU
/LWQ45ruPOyoQceh3MPUQgtnrlY+xaVTxdiF7DMZnIIBTL3DSdvBKyPzmR3K0kGZ
yd4C+PYnScZEvrImLM7RZMFqk4hF01ESU4L3/qmBgtRaTN+EwlGTbMOQtfNFBpuM
PVliSIXcWAloRVPX9R3Y4u/gsEvIo3ONr1wiOrT9qeHpvlfq6x9GImXXVArGObmt
ElQWGHTFW5As6cuUDc6i2bXf6OLgRxkb3DNT9b+tz7EA6k3+K67DxQqO93Nz5yLt
eZUYCLw3dsbHUPVFnStG80VsHu9EWC9I8NWWgHC91Vv0GkzA27l2Y3DhvLag82kh
8Hma1sKckt/kebAbdf+xEtO/9xcFEICFzADF6T5CclF9H46Rr/aD6TrDT6u7l7mj
ulhG4KTfjWdsksE89VjJcWxwwtPhJi1ZHNQrFVnnrWIJFnjjvodNOm5eHbmAfHW+
3V9sVBJ9vrC0rwtHPw/8lngwW+yBPCzdzEsyfUgsA7aDoTKNV+I54F6oy5LeHVqK
Xn6b72Ld9YmqZsDZTt1FitLgcvAwndUOlGYDe1yXKUcaToHZeO91zW+cEuFzs9oS
jTOtkI6Hvlkb1ypqqCgin6Z2/dnUBHwgagrWU97uYXdX0QflAm5abTi8aDzIUG6o
bTXU3ni7/CjNvLZbpSDhYDIMkeNwHKDs7fpOHF+zv/XU+no3fPSQuS49lrtwnJ5F
bChrD5ws4LNP9Pe3x3mBd2RmAkeCt2wOJWQBlj7M5VArbdVuc5UmgRXoGcLqiSUi
6qzS1Zu7+cqMyXoa0vNd+ETr0CEMfSwIGJUItk7u+t/OTQfD8nrrg8FoOnWJ4o8t
AS7hr4PLPj6lu8JQ8sv0mceKQ92D/YjRIc0pHldaN/Ax5+fDUFTNG5agMui72MQL
EPJXmKO6im7Q5OYSNgoBVT04lOu5TWu9xk4jdTmtEMlgnX8UYDwKbtdSonw4fbRG
XPVGO7d2E0crZoPSOWC3bWYkZ2RsUekbd0VGgBCiWD312S1aIuQM4MqylsHJs6lk
YKI/H3GBar+ej5CWECq4eLTYXtWRvtLvkDUL5dQHG5Ofw7isEqhJUoZgkcn551++
TC+yyM4TUJs97MfTJF3OdZVY3wB9U1H8x9GalCid/59DzfcLfecFbmAgJnPGg8lE
NTChTfB+PWSfJ+q6kRGHbUgpEEqg+o6rsWiLiUNe6KFAjCG84TeeQlU8dXj3tOex
KYkpPubZmbvGoIWIEugXCHaU7RKdjO3H80oy4ZKC8xsFPYF+AQJKqRwqhmWoR9Rw
FfBbbJMi4y4GiMkD15D/SIJHNB5SDv53bOnkOXMfYXbAApKDq9pMS9fj4YAslcMv
fN0fIIiU0VkoYRdZKajr4Kv51yx/l+Gfz3QguU5qW7L4BMYxFWcmtOUhiOraJHjj
ObGCWs3J0ORLJ+LiSSBZtKbJP5P4Ah3TT9Kjn6xrsAzvJieYSOjoryH1PJi4PKgW
6R00sha/DPXbTW/dmCVSu+dS7p86XVg6O2nSoSUw5lWGSFku+XTaqNoFPyt6VC9A
4TLcscCjUGZkvDGjrc4z78aHvGPiTI37RBpq+TnEt9hks3GN85fMgQOjqbjmZocw
yOct7WFuniZCJNLuAkYIuGsB4BB2nPRUXCiffyZ3w/DEtu1NSATKJ/6p30WbSz4z
jayQZ+B9ORPFyngsBTAIy0QbiKAgVSnf4UhjnEHPPc5aObLT94/ev8HdZdAKGAXN
W8aMR4u9A+pMl/zfYg+HRFhkyjwp/yqd6S/tXTPGaGyCNTvAEhtt7wBsvjxDwdsQ
AJ2wKCTawuDvwKtkTk2qsAODQG2z0WMSbzSyNuqc7ajdRCSc7JjduWLMdJfbhKU4
FnPhkIWSRSxJ/BmG3O+6ku62CAKblL7ybuJdGkQJKfnwi5HObGmAx+uMx8K/ENu6
j+m3L+311Cx3vtfvtKVbdvEF6mqJSNLv3DlBpEIcBrv19l+zuIqb4DXIeaecfM+G
msJ9dZ8J4Kaooh3+iAb5CVA8BLJAAbGV0P26wFcJv+IUE5cPXIb/6F22LNr95xGh
48s8a+89swqN4SwJu64TPS4gubcZidIXSyTZ8XX7pCHAJ0CvsKRTjIi2zDs7qbGt
JzuyZ60rzhQOW2fLha7xu/4iYcA74kGEK49UFH6s2VPXTdvs25SVJBKAqhugLEGQ
bHzwupX+8UVYQUkcKjkh/9WmdFY5hEp1ROmMd9rPFLBtnxTXNrfQn336gcf+EEVq
xLMVQII7kqQCM/hR6pKgnx2+oD+6IOSJhvHCokpJur7Es60SSU/C5vRUFSBwpNWy
a2IIl5lHbVdHpMP9IDfVhKHMln6Ad4ANPa1dP3wVsybBsqEGka7Sr7BUgAfTDP/H
xsDQk4Y8s11SCQPHVCKDMU7/wUroaSAKOZ1heSWvHy8YntaXCBXeSXmK26+gVFoX
2BpruiYKMCypBvxshTpd1n7RNrS1BDRyH1TkJrfnKGXdxyYZoNYs7Z5FV/ntxFJR
j/OpZLpjQ3UkhJfpMZJFgmqvkzULLdGQffcQlOMJfD5Jr/e2FgcM5REthk2HuvGr
Jq4QnFh1hAI7XWGDuVeqCWinHbP98RAXZTB6vZ4nE9Oyl4SISXdAdNYtUH+0FeAz
moaEzUskZoewOAhdpoU0uDVv4HUTt4e8SjcXlUsVi2Q0CmHODoIV6ubucqHB300h
3ZkBkX9niYsX5w+TuwbsdBWTeEaHbr25iogT41ej9aPEGnM86oVoZFfIdocqDx6v
+2INEQ+RaqptJJyo/43QQKp6GVXGXwqzlir8eV6tzQUvzpbdKFF/PWEQCY/VCrtX
cqs2598TdQFoCEWOodloJgpccbs2sC75tlYG2ZdCGOM3GUJULOU7ML/QDESo+JZ2
4sX+Dgkktt+MuxFHgWd+ZpAbtkaBJxZpVlmwHYq++lICGAG1GKFAP6/F93a1XFTy
0znv9zjkU54QK1sGJ5cz0KTBJkoVxnMyIsAn8i7NeGxzNcf61Pu7WmldjkI9plLQ
+mBnQdgLDDv0RYITpmrAB6Y9IbENzgoqGOhNo0FtAHbwmYijMNe9UOUR6c0JFYWk
udRSCnazgG6ExaY0K5LduZtorGeYDLDcjJTSgxV9AN0ju5PBcD6FypYYnyENJ8bY
oI3VgvbhE30j02+6jyvInqmueWmUYvSj0L7Z405boQdcigwWt6mReczjOk32Hcxw
VNbe77QGoqSWACMuxWq9yfWyCl8dPCHQ8U4Jv7p2sgXh8SCVYQ2XYVKT+/6/CYna
ai6H9ok3/ilsCGeyG+tp98Al9mIBQ0nQ2oeHLQslvSrSLBV/5cnkNiSfjQHX0cIs
z4Hkit0XmHHRj38Nnd5cJyADJzkWMC+JsOKjXvFJpt08mNlXRiFilP7A5UnyUgdE
ZOIhVPISW5S9JpP1oEEWFZS6p2dXzUSqm/jBbVClV86gs07xFz5q7g659I48p24E
GakpuCffk5iNZWfcRdEA4xwKz0vGHO3ecCO5gUPyhXH7SOULTCLDDC6F9SKxiEiT
ANIYGbILebNb9g5qe8EYbEPOqwwcCHJpbyfIF6MG4OtoqcSXhuH9/9HSgMmRfq6j
lTgbS8zaUisa5PKTJaV2CnKEbNyijE5LfveRmjqJhRire9sH5L5VYOvvnJ0HLPLo
aHOUi85+t+04B4V1RHoXvaJr6e1SR/bVpWHk0JqoqDShWzyD7m+SjzCbAeq8aEYt
wCMV722A2IxAipWpf3S1GHNJzP30Kj+Ot3TMhybI1a8O2onBJVilc2tLzH+wPBQJ
9XCtOAaG1T++AoWkyYZDObEEtkVZYmELH5LDgC/Gp6VMicQQHkMvBoFrnvnuM0zj
n4bDVKgUBv9d+b0YzZApC6/Bo35cagZ6mKMlxKSvb27GvKncF2tjGrvmOvlcpZkg
IWELBbmFGQLmRo6VlaVOG8ZbvOi7krEfIsMRWq5cIX2lttYByeKvq7UNIfho9kSv
C4v83wC1+iYeud8F9M+lWcUw8lqk8lHOZuDkhrnYyGJjGtGtoW9TrOk5LCoY1T9E
ksRft93lHm3cZOpRLl3O282elHwjrbMMFYr9YYY1I08YWHNRf5MwS4tu1Gw1jy7X
ziig0IxEHze4eYoRaOz/wB4PN6+rdKg0p/HIndesd115WiM+dGLKl5lDx6XDZoov
V/mnHt9l2A1oOKs8MgEso18BjAWkE0gSrko5Z5gmT0ke6IlC8EAEVtYTpavn6q45
tgNqr/k4MYXWiMcNhUaF41gJ/RjMAsrFu/9ybNZIKtNzRPU5wcWvRifJr/oR8Kdq
RInRpmpmpnoALE4PVPRHc1QHOGbKJtPa1bStT3VdiOp695CmiJ9+e++50lpRsGeM
5DAwHsupaM+KSl0d2hY1YL0WfwWuD6zeUrzJR5QgIO836riMZw/sURCkEFG12yma
jW0IH+xNP0Z78tXPYB3YMuRx1Ss3JJwantgq9TFlrdy877XcBV/dIGaujWEabP0t
snHDqjGfHatSZWM9YA14SAspiE99jAoi6qNrnKEKRLdWkFg2ImJC9tG2mOFNm65r
0b86zhzrlHtvcko1x7qchCLvLv6EA3soEm6+ra5M/VP3vwe52SW6sg7ca6tAhhZx
9AZdKiEzoJsIbi3BVgOVm0ESwRGwngCwvk5G+Y14uCdvHxTv1X6Grg8qqo8OF/aD
dStgF1eoBavT0zzNpdzgBTAmS0MJnQJfXi6F3SBC5NQwVRzxv3VQQabaWojpM4L6
GJCJokkuibD3MBfF6Fkk1s8HPoVfCXLup2WMRtUHRtOM9Dcjn5irmJwo8d1i4e/W
gcfxepdLT7yhUIly232fdiJB+zekwUmBmCVEKvUoupWP7UQZIlcijYuKiRvbLmYD
d+bFBY3/rdk0Cynz2J29Xo8HRuQkbvpXjleI61tDOtlSucH9Tn4rjwaPBk8wwPIT
pPSPZDgVw65Pl1uF6Fig4dpeBRM7nJkd8QEHwBGmiFyEfiOQ5Kd3xKQaYrEtu90C
ciVh0XyejqfbfZV3bkuRwUcRQ3rvTe7B7JJfIbuSGytwN0HPmt9dxoW3mDTsHZMD
8PvdhxuKtLiaz4Lksl+6lNWZco9rnShjoIZNvxc9tbshvs3bgAmSHWLA5PlkKzIQ
uyI2LzuEaLlatrSWncZ2KIdpUM9DGsyZp6Lw/Ql/FwKRX5t+gMf4bLMzyPHMljdq
nouplyNxz428NSZKtiBzigAAMKfSsr80WxvQmYR0Tz869hbCTKOtTyH4moB6t2pG
TYdwiAmdkFSQGmSOvQl6owqD1bYOo/yeagVlGFT5M7Sr0Z8gmZccRV7II+rRCnh5
gVuaf2U1U76+mCwrlyDvJPjaFOBafQzJ0ZUAn86JA0xyuaJt+IahX4yJd/M1yvbr
7Y8N/TifXNNU8F5PphAoB1iXZyp8at5c04TOlygWYBrJ7lOFny9DevcvIvuLYuyb
9X9XEJITzZrw3hIzAoVBANfq60NspSTtUOHT3qAz/kND5XUpat3SdKUQVRDYNewG
w+IMHvxrq+1z5FFFaL15E9p5tJQ1XQoPLlaex6pjW7LhaSV451Okk4n+mVIoyjuc
MNdqHdAAgP/GDKEpEl9HKLpIz4lJDVSF4kde2WkuGEiKsaM34fSsN4BDZMXEjv+I
TpkgF8aapl7hSulBp6jlwMhcPxblJ3KJMk/uvzI50FTWm6jlChzh1258uXVNExZl
AAkmF6MOUBF7bnWiOop0NEJU5gDoufuYJZPAMeRYRHGNbJHFlxVYAT1SBlxmrKtO
A7v46LF4YrTq/+R8XMR4PfBeBiKGpQKOlwJt5lE1RdDIVGp7r0L7FMko9hrVfMHH
o5EGK8NntluTpzm7JQH7WbkY/5HVV6ZWlkzISiEIOcR6p1AtrWQ6vqFRC10h+A08
qOaonD72/zQdljlMzHoICYQh0wkpywQnR0M3FxcmthOo73HbBC+2QaPKkp/A3lSN
iHLqE1Lr7Kliebh2LVV+cNZ9eaJihwxC0X1aIF1Ei3r808on0c+htcNcrcj61nza
TrAv+clNTZX+pjvSnVvrvbsyZMvqwOui9FGQ726hKxlwcjWqq9Qj9cEBoQV/yIyr
g/i7RYQvSeWHEp8jmTPu2sWp6nXXUkVmHUmm1Ri+1U+W0wRbSXWOS5zWkYr6KbaA
ifQOKvEPV+MOrNPInD6ha8kiQXqdOmeJf7LlflAgos4JO9PjhSiPjwmPxuRyg/0v
G9TIEeRitNVoLyqgjQW38bGulZbwENKNF1OLfSMk9ln06O6PTRy71fvPNlXVCl0M
PGSoCLxJsV3gzwb6sYVmUKL5YhB2+Gs3vf2+ppadGfpVjOEVaVAH1TZg2Twv+hEj
Vwn2WImy1f7K6eOyRmZvzXiMNh9fqGMufCyRzLGmwpNXnk5cr+DQ0xTwuaSEkK6k
y0RXmviy1scHVmSMQf8dv+c75alk6s1KUTKsCnA+EEAHp7cDgPqzOFNpIc3jhU39
QPYJt+aEPwlGjBAUpet7nI7htvnRO8XtsyJyYPyDiUbi7AWpttdVGLEXvpDlxkaP
LiXHCYYHQH4AxbrIz9K5j0GPMbcghwcUBL2+g8z5EZ5iDmdeIqSx6XXdTL1raB/s
mnRVjW5fAzA5JFEnnk2xKfBVjOOtC84hQcHGUVl+z8qQnTfTR48UWwQWl9vHlolV
zD0hfBys6L3cps8ZDsBL6d+DagNxhA+nTfN4VusyX/YG/XUbk7q+duJwH8VHTAPa
0KJzOw4Yw5SCFwfjy1b6zX1zNrRC9km9aQdK74qO06bX0KucUKCA3FWhjr3CSpQa
8uMALsWD4SXxLS8z1ZKvojQAk22KrUZE1h1I8k1wgV27d1e5qx/0e+q3O4M4aUSL
EwzDq0QwsYg0O0lpZiSx8lLFBRW5yXsVJzqe12SPVXXxFPx6DETuejdfcDGv1NBJ
lBge3bcopW0YEugQhtZ/cFuQ/EK+jcVTVg5lnc77H6MAsTMG4uaorJVcaGezr5CH
G2HYqd+qEh1kMZzj3dV9e2gwHldAO+Ugh92bPGKCCsetVbByOXawCiK5yjXFj6kt
Fr2Zd9ufubu5F3CFLL6V1lX4wsGkDtJf6HN0NfWaSj69HJxYV7RUVYESdoGovene
avDIPd8RLkkipU3qNGj5x3NvZKO80CZylTwWXyDkeYV/NsyuJgfPVM+tXlhXORMG
nfnsSbNNGVQObMG+dKKIqLhbFriXqsaDd0kisUMOmVF+jflzWnDHzm7zt7UlWFth
pLvE90AhxeE9qU2XyGqVaIfp89qIMtrosoANRmTZA7c5OQymcpRLJ0Al/4af60H1
huHEPcqvezbB5Kt59I3w9T9QK9jWBYeOnEcQhFNvF6akfeLdC/m4ZN7oRbmxQI9Z
+SFKKizgMXza3AJLYPfggm/XFa630bJvWWH4e47vCGBvDViBAVvJ34xK8wFLS3Mk
ULOhg3ac+CScWf5l8J17fB/0jYfNNlISVevWgzFDl2SGXEmX1OolSkk5SJhEs22N
Nmw8ig579n4G/4wjWJO4G7XKThwRZ/bgp+Yl9TiqmdlYGJWCEme4XjNL28qZL6j9
IWwAkacNZFDfIcRi+RLShikD+swyrXrHnyicHl3m8C5cWTQ2aLb/3QoAnsyZjQ4G
778JimChHafwnJuG0bRw+9ajAxfbg9GA7KD0qoz9O1lQWHV/TncHKsaPox6FYYWa
6Wp1oa6/OEWh8jlmkv5J1nfk3K1xSmXl3ozvYPOnLYOieAzdtc4EUzRKT0LyJhto
TKr0Al7ku/X3vz3MiaUV1x6oFJqUBuHnt0aUf8h63UySDUUCbDKcKrPNTe72n09o
utQ1pcPNPxrjjrpsfbp3unxj/QSl4UqOASzpZ3y05E5Mh5ttAT9xEXIAhckggwKe
sCROJlfzjg4bvY05cOrSJ/FYR6lsr/MT2sv40EDHfCSTWgdknJSvyxiHjgU1WJJv
zheSUH2mqVCWgrsJ/W8tCUyU0jB76xcs1Z5tfFm0Pjs7JSYeQWpouB6Ke/9tP8I3
UVpCqRJvlckxM4tfXpXJMXOfWVCQLDwnHCu4056juT5G43vOQNw5jGHB/N/wihXJ
c2cAYvSOSqgL/FjKvUbhqfvpLeRUo727kQDIQ5fRfnP33aqY8TBqzyANi/+5Y/TK
0GpkyfjPzcs/KOHEpl1nt2vzBCey9z0Mp9xKm6+rY2s6AiKfJcRu+IAvSVJMXanp
tPimeoDzErpDbFBiIuHFXt1iEUxPMiR4ARVR3ErS51kYeUhqpdVLwxKOU5srMaVz
af+Zy+qkH0PyG+FWI3Gf0Gu4FVPUHUG/wcainSW5PXISmL0hIiFwnZHBAqXWzz9a
xlUiaDvMgvWxYcYSoCnwApKZTZDNfnxsTYV7uQmsY055N2FrJgxBUS8dmEsPMnIK
6Q2FoLGeK07Zt17BKNCtRfrwKTl7ZP15FWnJ0+djfm+lYi/BOsFM6ELh7ncxKfNe
dp47/Y8qXsh1Gq8a9zsnJlok8O2n0cgI261ensfTHgRXIoCCh5QXhEE8hBybHvY2
tlG8Esvc8v5Sh59Qx+6HA4iyHWr0g0Uoq2MzXGMbR9jHlqFuUGY9GXDG3z4M4mt0
obyWiKdMOAqoZuedU8+YBO/hMn8xY0gRHXnoV/3mLZofIWBr+WBBr0KO9lxtgOPB
mNCQx4ReHRf67QiA+0j0Z9q1RZDE2Mo56cOT5aPSwxKiS8mUEKrlA5XUg5E8mzTf
beUrWpXw1pFyqVT1Pm7X99PbRlw90DzyyhupJ63Z8GYf2nHCyfJotdlZWHiOiBBP
LZkXTXj1fO2GUsv6p5j86J82W7th8cSWTd0uQ9eIBjDPWZDBBrI1KUYiqNPte1oh
K3wnuw+tX+bn/sipj7nohCOZrjSqKw7ib7Hdu7XlyXbUApF5BAe9WofZ2CX6W6qr
hgOJUc+U8eAeA6eXXeiAyWSRzoRoqyMjm4yT+3Jq4a2HaKbGKAceWDgInI3yGvqq
3tAdWqsd0uzO3a/3zkBWPmwSV8tSJ+ogxfGUtfOjTWzsE4oqUPplm0WPJUJbZWo4
VPQQr4+tij+2uMgna0ZTkzWAR4CbTNBKRsNjA7B8QwgaqgNhXFy68WuPQ7Lhsq24
pHf4gvfBiIti2/w8wADMXaOGF/9LAU4WQSFG8hHGp4qQTQ0g0hnU67ss4s5NaYKS
HowtBhzXYRHjghpSga0UgvxJDVYKQbVbwRYg8JW9ULTLWWU9b53zzSfGRnp5i8YN
9wiYmkxnllpLL3y4a0vth4vGCKF/76c4wb+4+5rbtC6UqJbhv7oAuHKfyLO4hSVg
zyAWEfzTzH8A8qcgSpN+khvEDQYCL60jKZY7toq/T2SSOVyIsfdh3A1f8iK17/mI
QEa9iP4QnDzFcvYphqrSd3CffLl1EpsjDUPkY18+ssfQjmIdgtzFCzaqjoxG6u6d
qToWk4I+jLUyoqJqa8lGC/6Ux1GlwKTt1OXDv2nCwhucmoqzHhSnbycHKwKZIR3N
Q7qujpH231ZyE7WMrpbt9d9Hh4WqK78Rz0iz+tawuZj+nGsElzld7jxmi+braZPu
+0JVRDcGIW4fp1YqH6b3We+w7Z9MHTJF0RVKLem+K9t2P27/wAITWRq13KHrlAPe
8nebVuAqEJsWgxVPjq7iqAFLCHuibTGq/ds72UxKsOYMUoVClqugCj2vLrznZKR2
gkKtwUrmf+MrP4blps6sFqWw0MvOYpn14Mp4TNuXnH3iLkMvhKdtyjGth6t6pSYQ
/RiXDo1Ca47brX9kZnvmrM0/jql7Pl7tK0UpA9qR6MlFs14xuo5fjGpBRgOFUpB8
+2O/CCLFadNf3ha8gYckCt7bLcTiAvZ9xZsdSCggwnMH8eAT2Or4PMZnJVVHZvBL
erPnR2L/BCkCevTSs+BQHdXMdopDgKRbUEU8keokX+0QjQ8g6F+V2Uv36Yk50buX
zSnqkZ0vVfoGsPlcF42kjf8MBjNxflV4C66aPs1chSdbGEYgBGUQAhKBD0Bjvk96
gjU2GjwlqaQOGptgDCHxL+6DK57Cq6kREF11r76UJCFBYwU4GhotaozBNeCNuSWD
xJTwZEpNjxxyBpOJOD66CkneUIPtLRY8tctM8UsJNZbOvdTHrRu5VWKLa1VKqnW6
7ch7gUREuFF1WGyPwwKeDqkPmoSbgna8nzXK/6RRbruG2eF6LhsJGYy2nfAeH3oh
HJ/l48+Txn5lWKGrWfJIX0Z1Z0BMQ56gaLMsvTcne+QTZNLTbowg7RqdFum2TFEA
uzu+A07e2qt2okDF/QjuD2DczpofaUd7AClJvmPkJpabUJOcduXMg3I8dHip0zpo
17jGj2EurejEIeij+dOYupB+3KGOjTuZE8IqWHhlUIBmQZvJDCXkz5xM01fReG/8
aS1YsFCi2ViGI8+S3hwETQhYL9npcdCdvDG+kkbp1j5IFVHHeGfCJmTXD7V2u/+d
IZe2UztsIB+qpoRMgyAwMU3gTqSDEfqEcVvLLUuF7hW4At5eJMqI4DRiYdaTvWOa
6Spdp9H1xyQoN8ad8Wy9QIV2NnG3p7Umdf9Igzp7eRPUskayOl7zwNXCKR7Mfz1E
Y5CE2EOLhY9UascBBAy3CPPy3bXDDGqZRJiE1Gv2RiujuYM0oP6b8Sr1a2w6yXxH
vmVg8AHBMJV5xsqcsLXp8m6M4BdQq1f0JBRsGuPILgVLkwV499ZMh6jgiyXO+zN5
QkrvDOoKcKfTjdlXP2KEDh9bIj0awab2rB5eecnTYy0lGGh0VKc5RnOR6lCmeZU+
XdKiSHgQP8wnDnUgSb4YHLqc7csOkWmFaY231rQTp0BhRKtiGIvbOC1oeAlJUd4J
le0S6S306NnIKvfU9Oo/kpeLxZd2yUmPfyD41HMuB43PVvLBP6b61Bm3UiDDlE3x
HtBpGfnXM7La5wk2EiNL0Fo05rwbD2K7EVDce53tPW/5/sgSpHG5WHDZZNl0lYjj
EWocxEEI2X42uHJh5/NxaGv/z5CL7Ca3hPATfVSTlpIAb767gEgf15pNL1E1g/y0
`pragma protect end_protected
