// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:53 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eW1uaW2ehODFbk9lwJicrsMdva7vcgKXjshSjYijAuLSLMrOfUzeuxxBT058hM79
Jtno0hngN4CPa9pdmd/ILj1jPeEsyaFN7mqxUjfY1iXozBqWxuRA/6gYIMpJSWj4
gDBhYKry09W0YBspuv4iiqFnaZnCL9DdPTXcSYLXomk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10064)
tcuh75lEb53VHI0YDouilowbtPJRItsBHWLuEq5PSCJgVfZuBAF8bjgLonkiu77F
UJBEuxd3CPcV0NE59VNfXrzDWV8DjCKjEATmzoGaE7dkjjuHFf+8I0B/KaHYXi0B
rrvQZCrrS7FymcKGyaZF0uLjAmy2ECMCDBPaMu/dCiYOgurp0oaShgfume3l/M99
XW5pKHtt6U/V+owbgwGWqcqekpqvMVT0cm0eBXmN8crUlmX0UYQns+ei8VY7VsPy
Upt3bkBxOYdrk3SlA3BEeaGDwxvbNLswwGMkAibUDWyNOSz4DakkCGo7BaB8cocd
5MyckcAg4M/QcDPJLIpn4I7MzhXV0w4llcxvgs+vAcfHaYlv5I4u3Lp9YTQY9Adn
fq7gr7aO7TdZ4hV8Aacj3out9/O2QB1QUtx24sw+xg2D0cT6wApHqxuqkciXziWv
pPnIBuFAV2qYDItN/4usIrMfT0Yuvjr1I2y+RKx7LMPGyHNNN23Ubv5xIAHWvi0I
v2TZNaHeWEwYDaGVY/ufx3mzGiKAB2pNHKrrXpxiAOhsoI78eJ0GrAcv96KKKJXl
HZQScn0EUjniwZEmfHJdWj57genWSJWecD5ag5KHWjsmH6qv/w/PUR27Lw7zcxRz
2wOaD4hCpLhotexoxggFtg16eLEAyp+S691FB+mO8Xl2LdtJakodthyIKsGg5l1p
REY+0pCbKkVsRS2+dJpsbYYy8QRwLbUzLLSHXzAZw5bt3gVZX+a97HHw7Pi2HKFA
JBchciJZ0Olaa9cDt6yFmvwUFtlklVKIUBZ64qQFPj08z7knq6rmd69QgR+nY3Md
8DfPmT8YGXzZWD5IUqGpvZ4klwBpYYejEP39i2scgnTrlxz3m3gru/CsHgS8NF58
wC0qhPvsQ8nI/OmI8p+tchuh8BKDfOzzhY4RPzobgdH0ZIGhB+OJq1bm0hT8Pm2A
OkH26fgQ6slMaZBcVsb17AYpjk2tv4JHPYKZJcNTLsRv9QOLfyf8wT4Ds+BzA0Fr
4EdaehPmXwFhtcO32O1nzaiRG0wWhvS7YTn0GVxPuCVZNTY2+M9hRWXvYuNqvZTe
cS9rHz5A4UePIDXtHOLG8ARLHObJHWeFGhKWcofUSKSj2xJnCBM5150a0SncTtgi
l9tcT6p7HDn+/h5z1LCNvk2oTD3GlfH2xJyF2dWwdU7XcEHVMCzratcICMJ8tCSf
UB0r8nNQ/9BqOwEXUJGG+yAcGDHHnBFzx0wVpdoCfrsYREjs/x09u74+pu3n+IRy
dhwAA1Z/3g7zC1bZMuxc8WkhbUhif/ABqwk2n06h/Alqn2k4NVAQzLB48gionRcI
fjocIJT/h8d69djSetN/z3ewC9dIZzhwJZFHOjd8x9Qaj/asjf9AWJEsTh0hNCwg
1oDK5alK7mfCB7trsRSFgNJnUdBQzxOOQluYROnPbsjlYX0kARfxgXhn3MS5yl6e
CwNzpW5IYb32CvWUYD8FlHMnimnIY5Ln9viGgBeLQLefj+j49abKtClxY1BQWm3d
iHZJgPIPS/b+YHaVZOHj4j+j+5UoG+sWpOlR1yqBMq4aKmPAuFnT0XqXV9BlT6B2
T52MsuHg3eQqKcfuH1LBHP/nTLOBSyageqtTKxbM7pE+GEaTPVBdUs9OYXa7vjg5
jmg0P449yj8phpbhOxKn4pi3cB+qk+Oj+ixBG0IRr1uEkifuG9rxliI8S8CbWb34
Gc7iyY628Q8epF5zyBP0yBJ6TXa0BVi9XVjD3DEmFNV1KFiBVdVens8/qztcQVqu
t5WeepxZUYz75P1inUE7f0HsNNk1r5dEKPfxO90VLsFmsQ2pr5D+8IA9FR78Em9U
HG8V0sbU6qOiT4hWtzeLAhuoahIcCvAATlKMNt93kACvFcHnaR3CzNELhOo1YoTB
TGVctJ3dqfid0i3kSjBjO+Nwy8Qsty0pGIgkeUwl0Oz1X/NPhEO+5M0RguwmXjj6
mgbmB1r7JEx6FanStBaM5i7F3DbOhLhGpY7r49vZhx+GuIB0judC1/9qT1eNJGS8
NZ38WSWMlySp1pR/OuPKc6jop/uUtYF4FzI5sWoOWz8Z748TOH9LDZoaBsf+dt/i
gOkRb095VCsV/lrZIYKKdWXH35Om66jBIyFLxpCYYrPf7VPPhLejV+AoNpLDLRr6
NbHh5hJbyKBr44azrF1yYRHXu/tk9YwisONZ5NT4YeFHE6BAPsW1smgzha2aWj1U
gE0xBjnPFkFj4m8XgzQtw68jMjFEswqjOGHVjHvFGFaiwRG6w2azZteEdSx8JKJO
yayJeuZz/abRJ/kD9ABwKgNPRvHYTkQedR6J1nCRy8IsHj5puvyAx4Z8YQUtaGZx
tydKVQK/xmrw1bNC2msSmhv8OMJZW3Ev8LWqaYvBkx5U7LmJTC/qKA1b1vHtURXU
D2kizHrN/+OHQnPS8z6zHstjk7ZFR2b6vQcMU4uV60bbBasg8+ttsFdDpFRsrQWc
2+vxtqsnNHNvPivu1+BZmiv+OypVQWPYz93Qbz39fH+fczZRse/Z+Flp8Bp8GHfT
XqnkvlY16uJg42U4OqXRfJrS8g8UHrj+s85eX9pJvCIAfY6yhYclt5frpHBURl3Q
2MILr8Y+T5CA6CXPsTT4N8iW0ULx4af2PDeADuaNcdboCAz9sptmulwOHthrBrkn
kKTTy6O737EC7Pb05y2lr1QGKhkGX7GS1qCphZplVXSWSjjZ6a0Ax2QHz4GkYEum
D0bD+zvJ8W7zKgoDD8koct0Ma6cYVjZIn8VDVLPuhxtgUgmKi/QadScxtOFlFmMM
BsYwSGfzikc5u1KSP6YcU5KJV8W2O4R/mew5mdwB9NBkea99+vVqrUqm4y35lJUH
Fn4DoRB55qSDk1vfwsTObRUtGgC1GJz+t8feh+T+fhntQWTTK0kKq6clRcNGxZ7e
xDfe9T1jVhVs5wVIm0FHUIYK8xuDPdHne2++C2lLG74tM4qvygj4VCxbFGHJwIYx
Q8GgUQevhXsebIZcFJLgzOmoecCVNt0r3OTLll508TyGQ682KCVCzeWqI2nxLUf/
tt493pY2BIapBzpQyP/39STYOIt4g4pg0xpOAowIoZdjg91DmPjj87l1YY534uSu
y6N/txpgaGg5RAoT5w6c+CAe1LjWUAM3KDCcv2FbVUYyF82geZoGTUq8OPXoa02U
QzBIC3YH7qfcfJwSL6qqgRd8p0xaWgV1AItkeI1a+zJaYBGbXgMASHl+alJaGaTx
cyYvjmu/aeA4zvavnTdtvLE9tYX2pgPa1PtClCpYoAI6VxF7lE2fPQmtM3TlR5Vg
2MIVUXpoYJwkd7LqBZ61zHu/Yd+d3AntxULk7JcvMY+zC8F+LTu/XUfgdCz6iCq1
GtxQZtvyGMywYJg8nnY7gqZFDIwlMpt6DXYQLkQTjdjrerAk9PenVaP3UU1xumk6
P6TaW6FNHwu68cW0+AA4Qb1qoknadjeoefX7rPVZ6iDyNvdq0MBZpaPwXUOkTJ8y
5S47hf+tzQkygRbgVI6uIkEL4w8zEtuDtOobmNGkRTQ6Z6DO/AjA1M7WM8kQS5Qr
QdWIVcPPN1zf3uDA99DQm2O6fW5zRtVoncVfJR07mRHu40m0QwuLWLxywiL/7NI1
zFP3YRY4CjsOuVAUxYkfr9VFXxeHT6yIlmZdQZ80NDOABcAq0QkNavne0AvMDKT0
R/yDAaE2nmSFWpWSjIm5sAOH1tv3ZTjpDxKlEoy8K61TsPtrK42yfBnO5z5FgVIW
uYYdLW2xd7sxfZQVUmYdsEbNtQfZJXj1nm5Jf5j6unYuzFipEWRhOlbZ5sX3wTDP
5IDaP+KCgUqcNlJVfIGgKUGBOmG9HqbVNBW+3j+tKrQcnlNTlCBFumvbzcaD4Tqt
AL5u4mjcI3pujacmxXL9eS0YqMy0B0LAOZ+jXpcbluJpLNimRFpCjK+FAirBFGep
TLEkedIwsp6HEnQltDmL84AwuLi434HgMrM6QN9kA1HntIAkXDaYFFhhGjgBhgLz
2vIAbawKw57PadCZ5lf77TIJAMj5pI/WtFzzh0H4CnHrnZM2FlTlKpsBdjVDy459
/HYRunlyUnoBLUJ3Vua3wXQkavKBRihSPLNDyy0ZEwsTr9xX6mvzQ/dXFCAGhL1s
GYDh8MY24wluLQ5Ykgb7SUOFXzaNKCJPNvt5HgRolE1dQ+dG87S0uw7YsG6u7Yci
xcIk7lE2Bj/VJzI+cIt0AR7lSz+5tAZLb/4LJoO5yI1eaJLbJmnPhGAHUtbR530L
KlEG/1KNRZyU9/6rC+9UA+UnQ00tccoWL87BH33tYnZEoPkXz42SC3FYI0x+9c1f
czhPlVWlf4Oads90PqEZiCbFsUxI1Q1nrhCtQWupWDptiOfvsH4pWQMn163cqbwQ
8YG5Dq/sZW8HdMaK8x8ki3cMGL6ncEn9fz6XbemA3LF04SQd2HYfWHeEw6eU24Y2
/Bfxa7aYflAGCmX6Ne024YypVE8X8fKD4Nbr0QIx1sZSJRTb1q3BV+IQJFT6T1hp
r59StBkOi5Oz3gJ0oN/M4rXtWuQUJG57pm/OspkzlbZKIAzUAbMDQJhIdLKGUxSB
/ISpERy4UiIpePjKAzkxT1dCyzhlRqKbwr9DU4GmHpssQ8ujWQJVbIrkDQbF0qZZ
YuQu/Kpl8aRqf98qZeFl3/UATTLLBGIBcUz3p5B/8JwVWObDOlUsFGJ5Ee7X63iy
fSm9VqVCSDKusbX2e6SpsSgvNMH5w3QfuzdYI2Yqy/rE8HyGGZBsm4sfkVefbACF
DdOa9A1pvlMGl791Rq7/ocwjBefGqkWgESJuvsITrXyAvgJXlPgTNa4sgz2AHESG
4t8aqxciDBLy6lF0cl8H8QH1mjWkNYQcaIgzWIDpJMVqJP++bUxQVrnjqH+mKZ0W
o3U2EzV5YsEphvPS60Z79ugGeM46H9pCseS4H0kCcGqlqLLbz+W5pgDT41nluNsw
E7WcB7IZV/5I2QSKJ+ajaXOIX7WjRXLX1s8tS49pJs1NatcxlLaaNVvmklwSiCh5
j7j6B+iDMVwrJdmqJ5xF6ir8ijrbzRaDhrJsIFsNA1WIXBkpQVGdzNHpD+VWleAj
W/lFSZbnnCJJp1vbbJYPaHIy/ND6AjpLHccyJQ8MlLmdRzA9nflZjmoJQPZK1XLe
gejNljShXYa0M3dCeUi3Dhi1u4aC/qn7mGBhcUKK/psQMOOyW2eWHo0p/S8CH4bI
eeLadfJ4/xRYTYl3U3EBnJKv4SJenE7dMejnRYYBAB1N/0zt87nI0/5I8NH9s8W0
Fx65mD0toMB/7xceerx7y1VrwWPdMov70NGMXNqCGOkySXRHLv/0URhRKcM34DBz
eDeR3g4llEcpGPVgZ3FZpvXA8PaMyJRSqKIh6L/EY9rWyup4HKEo2z6kXiQ3101m
G24gg9cuHfZSqYIHBcaEFukePRQqjrD/niiUiJwgBNGVH8YwemuuuSRq+CDddyKz
IRKY5p1xHVqwYHtYckNgJK23izVr8y33a5MnX0PRQDkBYp9rm0yiVpolTh0f9wZh
6cQa2eHzGWRvmRoN1f09Adv9vSjm5tia5BPS0tSJCzot869Df4zDo09aI3VBQLul
aNoJwxw7ZnqQVtE6p/KflowM/U1JbqjwEEpRNzbxPkq53Q4RGtc5LbV00PxLMlzO
5CUtrTxV/Ccsl1OxPy1mNXZ9ibWfkdc2FCXDU99JQqiEgpVBoSkkEnw2gPKeHl2J
DZPnmYsHzHaCL1Cxexq1EnvnZSREXc72VLAA0CraH/HdsfBNzDSB0sr0a1O6Lg9n
nqhkPd3aVBfGODGCxs+L3EiLxe4ZBXQjabbgy5GmE4evgBcjYhVNChx/Fs9Z/3xD
dr9ep7iPGlWeKNYkldTBugcOjeoIxSS3pET7xeCMAsdPcIJX8PxV5scsJUUdAzar
yv5SHpmprjxIrEqUr6oQusikD6iwBI33ghmee7XPNblqnZxX1gbZZFbeyjXbuamw
80Gh76zpr/VRPe4/fvXVBe1n8CpPe61/dZ9KnEd+mJgVwxJqyeAYoQOlVbZbAvrO
B8ghst70E6uIaul9Wa4eaHr2eMEq7DwsrOyrJW7MbOcQjCPdoRgAi/Hkk5KAwrBl
yAL1NdGVcYOlfWIp/8kHzu+EWakqPA6drNuU7dzBr3ggVMZQhqiZuqXjhkeHindJ
wBKsN/Zu5GR+l/4ISG1Kytb6k2QuOsNCQLC6WW5IyX4Nhd9MByaoBrvawSqF//Pp
MSvMYe9NHNQ3/jPQcALO3FdqYgUDhUz99kOLNC7CqbHi5Q5BBQbYnsBnxSxa1+R1
8dvvV1AplpcKvRi6Jo/GWCqwTWh0muxrNrJUL/5am75dauzlsDvlvWAbwoBvB/Oc
D2bYWqxRoWS2kvpWF5x1xmNf5Y8hgnAbKnrb+S2bTMoZrhEGXFPyaVzIfMlgzNov
j7q5fZM/vYiBqHTtOu3AeXdD4taA0qSoEI4KeLKWLwlENVs4RfSwWxhYkbpC7gk/
vzeOt+m1gUqa6oNC/P8WDo2XsyHPcY0mGCQnzbcRkndPpf+e5wSklqNv08D5OTSo
0VlrntIbpQ8rFV1QGMR/w8NKbcSeYWUnk4TSz5eKrVLSvHgaJQly3HjlEB0OPafd
42SHBEGvjU8WZtgDfIMPNV3ymsGo5auBmoN9nDatFdj3jiqyNBsDwZ2SopstGLUA
4WhXp3sUGkGiUTMg2aTWy1uS4KxWz6pWZGPMC5gigO/OHhzV69FOZyE7STIqUDOP
h2XY8+E4ZL2+Nq2HWI4kqrvvQGANS2plqylfRp78PYcn2xWePa31nIn9jr8Owtm5
d/6Kd9A4N5zvta1+5DxiL2KFrW3QP5KFoF8Lk2tFPHTAl0rLzKDuAlTCN47AsmJM
UlTl2NIQpLVtWcShi5/jHvtjsRbXz4S5f1bAVWhkCe3m9FIX7pw+srhvM3BVzDvo
sKBLPuJq/paPicbeqNjFde6iAOC6gEKWoTy8T3oYvfYw3+NuCerrKJ4N/J7VVqBr
W8i90CdEfR/wb/1zCFRhAd6v/HlR07ZHnvBkyiJHEgYiCn3n5N/lbow/Miqrgb5A
uQXQDIZL67Wfwm+uk90FRMa3Nuqk7AEeizc+FhuqpB7UhqwHDuRIGXLrrcFdib7k
3coCK/KmbJwRmOhcdKb0pOT4/+W4FYXka/PmkBPM5cyE8k7XUZyIdCiyoLLAz8Is
1ph1fXWQsxw1CjgL3JrT8i7EzoOlVGVSAvip1nvpGW4ZSFEOrXbwGTYQDV947kKG
SR/mIA2ARVpPPqbrB6MYSorfp26/FUbJ6vZ4nho0yosMZ79FCTvWOq28T2CdRBp6
NDWG5M9T53q+zkfDDdCVU2cYdDYvhgkda26wFDgq/2QLLFDxCEP0grFQSi8WPYf4
1cBcjAAiJoUepfitLowWKHhDo6QNfm4g0ZQIQvPuhec3DdBrg/7wzVN6Ugc2KCPk
aEkCMOXY97iXT84WekfX+XxXAWazHD8F9IrlVi/irq8QACSBnUWLmiqyFHcOXJo7
ViXnY4oBxyD33BmeTXpVkVBh5ayxtc2Y917Q4Yoe8uCglzJzPJSjjkZPuspcsar4
lhK6YbM29lWf6eSjqo8z35Za0rr4zwEHtO+sUaLk11YkwYQFN5UsmD5+Y+q9ehOO
3t9H9GEXoL1O9XPVJQ+Az0dxSAnJjTAYkvce9XghRuJH4BrGzqtqctkGsY7WcJQS
TIdvke/RklQMV3s/vdpcVh4mNWzZtFXkeHpa+vH0ZDhchBPHIgRGMcU9b4m2JRB3
DF/bKDErbvU51Ax7BKAGPhqOjSRk8RQnA+sFlCHmIHsG3ryv+BUpYAnAPYcNRGf+
Mho+mG0zqwIx4i3o5mkr4Ine2nI+MADtPaXe49mi2Mef53ADDQRNmypSNOCEd/3e
hw0WBW2osvYozfKjMVoyhB57T0gfySR9kfPPlmqASUhuPMnoWA5YiOIqSjQ8QlNd
EinnQN+dHKNePXv6lyg1ACtq6Vbz2G/mJneK/YB4joCtAigL5v8hV/egXbNm7G++
9I1wPSH8cB6bVmTzSTztdwNhj24JU1Fxmwgl4R2JYjX5+0Ee4uZsjkr/3syxr95p
tF2pT5v5x+/Jyxk7kv1/5s3izywyBfMMoU3QpF+Wx1litwZyONlgjqBnoXm0U3iI
BzmcBLdfXQ4CyHvKNXrY5EPw33JWEk7E+zxEy50Dj7rxKqMcHhgQEuGwfWomt8MB
F6fDQSz4lDHp1fZDCbmmBwrE38eNHfmGT7DUlDOIMniqU2wF1BoOhzWqHflKfi9t
HnzE7MB4jXl6W2iO/nKd8bXxZw+fX6+N7BADdtweWX+DX4HLnGt0MZ3D+zqKF54c
amYbCi3lwoLeqEFmbnectzVfnZ2yW2r45kYLgKguRBJRRQtE9hFEGkLLJQMxNQT2
zKU04eS9uO+txnULwFkfArkDQzmb7wfPJPsQhxEjXstxVx8XN3ZZnrOOgldH0mEX
EMOzoIvYqiReDFoGfU7KXY4Unemu5VuZNjYMSsIbGSbguI9cYRewn+kBKZrvlgLR
bLpEPlAR+drp4Mwc+qcNV1qGBw5SZjyQlEW7S9Fkx5GRD+UKYGScOI17W3H14hNa
z1AUwcICxTxUR7pZjuqFr9L9ZqcQUqqr4XBv/PYRyjbjIQ7AuRQ6B7OnqLfG51TE
LovkcWGJxLSZqLsPo7qlkXPxe2xP6XqaembEpTLQaHNQZgRfbW6++MmYUGCBi6At
3/0p6b8ljq3vIvWEQfXwHD9ED7ac4Gh5f4Kg36GfDBTEGw10QOY26v/LuJIexruU
4w0BTHR2+agrCiWp31yUpWTj2HWwCLxYf96SbWb+ovKqKsY/Njhv/BCIQbDdTUBQ
/HxQNZKjpjB/a6BoBP6YlBLY//XAj4sAvxhPNa2hEgqsvcc8CrIm0LQFdV/uwLPo
5bWB1c+c4NgzhsqdoZFJkjtGpgpMGzFurYpc61TW1/vAvK2Si/eY5M3YviD3wrPQ
YbwtfeM6J3CsJOWNhPPuwDkhkLhq3toEJ5tgN3cl/wFssQYWbiNOtvnE/zdk83uw
NXvIgAVnqHlQL1TIHoMs+Aa9IRLMk+dO5a4AZg60Vvq3u5UMVZ10dvwoVRh/sm1d
bDo0hkjG9hsz1pyOC68fGinuZM/9EB9BfUGmB3bRVhMm9snhzg35yKAALc5O5F6b
2HRwNTxArHJwnw36U2Vbbo3Erf8bhjfk3ctebXxxiZnIS79/q3jMOXWaGl5nxm6K
IV2vWpYnupEJ0lJGqzbwJrse03pwWMPrmTj8arG26SL87ZxyQFDwWs6jF+JZVh14
D1ptuPJ5HTSqcmPzUCoRJDeMq6xcLmJqhQwbPpVmb9CiqUjb0Rtg8gvk8u7c67UG
5oH7Q56+x5+WyqWc6oK4I3G522UrexXjzoEGheMABfwTKFynrTAsL1UZ5F+JGHcZ
j+SYkZs34c9s97s3h1+F8vnGQPysHGQ5njn8R4PzuQHO4/mt7E6HZocce5kYj0Aq
Ndz9izXtXMFFIDHqB2+9mys33SXV/6CjlIVy/m5k8vyTSQsmiLe2hQ1X50SPkHx/
6lk3JrE5o5lIXvkK9Uoal+svDJyuwDK00mFUoi5OlGsz1xsZy10KZhOKxCSTWux9
lnlezfHia1k0tUNKRfUdGvQqOACOUwXIJd9zUeycuRf9G6O+YfD9j7Ar8rx9HoQS
qr1CAgrYABY3y21Kw4+oJaO0sx2gWEjMv+VhsOt7xAI/tw/0ATQ/AZ0n+zBdpHDB
LqRcZ8M3dbcyVKM7WMbJL9Wg+DqMxSHtfb7Mo+UjA/FDHK2V+2V60CBSnMHge4VU
Fef36eqanLiC03yUaAUgO3hzGtQaIKX4eeasTKKu5BdsCA4JoPj4E5OKbO34Kcd5
OuRmcVM0jgPA44nshsDDdINKwOILJV13LeQ6s39IEarfNGEeE/FlW/AvgKt8sgVv
TPLYcWjnINDfyBRpH+tF4a4q26y9xBQYQnVDzbAYCzv7X0VFkTJkRCaNwQbL1PY/
YjddyL1JvsLHoiMhu5IbTSIE+iV0ws38Ply4VNV3jGr9MKsu/ZzYKvvrG26Z3qIJ
aEJiHuXV/lrbcTZomHJs8dfptSd13xT5hQfFWL88ofc5QgvkdBLP9spTDk43J26q
GXreTQN9Lu6gDfj4SZ1MLgEA1M9u0WjjTT666zapyODLKsh9mXtx61MVCNUQJD9T
1Y0kWpF+C5hG/n/9GFQjMzR5Z5d5mzgcQGZDfLYL3/R3c8y32PK2dZP0n5W4m5hO
fGf5vwST01AQ7ZVAPEoIN9EwKnqdktieE9ODgH9weL6pfuqQoccaxfSPK08FMlib
nS6tOIa3LKF3LpGuytTZnfLdqOgnZ+bFQ9jHW6yjkTk1cWcEsCIsslE4VhNAISf1
rDofnjqefBIGbp3WzjG69NVN9M8pCr0MdO2nm+m7+6aEedViTAq3ri4BdRgd2m1m
CdxchsqIjt6bSaJyD9TvXvlv7cNCDLrsrmnzlVy4dw/LlXm6+fymTuHH1DUC57oa
g/QxE8scH2aicTzSTSUhEd4pFbBnuJVzyJMaxRY6ghPMB0VGMeQC1pB71FzPofDK
NPRrkcoBtul4c+6wP2q8C2ExpcY9Wy3W+w3HwLESmf7wRsIgD+g71INLiTlTQb5p
5L+euD7Esnh2DkBQFNk1gkrHi0BM54Us+x6SGshSzizZwrh19QhiJrz6r8m7mxfe
4aJHOYyiwuLXtBzyujJZQIRVit9SctFAnSXN6bafsIGeXkhOHrrKmfWqSn/UYQ7Q
O/Z4evFTGiTVqKD/lc4bpbRL9Q8Y4wv66qm2Z+7sYixG0zjGJXoGWOOuS+5Ot7Fu
i70+k0waJ8sj9V8l8vPm/WBQ3qhV5SpdyjNdrEdyefZC6Se5GsGenWBylCoCyyA2
VCTjAB0Xxu3vOmkJ5k+6ZbSjDxg6V7sk/n2FJgpoHr13u8x4GD3g68sQLkHsmw5x
Cn3paDUh2ReaFYFISR/Svg4fTOe7Rn52IJdI1HMeiL13gTy27ZjSJ4jTsGAiQWCu
Tf0rG1O2P0eBkPYoD6r7lPGDvr268PC1kCXCuQm0sI0PlagMtD+XLznyZ2USaUsx
ThGWF0Odfn5LAESu1cIhHRQcFdAkWBmqRA3oaIbPS4Zok+99Uwbk4b66Va/Ad0Ss
wPsm9ly/3UPefU4gmqAisL+Pmw7dMK5AbomPZuIfwNqAr0AxT+33UhXUQkfaZUMy
n54s29xcIHEl3NnjAQSj1HopbHPJZ8ZO3iU0yb86zzgX6wX0nqNAy5Lx2W8wyCl1
v38VwV76vQT8xV7GlG1kh0JuRn7c9MFaR5vT2cFpCidBhtSZcZiiHsJufV7aZrDE
hwd+B8LqcR7oCgKIAYhNBwgHoeT4HtdlvPegPvRBrNMJ8pHDe+oxeRsJSmkZtnQh
AUbXZk3jDUxpipKHMJ+B1kFoqVZUSZRwrJkZDLh5S8c5Z//S3VYeVbf5zl4UaXCx
teOmsBFGIy46i94m50mAr2iLS0vnezodKvEppl/RVgSnswZhcVvIG9Pttc0ihPrI
b2qRd876L1glCwoGgN+nSiNQ22kCvPYiMKbQ51X6VoXLFGlnLFg5ijYopd9Wvn3j
EdtSLPAMNtvcPBeORkcYJlYEjj46XsjHxi1yzoaN9SRHQ0tpBWvi/fvM9ggUJhcq
Flp3Q11HbIs0kWywudgv9MwRgrIKJkZbxySLdQyyeOqNvoJFgcbew5eCehg9Qp0I
4nWSQyH8ew2oCIEjelh9sy6/qA60ZZ3JAHq6C1joWeKBHiDnK+Vdioiol62mrvAI
wt0aoBU3H2NOD+FSJWFnyg3D6swfuh1D6qMnDQX21yIEIqxPY+fhyKoqdSU1SIaE
lUs7/nFVmVl7EJUOEToUhbsPvpyf8Wg2U7YSVC9kziKRvIi8N1SBVj1CGzO9ZaZr
/RHhsVKEAzbqyvxb89+KMFtRmLTxdd48rv/Ii5+p2CULtFHgDdiISb4yZnLyE1rX
w9Rx3chXayl+zMYm80225Hgr8VS7O3aO+X7OctwCtoVhyMsyKUWbvEf4tjQR+vbA
gaanTPMqP5QJ2uV0UikRgpxSMazU1d146TMu4Ei8gEK7OuZx8MOmy4V3GMi4fUwV
is/QlFpYewirgsJLmCykBJTt8XExSVSTvByw/sQFHbrljXHmqqYFJ2r0w2eiqtyG
1lA3Iz5hmvfS9YCJ0mQCl9l933C5pWZbUuFIFMipvSj3kSeEAyJu7d7JHSgOyUI0
5QXJrTFiQMmKVATmZnOWXO+yNlJVwCbBL4BcaAMjxkfols+/xIZt+d4b6WLyGBhk
/fCYTAVjbsHlcbagQRWj4ArnbyGDSas1oKpok0EhEdVxERgVVdJEjbexeLJup5rX
cZzjI7D0aaUMoXcbPqQ67uShEmGtdxP2GAvIu8d04q2dN6v5zfvDJLYcjkRQY+9P
i0jKHtfFfPfreriRsYydQ3nEGy92T4t4z0muQR0oaTbUNrd2m8sr/o2ZjhLt8Fv0
H51qNvRjJ6jc+6Ln6u11bDxIcrk4sqpZmKrrkonk4mvHI59TV4iypZ4uok21Icl+
VqEtTdJCS4u064lPlkxq7P69iilllfnhxGCFlYfPpLKCniohdsBYI47SILNZYMzY
/my6UQ4Q1zfE8Ws5nNVOMQ7p4AcmZ+bMzcf6aDWH2bgpcM5swYTAHfV2zEq8mJ51
JJ0OUFFtEGGg+FQR/4KBonfuaGEWv5UiRX8uJI6KL4+xPX8g/wa3H6Artew/JJwg
ZcaXQAvlQ8b8BK+4/rQaS7jGIOC8PLuTkzkkE8JPupwbXRJfLR5IzfOw0F1LpRnS
aYJBopV8n6P4wQJ26nYwuzIgCbPtLvAsySoqDHoG+0/xmtxEy6m8c+xvu4pS03pw
I1ImyT4HlpwLzZMCLZIayYLctgd5qdyOqaaC+r3Aq/a0T38jm5IDYVOw6pPPi2Xf
8C5B8K0SKQlhfRJukuqyseguNSpTmy4HzcX2BZ3N6e5mOEKFJknN8gdySUjLHcOu
EPwfzGtDuyyLWE63a7tFMuTuX9/s6sgfu7i0/FuKyaN4WkDsu49XNyBPdIdWkB3b
kWe1c/b/Pt7Os61jpa+UXPu/1ne1yWfhXnXlIBUAm+MQZ4Ot/GU3h+4ssfCLjvp4
s+scUSlUaM0L4wgEK8c/+eepenXbGzJoZugYnrMbPUKwdxmn2q7qe8Re2fhknhGu
VTAxRU/ZluZhJlVHtsvsCBHAFmK6weXlUJcflJIJjpk9pvDNldsYEc+bX6ztfyym
VEpkL8FeCZaNtSq/2+uuRV1J4keDhPFsYmzxdXGHy8xke/hmQ7QTXCEy6Sa2OWst
NYFl1t6fyzyiSz0rjpcGCd5uCKgdksMSCy7qqElc0xE=
`pragma protect end_protected
