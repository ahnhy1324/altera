// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:52 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
D6KvfcyNHhLT9mnbsUcrDl9UpXg2S4BSDYmIgJR1ikQ9sbJNElQJHDOMUG7jqeqD
gM7D8Ay89bZIir0gyqDt9ANBa24WLxPAsmypiru1Et5+ZwuOUqkEqWz1pFoHkPXB
VSj2dgC4dci9ryiS1WhksHE9yMn0lBU6dcRyrNXiWxY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8336)
FjXI7yYcN04dsaLBWBdoIyvDSFFXz/XjvF2dar5x68oWwPRqv5H+5qVUeLoqJTC/
L6hkQyoJ0fV9vYLllDg53DKexwsA4oIUo+ynP1XztRilc+j9ZLgRjqLFtmJF19y7
k07wJAbECFbPOle8JKy1qRecYPukxZZddV8Wc6el5wz5esdHhKSuOU7dd4j/mW3W
sYkVQnHRkvDy7ciRY6MmYLILwSyCQxWlQVgTkSsMwUh9KkVrlL8QiqrJDfTHUPvO
JS4HVc1U6ecxye2Hu6uJq2ZwNhXmgoWClxoj6IUZuXRGUZTT4oNA2h/h9X2c1qcl
dSjp13/P9x0oPItQ2l97mzE2fMOksf081ZMysOUu7gibLf1VLHCz7FiPckvkuCZ3
xvFIlEiB1rTSFBsmfHUzhUo+q/Wb1XX/FALTk/TxtP6Px5ke9H2uIMt7WDKFtOP3
A5wkiex/SHj9o6wKUz6N+sDsxwAzP20muM6tykjhU9x5L+Ew9r9urDjixF5872xD
om99qZqAOsWn/KPJlKk8OP7y2qbkNTQSlui4oQAXjg/l529yB1MDH9UxDGNxQet3
9UJG9naXiXtubuGvpYkLpcv+rYNsUJklthoUZy5g2KSwT/lqTD6yLTSKGWoUOfSs
wPUt7t6ln4unT0pb5e0ng/WGtZZ2csbhrX1yBzt5p/XyhD4KdvFRjSVWKoYwfTaG
zHCKjQZSqDgmCLJBXqpQWq61r2yPVMi7n5tPN66O/oGx4pUorq0w9JpYLX0CJGE1
9hLucb5NOgG8M1KnwSTArHemsp9EpyV6QMNSMuUrPzkb3w35GauR0EtvxK5YKUq6
Beo2Dq+V28oetPyxV6/X1fG8dpkbijGyKRXKeA5zvpPH/ze7/mjgO0rlO5CPwbzX
PUAC39cUxW2thn78Akkh4dQQSJu1K2V4k/qu0+TpWLtVKyzSdZK+EmlGRJ/Prr1i
lmm4NSRVcG9V81SLcsh/cI/FrmaCkNVd3w/4w7Tbo17Psgb8m+FubA0wlxAPxpUE
ZUwM/DIEGlrcDZQ11Za7IQa2Irs7bkMIlNSYf83mqg+s4pUIfoEE4kB69loST+UK
hvjJ3KaXxpjXHqoZz/yJ+UaE1CUW+2im6rQArDFZ2gO8pmYydUjteWSGxt8d+4cY
lrdkBzTOpolA34pDlZDZdFBj51CE7hZkI9n7jv7Yfec+YC7/soLvVfhdKktRGfPZ
e3gEM4OzIKZmL914keLm4BWrWYxFk4D6YoE6NRrVZ7HYXs9fDokmfmtCtTawk3Ck
NUO5oOXIdTXYSLh8+KqiMoUPOSaEwFXrhiw4FKVkB7PsNeuvjHuPvJwyitSTNO8T
BfPsgxPgVwIVMy7as6wZ+3lzlxsY2eAjU0iB2TbocwUdV1GT1xq+/dwYKS/T6uak
o4zbg0pkaj+JZkD0uhmDKBuB7Ny2u3lTEhsCoDWTou5mAspKnwvYc45Ij4p3SVO5
MUGszhT/sMbdLHW6LQYvW5ZmL9k8vTQYj+1xVZwDy3sPuUYzre5w3pzVFB8NisMK
9BgGLQOkbE/HkSstGsMEjhAx5Nu3F1uzs40UIgNxu3oK2/FhZX4DiI8OTRplNZcc
CRT7wBuuKwWCCB+gUYy/1ZEcF+4ONrvyWhI4M2Mp7My9HQ7xOjbUUaxB4Z1ofjvp
7kqdGirP9x/VqpTgkIKE+sdm+8+Y1Rt69MV22UNrKTX/rY+xytltboULZcE4HCmG
GClEGW6TOjUDSsYW+3IUxF73znWZQDPoXnB4OCNAUKimBr+yjsvd3MskxLFbRcnC
WNH2WPHCha1YajsuO75eCuy7sfoScnKHMktqcSOBdeoug58JAPKkGF6tYOe+btNi
umi85RC09jP6aLX7RrcwVVYYyjXbHeBUFNNzlZW7dMbwCTvz3o9Wl912N7Q38u4u
nE9cInAz2lp+Fj5qk2OG5wA8TZbwsTi4t3gtTxFqSt63+JQJ9Y17mraaFCkQ6itp
7mOGGCLoB7kiApD3Axq7ZcRR1AIkWxWGvOZfoD63D4WNHRAp3YuQxRjU3lKELXEQ
q5C4uTFJngd9LQut2KuJo/y8zByiT979KQ8g7bWvnnrmkiBSpaXBR0o/ylhpXb7J
539GSzHKE7bmYyYrXsdo3i/J+NYQZFkwUDPJNpq7pKEw0nSAvWWA9ZVkpyWjG5CY
EWLSfOW7K2W0ihEW5r8AdsCf/kKI1qsILg2KyVF8uw7JM50l3LNo1/Mok+MhFkw7
epyIee3W2Jif7kxVYj55QN0X9xOYYweqs6jzmImNO6FGaUBcd5WkhWdbyXx64aF0
ifuLbPnsZXN5bStu1rBQG8EVw65YJPj0Eu3bIxTL8t/OU4TyFj0L4uWUDWUvkIQy
1XcI83RbhRW4vHcj+74XcNZ2ZA7JYtX9XuHCMmc5mticBLuT9aIBoX457CX8Xi39
/jEQ2b94OZwAlyyD8u8v4d+HFzWvxzeRFD0qcOS+5Ugq1d+M7onKSNRRyxts0i1z
XWFScjGUHPwvQ5mBN+o3tAz5N7/0j2CdPdk/gHX/yX6nTAG3m8jacaZAzlDvUxEt
OFyZWrhQ03j7T1ymQ+7kr4gS1h5llzh80wI5A7FtQTGuJLuwVDHwGKbaajRMK3Kx
DSiucoZzkMpMGn9kUPQl4r7HSi/BBIZjHnNO0UFNBEhw8QqO3Q83SDVQRjnrDF5Z
TP42Bqbwf+gwfakuEPk9HxPCxmpN4z2ojv5kSZdtQkG45g8yPsoj9AdM8iMnAf9o
UPCI/uf9stQJqj9PTapTSrUGn1C90AuX1TZowGzsb+ppdHWQwbrfwntg7isZ6wTq
utqicEa61IJFlf0cDGFXtojWW/g1zQxjLRVwRpCUrxM2RpZh06dn4xe3Zs/2/Q2q
i65+zVfuAS+GAodqOvGTesAfv+mz53Pszcv15Is6gsxkANZm5xRQ/OAhk9xT00Oh
lzLQmu2qCny0x2x99RSFnMDdA4nVhapX9R+10pkNmE2lrlyKWGwz5BAJHxRxTBWD
ixFD1rZrknW+t4u4E71KkqAa+DjLPXWbkp/tinvQt0SacEFSai6+dKDaS0hvtC7S
67Oa6Y80PtxQStBKlljnW35c/gRQmHjhq0cuDo48U0UqvWmxpBR+Jr/ZLX19OPrs
+t8LobMlwE0A0cgbiTYD6vxFV6FTL7pzRtg3AtEguyF6+blIXLDqnzVv8IdEZLpi
OZPQaEZQHXFSVel0fe91mrdXloiQ3dWhg3v4nyPpOTsX0vozWcCBBqvkmzqJvDq+
u23e/KFT3Zxy2WPVGdZ6BDUylwnl99adJXDjc2XBtnetHIHAz67mxrpHoum5phmq
NZh4DMmcFQrjKOu/7Nbk5JmW1//J5/C5AIlRYqfawDXGte9112XZEP8zGUrhlPhp
12JtuhsWtbT2/yOU9b7QT29+Ff99WGhNkdUmBhmnG3urkzPrTsPzmcGf2D5yWrao
jD1yrZNzf/3DrcMq/udU0HFip2jfaL9duISiljPRr9VstQMZc8NylaDapZayWn7s
D091EiCsiWInXpLWh6WojudthqYTey1GHvU3j9jDxuOEVfryj2g1DwmXsR/hgf0Y
1l0AyMEO0Nr6jiJJXXUE2pPrfYPe5rI75oheeLAT2cWw7EYaK4UjK4tOpSDPYH8H
T405bPYecz6bpql9MF7EjIrpQKQF680OpCKX5yuYPP5HSO/YWP8ZPo/nVqTaFMpS
G2w2U3YXv0V4GlmzDWaF31OJGgWigNcS/W315P1tWBLquR1XQfg9bjwzyZ8oUd9f
RtcdJwnJK8FOf8dRrtyEbDEdEqthovTAlqwVh4KAj+rYCT20610h0iVu2Yq2YOQ7
wHFX4u/i3gd7nkN18buBWtC6S4Gc44l+nCcOVUB0ITdUjeC+Or/0Yr7AiBT0YH7H
i2PkYEcrethHZick04Iel2uLVSDoySWsQrl97jFUnpDkrjqqwJuVFEy8KE4mt0MB
UUnzgFp5z3QSBIBL1WMoopWKKJhhLYbKVi6y+slIf23ilOZSIp8RItpeJmvnLikE
BZCBuSvAPOHt29kuKRqmO8CfWao7ZTqB3axaygQwHHP7Dl7ZRBM+inH8R98PKg3k
GjTd4OF3R8Kcm/TF6b6nxFq1U6acBfSGI5jeVLXDsrF/c1ntJ3Xcq1Ax1oeX+Vq7
MH4T1Uk2ULTKfAgfGGAEkGO71cKQTK4wqPMm+tFnaLCNDX2pi2h6WaR8EhFm4vyN
OLDJktS9ZRC+PyHCRtKe48lrmK7KUVre3CK30Nq/KtWQ7GYot4l0aXh3hdT84fPM
GA51gYSYxSXAaOAcgJHFTpkM6e9U7l9qiP3eJGJLRsOjTUTev9sW1KCOCPfSv/eD
6+JSYXmgrff42AuFfqEg18tMROqYrt7R6Dd3ab+749S6Al41qWOrOQlygw+pxSKY
V9zp1Q1hi243HzgMqv2tG61ThqsiyA1djDCLZqX8Zqn3kpk6BqQhVpDw6RPEpTlF
xxO1KtVBNJqC//hbOOIfLsEKtUfmPYVbrzIUKo/rAjohFg7hqVrLfbLwsZjs1sSD
vjKTrvlYY8K2gD4utGy1RW5WgjDuo4G665Slv1MHllKs0zMmCw4smeqSKcO5C7+B
pNwBirVYyTHawtWBOanJvprpHytat8oazrCFdu6zF2NbZSx587pRrZ2GXke5naId
FiH3MZR25nlEACGNnEhEDLT5nB2oQjMISOx9giCEXcMxU7IyyJ7j4B11U+4wpkmp
zaLeWlbw04CF+vDAhvnjIzCK1HhW2UK8tmTbrGwEPib9qh18ZZzoB9F3AO/6EpM2
jyyz0GOjJlvSk7/UMvRtSolk7RzyTN09Ad0sifsSmabj7PyKcxugFO/bV+a3KYrF
OXgDTXlUxMvIm/uQ/GZSEOrbax32S6WhLNdXREmh4Bzh7DmXu54YkkoFQke1Wj6X
HM94RymRObri5jnNQe7g1hj1Xuxt62kTkbrxdnApXhMHpp/h387ZM/GEVjIcj85i
ktPDD6uG8bMBZpAaMnFCNzpkWlEX3/QmCzD72X4twbs8+l1Ble7TO4nF2gVbfBIV
UepsozThVZKX3wifU0wWCUz1pqlUrN26tDrQtgpEeQ5YazpO6G2xyeDdB0XBv31z
w0OM/KX8NbmilmwPz9YMEQJrH2IpPRFmRoCdr+pzGWtdAOF9ReIX84f6SuQZdYId
t7vjSbPG5gKgIC1pxAj52XUSVjcPrk3xumfk5uY/8pvz2PLVTlcfv1iiTRayHLYP
6n4ypKVmdCDmI0vAKpamYnMwcd2Mj3phT+vaLjnqOM6ealViv45U8SZuDnq/30Pe
+0u1tqMHOmyNIS83COf3RhcR+RmUpi1NQ9NaxJeyeLY4y8IN7FtQWpfvyQn1FXG0
SQQw/3ublzoGYo44AEIwhAJh1wa+L95qvQhd56Aaw3SMRsOloK+vHEuqkKpXOaSM
c9E2w7p3Ugpds8/BzXte1qanLvFXBrd/uvfXlWe34JQV33CSRsXnw6F7kuzPhuKL
GNf31wywN/uxQAsm1WaBIwIMGBtb8kHqA+c3hWzTw1OjkV6AZ5f3FOT2FxlB97DM
vX7goyBxb+kaI5ZkopC0l3azXFZ0htVMbn8EpYiv/3hcHcfDYuGLgdCVPqlh587S
zi6YUCQ5OAqciZjYUoFSQrUwif7rjIsHLuBKhANcJOU6Jp3Tfp8hgvFuvUoHveVP
/J11BuFCcACTEFtg/YbwPllcil4t6Q3JnlYYB1U1yr+ETb0jr7Okdq3yI6VJTa+Q
ijzxAUFSw7PE/cBAi1mOZCiWGRfDAOZiKJazzLxv0d/de+2R6c/A1t/qxS1XToaG
Pw2fwiFUzmK1B8heQTR4HMci2khiOskvYG1WS6SnqdCaY3fMwm9f9NOx8KBu/sJI
jwJgoBqaS2bKCMTepj/1vRk08SryA7HQPAPiiqpJ6/29wblaIQVBAkniknwL8X8K
Bni3l5JkQksgnwBxFlvtQ1uPNwmjmNqOR1pItG86uTZRVfnOZY8rmvpYRpYg0RXf
jL79Cmd7LqLed9qZQc5+4VNILe4H6LVXXNznfAwBIsm0mlH/6oshPcvVdH5YfPzi
CRhnk2fZpVhOcrOASCGUCZHbJe2VNJy+FU1QVmNcD5JTMFc9jNb1/KF2xhwN6q/l
uwVUv8J9qSUdACxyu+7S3Xv1uVsq/HiVs/6YO16ovjCFtJvLRKQVi2EF97m9+zVz
Vzpg0L4wz3zl5wNxmzBhcgj9DxlGEPCOSrMof/qq78KPrEGTXGwzmqW3knk/EaD4
AmZFdMru4joDPxVJBNOYdJHB6Ms6nQEtGuAPrOTerklH4QVhwzTKiLJGfOLyhxyz
TiNrkfDCJoVhqPjoooAFiY8R7XpABM/sMSMPPper/c/IkrU3r6Q0KPlg82Hnd8LJ
1jIb0ELDanVte2B8foKnrPtqO8i+IGxwjT3y9ai+cYQfJVpLWt4tQ0G9hUwFaF15
KLhpSx+gPCIPVcoKDh/XAi8l8rNzYrxWa4TK4tHEp2rYZuMT0eQP0d/dKcxeVhXG
dCC2bzQO4NcElYVtTdfEbq8KIL+eekv8P7s2jQjLBWflglEZA1bptyO3FnK+cqR/
KDmjXudzz5Us8Sccz695ed7fadz9jEe0S1Fgbkd+4D3G9xZbtj6w/vifNg92WJCA
arvmjQ2IR+hlLcGQoRY9XQGy9XvwljH0nYZ2NMaKPhnO9cCGekvqhOv/gp+QJid1
xPyaeatO2kqsUzlCoyOf1axOaWrkLIbhPlrsXvi6UBHpeMWX/X1OnX+ZZiTeA4Dv
yeOE4Sfu5W3loVZLz31awpcXZIbGofBP3wAOBg8K4DbCkfv9el08gTN7AIQPzEWq
qu1Bn/n8O0t+wk30NODESjbCBabZFs/ufl/hZ4cQg9f8z69Of/VmYOOhEIxjrwM9
W6IF8VsN8iIvWrwMCanxenIePnuC3L2IwjICM7uXWZUqmZaR7n7AzA4bvER92K3T
7165iB5a2Rmt22WPdL0+vcMgy37IDzhlaAHtFBtTIncF3KRujaYpwUR70NVXD7CJ
FPFZ9vodZX0YyeGUCz/MiYXkxacQz2Mb6gwvhg9DI+bhOSglY/ZGVA8xSeMGdZ4m
Pygkk2tpSLRjusMerY3YgYPZ6rlx07lRnl2tZChS4RjFJ/4dZGXiwMouDLcrcofw
gYh5xqUq0MiXlbFJ6fR+j69Ow5G2buBuM3tVsNu1zT/1KkcLspDIaiEA/5yqKMVY
FbYbPv6nqB7KgMTJ4jWHtO/4L6IxhOPBtcMkOoK8zURKTvdRfeHfpMZnBQR2kIFg
wwrre+Z8zc6dG+qjxsyWmu9bTiI5iyEW63CPcXS1KMQTrLFBxCFmqEhvTHMVTuAN
Eb02gP8f/j+6GaXBNyaqX0GtXLV7OORe4RM///+hfIaCTcJSVbNI5Y0assue+GXq
aHHMfK3qH4vcXzh2ZzyQhQzQSxXOnzNa0mYpWsVSPHjwUbTqs5vy/slZJvLRkXvv
POfU63GH5rAyDT5VlVUeOVdj1J7aN3/C/W76MT8miSfLAUwMZRta5PRfrIxWf6J6
Y/6uEqfv/QDIpagdAPFygveP2dmcqRNj+/pOAZeQ2iweM7+bwy/ibb/k7yyfrRxD
r8K+lNCp/CqvcX8tPOUibFAhFTeY1c87Os48+yooehsx+K4hY+jMIBZV/++3cXs4
mXZw9B4Wr+UZZDlNX9GSG6KWh6tCJdPNn2zUaeBa1AvNPz9UuJOrVJ+NWmSdeSkt
X7BUmGDEwVbqu6QL1gSn50mhKlR7eC+9kBLXFAPngXMupJv/VZ080/3ZrFl/DZ9S
pmHYpf+J7LOyhZj8AAVuhgiMMyy6UZF4PwzHcwURvGR8YBjUsk0kzKxiCOTK+l8g
VGqIkASbEOA3GhambUZJjifNoV1KCceUgw0lKfxTXuLhq8pDw8gQL/J2nVp8aTcT
Aseq4N0vALCSfBlgMV0qw1w9Toqo3rLrZTgZxEWGpVJxUKckUWJvsBYE4rtF6xmT
1KlAB1Vci5uZ+cg89ykLIMoLPN38X37svzgH8Q+Lb4ggY4XS+HO6MOohl25nwroZ
+PgrED+Rmdw3BBiLcKdQLQN1d+o61oJHaPvHpYSzYsdqEPVtYZSCI96wwNH//kph
jzLnnBOfkEXCA7HbbXf8iRwxjJRDLkUqszmnnTC1Kiq0pren7PqLSdzPN9Ph8Ruc
leIXmBKVJ3bnfU/hykDBAZJZa76ZU4tuGVd5/W82I6mjzrocopk3MVrfciVolYW8
o8/ip/Apk0vZEmZdpYbhbnp8D28WNoUxSOUVnmHwJlMX3YN3ij6C8KmtxmO0ZQgC
Ma/5Y3NL/b/KLeyrWqrJHSqGhfCf24eUX4L1zdA67TEk4Pqzk55xc7DUGv7AW9Xp
qT7/NUXgMJJXdy9uVRuSnEbyUZCBjRZQFNpb1CZtMVHrhb5hE8+FTg4y3YntdThj
0vlgAc4csMYubzP25QmVpMA95L+wlJyJK8JncvgTbZ7utSNxpXzu8ELUO7+UE9oD
U4FhwrnmJDWmQhuo26YGoocLx8XJGoV4efuxCvZ+WifcadCtpJDdc7c01x48uuVy
VDLLiEqkbDRBT/pxk4cbGl9mWmnFNXLntooSl7b4lf7qyIlZMrjTNf90gvEuHXL9
N8PvkqTXzEKlMhjLl3+xevKih+d6CEXWpYHJoo1W7NcwFRgxGbadWgWAQPGWeHuq
uAwjzK4JbN7K7x4X42b/eSianNlUdUh/+dxa1Wvj5LeHrdweh3xPFFZxjGgg9DGE
G2a2c8a4aKFFTEZJFMklV1gwWT9l9PDDOy921OYAQKv/JawqmkH4pcHSejGOa4dK
s5S+r8/3m8ynhJL7ytX4uVQWco7evCc5z1FiOuI31cAFj8z01h7BDpbmNg993CVB
Z3p9eqYOSfu0BM+v50wdrSrUeuVQbyd+VXhV96FpY0LWAoDvAb0XrG6jplO15HCl
cqop1EnEryMiV8hBB8iKolTiHdY/Sj81kazRBaqffLzJzTj3IwcGlI2t3oOxqOVG
191qaZL87rNJWcQw83IZ2epkthPcqOcPFNd55IIP2Ipm6TRcVJx3MYVgNHfxgOY1
Yqz+hLRAnLDYfAgInh04MGMp2TngXSBj+YeblXuzgrlkNix+Ixe+VfjEsv/5kFne
yyjSdMmkly4LUYn4L1uB4dOQrkEJfViQTD4yPMIZQs1vq1SRDVzS4i8xqoWEB2V7
Lj8oPsy5piGPVWi/8NAtOdv1o7MSjQFIX7b/lCPtDJ5fCHLsdb0uiHPN8/Dzt3++
evDcMVrW+I6cKG67KcoomMvRjysBDaFUQc63aG8EU67KV2JmZ6meNSdxhIgs5PWu
eImKCjtkhXHRGhRuXz6ERQIh9lJa7HkJqXrgvV8k1IndArrPepnUvguf1udDR89Z
lTUTc0lIv4P8mXkpcLDznh3K2tdS1HL2HW36bbfM5Vl24eJhXpAKanWMdFV08lob
x+boHKs5TtpVDM8Okju8VH6MyohCMFJVR/yuQrZ/iQttsDOt1YVGCCbQXmqKAvjX
22HVdPBIy4niTGaH0TmO/GLefj/pfwZa3ouDtAOBpTUUbDwOMREb9mt5ov/FlWt1
YZ7tJYfUT/T7vyywSW1AB/txsSZEMgLm1Sv/OgbQK2a5DWMgqySkZ7WDUPh7LfU7
hCyyWpL699h1DOhNwJ3kVH5YeVD1GVfeUgI4TqWkfsCYYxBlyu/WpRs50A0bLkl8
gQ4SqEnreywAo+CtUTzl16P//LQrYgQmn0J66RCQ3dct9pGZn0DS0oxFWW7KlKkT
kYsAY0UpH4Akl1Yapfvg0aC73V0dEfhaaE+fZ1VcxF0ZChfjLJNTAMc2d5LSQInu
xnj5EstF0iIuG1bgJsqqOGRzqJJB7gy/36mrKPwUuJi8jOjAPsfDhxE9r6ocxlDZ
DIsw7cYcwcLhLqJVhl6hI1n/WrPQQJQBWXwwpCBNSrtlqW5/cHjwEgGY1viOllkM
gxroktq3YCzfSeoWaF/Xu1M+c21rzEl5jY+Vz2vWmHD+vMuEa2wIVGYFg0pZuU09
P/XD4GAnQ7rN5KXc27jdYoD/Gj1uJdLlvNu7AlFyFVl1fD8Ky42L5CbPweF9V+1U
5+h9P91gGJ6Zpu5H9So3AGlDEtLU1f/eBJzoIxBPpuemLEut8kuAoGcNUUzeZ5ye
UyylVp12KwQ+DF0nWwP5eMCkpyO8O3J5+DJ/3dZw2WIefxxGrwhlAr6DQBrAHJ1K
KQwge2KfHHOV/qgVlhIkHlfeDuxgWKaKGQIXV4xSw8n4ubHxUhXbRyaFVRcccX+1
L4nrDOOrGbeYrn/VRjY9cnTld8SB2HfaOoyl/49CfPW5lUhRFbY7x3R4DVTE4OEn
OrdVm7/46a7756LZF6zlqeSWYXc2fXPlPrf88AJr0PJ2zBIzzRYv4fBkUjl2ySsG
ZH8cJmam3me58jOb18YNX+IKUN3ad+xZd+V752qeObZaSdpfhOotfQ4A8PKYTNfe
1j3WIo57k7sUKkiPRZXMiOL2hHe1A1Tvd2Jd3srD20vgJIAkHzOTXr6bdJzdTFMj
SNuNWsmngqHzeW02LYZ/hK5CjhmGL2D++JEdbKzKa4qbqXL9aqFmOpFIFrMUszFP
tVjw0l+7jWEkTEH173ds+OOl7XwDocriu3OyXPs/EVqh1wY11NrWEhrQXtOlr9FC
ER+I1cJ9cussRyPriiY32ULo8aOCaQIVwvboWGLUx/74aHX0tPyGwVDGyAiMbu/b
oJzQ60K2Eijh0jJNxNltGpQN12h9XrFVRp4l3e//7/1AlNiOr3pCCAosbacGVkaT
v+b9xdRA+YvntFgXcIkKJs1hc2Q8zHGo1MLE228iU39omkPXkrV3xeyiNqejGYe2
Wt/YCz0QwDWgLUNAJM0RqmGJb14o2jEkF+52CeConjkGd58GqU9Zdz0mJL7KBicA
9uSwE20rGUTAViGmiiduxcn++ObpWyTnp88AAofI0BQ0vUmEYVqXdWDNgIezJxmB
qmwysI8JjynnmjAcQjoFmMkUX7eNpTK6fVMutR8tjlmfeAX5/r56xGQsKx+OBCOX
celwadVuIhuOBPKeqegkTaI6LQ7Fnl7VjsF827T7FUc=
`pragma protect end_protected
