// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GkMyv744MwGvSpSXxiJd7mPLRYiaa+i0/RrXeL7sXlgL0jfbateL4fzwTGYN1/7U
+5fAHLRiorHH7DlkdfcsLZLYAQz0MaYsBNkb7vKx0DgEZgxJFbISBxWfcA39AwQt
69K+/7K1TVCqXHh/MoaAZpnPooBGhBci6Pjwe/+waoY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16400)
hZ39qigvKTuwJP2REHQ/g+rk+dkGa/el+UnLYgqfO/JC52BAZdo3bzVvuR4ldLjB
aQnttKEFwsihB+3oyT4TkRVMj+v2MMLi82XIOqzPzFs0/Q9WKZ6fFfshWi+4JkFx
847SYp4vOjw/CwsUijweKM3ONSP5nMWEcqtae2LJhoZPj/cG1sndUew0FT3NbCYM
hCKgnUrj4c+/UFn1g3jN8rntlb6U7LdABccG2jjlUAqlllT9cdUm5jHrQTP4FdKH
+dTCMyD9DbKVZq2WqACNbbI893a4buM4JzFdzv1Q/z+ienFuTKPsUu2o/LD2PWQs
BtFkeEctfNk4L/0InW17osl6tnGwQrK8tbApEatCb740uMgZCYznea3gs+xAYXTf
pRG8bvRszrvFaY9o4vtmokL+OUtgPUizcaGeqooY91aZIan9981zkWi+b3wO9gAS
haML9IpMjmDsqmr9BEvEvGUChxORe0LLTh9pPkBEHFCriq1ZThmUnRZtjLwKYPBh
4msIYNIjpH67l/L0fr059rjbBhZ5Vs4dn4u6H1xc1vS9WboYZAU7DjRRHGQEsxie
+UNp0RAB1u0lGRC1lvSbFa+FFNgcLJGKqAu17RFxWrfwAcCIOMzQGKkf0biarytg
g2QjOpVk3xqu1g3N5TRzGxFqgb8uJ9tQko+qQje4O57oPb2CoxkMKq69pjuni+AP
AgCXk/bMQJTl4OxjiGVfuPB2G8FDEONWmCdAJxtxIUSoED3deOWCPsL992r//Ox3
JqjZHzcwJqDNikHbZdGxqKyCYihQgxpp0AR2McWXGnOZtZcVx9jXxME+zHoDSxS0
K1lbQEevghOjGvLuklN78AglyPoi9pFooYJtbZLqO13JI/52hRH1nwST+6TR/w7H
dAp4kS+o9BYWsdcPcbdfUQE8AHgmRkiVm5ziSQSQdjOkp1SEjcY+Oii463HjUCMF
CA2/TYjOFh+rPd9k7iKEe7F55FXLkyfPRLuKz+5JNTL2uliMpXDOkYKNuM8S08pp
6TlNQdHz+q/s46skNdC5ano0jXkLF/UNDCyWQ4kDrHwlw9SBNxxwSobOY9G3RHM2
Ng1eJ8fPGHtIixOJICNmiC5N3ebE7v7MzZfs+5eVX9GrgfQ1INauWTj1Q84Is03F
4QRn8GXKYDI1Qt6THyJz7MX36eIuLVl4PgPW4j1SqFx8RNHuga9+SNfJXOWB8DtF
aEn4JdNR/W/V2GfKivSMu+SFXHLtan+UPME2ibeq8WyhrQ1ibgWZ0GZQVmCGAsnO
I0sy2ycA+0OGQqXwh1fGUllvVDCijUSST89xN841SbONbMqi5zfMf5Zz6fKvhWNq
VpwZ9ayc1UjsDT+j12/vPLtB/VXyHBoQCcU7IjZD5oc3v3bKk7FoODjnSNxR+Blk
Cat0cNfnVwSapK2qMtPv3PbGeIYlZQ/DGUwe0RhON6NXxi41Ht7cYzWHtrbDX/7g
SaGjDS2GJvEVAWzuzTZRi9N1PI/xmcXGoFM+rolnYvKf6m+d1lsiT0/+WJCGMFSk
oev6zUfy0UW7f0V6Ib4m3a12WNbddz6NI03jgdYbAI5OEqppJLCukXBpYW2SFayD
YE5npht1XjWSaPTniRHpAzALrMjkyiN0rP/YA0iYXXKIGizvxWbFpe5pSKjomPQU
FRbN13WssKVxzAMajur3/Vh8yzILUovzYeGr166D8tUZXNeHPEzsV99MmJxr5W/5
TzY9mM0W4gMzVaqoGnAvBDloyohQzGrkqrjG2PQpuMJm1irlOY/7sw/pEW/DkvgE
IPC7sXkCV+jEetVVTJXYwBy09socsfwT3Q15MJkAv+mxnjW/CSkecaFRINLPPVlN
LR77RmO/B/5hXCl7si2FFqQjA2Cpm8dhU+I85kvLr9fRVflzWBoXpj2bPDri+vHW
3M5CN8JEFP0RIwnFIyzqM8oUGGVvtdLDqCc0clu785/jM4hBj5VhozbBydZXJUfS
7Jbj7J/10iNTIHbHOeAeE51/PppWpUdN7VamNHsydBzAi2omEyE95kXqFM2soOmH
5yncoBBD9Ok6mLMg7u+9w4FP+6LbzieQteUY2er5/8d+MlY9r6EKg+hxNbqbYmQy
GeMRI0SOC9CYU95/8MZR5a+w0PhCoWwO47d7sqWiHIh+4fx2mUUfOnXF9EGMhabo
YtBAALDhEXrBVf5KuoVnzpP5QXckEKAOwTGZV4pJ3JvCrRfgno58Kstx7Dk0Mjw3
pGt2h3a935OZc5YEsC0DF5q+vWt1NY8Jhz6qdl54crrzJLw1k4vNXC7IXQ8Ijggh
ViSJqJTF5eBK3Vb1Dq9jJ1KeNjB6PNcQaoVbCfFsGxo1pOQJtgdNdLLRgBnxhbFl
zgCOOhJ1R+MQ4ZwtqYMviFvGNzU3PL2ozkh0TCb/OoCWHq2YCGT5NGOp8xhEHqkN
92iKjDaMyIqFyx0Hf/14mUaL1pWZr0iFhqpxMCUvfNlcgtPhmi1BhNa/yN4mi2N3
rZbUxw6O6Q6ODYhP1j3v9QXskkXivqQJ4BsvyHl3H/5DOI6bcUVL3xWreulTAKSv
LCPBLpOid6CsTUw/70fzyL/YUxlarUqOQ2A9LsRp/vO5q2onSMTOT/MuMMDQxmXt
sCyVuMJHoUmp4RPlcbmRK2yq7eeR4k3b+omMT0Eb5szfokAsrP0v5Le7CJVZ+wWW
0OqlaetnA4nizLyOMbyxVQ0Qf3zCxboL3HZEbqavGO2VJbqW++wwpNdcIOZiC8pt
juh6yqS7cfhRY0b8kswtxtMX9v2ONDNGh2Nm7HU21laiaO39Bo0kpVlzga2DJGoP
my7V5iOD8M7+xfPhl5BwsoIY6AadCeYiBubCpprbEZluDhDKT3DouuGpMD1TGms/
dqnZL3JtXEiuQE8+itFtQgbsg7WVeITCMkTp+hLCKKjlN4BNwXlY1ACFBdaF+mJu
GI/zLq6MG9IPOpj2LoOst5J2/lptEwt8sHELAe5QqzCmCLuZQEcjVEJH2bbh2m6r
iSiGLo3Us+i+zXz5B2zmwpW90DqZiaY5Zxde0YCMwn2NnjCFPEPoJCJl2t2KNGvB
bHuzLD6cPbt3Y6HxVbBqYXnEumgkN8+b6jeBhFBsywtPeWRWjJltBWPD+xkQLUc0
wc/qulnOXNC+LE7rBZW6+m8kqgZOiDCGCU7BxPUYaJ+OHEC4SYz3SZQZVaDPrAa4
eSihUpKgKGnOUlOm6ii4psrUsVJMCUUm9cRRi3AMmtqm8T+tVihMGsdzgzx/RJfk
oPT3tv3IFvWLgfvPnTnBYrPSKiEF3c1bFF0tJEv6Wr+PyWXQKL5WUr2790b6RKDd
5Gg8BS6pBE7YCXjmcJ84G4lkqtsBbcRrphFZgjpDD8cwbWcMDnpYC0v2T+ZCZWxN
07s+pufh04AD44xfp6LluOW9x5iu0hEtL6FnDfrYUQRN6W8yZ8DWA6wl5zqBumSM
djilU4vfsCVuNYmv4aBdzkau6l550yFk7q2YJWQrFGpkIMHU3+ivnb3kywhKFD/J
rnVxhHg6SKtLWRIzV+g4bkenb1kviOvyuWONx8Ag9HkGk357R46/RfvYUT7P3wxR
woRjWka0dHFqKK6/g3ZuTEeFWoQMiXdipV+5eMHTVhTNr/bbaZh7tD9HpfFBSGLo
qTj5Zh771tg/OqVI/px2ArxK1FgizN7o3U7ET+7CwIeCUa7ckQGBTpsYQJLXGe/W
fGXbYXMZXFcJafGQ254vfGCyxrYRUqz+xsgM/LDnGrMV6ciqe+Sb9B+1797QMYP9
w4xNdzIpI+90JpT/rkJN1DKv/EJSH6uyCjcLfCIsP+OzsOJh/UVuuYw/F7TQfhBe
6fQHklakN2OasxGoa7c0IewoHUIeZEJmag918Zar1VklcK6VBarI/PpcJhM3G9ui
AgWhlNjFmEaV7/fVTdaVjzYQjacq2Ks/hkaGfhbU9Ww3siFQGZssKpR9QVzV07Cx
AeHwO80yKyyNtKHD1DeiEhn5/KNmayquvqyx9IxzFNHijZXAegvIOlEXGWGXgpKb
+uPH6qDu6TLE/+h1Vjs4Xr1QMNg3ooITQd/D/4VLGwFSqOSuGqF69184vyD0fIyj
JixFzcXJOaDEmW04OCYe+eMjgr6QU4l7p/wHPIyZNrQ0xWcJV0jmsT0p8Nop4qBg
EVDCaN+SjBi5hJuCdnjAkKwH8Qe6unhqSTJqbHh9FXDI4EA7xDRbTIZ3Ce1fJ5jO
B+NONlQuX1TiQ9pKIdCVxVkLjM1mjZpbbGNyXOf5ITEgi35lW4rziByIwRmFppS8
i/A6oi90u3BDHVATvOwDVOGtoElzezncGn1b2N1ePlaBz9lYsE2RJg0ect8IqCl/
JYTop/u1u38XLG1lb4/uoJhBPSoDNYKcfgVF9VC/UtKWBiz5PYRDUaTsoBWbm1qN
FkDzYd405UUH6XMxTxd5IizkO6iXjlkJvg81ezf42JdkCPUcocTiDGTpoPOYzVRE
yo2wZAW/7XkDWDVrnciIJsUqCBqIH/Em4dnMxIVVqL/4Yq2URuGHdtEVQvmrrhVs
zIgA/IzH/8i5pJKzzDr/VEhR8avA5NDpLp1D7bqtZSMITvPwJPaaIuQ1lgjEjy5t
HycpwpJcZEf7OwGoyTtGotY3NShdJ/GRRRfrwX5lpjP6hhQbE30C0UzEAbRkCpDG
mUJWhb/cP+TDiU7N+1fWjnT2yedzIXmUK2ngFHMFvQFUq/3ajM9k85SFPq6g/Zny
i1R7qoGfKUfXYr7+tqxgTOFuiZgFXavdwfAMvwzSht1lk90xs7cr5sD8pwYFBYG6
7v8UQtvK6WX41yMBd5637y8+mZHta/Lg2MDcA6yxdsCXGQJKEi1PSV4mBvBsQKyC
j+bvrYDoxP8LkBZoYTkNhCYLrYckenMIppxCiCRcyKsn7QQk8wl4XxH9ajFIjQns
WVNBYn2QVBUp7xdP72rdneq1BKhF2hG5Qdbl5uRuKtbP7ReYOWVj2PcTp2K2BZZm
k78LGOyXIh6VkNJ5e/jluMeznljmdViKfikWV+0I4kVs8eIK+WlD6xP0IxanjQKJ
CYjFzBz0460TRxszb0k3DfhhcwkEHAmgYYQ1g45zKOIwrHbPNSyHToSAuqk/oIOs
AeGygbN7mWrmmAuz2Frjw/UIpaoUZRuz+Vh0I7W+BqY69PXRitSxVTmZ9VeogXQV
pz0xh8pQx7k043y2GLm73FesxRL3z8PBaoIwtT0i41fC0aMq5zbHbOuEyVvp90KP
YNT+O1M8vE2vfCtU7olzxI5h01rf/V8x7fgtMWMwzOB3DAnHFeVU9mbGosx+ekif
cJWni/BD3/IPKxU+R4ZJfflDALdznQ3rk7T5rfwwpgnJC0q/WAcwClGDr3yHvU8A
ix+/XGM+VaoxUS43RYc4YQD+UYnKPOreB7z2OEzHCV53Rc/FVIQ2TVA2c5Rgn2eh
73Ay8BXNxjYXOqfPa5uWOwkRx1t620yvTeaRMFWy8JlFAnZtnj5/uSizONSfN2xG
/DjiXi/q4Oa05Wzn4VKeux8ijPMSnpNs3s/biBuIBCS1FA4gWNx7nnPqU9p+G81Z
GtGT7Vuv6P5aVn7MxRPNiJrSJ/4noGqOImoVYPeCh4Hweu9hFKY82resKt9vn9wR
JS0sIhqfPm1Byl/VPNPqoCRMlq8WmJdrea0Rrg+IGgqOlEKf0PT4+63LelbBO+gR
wNj5peCBCPBmXYmwJvIoc4Zbzk9a0BtbESnC2aRtb8cC5Asb+wdvGnHRDVTFoS2Q
q1u+St3b6F+GofEfNTPc6pjTqBsq307dqzkVIDXEXYqsKjf9Xe42DK/evrmN2TTz
fkZyTzFVrk4YrVvz3/BMjqv/0DEAJyjCUI5yKQZ5BwFU7igk7yUm59tthAFA3dlU
MruIx+IY1olzXuNmcGU/57VB3ZdE7LE4nwXfCzreRwhFXaYSYcdxn3PSM3aPWCx/
VW8cMr1lvXZSaC8SGM0AEsEutO8PbR0INxEslle4vRzJTGjcSOnbQyoaHyRz5G3T
B/WKKODYIEGr74mNmKuSNWy8cLZ9lTCOdOoy5jYCnSYWGfBIn+4mgtkpsYbYWS9N
x3ALxmDthPdqz6n613g6yT7CHx4Hotmn5NIoahVNbHlqXufV/iwcA3GIaFs0m57F
ur7DT1RgmfOrvliSYenBCrYU6KMCewRi/txUjoBrnVLlw6ovU6c8BU1oK8QDv+KK
gO9UhoFiUpqy50QaG+/sqpUq9XBQSIc4chaqO/9iZUVV9hrqKzhfLY4BH1/+dlh0
PNha50gSpErDYzMwC8SucIsTKquK8FPh3G40YVzXXepEtHgCFaxOd8cf546kUn3i
/E9tf/BkmH7z5lK10nHJhrOFYyhWcGtsORRS+vnR/oQqjPNMEsx/V8mUOeduhl6L
e0VTWPKKnmo8bq/3WXD+CR9rhCqvBgXfM+5IrzZe4tSNCmF06VTOUWs8s2PYtHx7
TCRj97I0qtGCWxaVgRX6/q0QXpZYbOwVL1dFrHj9yKd1+JzFjaqopMUBmpMOSUYM
Xujm3ZenQGmDyVPVczrh0wHlA3q5SrFa5nHMwBFfLlRVN6WO2uhU6gX5XFKvY6f1
KfLdeMwnE1N91uJaUN0Aji0XmyO7qVBXUt8Z1zMAhhKr8Yujrln90MEDorM46p8f
BmM/sqo3j2wHa5jW2dqWFi33mw/HObTxu0WbZLmE4rmFJfWr2QKerZp0T4mZE/ev
vjiccdjktJp4xAelXKgoK1Y7H0mYysrNyG3gWqxoH2yHjrwKqmtIFK+insbPXJOX
+5tdlyK/F0Ld42Ob5Se0l0UZg/aPn3uaOdWSxCuOgoYhzN2cLk3jJsuWLnl1kXTs
dbiyFH1k6ME5jwkkuIaamgy8G9pkoThqS6bEePxVbYRZbyfp3JMnrfdeGIMz1Tzr
hKx1s5Tq42Nh40qB0UqvWTSK9qkO01ASHHel4nq3VFTVaoEag+CrvCe6+pTadqQg
66GU4GaGLPDWxzZ+bhzgzyWCYr/d7GidTaAko24ubn8CAhp8UaN+LIxh4admSrgA
q4YJUDSMdY1EncZldltuPzI7JeD+4QcMsRITMpB1qoH9fXNab06nbnsaqYJFq7Vn
A0SfUnV1CBvPty259RvKwe5tBlG0LVxSpY4x6sTl3xcXBtSVk8YwpnVzB8omyg2z
WfBozTnXYdOGr3Y4ldjoN2zYj7Ihauey4cSfkSlNvwxRB6AeY5taBT7g8Ug0tmPb
6OOfH40cxnU7HHUwt7y6Zn2x9fgunv0ECO8V5OjGzMzs+UAOmT5uhY1Kz94IZpBN
4xYUT/joL6g/hVEdnnONsmpncAQ0hhWmDEc/A8TmuOC7S61tLuSJ8iAfXWZHxPNT
SAx2grW8a7QajVBptuuXTJebw+jhHLpcaOYhFOumrVWrNYZBdnJtVg2d3k0BlAwX
FQKxejskShZbowKVGrz5dGCwrqJRDJ/3apqsY1j8NwJzvUp8L+W4pl90jcHVX7g/
mEufGkPAMKv6OEww6W9CmawwIK2KRHVGltBn6NyGHtwB1gkJuaMGEjyTWkQo4Ukq
vtSZ5T5cCtGHOvTeAFnzfRhpCDEAcatIx29c49A5tD3MAvbhf8oriOB9cH2xxj0M
JRf+q71d1l8Zw1sinrr7pPEFDi+hPJNL304bBBFK8nTZti9RuF+BQ16qml3ppJaQ
AsE4xey/dLAl9vZ90eCoV6ERJVqIcZjHN5cT4R7hoCCFT0lvkE2lUSwk3W+VN356
8Co12/yDMZR8liR8gerKuKGyE7626fBQGN5ju3BulEscDu8Op3YIfLHTZhv3qlsQ
axOlCbl1letIQR9zLvRI4rU+UFR42LT2qfirtP2stSuXt90qdAfVz6mOVqtcSF7v
3OqIYMS1U7TNhMfPOAOxuuToNo4nT/OJf9ccWcrIwQ5WW9q/l59bNehTzzTuzrue
+2dGrlRSYbGthyKO0k97aptfYs8zAW8xhQnOK/SyzXIOAL5vaRRykVyNPk7zQMVO
qEili/rh1iMc5DbVfuFVQmahjZxmkCveZMxl0UlIFBSJHv1fJFZmwJ/AtndADM3u
t2r07F3i5ejKbBOfpxO9+osOBxRTh8tWo5CPEBZrItqsSJHQskvnVpA2VNO37kpb
JKVc/O6CpPIogenmTi9jttvc7HLnQeYMClXwOwrd1HboT0sOm93mOatkUSFSY/I5
42kDq6nYqcNPzp5+6u2l8JllsVb+x9KCPrbbJ5oJtw+KH5oPm7jhUBIr7BD3/1tO
stbrF0+GU5Xi5y6buWtAnjOKz9ahOpwXAPUT/lXchgBoixXo3JdnSFwYva+kMVpu
7/aBI/erzocbgV53FmfIZP+I8KP/LNlzGsZmUi9gygKTBizGQYaC2PHcILVpODQB
sAnZd6bazBGOYf4bbJ9lh47LlhNDM/8LDno7TmKw5n8x19KWfR35sE+MuXGLTdGg
3i+vrYbdBarjNyNWDmz5q9x/+Ei+ACENxvOLakLg6eLoSwrXCz9cyL/oe8C90W/s
w2ENp1DCTrrE5rtUgTtSpE3ekDCEs+Gbp/0Xhnobxa3Un5V7DX/BbbabYT/fZ0OR
Rk7VjpB/12wks6Sn2KPAMfrwcAht/W6vyaBNhoLOzlhhZUGBQg0WHwV1swKfh1b5
/y4ZwznJsuw5o2rn9cgPz7+73FTWY1FgxsjAKSO4pS1u0/uBNpAYghNatUow2PyW
pY0qrfxTw0+U8Goot5QOQKGPRJ6s+ccw6phDH+gX+ZT4ZFsUg3xq+9gdFmjSI3VK
cZoS6gJESG87hQkwshSUZw85GI9Ui4qtkQOVG1d2GS8F2QbDcg++5NMEq479++GT
fO/8LoXopewlKJRBUMWDwYSUJh0bgKk/hPk55U8cUBLSNoA3JScpVDn26a+1H8xa
AcpPJ66MdQhVbY+/8oS3hBjZCHwVQAOm/g8CtuS+k7kpNpoFqBMP03N3n3Ek9JJ+
e0GLzgGTnQSGHgSmmhneqGc+vbYSc8TS99VjXSD/UfLhNaxgwnLtX9V73Y5kuQCS
jEG4aC75AouMpme9rEN/FrX+tYZ3J2v92eA9mH3WAmjNfQ4vgvhpM6lA3wbJJlh1
ycFqSmRj8+fkbYR7VXFkEuEaIObDPFXe8IBhh7ii2qo15bX7ZjqFgGPMecNHYjkJ
oJdsYUyXdVq/reoyinFVuZAKQPnDH8len5zScBXv2pIJzj3SSCwhQ03vIWKm4NLH
80FuBqjwcYPpx3wKGwnaDYShLRPoXRQTF1OPrWV4ud27vKUbhhDg2tDYB+wv6mlE
UrhGAwUKADL9icESkwWs4LgZNBY0SMxMysd9jhu6WKerAsnMTm1XZFWPJizDUqZR
gknWauf4Bf3LHZr3iEt0wn2EDKO8BAR4ZH7KLZsf41PlGiYXiAyKS1v4o26pEjzq
iTbQF6fdKVRAyWwwH4HeCMOb1nnat+C65oBKmnWdmDTdgoUpyj7UmVmg+tDHAS4/
RKEb51D92pvBiUrjPiJkHao+7TM5nQOUKVn6XLvKLKar8W3U73+GsVamVufkhx40
PN+l83DF5jb3yljaESOfFPRkjRcse7Q4n1iStTUledFpCgtLoBD+cQ3ogsmuVX4H
+jd8ANKDfQndlqhdoDbwcU9bpo2YcgVrHRdSlHG8+mF6ryUIQD2/dMBtObEHFeOl
6JUFHtx/iRnvIkwKnIiei6fMzyFKwBvCk/LQz8b8B4Q9zIZTEonyjgGgFEpPwpBd
xD/KZXhxOVcAQK7/rOcPT3tNY1ZFuzqqJP/SSph1uLlcsWT9xtX6wClrsmNYkiqr
PcVNgXSnWWvL9fak+BL+dL8nRC4RlYGFxiGlzcm12qBc6WKI408Uk1uPwBvBALyV
fiHeY7+BL6jU+s1x4RS/Ultf/O/+ShSOMzF/zx2gDuFcChjBafwQgDLfin6BSDVY
ELM4Ljonx13rYXMFBDatbjktnaUdvtHC2J9F2N6uDwMltqTxIWIJiOSZdmTtKg4B
Wb3i8GPda28B/5fIDIuMtM8eGOVqpAIvbL+ZRFcSB53ulMpS3SSqNqu0Rd4+2/xU
sYIOyjzEgVmrclkuL6c7w6yblo3xW3yENUdbqTKo/Qqpl9LJuuxiiV1YSsvvvY9+
5zk93ryxAyio+7dU9ogZvydk0CcpqLbm16YQgDM23DUU10ZSj4rOTZKzefgdcpMn
kfEPeTSMlTAp4ryOBWQFUF4Kg8ZLwluT1Zco9bAA+VynSEsXUwK0km28rWI82B2D
yyL8qS6ym2noBWtqcX/9emoZadNpn68sNIcgLUuHetha8616MzDTsAy/FSyJtBVM
YoXMIrFl1itYNudK97KP2p+i3Y8f7bcUZTWuwcGwCns7+3zMmpl4iyFzr83gvdm0
UC3ebeYK5ltoKQXX4g9YbEE0wTSUCoRstgtdCiYi+1JY7oC8PNJg1u1St2bCmiW6
rHlTeZ0oUDiIegdJLte9QEDrlN+yQw3bxeoF8kDYHgB3N9oBdWey3tKNYfVeEBLx
bZOxrjE5MbZe27ztbXdQEGqu5tGOAuJ2KElqNMyZnhgYGSL+qGLDzpXbNvpuCVz8
I5w2ecc+VCglYOxDklnS9+iJZ67/V55gc3cNBXWd0KCvE9+DrIO91c1LGoOPzS/H
ILAqfhLf/eEI3QvQH4MAjyvnqX1QGb/2X2WhLZ/IeXfs1+lOBWZ2a3tkqZsZ/+mu
kQsVV5qLu1Ze+L05eB03j9CPpqFwEm4gUOJQ9rftg2lYXzavnFXyqGX3qCTXsxQE
wlhfwDE47nZ4DCx3y8Slf/EtuZg3fXFqKzVkY7F8mv8YEH3GeJBhHuC1aADAGA0e
/LtxELVDtt6BpfOVGjf4MMvRqGy5dV/Npf8IFGhwVwNkfLbX1ihn39GVcCa4iHAs
44/nSxi44QKbTm0UTrQ1pWwi0ScQA8h6yMSZnIpfMjjb2MhVKNmykRRfCyRQggRq
IJYg78yYa+dADnf5bhrcFGqFXy+s9+ukuKxDLP03IZNzvho1t12GtI52PX36ngtz
oI4QKq5WTX+NQUMfchZjpu3MO+SFcwW+ic0rWEHLg79Z9PrOQmpgsWaZEH6lBHEa
T4hUxMfrhWY3nwU7wVW2DMndw31xCA8YnNRriaEbcx5lpQ4LJ5yUcULPhvRwqp2l
C4lnW6f6Iu8bvewMp6q155QB1F7abogLzSMb1JQduCKEh8FTKnzaDnHb2L4go64W
9Hlk+fqSrTLNe9mAcNX7hTyUKYkBXEYaw4X92nDpl0uO78u3F7wgnA91j98ECa32
NYTxiyrSOwxge0w6qFfvMXsyZruTgPI9OwdUPUZbVH5hi2U3XN+wXgcl8LdY7YUP
iw/sWH+B0lMR822SkTHcMUjA1DR1wyOHcZq9WRlY9rOrerauvISzH9pnC1k3v1z4
gjoS+R3l0J2x4PPjnl0oPPWBuFmU9XtdbOJw0Mhd97sNt1oAg91dWGVlUwWHvDHq
u84yGfEbjyoeQG4sCilZF/JHzVOCxV1mpDBb150Ayzg7dgw5MzuKpyJlF7xFmBVb
mbfZtNV0lnQLYyseobbglbiFqp8e92jUDPTW9fiqgKFET9xHl1v7BqBpfEL9Y7R5
ZPMOdRpQq7vLHCpf629DEkt4IJAka1Z8s3TqJIVWRogr6HgZYnG9Ucf5PP4aIyjq
GBMf1h5BLWUd5WQAoP0HnYhpfJVQQ5ZqPui8frpcDS7wG6nXZsvDzQSWmxmTyoph
T0pNct3/QTUwc36wSdNO6OrtSBt64xped47CzYTsXKEB3TL9gTBKwxEfAu3wR4V8
nFMjmdH3DY+52mywdms0YXKFmZ2vyyB09gDEe9gcnCv81J6EhLOOj8tT3WaF7sOb
4ZTPahpuvzVpKcv+zgZAvYqYP/FoU8AsgiqqOiSiqHPVok8H9YbAnwGHIy1lwSQZ
LyZjfWmi72uWNP6JzNgiHpbwVruhbNqsDYNqA+uvYlHuA/irplM4+GOMjEMIJupN
XTLrYeydVk489u3cnOf3iMeTQpg5nDYXgcadjG7LzlB7tG5tBt9AlV8pIMEeCrqX
JybYXyFJE9L1JhT//2nHfaGeXf30CzIfM4ByXGbXzc5NFj0ffE3C9gMhlNraUfGC
MytfIuEy7HTxRt+zS9INl4imMh45ln5lKhOZBHg43RfqI+TJQP/oL7QNCixYxSqR
C0xjt5rNcB+BhuswHtH772TyEe3gQ55JMTW0AEMmV33vq+JJ15Aw5/GZgFypIlgd
ZpD/XYdJse0O+SGcUJUHw+Zb96AMDlYplOySgJUQMmjE06q28ZdpvP54IFPYa16z
loppOp3ffkZd2bTCmtWLQ7J9kxCsGtZhQil7tIoIc4d6gPyx1Aaf5sHkbAYM8iEK
5RFUW/lUqW+eDny2FzJhfW+4vZ1zmo/r0xWRpnls6DG2//+b/eqllsduHb1n/38Q
YCpFdaVNf2IbCOvQ4ZROH04FO80o+ddoa9b2y7W/wdKzBNWUTCLa8eiQPl8gdz16
rAjXbiXDy4qeB2XwwJ910ViwYV3eJ9Pdb7jiwKonPIKmiPooP/F7MVP4sIHjpy3Z
l4uefwyYdTZ+sR/ZosDQBx15U+diOdtBlccSSHAYksPZLVu/TguOLzl8HMtZELNL
32dbCF515445nhP7NAYcVaxbCWj5bX8Ta+KXrgRs9WaiRbsIM42h7dFA0TdhadIi
qphpYopbM2ro2OJrmFXbmKMZksP2HxwWhgL4jgRy1A64pgEFjktO4dnLMOvJh8n4
NVdN+l0J1cFTeYMCWJ6FKZCU8xrEETdicefqTfbPlgZwcyXCfLYEWmrJD+R3rLG3
uGPoUZ2YGJIXml0ZWsQ8a6o3IpGHbOuXCHJfOzjxvzQbCxx9coz9miv3wSLDk1yh
ySVwMcbhGRDlBMpzYXrkj5JbWJiqoiSM+/oucwCCZ0VhryQoMfe33xCT4a+AezkU
BPNMMcwUq9w/4+JUWQcG/poC0CDobnR/QcSmxBCP27rRv0AoM75BMtbEuRfFgkd3
jFsxYwKh1lW6R1HPGEEyboByhNcQU5W95rnLMe4EVixcKcjBT4q2lG8fYJbPSYki
FGyaJZvoMR2uaIOGa5SXG9fBxB4/cyDHKyehyza/S9oKC6DQepGUC6gqYjivKoL4
bTsgOkGJYK3A8i1J4l8FDUrxyEQ+y8ay8iTebenfsPHo/y4YEnO/QCC0ozab0ykZ
XDoj4kwT6t7rwFmiZ9gE3h5WpRt3A5/DfTaAONsf5MzpUQahdCQbne2rY+v9M7Hs
Qm5WBeJK55eZGIpy9YJES07eMEEhiaNoisDvABVRMEN8x3+6+TsTJIIe6VAVrqMO
UOX31KE8OMCsU19Sz0nP8BvizI29tkgNLJSm++ychwkqpXNPbkgeaXtaxAmYQAhY
thhNjfxGvMB2MzmRIdvk8WY2GG6eUaJ0eXznjDrdQ9FMXh43D1z9IEsUkeUhZwQg
2ZTa0++tJ5a8zGJaEMqx919tCn1i2gZg4lKlvIBHDhkI+Odq4UeDrwMP/4JEpJ1n
rFjT4cGur61XhEyfgTuo9ocUBlFusHAEy8l49zTdl3t1UfuX9I/AyAZz2MeybuT8
N5aETi8I+R6TEGX4qlvxkVnm08mwexNRu0359byOHQ75HVfuJGMBceD45OlFKvqO
HCXfmvHVvJ5CsMurZ1VAwcIhXnVxx5NrfulhSaIPl/KPaGRUDZdjnxDIAA8YOtoJ
AKuNcNPkqkEm+oe1rUHRvrs8y03LchQowG/rdHGZ6oOCo4UhzVswxvq7onNB2oeL
xShda1MnjrLU802b80AQkHE4vG6112DnVh22BasZz8QgzmqSzt3EIg9YJZsU9zLp
vqc+CX7RDk5o5bsn1b5qJjUiQI4GSUB4eOiLoWHPo6NT47Lc3hsFsCfRMh47f2Gh
UlnYdrkoZgUy45ZnFi9Oex6+hGc2QE9N1r7JJKJVxdDB7GdzWqNIcjoGTMHtRrgQ
0yMzhoO/ZixaqGNf2px3XlZ8A9EyfcSjif6Pb/g0jk8JgiVRlmEMVIX9So6zuW8K
ZjMCCT8JjjEpetLJ7muSLZQEPY3IWO3ViaVxEwH11jKLu8ixST5m++f6tNvxkVFX
r4UsbXsB9DIcOCgM2fQI8y9OSHVphME2igh08coZFkXsqxi9Q49/yPLlOi6VjJ0Q
BvubhcvXzK8A2DMR4bocCAFGOr3nQdr47vS6BZud/aaoPoH5GgV0MiyeMUJWJSzt
FF3FXZDsSGltQ3N7Kh2BuM/R0/0zIq9O4wO1SfUIxyGDgQAtC+gmhvTjRa3+w3kK
8dLk5rKeSu4480ywKTl5J4SNdzGxvYKlVG05Opdu3+LDZ31wlryxQHYbg1EW7BeK
2rjCnjHE2Y6QY4LMWiyZWAoX0daqdxoHdUehNFo5vxJaRqea6eBoFUI9h+T7AV8F
/JtCb8QGHEAfGbo1STeHfv5o3CzGHn849w3JBX+kmWSyUfRI+DMCugapidcC8G6A
zG6StrgUEQ90BS2BxQ/UYYqSwo2XPwQtlhnzBPMy8BB3utRNHnmrXq+krSH0H1BL
0QWc7qEpk/ddnTfLdm31PWpvOIBLrhoBlCa9NJqS4RM4NiUTqAzwQHyb6K1YgyMr
VkWe40+U8f/xpqKz3H6jeO6ZUTUAM5HrH+k2lpxImJ9KbHbNF9kg9fsXB2rd4jjQ
TPC3XBcrkvgZWtQ/o2NfYUS3UYB4LKU6k5Y6jWXQF6wq+xYZAWkD9KJagQlUByC9
9nCOH7DHIqpbwi6P1hGsQXs/PTGvHcWOt2XNtD6wkDs5LCYqt8va1Jp+j5opae1s
qXYH+jWoSg4pe7OLM919yOTPZmj+eHS4fDk+JbzPMMSTmv+NKGa0t/ym3ZXdh2Be
W/IBbRZJace/uOF4erLtGxVgDPw83vwX+r0f1t5CsBm8O/WhRiyk0+fv/sa3A59Z
AtrWza8IqpPiyVt4/KL4bUljAgUTAe0PeTJzwkPXEbjLwrDZ6hILFW4MXIspCJ7R
yRQ1tOK7a0w3AeAFonVbLGbI2DnWvni2sZqfpsDY1NGb00J+hGCpYpXl5Jy3nVLw
+pua2UGBlVJX933RwuAqfQt0H44r9SQVLbyGFMfEmWl/vrD2D6IR91+LdFGJcXny
VBzl+gT+/BEhbQ6+R0AurAtlCTxZ9aGktIQGblGAgFX+pxgnQm6peChspFidmeyu
j9T8sDcPmlk3P1PcptZ8iBEEuNAbIi+VYAw7IFDHKbAOUyFi3emAeUiI6O5v+zgl
aZ4u2GhUsDNrIAFzwBQQjWJUwcwfaSEY24ZPw0AiNQLM7nxyDk5CLarF0LjzPbep
DjBvx8nzyi3806wjm21LyZPGYoiBaHX9+55VV0lrROzVRAYTPvJR9UeAVupCBBs3
YO2ZldEP5jKGO+Y5Hk5eAtyjN1odj6R0Y1ubPqd1oLs0zEb/NUrRJa2re65dS9Fz
9HD9bvMzMqimRy31mUJxzzyGlKoXdQcv0QWiIZdN9ES3tw3Esr9RvTgsiZJ+zajL
TyxCWyI5cfBP2HCGTR9DZhl9lsYwb/d6uhpnIubniJ2/2BFLEQVAGfUaheES1LjK
txOMlj3Upimhk/Y4BWTZLoZqrGqkrNyfKGuX4p09OnOK+7+iAmBiZm1Ix0PYeSAI
sJcovGdN3XetP5GPjxasKkXJ4UJyB6rQM9c0xNvOjqju8hmT7wFr4DSNTwZX2pzi
s1eDnHhjK7TFhq3LHMcwRU13LxMBuXnaz03c5feKE4mv5xoeCJ2D1A6ok5NXyGu8
DaFuz+aAm9YQdP0kvn9WFDsHug6lR8Xu4Z+j8TD5mb3vzjscf/Wk2rioiNdBA8ba
BwyZ0sKZVOwQ8nPiG7J8zoBiIh8aoqE7+vSMRayL+6zf0+hnUN8NPQ8uH+B5YHya
tpcwMqrkIFUn7/TCdpQNfDB9iHLX226uXJC19mE2HQYOvjjgF5admNxBYFEJ/jiW
EZOwaAT2BjxpggZSyBRrpEgaCyZbgzAZDfr/Ycyn/EhB21+nUvOuYFzrrqR0CxPD
U3hJ1WlVScyiC4k/Xwm5+V9huOFXg/MrepN/oFJgI1CfLzQ70Ri+4s6XMen7+4ef
S3CEasPMxKz/YrKQ6etpX+XQ580Q5vp1D0+wPPCkOQOquiDoV3I5kW1juLGkV15K
qyIoSIMZ8FanM0qkWSSoYdLyx/gBStutJRLwiIMLSSlPG7dH26iJJhTrejA5FFr1
Kjvh748tmCW7yopJfni2LybIaHXuB83BA7uK2FMFnhrF31r1P4+WH6CKw5l11yQ+
zCz2re9uViY6r7BcFbiW+kSwVh2sn7qCuTV/u8qr3PEdE6Pmsq6oPME5w7C9MBL/
cAOobql5GuS8nH4WpTEqjUlQvQ3DAM78tYpiiv/ihmRkor0gvhrMwz7ImFIfTBD8
ig2t+zOHAjB43FOD/Uh70+jhfJY1JY4YnbLpMzUBwNx6liPPJDVh2u+6tWVQAGxO
BT+AF3uRcz7mk7vyVnczShSyn4dICmzeHc0L05efDBaDoXxgu6MuHi0wIn9bAN3U
aX2u9qpfeys6tno8YEfqw6lLJvhsy3mVGM4hzuslxqA0bEUO8IQf3odcZZqQPUmX
DSD684Nhs52buuWCPCUpSawi4BsGYTdMmRnvUsNl3Hl/p4+JQBUT6ChNulKNvG11
6kWgUGLy5bxKsZY4ODUsdFitOchlcPKxHUHj7hdzcIRuW4NdDNXTSdIzVm14e0lA
hx2rh/j8HYrUxgUfsYHK8fUngqHqN57iKlM8eeumLtsc2OQDzBwEkIWbNwpuV7ai
ttKmSCJSctmkG146GVdGT+fvju9HCSUNpfx7Mkh1opM92HYultSJLdjAj42dUOoN
xOayDoxPb1PXKaZ+Jm6GJgYGHx1THlDkInudP3i2FFbzgJ7QyRJH3nI/afi9/qgA
puiSwFcxsURkYZc3jl/8yRM3OfMxuSy70Bs1hqoAxjhPHvjI0g1RYwRYZQsPn3iy
DhUkf/GTAENnWyaCxR8i8ULAI1YB6u7+hXp+x1xuaQzmx5SdsI2SSdBdC/HaEjiX
GE841mHx94WwUciqLPTGIByxovRTZcZ5+TPX/LMFARUDzCSBMui9YeWL/V3ogeqg
47ceBZE8JGbxzDiDclj7bfe+cs8ll8qNeppnWEemnRu3ILVFRQ5T0Fnf35v5RDU/
eEbP/htlYmQxZovAIr7BGOmKg8LUrNf+iFOu8NIM7y04pWI169VO7AFUORAZxgos
bGX91l8X26ueMiRGMlVx4ErIaWzxabrXgJ+9dzTLRpbfKLcXdFjy6M7LGJVGo0N+
NrRv6mFrK4amUY8/In9V49Tdj1ea5PMmt3zJbc3+TkuJXF7QIzhGfiGd9fuQePOe
14haNoigRGzEBnB9NMGwcEDqFMRXqN/y6W3AZpGBy/jUe5Lo7OyEqns4gqejQVf8
wRUhC/ABnDbxs8XsgqNQBaubMDXJDDjmIGMOuKSRVa1YmdsgdIQbYK0h+Y64nQY4
FoNLhc7jziUPknGPPZpUq7YOXDvQcNpULZNBg6hykK5nxJrRSi/90fu9jYy4TOeC
diSouIxZzXIn1Apt59L0qkTPCJWmwonYSOb974hHdVJQpSKURNdDUkbwIvd1gP2/
HBBAper1zNIucSsqiEgA8Zs6qar7W/A+dp9MPLDXkdpzRfC+FlUNLk+znFfWO2Pq
Ghmk1Mjg4g29Ek+NmFXxc4T0IIWLktgTA+wykVmTNfzv/DmWn0SHFWU/9ztTKCQl
MWssuujM0kG4QhFFJFyMYtT5bjcIdC0EBrvqhUQXLyyt7LZf2keVZ/rgMcwJdVYW
2H2lm/mREh1O0yjmiDnPcDy0nPSR3xED6Wp9+G9pfONA5UIxgCRGEY4cA+6HODIB
CLRLrTW1xpGpfVyV0Iuc4WWmehNQ0+EMz5d5+l/8Zc6GNI2DHT6qrGaY19cjUxqP
tZ+urRmGC8k9R1cgo07KgD+KnRP252fZVx86z6/kZ7NkqOwr0MUNut/EusPHVM8i
naUuxwb/wRl92Sv6mAVQ9FDMfy0ZJgG53VbIT+NCLOkf0mGb2vpqdXIytAK2RAZC
LkE7M76b58KoL7vAR6D86o2OQw/9x71xANn+IymLXxXXQgtrIpF3w4oIXLDFKqsp
Jlwvd4edE+JZzng91OLdYW0So08tEwSN+Al1GaQl2I2jWISqnumVmgBLVsUF1qZX
b1jQ0QAhQ3+2g2pWrkFXyJnbILj50VNXWSEdgkZPljqlZn5aEAplEo0ue8T0g+p4
Z8EHnkWolNO6ma2ckM+NkFsCZBhzNNGrJaL6cgh/2vhhDptgSUeUga0TO1F6aNYF
FVkHO/Sne6yN7khv0y8hj9ImtOgqdmVeyJjSKpkS6da6LQR9KBHPHJ/DuAwUBpJ1
cmo3LY9DoHt5kwW5ClBC8cCQ37fEP/7J+5SEOq/k34JbV6XNHBeYuekOPwOAy7QC
kU29qVAgf80MbekUztrIxnto9qur3TFmWKXn3SA9ShSC/D8niyZAOfjgqfguUJU1
Mu7+gh/YdQb5w/nUioDQ12pwdNuMSX0OCS7GHP4QU3+pNENGO2ADTMrQ9nDfNToE
Av27JXwqCJN9n0CfBJmymptIKQL1zfKi+4yntyTKH95nKVJp1IGAPV5tbsDFnq/G
Zk1E8/AI6Qxmk/5oqYIDCLBx38PHKgEl/el+T4AdKMQI9ZEj94nFqsx9WoeUTDKR
obaiZTFxtYTOVuPwjqR/zA9xeVu3hE8542K2F7NpZL9J7BRnrBmkDQqgw13+3hD8
sCTw7B2iXtbrXvXxtj5WDOnMspnpg6i1BlO8wRa+A283SFt4t39NvjqXAGWBeQD1
8IM+6jYvt+6xWlu9CSXdNC4sx0aYsuaJ0kNBrT/79/Rtnm5RXCdYK3Dus29hTbDa
oIEtKXvzXb/PXTfGP66CEgZlE6SKdl0fpxf5lT9GlyR4MSRhuF8XBnCzCysHe0NB
bS5GXH4SJy/bqK2k3evi1Zx+9ZQ4yZB+S2g6avbkRHsumtmm+Q7S0q94Xp8VF6jV
l75/jiOzYwmXKwCq8/gsHFV3CIaPqZfGV3RICLFGfCJUt6M++xqCoZ5J5cQTbCBG
2MHkEuZkWgyKFK80smm4uBpAoAtdHtwE0IKa/MmbqtXl3yfY38fBU0XkB5uSLBPJ
UiGWOcYdP3wNY/3ZQHO6kwCLSCch6QCIRy94UV+JAQlQeqPK/nwFjm1TZXv1Bfjt
dWtg/Bsi8iDXu3xAF9/l2KMfU8GgUrdJvuFpgbsFgFGhBTfQU4bxEyHetRKFwY5t
dlCAqZ992Fq06z7HxX26LCLkjX91aDr6TwRp9WA+unMrMgRXhwQ7/16ldGk4qEV8
u8dmOKdfvmjtodNDdbD8Mv9TLHsW8A3AGVkNhc92foRL3lHceG99uPoFoaF6S1J0
RNDlCTuXL8dwUoQbU8HpuwtMVL61IpOJ3Tax31ZPPWR2GgQa1MHPimFSk4z6ZgWJ
NlRTz1xUYRt3nZe+GOSAcfD1X+WpeWxkLr0sHJLxRem/2iKY6Q3LBWm/rsfe/56P
DrZZX/VdQe9kOm9HusWWkQcZEvabpwAP26nJ24vmxrlW6nyLRC6Eso6P51x5edcB
J/eJin0e7uvo06QhXFUjAchzGR+385qnSFY8I3NDR/add8Eve0sTvY0jDIK8VICA
Yd4TO6+7keprWI7s8fbsmNJ/uNPUVklmXXaoHiXK9OeowkCOT+VVSU7ZgcwEI1eW
l0iau5LuHQx/AAg/TIpiNBF7zTob8UBLSnpPye1rGayvbyiCG0jJVkVTwKNos9uJ
gb5W1TSVRKkziub7rN8Vw8Ys6/gbUR4tTFyjrYGnsa6d/x0te/yqRAXzdhXhXwir
cirvRaovdwpiDYKjM4UJmYxJ3vaQuSn0AfoaYa427zHW7aHTvT8L+LIVLMdq6Vsc
KIR6igkNOCXETUHQ9SytmbfXifk8D/LeKwlwHg1e1QSReLvg+1A8r6losm/o0oFW
w/TBpgL9BV+wWfWycsvMbQ9Uk9nS0Los8Zo2AobvAcPHdd5hTgoXt+1FeuIWD/1r
/CxHCorN6IhktQOx41P2szlMsThgMlOgfItlpfWHROf7FHaIslngYNcU3MJSm7Wl
Tcwo0Tk0ZNZO6vusVNey2u64ktByqV+p47ejErtQNBep8d0MOy9I1/4t0RZU1hVv
CqRJj14gnQuVZndWLLHc2hjNWD+OOYbZVubQCGKVBzaAjLlOd0aoiY5VE3iMsFJc
xxvbQjYXsd/PaGq88FAqN/c2X4Z56DUYuH8MlI4GCun7DBlZIKwJx9XYV7Uasv/E
0o3bhgrig1KVTOyv4aBM6+jtFYf2WqVG75f3COMU+x3plmu14RVMqdNt+e2Y/7Tm
NIR0o6MmdXVaJUvTpSD8g76Uzg8kWtvq91iXZBkCQC0eMEPIvr86jYim3osl/Kor
XUD6Rh/ehGZZJ5jX5tx9XfGDpaaZ5wxuUERbNQ7o1GlXKSyOXUOnEWKTeZlNsq0X
VjqzsN2Eu1U0yi0MqIwneJD2CB9k5kQxy8NQF5mOwjF43GiRwBzsDp4ZFAW0GO9s
Jram5/E9XTck37pyhXTCR8FeGunco3MOakfoXXxh8xJqft0wjAhsK6OIDPPm0r3o
IFV1MF+rWgG9yul+o+Hj/CloZ2WW6ifZTXkMRhQM9snNGPyH9QROZaBcRVxsO3Fy
ayB8Te2zUMrr+LCwaaJSzZdB9jSyKc+BVB8ihE0b6JQHYmTiZx5X96qKNgBRFurG
nEkvkTI2MkFvzcdBGxfzubBcnPYNw1jHBnO0T7gD785ywSPjXgsp7yEW2n7LPzP8
KB5nq/GaVB0ALYRQySkzz9uwJ4eocZfbt1VjmwYxlf5+wStGjutdjmiRu1zCVNVU
CcPyMKLeMnTup0g9BCJAOrwM7atfNO+Xw+ZZD90Yvk6+CERqxk1VaeCmMMD7yPTF
J3iB9rLVyk7oUFWGwgr4Js/+smE5nROf50ViR9UEUYCHidiwu2STXMNuJZCeCzvr
w9KEd3bDJwVlXtfFhnIJHhYeESlpoilg2KPaA7rRHIe7EOsy8AN6vXx127AXccpj
wXusQNv7VcHD4nzMwyG6/5CE+QFamSeBVOut9ed6kN5SDz2CH54O0w5joSbVrLtM
TQhosr9UkDPMcINHezQlrrYiaWVa9Oa1ZuTA0gfGvG3ahqUrHn29h7vT5r9FrZpw
xE06sVsbMHCiUlfYywCIWyCJfZjLf/VXmF8D1+Y21z5KCCj5RxbXkLefH5cAgBgx
zPmlINDGY8ZZNPaBSVH8wzfmBufvEgWH0MRwBvMWSs0VuqAJNNhhPN5c4nga06JQ
bXC3zTRSCBFtpv6hDCpbnKM+lEIUPnnZv9dT2zfZi5pfnrCZRgQ/SQ78BAis4H34
U0r4l8Djl1+7rqsHWcqErLT4IFsB2VkAdePdRWSxI9mBxOcWdeRYhvGTThcRwR3K
SA2QjZs6XjNi75nk/3MXaeH3IslgLFNtwBiCsbGEGcXdKCx/K7UQUKv3F/dmOjRt
nUXbsOOlamNFv31iF/47kyBjdfHMDOe5dv7znPqGWeHt29/6xce87Ze1f+SUCLHI
M7YPbHyv4QH0fpr4fW8ooll9fkEOIcgPiUwe/55S19YJnEJ1GRdtfeicb2lOXDOL
rdIXCEvu8Q6D8bkQ0IMyGVBom8UQ+Gn9BbuW+koCVeE0yWA1fRWEdHrXBJjrS6Jr
kRIHBsHVrKGpzjHne1UUmb7bTUfdecxBO/agOHWS3hMYNwEWQ5yoCCI1lnNszdIU
/cfYta9uMrM6qqtp1NwwiLr/Wez0+gDAM89AnIwDaLmGTFW0LIbW3ctfmwPNvhOh
hK9xaAErjC60PW93m4W4caLQZiD+ByUzTNfd5yW9PTo=
`pragma protect end_protected
