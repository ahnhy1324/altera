// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ILiFbgN315llLjK1PVqxYfUgTGTKoNOERjkKFci/VQCN6+vwlU6a7XwN+yDI2yXn
SuVeB+BC36QNk9x0YQu7yakGYGhAQM3GToF8f+W2gtG+nNNujzSG755vaLUgUnFZ
5hMUEdnZ8frg5I05zEM6ZO+OOvmyKLkeLh1FTqkELg8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 62928)
vVvyOegolmAyPm64AucByLk4HKgrp/DxKXrUbtVyfBlRcokstc+aNLU/ijqO1o7H
iwVXxj4I7SqrzytWHOsk5NWhvExU6jmWU/9MlUmrCRoTjJqyOnzxqHtvJKaUdoGu
rZmfwQg1vqNI8x93BRMpJMRlhOsQx0Mhpr0LzhLHN1H7MpGPqWbwAtSjV9UbDUkf
Zxso64J3mPxIbPK+MdkR+oZ1oGcY1A5FZwM2bfNDkdzNFC6tGWOFiyzKbEjPKhBG
/dsXPpH7qjGhsFX8Zz2aCFtpKbYK3/iCFMyTqo9juaNfWgU6sCsKEVD924/OcG1B
1wU0aCtPlzQcfW4Kz4kHQmagX01INfunWajf+hpr7sM4HVZfti4tsImgxzHByYB1
uHqzpTb3WjRFEB6Sab3mppvYwbD8HuY6JYJ//6UTFAdtXBVeAzN8BcrOD9H1sYd+
IjBiQ8VDZmrqHFCWRkOGtrNRbZCXpEb22mGfJG3PsEfGuWLSRdZnjlqKH7PkFQIt
r0nhAumqaBODfKL3cPV1cfWg0cX7Jl+3DVDMBdSLL7a3g/RfJV7kfbn4pgQCZPQZ
TtC/QCXKI0HWw0+CLW8gp8TPQiTmsBRlluk0qTpN/aSMIRfWvxEvzAVq418s4i1v
BFAiF79PDoERdWf9Jw5VHepERYxtUvlTo92eMHeSie2+fq0VF9B/sRMph1CvDrhU
SV9HtEkj4C+AeI0Cbnbdji7KEz+s5gwZS+vHE8g31HZ9c+MxjEIIRaD1fNOOTmvF
RULccZqwAtnDPpDsp+4cfmluOAlvco65IPov1SKaqMeskipvZFp9zgDZkpc68+zk
jGXG0X6JhwWE13q9t2pe2owCkLyrd2FWF5/JPIMGwxtPDgBo7d0OOU6Jf0iQiOPr
ctditB7hZvKadNN8O+fNPg5DwECsXbCmfxQ8rh4fJaxetydyELexq5bYLIaGGf6g
kpZBXktO2466TSZZSN0drkE5xlKAHydPWZHh2Ktqc3WR+rYyuhiekzXh/nUtfs3O
8jXxCO73XwhfetD2Y6idBqzcdSAX6fNo9Sy7yIGaW4zYkxv/zBQGiLcKE0SvaKWo
kpYs41MyjK0ehf6p0BEWdRQOsMH83QLpChjh10VMpp+gJ9bfsvQ5y0M4cUn5egQz
MXC5NkhlY8ycYeemCoBSpG2uuuEiOor25exi+VGegL9Tr5qRKbWVO2qWX421t0FP
4EfcjTzkk74sSvz3RG+rcb1kvGmfwYBBABGN1Qtk+J0bbJANti6cXxO7jyfCg2jH
3I+GjpfmuZXpvJy7nij2GeE+wdNj2QjEKg3Yq7SFTLSXeDcOejHGq0WHx70VpHRS
DZ1ymMXFdOX3iJXsJ6rAoOU9E92TF5zpFYPaW4eCcbnqTvtTbhjfWcPhdvgGVB23
s/mYmXN3rnaFDwkR3Pmr5iTCoO/qgYiDfOqYEEtxbzIp1WfR+9gDXJ/nvVDMxGxa
gFexjC1Rf+tXghZCxlB+0Mlk3UziPCbS1W2ss/LUf0gH0cjsmkRwVOUkQZTNgFrs
ktXVxM38UkCz6hPmtQfpr4lTYNnPOZ9+EN4LbVaTGCZqChyhuPqwEeQHcFxeqsd4
GZsjetiJ2OLSB6rZmn2+rhVDLux3DGvFDFQkKppGuTlEjQ+WKq0Awrd2EYeRiD4J
e0VeErkE6YlCZzcLJgDvxvxp38DiOl8SqMb9M2fS4VvvMJ2Dc8ENMgZUq0CzBZlM
ZQkumSTXGylcYmLiALBmkcKlsQfu3KIu/hQul4PBYoUpQWIjRSy4uAHb5SBWIKyt
o3FNsu5DyN9CaREYdb0qpmiqNleH46CRNRtKJddu9L3atrH4bxCG1n6oYwugsnzv
2wYwgLF7qPhV8Woyh5oRUbQBLpP+NakybaAx7jnuffAWQLZcTOlT253QRfdjZdzB
h7JizkE+iN3fQ+ztKNLsIA15CP8CdqlRmj2h55PZdgjAtG/FefWGIBAbB5mC312T
e+2jwH8+dVGRGoKs28cw2ThAVwJiJ4q88D4cTuY7h5LQEH+M6D5AdQ2A+YZR0uUY
rD/dR2Wzjc9NPRwrjaArPchr0ghxqwJ9tv49mTPWo8PXWtgtzAzN7LK58h47Lp2R
cUl3A6LPgMlEOe3V9rMeOPkThcvoB9SFE1QKV2Dlo9Ueh8vRV1aasuany9vcZKHT
1jWnsE8VS7yXbaS0aHNXAZ1VQLIog+TiLO2sjNl4ZD3sMoP/Uire7812na8llCu2
8dAIQSW1LGyuouS8xJYDvM7DwZmhxSwK05NcLynZfAsSucGJhKEeh2V0p/azPKyK
lUJosZeT+m2YSJKmh8YANdYRCAF+uYr9SLrZKknBPZkukgTJbwO9FYuJIriesvDt
Knap8S5qx5aVB05lLhZKIF/27Hr5efjADswTlfQautwRw5LWFTmmmXFbhS/lHIJz
rVQhS8aqp42Z+DNqXCbWVF/ZT6i9GQ5KDdrw33Zqdza6qqg6M1HK2a0biMQOTsBJ
PVotbamV14Y3su6M2OXxd6KOwf11uh3BEYDnimgu19TTimxd+/Kihguf9o60emxG
7xWdH/Ilqh25mFn2g/X8U5oroOCX4hzprRRywz6TFtqV002ZFFmljo9dAfob/3Ng
/scD9IKlU6udEZk7wel/NZoC9Uf487zuczA/WugxX+vwUm+P9VXNUxP5lFq4kMKc
G+ABXYcnHAJvFxy9RBhkCoEJbo7HSX4nlgZlVfa06XMotqd70IuMGhCXN5aoaD4g
xTkQPknOSanHNCevyHwItL8PEQ6lse25IXa2djcltLJyAYegUVqwqkuTVvHS3ppe
Wz3fJCEWbfx3bK++mMRAKj1Ven6nchbvUQXkQI4a7rqNTpHvnMqgkEf+yZZObkOR
LqLkrwD1723d/5iNlWcwPV/XyOB28NGMWe+7gohRvS3TGHekSEEgiD3701ZF+1oc
gbFqrrsIXDGdHScUabRCf9kOIFHUrqAVpltgE147YwB1FAEVHDQjO6ryD4+GjA2j
6jpDB6DDkrbibqW8NomyzExdnMeV8oRlHCimrSCcv3QiyTn/noF+78BfTmiZYt9m
J30UjVwllEG1bUth/O8G7DAIIGq1JqGAsS9xapIGjS6cyyXaN9WqLtJ+ukGQ6Qlu
SuiwJA9/iVmhb368VroiieX0ke+tvTCN5toQaEAOHNgwsmhmFZtkoh9OrZtg7KHu
vcUU++z6LiDZH2iYDwbS3IeGqVxv4RGdEj337KFTEyrBkOihCrAa+3OLk+Qsx3qM
ahn0KG6797h1RvfifZZpuepvjw5db9nDqXdmqBAN+n3NqzfQVlqjvNnQPF8Qdw6h
fRFWDxNpubzFCV6eaEkeNHpcEV+Tee59QA4qVe5frQDK6Bycxf4L0CAD5KpJOw/0
AXSQMBGw3qfsqDLEQNAaWB9tAma+RmjiAlXip9x3TZY/0iKTUuF2XyGXCo0emYY4
2mbtlUsOKkwu651EdiQjSrsIlkybwaqIMzY5q9Ouj29DOF+v1zBz9N+yN6JImMve
8knXOhnd3DxsEnSFAKGgCn/iNqn5RdcH4dmHyZepxjsHt9Hz6Z4rDf6dutzYHQTn
3jdEvl87Jyn95bz5x3qIMBdKHo6ZgcEhEfvVHpQaubZ31w26O22Vmgao8VJSI0G9
fhja+ysJeyDh9c5TMgAPvAKrj6aqQnoNe++nkO5bxbGB+wgAoW7ynHzaqdXmSF4O
yZBYSf1aGBrEtaDP1Fr5+Wi8h7HJ2TthTCOBxnpqP/pFRuPls3fd+hhZZrIpheug
h5YKGFCkG6xWN6Gg/ehC7OkL3uVcIgKLe4+RKWbE/8q0dcbbJpiTrpxlgg41IN44
PPErY1Bgouzli6YyohLzLpJ6mpEbuhphasSMr8Ne7ttnX33wO6TvpKhYSzsKbhNq
fnzTrL5HbQTT0wpP65LYtf8Ti3ZnFKrqC6k0/Jtu3HaX8sJYyvRIhY92W9lndKr2
58R+YV9HkNBR1PBwP+pqXLf2N6gNUVNR0OSDC5JXHNIQNYJ1tWcdu03RcXqPWKoY
tMroXyC7yToH9+D7ePu2qpO372QJU5uhBgSKpEJl/mwiFBYZIXWd905sWFpJd9sG
avh7T2SbQflujIsikJm23x37lfPur2i5Sdll1PUt4LGJd02VyE62sRhs23t1NB5j
CBd4efQ63bY+qNfOItsK+hEN9j/Az5OzAlq8oC1cxmLPHFk7lg3rWBuINCFfi4BN
YTmS6FW5E+EkEj/bKlBue7xw0Z4i5oyTavrli1yf0smG8AtYJ52FTkwckGQ7uZH7
u73c+7eiJZz/eqNr9LF4ThcLWN0SQYrhf04tZ28hSNcIlV4lUJz7Qtp9jQjFPlYO
keIMJD/+9iUeW+vefl5IbXgQiwoLygMZbtBKN26hOZYiTldVpoQKxIYwlSxs8nx6
byPVfdxaWGxtBaQZb+amdPiVuq3UH+b0KO+0u1oZfcYDUwIx57VfHwq2EXNI5/4H
gGt2y4hx9O+3uQ6QC/pvsrwF1G0b11f/AshVpZ36SsXKkT2GNlyHCPoRrCH8MEf2
PSSnNjbnqC8vYCG3Xwnn9ltMiuUuvx60pCcK/+elvcfw3DbfZbWZRhACdqOR0tKJ
GwzJABPv80tZYmPHHUZX4xCq4hEPr1EKVt30LdfkY+pakV+r6PLoxCRm6tVbmgbz
GhkNj97ParbdQKVn9Ft/icAnwA+ye5/xBOQEGXeiHaHwp5g+GEKksJY5FU/To+4o
Rlhdo8EyPy7AddI3NHLO0U2Zkh9ylGeR6JNRH8P2UigUJFJfH08hvX8SoqlIVhGr
9vmh0I7nq2X0oeTfZJu6iSgQesiZXuBOQ1nCM/zSY6G/el86BIoOlTuGq0ybT05u
Xc16a78V5oRKzD3F63JAKFCG5AD79jcyAxWJRiCQFW9gmLFoiRKpwG+VaEpc5ZBk
0DYG+ZmEGifOIKQIMk0EuVqfFbKbV+hUDnUg4UMxvvKbhgB58isf7awOzAG5Zrkc
47vQDbwfCHFi48V8ncRpjAbX2J0rk9jSF2Hq1XgW7TjSbNSlkRRcxkUGptlSAuy1
/Fcup2LgHCB8bWSh6msYw9RsvQ3hf3tj8Rh8lUbgxuhaH8m5sjVqZ4xXXhgtuuEA
lmHpCUr96+TVjF8XtLNi2Q0Pd/ZwFSUzBqedRZHwBvhjCFHkmG09nNqKkbA1LKfO
b3j7yO2llIUDNjslIdo1DUX/dApnsgPY6PKftNO/TgmE2SUrd7zPGcMPm4w23s49
CugFU4BNoMLb5EcqYRfoCG+wm1RkCRVKRvmqkv8mcaq4guYJ2xDngVm8u18gVBcU
CiXNziw6jR1DbIqWaFqtlYCCmPLy002WYeaRqURHQ6eryk579JEEIQg/GEaft2cB
wsLfqmZHHSftUHgvxS2KKsHm9zGcAESsiazyefmZJR6mHGHvMr/cI6nwEPcLm5Wo
qCnl9atAX80w5YPDCNE4v2CEMceYoBV/J/IjckLZevwPQqMt9DAJaktXgMR8T5KM
YAcmUocd1wF6d/Z3PfhOqBJs8A14PaNc4LTntiQNRXqec9xnR+YELwkdSNw2Rxo5
Z63mKCUqTSOqvmXDQ5bGX86ABZJT4T/01nOZQwMkMtWswrh7T05SFCo6vWtqreCX
TRBmoWryGOYgt+O870Dvh/8tEb47c+Foq/8BLendqlcKxs2Q7Lws2x2AY4y+N1t4
8p2wl+rMiJML0/JKOwSPH0iSWkwObAEUpQ1CaMc6xlGncMDLkqM7ahZxHnuWkhHJ
J5fbvepcdI+T0keeZ4QoVxioCj8GoUex0iYs6Uj5PnlsTn2tENR7zQ0VLejqsp0o
XuGFNQBa5QLg/2zsynqag0umy8uwFeuflkdDDmeiOEPaeu2PEzNvLImYdHiPosIg
iPtVj/9mEw9jjsKcQ5/nzgKWcgHac6H/KCBBh7HEVHPbf9kvkROxkbOc4Qp4Rdyo
8yseEjMdnsrhCkWLV9nWwNbG5s/YQxwNdRF0uvY13W+qVQXm2CMd0/SxEDut6uuv
c6PXVCzPthvaiYE5j6m/0ChoDM18FKOaoxwv100Ct0FbWrURORIB/ITUZgEBA2YR
hscKD7vtMIHd6aeZVihFbUmzUZ21JN+oQjYBZ0oh27RI6M0AakinVWlR/0v7+NlD
f1lhrx9z1BfTOeZ5RiyYk+nWGQ/mWABohZxNME5OW2VQISZHaMyzBfqkz3owPHHW
spDqUMqxbbaaotUKC3mZz1kR4RFvUyIhOWq3LXUxyEKZZN9nJYpsBSqcluhtsxq+
iOCSmmRW55iAm4ywXEEs50pUuLiBfEGOCrL2PqIiBnOeeUQPAR17OCt7oeo9/vWF
uihnX5QtJc0OvxN1GO2tBN4IhXo0Sb8HrwL11kQzeUTZtYWIr/54KWOfyfWBYx7S
nIqIqZpv33qbW9l6g57q9d0QvtFj2dw3KDYUi52FzIT4rwqjhRHROkLrN7N5DqsL
xltTypuybNdu9iKbZddeN/pDe1uzr2qjbPI0Vkds0urqIywn5I7KqzAOUZ7sGJTv
UXMDEHV1CMJiY6uZtvb8dURkTFbYe02uBbdd2pdfGStHsIegMu6DZSB753IpyXZ8
qGdHtfhaJX0j8phLBs1M5oactkeXus9PMygrtyn7IIST/ajZE1fNVxElmHEGYSkp
YHiGxVqX+PCeEWdajZame6YZiGf0sW5Hnn1BL6a/L5dgMGft4I0nFAYdDWPvtWaq
/9f+CNgUWlx/W4nQ1aXadpBwef+sZCh+3/pR/Q3qCoSSOMrsEp/lB5ark1r7z/KB
mAB+AV68Mt1J33aOrIkgK5VKtnzeElOeivDAe6Rq0RHN6XPw6vXw01PZE5vYOsMu
/IRglmYbLvN5/OMuPC8+37SZ/rwIybr3myn5bYpeAURBmBOZ7vmJ15kn3qEDGh9t
lF0E9gY6VNCuAj9hVXYFAa1XwRZQOFMkpDayRF0LqHhJVSXJ8CYZ09HGsd55eQmJ
mV+uars9RZ64MjUo3nVsz1Iah1KypDFjOwAtIM8z78JhS+sDP8dYW/PILtUQqIUi
lOz2EQ1NckIP/8VV0mj9P7hI9nY9Trg3hnotIH2wMtY3vo/4qzoVzcotN14+989k
iPlhlrLo1bMrW4PjLaGmplJ8koor1q9s+d1T05ziF2+vAGkd8BYmhD9sf6uPxEa8
EB6KMPcwFOWLZll/4je2QPbVD1xGllFbnJJClUZ6ev74aniYwa0YVrie/4UxoFcF
BI9FyBXBnTUIeW4nvzfYsdhQvFHm9ySvrR3iiJ1xUdFr2yM2uzTqgLVBXXQ/yV8y
g0yCpjF40I+Kd0W3VIsr5M5v0yKZYY4btSem2OqUk83X88HWXuWt60Z8K7LBZrzK
tcth44aXm5GuT7FtqTpoeZg+Ti3+sH+e6bAaICGX6rZvmU3Gq9eOfwurKcLWxg63
wDjEWjVdDsPsLkASE5w8Ms8hJEDlGikaB6DOzFkCV7Ej64lomgGFqJHgAmdCQHL5
EiPKsJOKGtJSOTlJhJzyGC14cAlfGP5dycPpZbirt3YyDeiWh1PDgffr59BTnM/H
c/Bx7jDlpd0wiLIP+M9lx/cPsfZUpFeKGOEE9gS6J2dwgGemYreOOtiGFpzGsL8K
hCx1fCfDLKVMrITwSpqlJm3fgFWZgpcXGc22LGb2SR6r2VxMB/5mvbOm1PYmFu7/
3b99lHJUwOi+KzPBeRa/2ccdCEuFxbMY24sWLdF55/yqqhDNzvi8keFSAjWg2Klf
512gMLmxf8MhE3Rjgoej8fG5E78Z1m8pgGJI92rgxGbZYVlEFobo+dAMnlwGrNB/
h/dn/bZ27wxAnTnPf3VacamOLlZXVozyUbiV3Okylt7wjhau3ttsGuTXmS4q5D1L
IVVOqzwhb7x2pN76jWSRw5g5JsTSaPHtpudm3kb1QdSJ5YH+6R1UtJHMFsAeOtE6
qsahrdO5SF2DvVh9yCqozDho43rN7FUK7g4jffBSxLYlzhYahQO8ymjmAsF8gX04
7jR0tz84RGXSv+t+zipD6NgTCZVADtxgKlXNJY08qrSiJldLSPo8r8X3Qq2WSrWQ
t3WwPC48e2DAemeur/xXoHvzvGIB3kThHWEyWkbZjKrdoQT1iEN1ANt0ndcC6V0D
t/tg8469dwgt9fgG94PmRZFfJV8Uau7LHwnugvwb8qJ4gYh7pvYoiq8ttBlU6w/A
6Ptjs8Txdr3xyd90ReNmLtJU4hZ6aCGFdYkSQFgLEBOiDDin/G0dsII/et8lRo6v
oWURL2DuoxEh5bsti1G1/+N/vSVO2TPBbfz1SX5avlOFIgYhaP+xVif7AUCghkZ0
WwxKdLDDsiEnpru2bHJKoz5oMbeXIsXzutsXQzh7Di0WMz7AY1pI2B3q86lIynT2
tcY3qRaL4PcMoQMM7VuOWbc0UxJje4rjlcMiLbaEAX55XSweEmy8060my9HUjPZx
Ozi/9gRO5oNRrQ7JyWtdes66y+L/ZJZSYxnQuBBeFciy9o6JAlVFg5hamNJvwnuM
yajgfrglLx9L4lPkDjCg0TOl4yRIsigqMF5LPt5p2u1Wa4xq4YPcCj+gnprGcQma
/DfVq9YIU4uv3k9ElGR//xoHVgRgTTerrh5f6l66KAFvyQzfPs69Z+zKoCw5HOlF
7hiFsNkgNA6UZaU0g0ofXguA4VCagjsDWu4IaE8ZoA2DKnoPXg6Opi4Bos5nnbDN
Cc6KNNg5x15erfLFym7d/MMOoYoE9wI3L+p6FNFxm00//ctGpwDG1kiXVKT0EfUk
GYyc3KZiMlQTJ/OPJRqvbnmwInkatJexh9oFDQYjf+gXo5O8ByQCKa+hMUz8Bxh4
ldOxttlv7E8dNwaGlIk1pD27ijWCReZOLl4QCiz7GTUgw5Zw+pMDC8V4vF00BNWa
MovRx9n0iUA4k6BX7nUdaVsO93lnAcBS3+ibHTa/ckJirGPwnaxMI/6bFTvV4gxZ
tp7xHzl/qCoN3XWaO2ZEoqeBPYohb2PMFG4JzXN1cVNTeFoQNKgc1oI/Q/KAXJK7
55QufT5W5xwW8Un0W/53TT4qVTXnMTFufM9UPwcqmDK2AYwo+Zbv/5FrmYT47/p5
W4Rr3d/6Mx9STMgw3jW75YIo9dKHjVA+8Hd3rk6MZjwa42FvtAEGQs7ZlLyrkpo9
LAiBykoRKtZkdJkRN+ALufJK63iZM19q8rCfa6AdT71JJDyeMW894bl5WzKe9mQi
QZ3oLTJYbDhs/o8Pr28icOXnUfcwxUAvJeCOD/zZM6klM6ETeyuvjmXUEmL7s+KF
AwGOxdWeAMos9n++XRk1lToIorXWccg9IddoVjSP80LMeinOKwz9rQZTqLsqVx7x
UBcBzofActwQk1aBk/q2WQQEq0Y56TfY3bTHQtyT6NPh38BrlStXgYlIemD1RjHw
ACV2cO0WiwUfxVwXkRXHOPq896+uq6y74+mHK1RgD7d5dQmNo9qrytkxrNDCRdMF
1fxI53L7MPWjXeQLjwMnSHizYb81XXk9y3DP5cSvCqUWH0d5D6vng47Oo6iFAOhW
frmyWv6tTCtARZIGHi1pY7wdzWqu5HjGxp3huASzk7/HjWIqLYIFwGDag/7qcawd
TRCHaUSJMuCe5ZSDCJO2f8fdteZntpbR0NpVt4Mku4Vawt2pJWDuWT5MQSMOkhZA
4gybITm+LgdSOF9CB1ZU+a0Ek69dFJTHuedEwh7rWekc7s0KBQCGKo8VqbA7JvK7
HXxqiNo3a64YtwD5ia9UsH5n9+DnNpwl1H1WSBfz2q87pQtWTxzAu9wg1JUT54F2
K28VpSpn5W3kZgd+uEA+LIuqS04nNpRZmIJziUrphvBIIGVij6gqabFGW+XikMBY
FohxiqK1y2gmfnBXQn8oGfC+VBEnEYSC4mxxTlkXmtUVsIurOgWa6CnX23oSBv5R
QWV5AyP0cyuj5vDjlIP4aY9a512MuVQuZBBDXXyS+X6XHwL/AwxRllR06ms66jnS
rKn58F7BxCxQhRk5ww31LIbWnJm76Bp5Zg27BvvIAOEJE8v1xrMD7QhxMyBfFYaU
KQFRX8BgzHB9EaEbd+cyDMGE5qzl28OByedqxp1xlRsQLioR50K2Jo/mlZXB2Dz2
HjoPLBJi/cdBRJ1DzqPIP9nN7jr98OHtWuMp8UvcMQTntq2EPkOjn8pvNtDEJbz7
nIlf608tVzgasXXtzXIy5RAcoEl8czFIrnT3zWvHMqOdEg5innbuGrwLCBhgpkle
GATHyN6bIb1lXuaqSyZBMIag8G7JbM9G0+mj1txuhPvCrA5mCXzfBriPCAPJnGZQ
ofB8ck6RefFtkuyEV5RYe3GZ5yPNtCjK8jzMGmP+Bi9i/ipvpQKelKglMiAT6aP6
F8nXy5OqnegZ8pRjJJaiUkufAAPZHbGL2NaaHR0OADl75gpoHqEgHBeyXyTFhhfH
ipWhqMD09WbhdCmDxBJp2Ngcc5F/lEwJuPvK8OstMpVB1ON0cCsyIQa6jdBC/KWQ
Yn68JPA5y2K31btfhVIsu2N0L8kT8MMFYg0D42Mr9Uq8V7H1AE+BdhgRvUWK8qOg
p9xHMRNasNctkfWUYjEOZFB7iCP8Lqb9z/RiUOWoO9KT+dDPnJXJ7N773zijZdnj
DVPfvcR/rZeNhFSyBAxRa1/JcJ4JN8cqs8B7Ju9EtdVwHJDxZEnNSsJ14RybAt6l
05BbO8XV8JaBiPaR0bk83rFXxcHCzSd3WMWxDb56bHcptyCT38Wdj1bFJL5raVGM
er6ZFH5XzmBE9a77M8HgUR0ljwTfH+yD67V1WvOWqRLxWp/a4BSIk9iPBLwsLG0C
aMFDuDkcm8aO9G6kNJkNQpIiCmFZ97sY0j4BJxHt/zhorvXK4PezyuxIVPgozOcF
h94pUYq9zBuZ5jHrDl+uL9uGhjDKiRqfCGFwNL0hLWQZ0YoRHr/tP6cXKMbgCV+H
7ITpQ0AEBPqSmsoXbh3WuFVjmF12yzBBAo+qykrLBB/BXr5GztzArOB+fKdFrBXd
LjK2XjIRC6/mpXjNjU1sv++Gf1pJ+bI2Py5LfpYBs7ujfKKL24tOmzttwJmtWtl9
FockBwRWhYuf9QW3iD9y7BCJMxD50LmmSxfxAxL+pTbAm3ssQ5dYA12f99IJbTe/
ZftujDar37pBVKfxrSKMfWGkt4zxJvUtocF/HYAnEAGwz4aOeQhb5wzBPvjF90/Y
1kJnhLA6LkVLqlaBTNqaVIV7nNGaSWc7Wft8CTLBcCblzTYGTnK9KiPZaQi2Kcv2
35qFn+7XzYZMSu1X35n7LRjFRYnkm2vMGDb5T/48uP6SANk/GfcQIR+h/2YEZ43u
6CTi/ePyuR5iP/TlCLwQ7FwtXXPdoJGIvJxxmFACvX1vtd5BQ/+jzV2N7ZM6nxdE
hbhkqDQ60Ij8zzapgpL2aC80/XvAd74yboiEAuYyxNwp8WGCczcLFWx0WJOb+Ho9
uAwwjS5HIZiY0zckjBsv4iMoZosCs21ZxyflZNMGVKAHtDPlZH8rhd+72v5wndxD
0aWc7H/yzVSGL13JC0RK4uTTa9HAVEry85k/QhuKOmUD8Kn14+gq0fZl8j59qxFh
QrVmFzpgVWJTH9NhOyrnyptpIiHuWfNaJYka5UokB5X6dvjRRyueq+BRA8AA9ULV
HnhfZJx9GvZAtvHKTqY+cSpJbkTQWt/E0kRTTaALguNgQsbq9eQfhTyAPaS0qvkL
/S6EItdM/k7qf+DbiqE2gEdY6ShSChniUMRz0or7qSMO+YxLD0QSUeDguka2dYqA
6tvu8GmEXhjzTqCCI7aLFMoQBrTVS1k121dhslbGuE2tfrEw3PYezboDbCdTTo7z
McIYbOGeVJfNpeHLUp4aT6tj4YjXJNNgnHPifEWFrF0w8Ga+cJL/mOduiuHIrBAo
zC9m3qU32oanXk8O/gyAYwc9ZShPVg+3kMD+h8fGIUPjR83iESneCb7ng2RgD+/O
aJ3oezZPKdHgMDh+QvcMgwFmeSeX2E/UL4Uk43gU792nIsbIaHUGMmeMuj3d7mcX
z7i104JK95k+Bz+FJbXdCYpqOwAQKZaSALjGO04meq4M/D1PZv6WdIg3BWJEZikf
yfskoGgdve7PWmLGmuHkBdGkNfER0twCdxRt8AWdpYDgpEk1Te2EFblKTZZ4Vg0w
an2wCfNjFmLt/DVW3uQi8PnHlY49qyQKhBXX2Ayt66k/J2eOszvi59G2QkeXEljs
KNRauesXUj1/KeDgO0gRA8wdk16dAdMi+6+l4VCVw1Kb/rf4FhBQVAXlk8aMFl0d
P5y+sa1Ns1lCAdncIs8MTR+aZ7IVsdcgOnBUGHwE5PSgjgBjbQ6sBHc8OYgZH9j0
WTm2k75hU6XvG4wwqm6uGABaUX+9x3N97adLR36pflCXTYtIur5UfEkOysyGb1yo
nxYNih8wEo9kC5Nq7ifpZnw3jGtPxlO35mKLSVwZV/WDU3dGAtyKqxUezqwGP/85
AeglxuUyosdSHHm+rmYAJLzzt/wT7W/5atLWoVClAjpCuB7k+LXdUQQs4+vz0qX7
CoErY/Xvb6nQSfG5RYEQ08BzQXV609WQHG4oIaiQHcZPuM5m6SZ4q+UpVp2XMmHm
qHmTNypo7yv7AZ3J8fiuVLYC86/5GfzPUBE0VlIQ8P1MK7tLunY4uB2sGhGgQ1Bm
LoawcZw7iKmXdX4vIXSJXxPGmDx8LlclT06BVw1+NHy8PyhU65q728N7MWl2jNbL
UTECRvU2D4kRUf1zt+5SRAbmrFCsy3wjrYXFTZgQOGKZ+De6+JyRI5fT91X/Sex9
TOBQjGOrOcTe3VqneBv2QL3tQ317VkG+godd4V/3s4PFzqSnEtfRgZQdFdIlBgL/
1kL7ke3G7in/F2wCBXgYB+dJFvYtxnWsra4JnbThUrIUaQ0bXWJGpvWdsTUUmhKu
Ka9zJlWniUaaWumPRCvE2O+h+igSGN+ut1WIN4NbMA+WYAL5Gqu/Yj54xa9lb5gN
3MzRcVz8FincL475e1BRhRcEKkUlGONT3MHxu6RASkT77C6MlhxUGd4n19bPX6mW
WfY17e/fqXXrYdKC6UzQMXD+GntBW0AQMnsQwWHV9oFsnkG0Dr70RBus4AzmelrX
nnKPuVuovUUSomB4dn29G4xYNB+EBAjm1rm9zgSW2g9zdTUmsPdO/9VSIlDEQkZM
zRAAGB2xUfarTNcZkWJeoECWv10eMUPWrEzeDyIQcvRO4EBMvFXHUpX25D0g1utk
Z1htVGY6sfMkt/kRrp5ERA2WPsQG91SDZZ4UK8E/qcfE+w1MWyc9veE+FpDIvL9R
mE9BxCIoJRcZHEq/30xTMoQ6aB+LQddW7rGSlCeMFDqXiFAEn8H2Mbhj+1QDR6OC
t48dIOnHWeDGspToAsv1k9tPiZYUtbmLxr6u/bAC0l+DsyQvIrO9l4JqiBYEXyu6
q/JgMvWF7iqqqkO918maAAt/y6Oz/tYfmN5MNNf5xdAGl4eMkEk+Wh4wj6kktpgU
JX9rSWBm3KzkMg3Xt0AS9wpOb+xzEpLFYIe/wIabHKra44RNKHmnv6wq1R5GDj1F
2SPKN3/9qMDHiZUA9HFmKHU9ozCIC3/Epn2RY3hXgq0byUWBcCnSaVyD7nO60OgI
tOhx3nrQWJ7k+IZBgzdUpQPFXgoAw9kxKwK0VyLR0QZ2cG/e75PQU7MqPeho/COb
8Rg5SHz2ndLqOpzYQpO7H9Fl0uWsRtFLcllVOstwa+czd1EnTw+DSkltILCHAsAl
SERIS0gkW0+4X7AbMu1TvTSIEqZ8KhbFoBcozxp5QpyASZNFwXd7Cbz8iW1HWk3p
0bCh4yw2kPTyCDXvIUO3zh+Q/Yc4nLd5gcTaA53ObI9w8FNRGTA+62MB33VWEcyk
Y2n1CjHBe4r0gYSKfTS1YBjuA5hJbjv6vepKKl0uCSfmj15+gllNASFe1Yf8uYCI
vh/1/2vLd5JTGbda11X6E4v00Q8WiJT9QC9xp62s7FRmaPPcudppH26hm6HaG22P
jiunEBu3hTD6ukM/VBSor9GlWq1ae6lLXF8q2KPmt8MJyhmrR8cAUsmUi36nPRbp
tI3BusA8tGJ3PLapLHUpk83NLmQsoBCRY9fZ8HFT2xwBmoGtaVa0TeHHB7xqsHPh
ZVsKaAv67o1ZBNs55bKsnoFv6eBum4LTOI3hTraETinxeuWSvcqqaUzGeVv3Ar65
DDsitpvkhypD1GcWtxMzlWAIss8a3CQDCmUc13NNyvRUDqbQrdeQ9i6CEJ3jxaoR
LUcnfGTCIuSSObx8sulOh4ys5CwsNORMu2EAyp4w7R96Uu/d2uLsh5YLI3q694oc
Te/jZB/LMocoFy8e4EszMokNO97N4AtQNeNpCHOy+AWyxWu9kRZthdAnbKTsEURK
DJAbOeTdLqOlbg7Tg6ee3l4dLsdHzsib7DBe/XBs/jZsz5Ufrl7s43z6f785O8u5
MU3eimOrqBPdhUeQrh/Cfj/iEmZorsBwgtbKxXXkkJL/ryheFlEIr3u7OV2VlPG0
DhfpLkhivYnDeQmXXNieNEypDg7KX9zX4l2JPJOKJlAPlVWiKW3Ij0lgaVrepazp
zrSuGjpSl7V9eWYabCH/5pKWWY3vOpyYCAsb62NGQVWyd4hX78Cc8zBuCB+0f2qg
SpI0y4nsFKFoZCRRuIB4S+ltspgQMfSMmEExjdYD6ZnAwd+1yWG32Qtnkz0XsvzB
iicuPmQkz7RNBthq653f6t1RRnZfS8DDmmb+olv0+VQlfo/PVcVe9ShSZWNMQaqL
IvWO2bZoPXU4yOcxNtv2yHQv8nSvyRZ+HuYrOehD3mNn7ut0AU1v/rOClHn7/ZJv
sdnjBWsOwkHav9iR/vIpjoLvRp9qJBrGZoa1qdnQJ8FovlWuEqcDWtAGQbQTaFNR
UQuNhym1QsiEUlWJZt7NHQ/dZAFmbFjHEPMYNh8gbcELPuOO7sUOYUQYyx2miPmv
ncc9sNKOVCxY0g53bbdFWcggsMmOGis6y2uR4I8YHHJ5xuCvov6GaLwYX7eaV5WE
jy2GhNXGBI6NcBpxDitoYy0UeEwqOZ3RD4OdeANpXC8KwYo9Ak40mFOgOzmKkELx
mzzQa+yjSBInhH69TK84YlUES/K9FhQKYEouo+8jD5J6S0uFnmmPvuci2USpDgM7
55wzLdkp9pKAzXcTC85n7fOKXlLXQdj2J2Lq8CdDLDZprCAwmRp86yinPdy55c2y
mh1bWg2OzKwb0Rp11WlkpxO/nragueZaLqTYdrjZeYZcmHpd69wL1VZzcXnazFbi
4SYn5o20YzGswD/f9u55MIlyaFTw6u3Xubg/zt6eW3yeTq86ANV5VnpCfyVyhk8A
H6YqFI79LZV96fhhJC4WpZiFNkaRP+BxwdsfzsoVzeZfCk6cu8wR7BGXkf9MkKE4
h6pvstHSmAVRHkZvjbxPGqS7tX4s819w6qRMcFSkBOcsWEGDJYPRzE8YnOpHjqlm
PRSOXw6WxcCQcqadVKp0F6qG+b04wb0N7I12w8kXEbR3Fh8omDiAr4AmDnImE/7L
0LD6sRAmDCpMGHEepHcCbE1yEnJk3h6usJ6YW5PWQCWVgOAOJytVnEKdJRwmdma8
hVvjTntvY1CKQ8fP5YyPkoVeBQxS9ALBmuoIRVzDFHxguZbF9WOgfMwPsb6n2hpM
x6d9lOWkyUMHDv3Nl/t1lIzvXAH/vlk8BSuVjvE+GGljPzXUp2Hvwjdjc0GOzNRw
XExOqHZJLzSQoEJAGxwoXrZoZ7u0HhI3Tyx8VD1HcOoCb78hNzjvQt9gBq2nlq9b
sumEU+Obkj/N2pNHBVGt765Ktu+kgrqBXgMNnjoJ+tp8vvewGYdStGwXJruB090E
QJJkTBALm2VzlNyQIFMfNXGkG8qDJriwkTOhrgRai/GJqvUF5eGoOPTFFPfBi380
Q9gKsVkVdOvi/3oDIRtWo9FVRAM/vRhBpecx9lJqfhigXFzODppI4FSX2rvSCRvA
sgE7ObpavAejvgojGxPIhCMZq9NcOBrQ2zyXgvRDB6DThLnmeJzdXnQ6imlAs7HM
aeFWj1ufvesb342rQniJ/8VhyxgSVY+nbpVlCLG8hphLLhDeyVsTtR+lvypXCnqI
YbWytfMncjnQXuVIGOHd6+JEZe344Ff6Rt7Z/68FlylpQamPldPh/smoP0W+IYr1
+EZkzqQmPsmP6M4s3ET/MXgNSUDf0fnhDLHj+9//TWgg00wvlXK7f4PfJaMgT0OT
wscyVX48QcZ5SLCiX57Lp6uJq45t2iOzq2zwR979kF9b/BcbNJg1hp/mP8GktLSq
J09Opz51TE88Ukc4VRDkvNyoYK3Ke+GeAefvxoAbsfrrzZncCmGQVGeQv26BTW7U
+0Z8l5fTa8IyHGHEcEZtEcRmyDR/uhJhIEWPgZbRruhQ5Pg0shilzujHDeWgghje
z1NOxti/fcVNKVrfqj2LO4XGs/gPbSBD3Q5HFXtjyjeZ5Q40r6U76OXoD2Aa0AWJ
9SDAnsaCxWoYij0A0Tqtg5SOHwY7MQrZcJG7YjrMS6oz2xT/icIzASYFtmAweKVE
p6UxsOv/HHWic9G28iDNscWaFf1V5/v13XaibTUzoVErirzyJCwEwHUX+2JJdePD
6fJiDWW9NyQmod6B1F9tA82nGOKW78G8EF7J3HcwXXEsnGw1aHIDTj9hkzlrPrPJ
+CsYxpfKKYxX55znQhrtF//6Wz90J06Zp+mVkMNpoIx8JQOsUszZvGTUAI8oXUPV
uu2am8lO5gze0uj+N/e0LzpeL47vaLOkjnFHRxNwvuTurzonfAUmfam6QttAmDQJ
Dam1YyoquhY4pBgi1ZeRQCtxTUlSyES4qWj6HRng7wb0fnlYnRohUIGcx1sbxSje
F0yj4inuJZazo80jIYrGWXao/WvzYykxxRY1kIl2Gm1Z0XsCIIkWlrGKu0z3fVi8
/Qji2wOKkTOXgMS29PU81Jv49L8OPzbF1t2ygtCHGgamDGnTVCAtP54vpFmbwldD
X+wruLm+itoh43V4ZVlJIGKr+AByayBlMW5bxMJToXGntZ/mjOHc1VYYfsIk/b68
fAWP/KGf4v171qEq47xt+iaWGrhvqON0/JSoLH40s3e1+gxhW3YoN0SrLdJSvHsJ
IBwu5F1olIl5LI547zkPX1to7NpcRIe4TPgBwOB9L+3EnScrOZv4GH1dqhHW6v0f
LHkPLPzNo5Fz86RZWRIzWsRSIwpS877FN1ndN6qJrTHbuhtes6E0N1lr6fBDjgG/
8DMTTqmaxq401WUDXQ/o4W9kEa1Goun3YJs+CG6FbM0Ezc2goD3JwgoM15BxSnPT
lpGfPfKrhuuiXVlB8VFc1bTbPpbr2wvyq1AIekeIFprcyE/9PKzIYcHCkLD5v7jW
iqq62VUiB47t3daIF3aSk3PeNelvUWyJkpLMFNppSxO5hA2qdGuPoGYK9/n32LEw
tEnQdpnUjb+KxBlkU3b/SpBfQDEqW3mEkBRhwjg1GdAZz5r1UVgw7TnWWw3E/Gni
fnwGwUWD6e+CdMj5jWeRA76+kCkCgMMsK84EIcwl8mK9cNrgrBZIW08vSuJSNcBR
kjD5rLU++gf1nmylXt23Yq/l3Or/zzZ2TzR4pUEwKmQyImCmxXdMJwjkBLfFUEN/
7cPHe2OlhTIZVQCv2Oe/N8qlU2RofxxMP/NGKO5AnkssH3sHZgArFDsNTtMos1BU
JyLTaRInGzO5sCXCxbge3g2vb60Sekyk2iGAMr9AOmzyYs1sDpslOBzuPFYDKdP6
lI6YfObMIsXuR5YMVWnTVVBdYKRt3ahmkc9uPu6Bl5e28hgf3kdlhsB8pX4G3472
ln0WDk5mwCJmal3GWQVKAe5rb7RFZuD+wzyfUePsIPwfWhhNaX0FxLcVjtvBVp4p
CyHdvnGyKowH6S3n/rXIalP7/I/vIQmt+vJ/5j3VJZZ3gh6arlOMZvPRahY7Py5D
UwEACz009ZInio0U9Io2HXT4K2hd+mwJ2y2hCvtnih7oNEPD9lR1b+NHlqFminAQ
NPEFK/ee/K+ymFpaK+fzVw8kUcA515Tm4i5ibboJCbhLbLtQXiB0cPN5gEehb/Xj
+UDGd8SYxE7GZYIIvTn+r+xL7mTkQCWNABi8MH0N0+dMU5VnYdYVWEj8hVIDeMQY
cIfyZ9h6is3/hknf7SPQZySVotz6FQeVDq2HtYgscGc3VrTCCXmmqfitBH0rEpy6
+zaBzNCquG73kuvZ/DcG9OnFWcddfhxI1yMcRZD+Z/o1RuxKxllJEHbVy2G+hbr9
Pl5WuyYTNMIx5gpdvr4E2J4pSTow16X7aOfKK+NnZReEmghMlPthFVD7LLhmgRNe
as9Xp0UFE9m510trvnng30VfXROBVw8Kx9A0k3FBxm/SgDkRHQUTKcE7PVNz2wbS
CBNTS8pQQ9DbiTgbJByWeGwZxpvGQrcBthKrzYifsZSZW2jHYJxgvK38owqRnF99
umDABzutr6pCNQUfoZruqXxkHZWb1yrX1lzHtTRCi4pyxDCOD/rDCMg768An7R7B
BvZiuKL67leeJfo8LQTPkuv8ydgSArhyQGLWIIUwsqdUzzgmnPikpFV91JmyKsKK
yikV+WoivGEIfYoowK3UI0A+s+jVMb1b97wEeJGwHqQpJb6MZ7LI19zLMA8A/kQA
Ga76BXrVS1kG+RYFoUJenqIoLqqjHUkSHRYLdgOfbouaIC5la9HsyrMthwFqF6zD
kOgyDWMFriCZeMSuH4ODuJBEGDKTKBGJGsIyJ9z1iHUyYjKtj2S7Gw4gobi2seaL
t2Sk7ky4bDWun7U/u3nYUFhtHJQZ8lU5evw9phoS8ln6XR3+XvscspkO+xsjhBAs
IJf38bDtxcmKA+BuiYh//IHwpYl0e9K0HITLbBeHdJtYPuyGaCCl5bi4g+2dsQkw
dfFOLXGjcPSpUPb8maOq/W1GG45+0V7C7zQAHFNoNmHCzD+7xJfYmIEhJR+GE2r5
8/NNv4fGeg9/u81fZnXcWqXGM3LfdL0RQMU4NNXEyI8vAxXghIWViBPNgjgYphnj
dhaiSNqImJuwTLKP2L4YJiAONeW4ABpI6LjBiHpgY16+QkuxG7WW9ECtIBcERXOk
Ay/WIZpTdiy4lTmtTkDx+RPYXMQRHDO3UbHtDoWWdeoGBVDbpwZHTSe0nPXxhfFe
VxSZwiUCMv9xh99AQl89SvtCEG863drkxA7UQSEJ7tKnu3SEbhazjhu3hDN72aeo
eyeiJ1JqISMvGSmpBN4jjpiyaFdmkuAav9HnHeR3loxpPfF4c9rNQfXe8Qyk/af9
os/tJmrb0b1ETnFHjze6o7uGsCricaMBSC7cyqmCxSTPCfLgXAzqagZ7ZgYaAadK
e6YUUt6DsO8k0SHaBH3KPabuZ1cvSeaRSWzkYJJE1oQjGXrdHUeAmynWUWj1zQ41
OOhlG9v8oP3x6d5dvPHF28+JGrnASZrTQ9Mji12kzSrCMMkhnFFr2KHKi/Tpgbvu
B8aOZ8LpHraN6wtOOz5miLxg+ARLURDhBjv06fSI0AQcB1kU/VDiX/O+g4tY9r33
jQMlX7k/i8ynhX7rTqmkbInOkfeMYyMNf5KIiWgqjgsqumAHJJmJraiT/afVjTIF
qJriuV976DKQ2K4s5u4IuVHTEtoN6kJsRNBG6xSHuJq86ASt2XI2VeE+F0y8So1z
wqZ8P4VydFBiYTruclNUiN8C6Mn7GYp2qCzsEvMpDd6+jAKS2axsb0Ax+C9ItXL3
cZHiWjuTD2A39XGwA0mrj9bOr7VttYvD+R9SIZj5b9a9tZzpKdozcsTjzAQeffBi
21ffoYbZetmwYfuVVhPMippP71hlbxlsjXz0j0buW4pVWU2AZoB8OhXfoT4BoVYm
s5dqhZlx+xTTijWNFnINlIxLzAeCPQoc6Lzs5mpIKszqHQp06KrCQAFgQZYBcisg
OX0OJB7VP15QHlDltwmid8UCAjvtgW7qbYGFZNnEw6pVV8Y5cTGvdpS94M0a9OKy
hLFRg1bvSqSQdaoEdvynaMFAzSZBjq6K1Xh7m0hn+7YRT3PqU92E7bEmgG6QWQrF
Y1XAPIbqCD5b+EbbMzXad7pnN2QX3dtjfJTeWF8Dz9eaVrm8e8apRxBGo4keMkyr
vDQjUEvadg5I9w8x+RMUb3lkfnEkHonBejmjmzpv2po6OXYlbxAjkeSIxa+8XrsZ
vbWkYCbUW8iwwfUdVEJ4OVF0KwTrj4bT/40X0GD99rFHY+pWoabrCgX+0iQNtWDT
hc8wPlStQY+2GQoFmshmaKKUIoPOmGFdT9IqtLJVUvgCppC+ErUfZAv136j7TRAl
89dA8RPdOuqDK9H1w8mI7G5OmyYhNy6YpvimXgQLqEDnG9VV4bCBhD1zZ8RkkuIb
SdN0DiEU53sFGUUUb6rhgrWHOjw7Pkb+ITmEFFgyd9OWoq1A55ZCX2xObdilIsQV
10scHK2D3wgPFWSscCxsPodVIalIeE1hqi3JyibFgGpKI3hzC1ie1g+j8NnO0Pun
xEg/GW4OOpAvz+F8Xz7pmpHrUG+DlVd5iBxVN7zHZo8scBH7We8MhIkoeb5PYFnI
ft9pSAP2T+v5KLlkOEHMRq2Wwcc79hh+rlJ++Kt6vC0uCCaoQCoUf/6jcg6jkeZY
uvkvOyLEMeeUgLW9p0EnOSMz1Jdta0KoNrJQ+mJESwEjSU+l+fIXXiM8zMFHIvjy
odGpYddNVkKCKWcIdgeTSX8NqPye9ad9qqPC69bXSG/OQJxb3asdokYEZRVumxxF
p07ciFr6RamCcTEZbGczl4jgc56CIaN1KQpJwSAAzRz7gnRD2XsbKY12ieOcXrY3
5WfiuaPdlZD0IFwNCQUtrQDyE5Y8g/Lon3gBS/tGit9MCChwTFjiCq86V/NKe/2q
P8foYkEUcqTF6ySHpTBEUsk/zPxRhYY448tvYkwHZkqN4+dZGF3pTV6Y58nismvD
UZfbFxDE0m14Z6tSlMj3UnxHAEycXQg+7OgxQVg+BdHmitYdgLGwl1goPCVVWi/0
Y3vJi4nU5DNpAMM2FUdGibm+80WrDBeo1BXMBREwFOGLJU0GUoqZO7P7vuhDk2Ch
rCbIgGMXnSZ/qSVl3QUyLIr8tOlCVeITaxAog1n1C7iI/qirBHLk1e0bu8AsYJpf
/+SpXNOzidOlF0urEXyxD0agdS8xikCEVgWSef2DUU3cm+g292P9TKsQdyl70Hvv
FAEwNLHIPfB5OpdNc7pm7uCMzgX/Mbe/tczBu0rmji1F1/3102Xhadj9EblasBnt
x+LoiyrV6HbmspJlDz0w0VdAA4/Md/Y3sEObKneonFBJaP8z0mrWoAtdehMdvkVP
16r+8ugg10wSf3Q0n6ojTSP2ASLs1UcHCWIuPDFrwLyWSqty8mPirzyRcHJrPzhr
Xcn4hq+lsxsPrBMOz9sb9qNccbnByvTi0e8dwjlB6N7QCskOSI+No22rN9c23H91
2CgsqA9AwPEmXR/LuOVSyz7xTMrkx6M68Hby4mDCI/NE9kr9V2KcmkjCQ9Rioxil
HeR0OHHeyzlnChzMHVm5VigrTRzyDXhRWj7sHUnJEom+MMUv1Xl+G52mJaYXOZkZ
1PDs80ud+A4n/YXgatiydJrI6VOYmbonVzQD3UhLHOmruUA5TZ/P3tQXDBUVS4Uc
z9y2JdZmreEc3/IPQUGT8weSA4e3B4RwjaeYLFKmOeUnY0y0OLu/BOzxADEgWrla
hD+buPdyjEYvCqGtkYwf6DeqZ31SJgh31IofbSaAwwJ+LdAw1cxpIq0jjfuOX1+4
TqqpVG87Y9CLgc9LCwggaiSh4mAJXJ+LDqjn/MYh4cAwx0ZchczJGNXJvwLQmbIn
iWvUwUtnB0alDZLIIH7my6hYgycKqdidlvkBAUnHNzA1r0QT4sGOnTI6r2O349N5
jCUO2+zJb27FhrahWKStTqkkjKHVvmnSbXuhN16rKszniHvyFi8p94VLwcHjX9/9
sur01pabNCxT0zJNiT3sS8sqHGMz3sGIMy1weERzzcDFg+Jm2K7k02TKBd+Gu4DW
VESrW6OOOqWLCjDtSEvXXo1QuXfqfYPEbQT4YylM5mhmbaJCNYAD+54sOCnc3V5s
k2foaZ6yzWdteNhqYlKsetpN6z8VDUHjW91r5u3j9+ef1xBDG8QLtPW6cPTmcas5
SWrgYJJnPR4fIs53mz3sFhwaUpEXLRB6wSKX3x002uQyXlfWXaEC77T/X2d8tGUC
h1TCua8r/iek9/WTlYJgNLHPX0mPGlwr+YPz3hvCTtOQrhV1aNbqESYjAz3GYf0p
iCcTiAQfXxl9MUO/UCvkojEJCVuHLdvKsyr8vIWA6ieKH1qJwGvgkirQ2vREtIE8
zfK9jWKoAh8crZ7LJcFVr8rFnVz2egBZ7z/7x/I75ZoWbZHU8Xl4mvyCjKtgAlY6
7oVhfGXSR8IdvYicFFnzJIIJ03Gj7lsC8G2jDVjRTtscvQGHC5XnbUNChqrHTr/7
wMq/2R+MNAn4W8/w8geDAuCckLEhzAxPx3vv+QMExkG9NCoYs13zDXvY4U9VHL69
46/XkdiT6ESqbTgCgN0N8tGfKs1Hgwct11G0aKff3FP9RP4a66+fZ/xiBroql3S+
1uXMCrlQxiQEhLCRCrpLA5FR/zwmladq2K1xeR6JfAgq1YVj8jE15HDjip24MM+g
PyeX8Mz8TLzc7gNExtSsJkFYNyMLL3FCHcFGLegjjfNU9WLJEvW5VImHUXa94u/V
3tEtrCDM7pFweuC9iAm39a51DQ0nkSS8BlZO0IIm1txmbKcscZ4reraBfiJHR9h1
ClLOD1YtZ7ofFe7wipCwaawtHhj5vvGgrgwKIVx35HZ3+QOJyK6egZGl2CHBg/iu
Bupt2bW/8u80o7LxsQUw1WlvHoSYuaAifpUJ57uw/YkCn4ZcVNJ63Xf/tiTMKBnH
3SEhygE9vpkuOZWPeRoZvsx2LqKDH3M0/WiC4Ode3CW5Zmq4V3FWWmMIehWdA0VK
jOuYHcSZE/WRTW6HbdZ3gZu7KfaCwHpcyrLiRAzn7a0VEssTPJLwD/bZoWBB2f6D
4EgR5wkAuXb+UxzYM/5d4LBJrVlvO88cigBL2bVcemYlZRQCz5BouujPHXcq1dha
Bd7aLbvMUp0z41ymGADRUfCxIhcwVVX1H5wMAV8iCrxqU/yNO/huPzEY9B1D9K6A
TbHbx5xNgokwvSz/aCvGGBN0WdqNEQLIRQnKTD5Tm++gGebyQcwnYiXXyKiOZND+
aLdwfL7liIRK7ttObycRQPAQVtZBd6p/T8fdwjb6oJ81JKg78u3caG1TLS1Bz2MV
UK9x4v8NX3LjOFFdJuf+SHj1+bmTBO6Nnj0lbpEmKqUygG7GE08U3UYitZocbzwY
py3oKkHUBSV5aqPB3CRjn2n0QQ7G4avtgxiBV8VpfdcY5tY2DHkYJlF8CZQNJdjv
Y+59f3rNMynmwUlV3o0Alf4M0Qp5fj6RfKlJPTjgOAi1sT0g7BSxOLguX6hU3saO
p0AHmhQJqjpJc7G25ooULwpeFRHsOo2Nzr99slfXJDmzaz8jZi2bEhm8YXCEax08
q8loF4efPSDztW9mnagLGG079z3X/e+qUgA8vDj4IKP4RsdSDYl9y9cXcLTovffI
OPOYQq8T3OthwY/tkeh5gZhTXpCqTsKVboU7F4GckLgjGSmgGEnMTWSSJb2Do6OB
GbuMxJT/k/oCiawF58/olbrUr9DkSomeBVWr66jCYNBVPGcxsBt/Y6n5fw3W5lNf
qKhAbdY1tXQG4KPtIjIxthpXqoZXlAU2FFwGIx0HVKQ00x7Ce7ecn6NoqtIV1BMA
0WpFO3tCQqcoGtlTqN5NPCUdS0mFJnAE2YBne+Lw0GbmfGkSqGwnGUmZPxgsmSh8
gHuFm7L2V4bGm2QCiwlWIIPoXxTsDDCwvbsm/ezBAK8fhZr57ahjklKX3wq02iSm
SFGidSkJU5CCu9E2b3EhWi6FmhotmmTwYKTBXnnN7w3hdEok6GdQoCmM+VVTYq5m
48hcKRWifvJ+RSwx3DEk9p5i8QEzTIDEOdB3VA3XMMn5m+A2BzXzByxMP3fwuy5r
pyjuEaCOJKZrN79hKe/ZIpbjkAhslVm4v3UUuBJ3XKIq8UcSusGkV/8lcfsMWYoc
HDxTdJAWqWSu4PBlCaiSzkFoBvkZ/NMzujQvn7GRhgLJNNuB23AffUiKjAGXIn64
pcpRO3H3GygnEbznLrPPZoFRelYky8dCNfb7n93V6wSisafZbiK9gdVWbPrO8hwU
tjqucwbAAOYPossD79s2714xg8vkD8o2ZB7+mdVmV/pIRQ5TX3OxD0f5Hl1zL2wL
m3rYgm23mNRmv58Z904uIyEWu0rY3hEPjkDwWs62c7TZn4Mef62xdRh0FHDIE6ly
eOCRomEfbfb6WrVnZLg8z5ApUyZ0jUusyfFWptZf3h4hn855mNJlFKi1mophM4uu
ZqCEhROivuvHlvZ1dh+3w6P+GoxrKOxTHHyYeJvdUh2rR7RqeIhy8HlXcJYBWCUN
FcFqRH5QB4H6bJJVEuEraLGHUp4BACRHCMz1hqeJcNy6p0TUOwL/klic/Xybz/8q
2b4xiVATbUctxZVrjx9CFk+f3zM38QTqQNaPsPjsDwbhtcm9mnJUjNQCdWZ5tQAw
A4HkZqecI1b7Bz3jVseaSwWdCf6Cjl52dLgZ/L7EgubLnKle6LDffoZo9C4mCQs/
3LG01xoj/NQRtPgoGDmDpVJI3clEN3bYtV3jKde04V/1mXKziSlzhQdlP13sYOKI
JMGg/Iog02Fyi5Q4UJairjXlK27lhgznESEZsBcDUQhSMUGUTo3TD6UTaOsC6HKj
zesP7OHyKGb98epijHYEfR1WbgqBhwjPbyC6/roysfbNidjqROI9PEZodX/3di+a
9hW4wBcHwvVUSGUcMhpYxfnMabmv7jyFUFP1BXKlDR92GziQE8g5p0B3dyLGdkyP
71XnPggspFZEIzXJwmQ74CKV9+CFFIHSDilDiwkOV1boLs7RXZgNtUAjbB0SGxx1
x24nJhUGUAqAOY+R70XIc69q5v3h+HEoaL8mt5HZ19Mgnn42PWl9biyki+AtEbl/
eQ99G7vD2mG9PhZ6OysG1EM8EFjrlNQCk1dE3Z6DXHC0JknCcYv+1OOXUG6qs2Ar
t5uHNFeFaGrd90veKfxINpf+llkaSs66vZNiuM+KikHRTOV1J3YCTKA/33kTny9J
szPNexdpUqpFzc0aIB7q2FxuPX3honxErOJRqc1dDvLDnSEtAuSfyI9lOlFglpIu
mPE3MHhTX01szY3CaUbbBX8l5HLANP0i5sU/CmA9qp9As+oawqXxPGz1tDImaD4p
5AE1hAR1gzH3IkNR4oOjNYjYwbaqwsAr3HAFSlZqP8uO/j3Z0KHbBk0f5AfQYwrW
U41ggYyKB4jyBSVA9G+YxdIchFP+JYNjMRuh5YdbFBzHNFKL6zSPU5s3bwgdhPOP
i/+Dz6wOAl6fJKvVyerR7aJDCUsmxLHa9bnqT2kkrMSUMESeRG0G3jSmMh6LgTH9
fWTMtw2VkV8I/QZRukVAVya/lT8KLIqdL1rqMJttaeJAQYz3sd0IIEUgCZOAL7eI
l2q/yvYb9Acoz3WQnnonXkk79CGCugPIViPHpkEmE/SD9GSX0ve+2fNFEC3Baqez
zTcd9cGuMSxosq9SSMd4asU0ho3GSGDL8CROrUzHfA1Tz8l4velX0F2Ws/zgdyoT
Upe/BFn34WhVK7d8TigC2lRscKVg6RZsMTyq67ox5itaxWeNGUdAjEmrF/LPh1/e
/vS2CG9vzLeJVyzLz928fQ7iVQjbycZAKc8HqEXqgp8BPEmpq+0GBYEdKApV8LTD
EF4OwPrhDoSTiYMkMvVcf5W8IjJAHamTLMqS+LeHCRe/h3Bdk9eJsctPw0/cQ5a7
zxDZDfLiYcvtVyDci4EKb214lFBdFlnVusSkBsmWYwOEL9M3PKFQzCP4x1JlIiif
WxnB41BHo5C/nWdxEheyJqD7Y6Q02h29+GQTXhypcbvzQHlzd655qzjvfLRoJb/m
lO8EgcA00rMb3+DvcEhBtO/LD+aVYEjSHifUQ1SUrUoUTvGp4gYv1YyC6B6ijr3L
lsPv1nQlu1D5HvQch9YIT7ofYYomBEwuGI7my5I+kkB/3+fVHuTds9L9G6Yn5OUH
hXGaBvnSFoWFSVlhIYm2fN+xDhHgvbk2sfEYuVr0+BiRfM82LRVM2e6D5fTeFPne
Q+OPoEO9QzH3QwinbFG2CzYsbGJ8IGLP25vwgfpel9+DiICMvIJYjBbVrPTF5i4O
jSs6bUi4fMb4o83K6kohhBhChSdmnjmMePKoS0jPgMqOq0Rs/NSVHGFPOBV34BiZ
phXxYqvM/B7gf0DulkqkAeXgEMNdzdmpONTWqinVmGNsqIv9CWHZWsMLM87Hqnrj
HN/b/fBGOBuV17ivyx8Vw9ju9M7Ijt6bv2spQDoF3/uoksxT5pYmf9g5ap1MvXdz
CDEbB5XNJ179MqpUwnv0cVX6AqyOJ4TqoNvnMDIexrT4K6AnjK7gcv3+D3fIh4l9
4L/uMVDgdg6RgJIot9n385uGUhYMAwKTOTRhtT2WWh1yxPlacYz8L+ZuLmpXCVYo
XIrXDpHMbPDkFaeyyDxkuUS+8KCqbicNV6zKYnJKtpv//S/jKbWgWmjtnclhxa4F
G/53TpZRF3RV0kpIrSjaTES4LUq2iH1gpB37LC5Sh4EUz52lHNpKw91ooK5sHeH6
OCswlgG2jm5lAzjQGhYcg3lOz76H5rj6KzqMcdqgI3MpHOz7L721R4yc1KIghwi3
IAIguczIsMo3kHYmv4AZUNo3x9ad5tWMnsgALyI5TaqCJ8eRlwEcjtunA6SeJ5Ke
fhllGuWldRgQAyPNVGceXf95lHLvsAvqwwNFBOLTw370k/fwjooVhiqTvM3tgBVw
PopXM1VJFG0xO5NWAg8tqAorp8kRII6SATSTwsaeqRGlYteaY9Jxy9aZk1UmTzD7
av4Spx39hOlisjAULzeP20GsvUOnH2il9KxBYFvEPFO1Cqga6EmaZZ+Aj/VR4TZC
0a6Ip3TC4pVWawjcJKlajw5qeJyWDQug8o8NX7YVw6bFO3vszXOtcmaMSbHUvsUs
PgXl4URWqLqvc97qrRHMweznKpIHVbznJ4Cy/Xp5C2V3maiwE+bbUFgvntxe8x2O
FH1ul+iJAvYI2RLh+rSXDZvGOKtvObCk3XvAgGlz3cALDQP2jVQ+DowdWLPYop3X
eQJVuZAZ0pTHW9rcBhevcsWXS+42Ubw54WyVduqUMOGtgfyFy5ayqZ2/3cC+8Kqm
06DQjwVvzfUJuD3+lGq7x927x8epa2YToPXTqKJ4i9wJW4PItLLxc/RXZlWbRL/o
dzzaOCdCHtwdXPCDgGIfCLVlL45IACvqKvEI0r9WpuiFUI+sGyWoPxXPZyImbBtK
b0R1Xe4HGhrzCHk9Jag9WYpTYZb4oAHQgOVfH4HnZXdVwhUOnp9KmlfzLV09JZaE
vyQx/Lonz57vda2Ap8VbfjC3xY8b2nubML6CHQLUNAbBw5lbumuLpjleOnj+dxZi
re87s9uAig9IxjzQrL+o/MQSLl+zu4YroWt4p7tdcl9qpHXwln+D2XPsxtnArJ5A
giwODJPIZ3OE0NPQ7TZgL+QiQb2sSAk0kuuk5kPti0+cGmOtwwdLGwZkLWPRAIGn
NHrl03tdyv3Y26vjFVHY7UAmmLhxKjIWMNy9D2RhSz26bZyAyoI7/JDWJiBsFtLG
Xg0sexr2Vp0N3qNkmbBCXQAl6pu7qh0Izs0CuzMbIyU4N5GBT1BbwTJkMyPXn7qb
4U7UWkVBpgqVQ+zcrJuNYlsssU8gasFVlNB0BgYTBW+Mrr5+PyxUufI69uKflQ2A
DjFUI02Pw2TDe20sKRohJzQ5RrimJUvJg1QB5quyaaUwsAtnN8Rs1UVURFtXyThn
8qvjHl6mnuin6FqrkP1eJ9ztqyTwlZ/WZdHa1mXRQUR4BTt5urB8+Hx4p9mYPDmP
a844I4knuvdK7qehpGCk1RVP/lBbH9+EwRT/1DYx/HGR8zz5o+Pxl4uYwjrwjSRb
hwIsUhwKVvzfaZJoYiNUEXV4YKmStsYx7/Ahq8lMqDXtx9T9JYA9iviemkHBsuVn
241Mh6QA0tcpT1Hr0DxcFzq1Xmmy9SV+1boLWplyAYmXxMUbRkj8D+AXWt8j1zPy
ZTVCOazeeMY1lIFPuPeX6ttfAe9fizIw0sJRGeNiGN0qKdG9YFetPgh2YrquO5G+
qTItqHJ+dI2a1eNBASa4L5kW2Zwq2DJ3FBquxBgIa3QNp8UO9376X/U+X9mQq1WR
BAcQVURLKPR5Ey5Qzae/RKc6btGF+jEs5DjzctI/ICI/K/VkUvY4Vqji6FvBBYuV
/t0CwzvGruNLlJeQ6Vo+GhJT0oZQGo3JRsBaizz1qVPxSdf5Wur2nTknpf2IzSwi
SwGISEVR611MfW8MBYeekGR6dbN2ipfQmLczrZRQAsjNYWNfbsN25ZDw7FLg1z2R
Chjprz3MKXx3Sh00HhnTC2CeocAGM1HWQBF9gyS5ZGP8A5pBcPzE4+1OUnpR6APc
T9TE9p0W4fRTv9Z+CeQ4G+FCyjRCfq0eLUoixmWO/UGQlTDGKOYc3W4U5bqB3rK6
9NaopBp54oKIUdLLBWxMWWfW/MZTeq2rauB3QuudA6QTj4vm3sMbst3lV2ZiiwU0
J3S/O0xVCbONPsFFIQMoP5W5iVFExEmhv7fPI2Afbqa/vprzoVVZNSdEkchtPqcU
jAH8bFvVfHilth29KbK1LhRldzexoUOwIjk5m0fJWb5w1g9cq89X9ZPS6elOvpBZ
4gNl+ESPIHhTAYvAt+7YVlxLzKbfrZdexamVoBQF5IoBVEgoIFAJnj1otZgsIQM/
5YFXJp8ftXvQNWNaitcZjWq5HiCX87LF2jPoBr9UyrVIBx0JNI9F+002LqgE4C/H
Qs0YTqwS3p1wwwJvBsTwBtI/mzez87nACzKxAmyjMmvjJMHe6WeNbg9rwIKTeUOu
Punr+kmchrJdXsw5OTEFSKkCiJ3OA+Doqzp8pP+9IAFzkr+FaqoUQWJR1s7EGx3k
j7tnnnKbV/Kg3c4RknAlgIQAAfza2J/+0zcv2TLVONgsuxUijvs+fwo44egiZAUG
P2OjZhB5Ay98kFBbTdpUuj3HzJvCpGnuh9bO82wm7285PGjsKx4rkjhFQzmZU5D8
GOZfeuYrB8aaaZNg7mjGif1brKXbGH3a/GgBWyf7/ffEpVbPAQlO9w34fggEFV11
EtgmAriZSBxVC8XCLKtMrQa7OnzYoGGJ2uRGaefCoAd+QqX1iFJC82ZKgyB3n5ca
HveozSC6a8byMSqkbUdSoOkMiGmQtnR7LbwjdnfNRMC3Px4GIXeA1ZLw/W80nafk
UXD2Ma0aUK0udD98MwUFDoQSb83YLtHXA+AzRG3z9L7EFgGBQP9nDj0x0PoXfEp8
3ASoD0khT2k30aCu9EmUnDibRF7GX475h0MVxOvDgjAFQlxME1jSfOga3O3zeVnj
pVuagZv7uAA7L2zIWNHIM2GLjFs6QFlfc0aOd4GpTLfNMrNDFQtD9CsedXy/iyjC
ofFjxFNfgTqLuGuRHzCkdb7/dCfnHZ3mts6dke+i/wVd0mKLaPRRqkYxIsNSOToC
+ZkDT3brpNDK3ed5mXPRjVS2xH1EHmLjCaXKIdg3LvRsPsTREE2DVOnqRc9ijDe+
xWMJIhtMQV05D3KOMCXj8swhVBbcjcO8R5jRy6pQVHsaTEH3MaDVVhA56FF0Gxto
AEdnge2OAhsOMbDe3Tl8vLa8CJ0cMAp4GFIUJ7DnzpReibeKDacBiOEGSSUpL2rN
n5iyUbuJmLm8P0J3zzn1ci1wS7YfssHbN7I9GfFdK/Ox98G5N8PvMwDxpcev40Ua
i0eEvDXnw7K7nBGAKJnBjG89sfyBrHX2OvITRNNNfH0a8VklQ1h9bAsBQvqH6EQF
EaaaVx6Di/BVfBbZhjmJFsNuSPlXnnEUQTFoIli1cj4TO46vt/hzhBGyqyn48dlQ
vdW0FYux+Zusq3fz2DoyMLmQOdVNhKWdM75pF0mOUHx8OXtata2IhwBrmVxLBtZF
Qe+8/kcz5Z2ASlPc85Rvv/Qwtd/9Tf+3C60SfW3v7rqyGqjP1hApG9EiC9gayhFe
WOhdV4GDfqSw6zbX6v/YhpafSesHYgnr78FPtSbxAXnHJ3iJ+XVz7L043uDlajXF
AQCR6gtoxoylZKhZzonWkSJ9IK+SdfMq/gaICVAMERmzu6M7+d9NLxS3pSL0mrjA
UkUpZtOQ6scSkVvaeD6Hu2xosRlVEkd2nKALy9aLm6l6g6w7/zjrQ+3m0xXu3D+w
wbaDRxQAEgFmLEwl5zFFgpymTItk3SfXk5iLg2sxe4a0T12wfXzRxzlikIMFmEQ7
FI+5gWws2n5QQhMcocsHmeoU4ruQmTbRKrWFaMApvF8kuafW81JOS0zhA5j8vAHj
6AVHN/zqEiMH1MZFD9UuqYBQWQxjLo8lMGsT/J96vh7LSNepD0iUz2i9ytVZhuw8
xyU0tstJve/ql0Ak1ljX2PGZqFk50jib8JtJ51oYwal1hnKCD7gVzPGLWyhUZjae
8aM9CPO2mYteeDXdWa+DNkdG5yV8NFfrcBL8c2mOvqIEotTLIK9uKDO+qTViAPps
W6VSg06/gtb/LGqXTyT9xw5QOeHEa9wE9ZN9M6r6mJSQOSKOUsrkfilglkD2DxQw
PTIQzASgMk/LwtJLJMzR25QEdIr9o5x45sSEDC5eqtJmXzh+iVi9MxsrzWq60Fxa
V+fNyPgnH/FzENWefCZoWIZq4qE0LgadBG9+l6wOH82TyWxZTJUOgvi1/AixM6UF
C57GfTT7r+VuQ/ihE8OBV0jdDcSE62QTStlOnmhfKuS1sCP7Iid59CQN5mlrnzYw
DEXRyF/wrHor9Fpua9bDU97tEykW04KzYfxnPGzqthiHJ2Vy3CY2sBm1SlUBz8D7
CSm8dB2PUUPD+1Krk2bBX89wXqDx6dlHsbxpmT5P1PHkmnQkG5E3DKm6anoOKPJT
V/yMQzthPL6NeBTWaMV06FKt/OxXsh/mGneqbCNnVytIXrhwe5bgZ5lYjv7urjqM
LEBmGWTKMJH10HhSjxY7wXLgBj/pPftqksJZa5hI/YWGje6nnJH1vWKVfsEunMD+
txAKT7ypQwiNFXLS2sQpheKG+HnneIP/oBkc7AjzvTI0lSqik2hOP3N4su+oADjI
H33iD6exWEBA4ukvnh4ODGplDUHO6z1/33f7qtZKguTpoSVW1QZRXsS06ftiUsqd
ld942hlflR+63pJjmru8QLC0eEmXFsRrFmpNoQjWQ3pKK8Vmhq9TjATXYhP7VyYv
dQV2XboLdSFEB/dgnJNcOkJDnbWuc9B6ZevZQkZvoE28FU5y9s4JYofp+vuR3Xc8
2gQ0EhGy7KDGDvxuUXyr3qlN9gbQavt3Nlom0/GG+j649/GZ0I3PdYkOorJt9IeI
bkiPfuz3vE1+OKV8WnmN6PfG3QHv2RJA33gDBGmreplRty28OU1rZVhjFx+U9Sws
D0tOK7keTYvvwQS/opmvkuVHoW/T/y6froh2ABXn3oqelvwNMAcSAfK6pM8L1gkX
VQJd7QmxB3NNZYTyBp5cowqVjjKspFTrt2x0toICnKB/rqPdBcTrtJTRexhrKMqA
Tlux/qGBbOavenK3430isGQr54gk/9/6PFnDWxDB+RA5TNIg1DX6jndWURwC+u8v
z30GkSZyeE5nLh009lfAkKIWi/9sffL1ybYbdJ+S9riCYnJDwW4UuXI2QyoS9YBU
dC0l0P0lH4/XNLucQ9KbNG+0c+GN7YxwtDnxtz6eWOZKNpY4gYHNKVj+L6pKXJlX
H+S3trh+PGbkpPKntvG389yQ/9js69grOP9P5wRslmsYrVkUBac09Q9rQhv/u5xD
OZOsm/7FhdwkNmKUDYiONCJMQbNbkeY7xDd1FkdFZbpbBW+q6qZan3ByNkoBAxZP
aQs73M7kqMiO6uA5r0axVvuGFRpCQAXPbj0OyO9f10FzJ2Z9aKJHw0H6m/CqQCLQ
sQEmzpjcXWc3KI/6ejkZRlIxiJaKkCuI3sDs6dQxNVQGuq9+8WZgzTU8cfWZtX4E
3zt3DZoHexz4HtKaU0UIqvST8QoUfqKUFu2HX88jiG1yoDPfgk/S99IqLGop9HEm
asMs1bWNxWTwQDgJEyC49QEq4r03te6KYj/VizkbSoCLlLRZEOEiUQnEK5PE1tuV
TdsCysTIlWfnAbEp/2/o8GA5XMfRgJoaA3E+ea3uFkpcA8Ac+4bVmnjxfvgkig1n
vS+Tx26UgMw2HkcdRmfanQqsugArN4oHdZtFNg1UeJiksoO5E5G6mbKxEAf7Zsv7
Am9cRFLRAOvdNdc90Eoj6an541ikVG0HNNLFzcAamH/GhHiS1eTEtSGeXUYznS1a
c/tpUSMJVbzE4TKDR61iVq6vBSreIaFzY7BhUgpocl8tS3t9YTbOIEoKtro6v6mc
/qfoc/Sq3j+/C4KWu+mH8Ep15tfunGbAlKiH6wXDUs+sVWsV55a9wBG5gPnIOyV0
nvTWlQfWCQYDqGtMXh5HPUdvCs2vOIxWP4yFcOLyx6gXp7GFftqVMFnXcSYtduKR
dBpgHsNAjmwH6P249FHaKcAQOH25Ymln2A/m2g4/DleCN6fYMNAZWyPgPZx1yBOr
CP3HnBqU6r8jhbbbBdgtQFgfrbd6Jc76r/9K757k1TdXpbsN66iyZ6RmmAKWVaq1
va+hocXbjOJS3pThfHY1OQIgPbiXyNSEBK1G3ef+Odxoq5DJjejxxuIW3s1ayWzM
JBIrGmNo/vmzlYraNKDW7CA8rRE9IQwpcofJsqRriy146GyEsGmPGK14K3O/+Xtu
/fky3dGFyKnbKH9MAgTGdEtSbRcTxdgpjHg3zf8EhW9GEQsIx+se89u1V/vqA6As
yNboiQE9ZqQApF/Ynno/zXm5oV2eQtRvD2CxnlpPgxmZbXDQfZdxjJoxD9c10g62
ruYzDtZEpgL7udHg3r+3f6IP3J73vvD8pcbDaf90nagVSupHvBuAboSVLy9gmqqE
UpEEDw/fFTj9TvYLpdJd9TP0BN+7JPp1nhUbX8RSZ+slA08uPr/sXERI/6PQ8wXI
p/JbVq5kB4fbRwgy8u7YQG44oAXiyx2Bh1Ijkn0jZbDEm2m0ywSvKfNRJfzpionn
mZaQAdo/jetZIv4Jiz/jTRzw3J0GcuZEYOxg0Wwtj/SaQWB+BKTxL98pvgEn6NiQ
+coUsyFN2nsROJOWhKTeM42HRKgOJIYYf+NFyL8giBg4u/1zc2TeMEr95rSoibJC
c1O2MX0vkKcW4vEW3877ByM+IZZb0xU59nsWl9TsNfmPR5IqZKCv+7+FGLp4EnV1
hVOmVr13yPJzc+r79UuKlcSX5UhxW2U2sS/3f1nheixdVIRvW1ih9hvESaGX8YCG
V+cAuH3GrGisUFnnqnMu115ADD5DRx6pkyaRLQ+EBNMc3hAl/0HxDj099FCQhzVw
3qUbBw3Xz+RVe8ToAN4LtgDODz+plEAF46u1Rql8YtFy7CJ/GnsSkJqN51jfAIfb
44cZ1ElMWPqn9mVyRYjTNICLE43nsC21yh/iBLAvvBdOErfC+CAGj96dYL+eg+MP
JJP4bNcBO20GgUWBeLWJ233drt6QwwNV1qMqCZZ/tXSrZCKzH8Aa4Rzm1TJDn64d
U4DTQe/qCVDzPh3QYHgl8wq5BKzDYIYA5EvY1mNBOcYTTMMm963kHHMXv3A/tzPi
lc74t7Zs6cV5iGdLxQkg0jskkWi50zXVl1aCzVo9ZJssznTAcaEgr/5I+LraUawR
COaVimBy/41K3xhwWQLFh7QMdynlFhlbk4dOrVVL0S09smVew58KjUt1Qpef2cB/
hAsZ62ml6q1foG5fBlOGd+JBUJUe5MtYQpRWBxyuZmWbMG3SmiC5QhrSWPnHVEZW
ScyCrWQJNS0VgkYkVFjYL5Od4rsXcyQ3tZTTAKINKee8XG2NFG0deMXRrDK6Ly6L
j0LhASruT7MAa+NtGEFfCzU0gtW6Indb/QrrRnVXRdJM0Wb0SDfeOYSmGLD/gugl
UdOp1k8kt7VqzZ4QJxw9UC0nKH4jDI21pvZQuqJL7/3wqk78O2WHrMNz6OhdTaSq
OQOWLfvkpNCjWB8m5XfLk5e3AZ4dsHROVWFrZAQjRi/7wyipwaTc0XQMm0A3UDVR
69HuU/sWWFBQwLoJsbp3otwNGQQnXFzXL9Yt1QWiD+yltSDOpEVng6EBaMftSdD2
Fp//ViZeApgTv5kggyvY1lXHB0+UBOHe6VSNjjyz/YhkW5aNh6s8XdG2hEKGRVJ/
9TAnzScFTqeiRMX/Ehug7eeSjZETPD4woXWGKqwI9RQ43xQlP4IxfKm3Au+CdfIv
0Xsbn0bYmLjY6rJXyYImQHQNzHx3QnZVmeVhdgG3rPamfU2H2Ml/VC9sEpi7uELd
51q2EtQKZG5xkHOH1McLc22A3M3RZZ77Bpv5RLf4AodXFp9ajAiE3A4jyt6IyyaK
eRblsm5DWvs56fkkRkkl+bJJg1TiCwHMcOJHjYxHbUvI8Jbx76FMz1HX8FkfN8Wt
peJB8IxtDxhZF1vw9rEjHd7HYV/hLB/aWP9b62c2Ogz2+udsdGJjqIqnCtwyp6LC
eEU5Zl1npvNrHsgxhaeevfjpajIosbikE/tu5EZ+bABGWfsYEyR2yzJZ/4q2eQga
Uh6zYBn/Tw77l2w1fc2h+fbJc31nx/9b9c8g4L9CP7CrTFXKFNcWlS09qzPIk71c
ghemaXyL4V4LyNSFoOh9qLIXslVxv8ao6MhvHetWNNparXEEJnwlO4U+2dGNrTsA
631fYjc4oSRPn3z9ER0RzOm/Han+veY++IMBO3Am0Grkg31pUGxc1TudE4cToZjs
atazkm++ciNphbnigujV0z7Xheyr/iPrJa4V5YfyyBL3Ppm50WigI9buxDAK1ii+
9e/9OFIUYrd6QNU5QpQ0N+T+yYIR+008yCVK/LUCcGf+qqimc3BZ7g4rTk6PD72w
BzNfpRqqyG25jK/LwB51HATQf0oJKrvF/D5IT3AIREUwTYNlgEtHvIMTxnJRWFyW
Wnj00gAOLCKUecCIAtq7HmJSOKe9gI1wuECGmpAlZWq9K+jWBuOe65tm2dNn4zWu
o2Q2CQWj3efx/JQQyxfpB+qoQux5+uGTRMnRjTuDBccYTlX+icfFMAjqrUOQewvk
kAevGEyPgrqfXsjZEsID9ev1eTkeYEilz0xFrrr7bMvyjV1pnKJZzOcXbrXtThGL
lYGY0Hn9UPnVW4rrhZotLKjOMcbcgMKW/BUmSsmPVFUanA4qLr7Qb1xr6oRuHhPZ
WybxZljDMBmbHG5MKFpqDcnSIo0et875S9zkzTHn8s6IBwChRE7K2bvmrkIJZgHN
ZHxOyiSZZqNhEgEje9OGxbVt374TLbUJwNApAViV4ZA3t2eKubnEvqLJTKVcMRAX
V95tYj1Lsg+VdUp27Nmj55YqBCkJDkHxFILWklI92VSNPdo6xUOAfFQmaVWLvvyn
DxWK0kLixZK4qnJ4axYZEIQZswFK8dJfXMxjNFS4TMIRvqCLj/3SOtJ0zI2nMI+X
wTa450Ya6i/dSjoWoo8MhxW0wOqkIwg6V8Iho8av0T9oPvXmjLmnQxnrItSG86il
11yR07dQfXp7pgo+I24o9gbAE99oPl6Vk2CzpQC8TdYAzCfxJCczG7QRZmVRmiSY
jpMeM8ajMsMoINyEv7m03xhdTjFt47xaFpA0pPYGqkUNJkNvlIUiIBIS/r2GDFSs
BKoULzgLNHkqX6/d8Hf0TtrbLw6AqWflFijIreVzW53dqQJQrwz3YiRIN28jT8nT
qA6gm56MzLKz5k5b1d+RvOaLXwMbzctdWzn9NY+jb797chbcvTVhSUXNObpKeEuc
TQhFTFjSJhX52ZTm54iwGxApEdq2py7/pLFSmjuAErzYJrcdCCvYbdcBLVRj8LlE
XFqInKAmUbhO3GHHC2jKonVyq2Cwn85FzoWwqCp2jPvGJm4N/U7FRS3FRJ1HHOtV
7hCUEoOhBsSk5I5UfTcMaXWxptr08MH/TZ/e90Jg+YvQUxJFw+RujD9VxW7K6NA0
M2wCXRzH0gfrrZx351dHyHkvtpg90sSRbvfwANw4p3O5G3Rr9Znfb82H9OOK+X3t
xwXjAfHRK66EbUiQ2Uli57MLVJiC79WUXBnZara5ZXxPl0FmAtx4nBMPKkF89nIA
oCapIKejN4+iXVEHFw6uRTMJIr4bQIP8WvrJdBACSPXZop7etM19Pzbr5AAYXxsC
9Hn2oFIz7IThp/u3W2buJK+0f1tBIQ5p81xMiIsRAlwTrHQ4hh+a9MhDFdtPbuoB
3lacxzi8NJsfQrMunACo6sX5CTKlTLi6TwVVr0Mpkpu9T2DUoG5ooSPd5PnWyLtB
6SyVGysW/1nKNsSsOQvHnj9cAB6dVJtCLAHswdYuepcwnlNr6YZ0h3aCGpe2sNJM
iPJBO8H0PAbz3qHsjzQgI/g5LqCkX+tQB/yqSRrFXgI0wVCqnXmSbPLNWRb1Lgct
dHxitki7w0KNaB5/5kQ5qR1ImpNGpaNIqli/elxh4UXPhb/Y1loqIboAKy1dvnby
USytzzmrUIae1r/uWJeY3Mt7wEnXi1ICEPAkUiW4qLzhKKSQ8+4h52hojP7ENBdB
vfotQvgSCP5TmRMBCfgncY68Zs4QJ4JzEGcQYORrh16vGDf1oIGaU3uHuDh1o15K
oTr7KAvbgKjUJgdHVtKohbWS29DqX1UlvcT2cYb6p52tY2s6EYFFPf8VOXuYQW5b
aRs79lfVgT2TH1Tyf5Wasv/8iOmuhF7T12o6L6CjknWUitfIMWOd9X3ZszyQ5POe
1o17q/km9m8CNdtJB65TXvR5KrFoli30Sqnn33s3ml40H95Q1tDda5FKg5/bPpEL
6FZV1DfJ71XDH7qnz5g5d119HQ4QpZhM2iKj3g/ZvV2RinfUzO8CLSKWnGuDA8IH
cz+o+zTFfVskZqddBMOPGYu8harJ8Fmf+Xs/SgGUV9HfwkXithwGj1pujpOxPyvm
lQ0G+BK6x6NdI1QnJTurP7kuTgJlqOyzqaFWJJm7WCn1P6ltgqm/nrjyS9oks4jk
c0Dro9+UFaA5+gnmdWoWeU0I8l5EkHUHYNJ1dISC/ZfI8wOmr/hk7i7zKi0OvGl5
R4LDC8bfbG3jD1f0UzrVwrCG/P2kp0qJhVQBrHqpglDsSoHa4xGSxn8tzODLSivE
nI94Mjf8QJcdnkdDF259Of81GbBnKDvkr2SSLfRFlyWvrL3J7OR01nBrwpjqmnug
FVeG9EH0E1RsW8tnSdyxnQaLJ/ybXhUt5EPdG8ieu7iIwscoTGYLzdvyQN25tR07
UHQB5IsVIGfurvq74De7ZG3coAHqxVJMFFZTokXs3MKMCap+gT6+szD1BZKGLLxb
FZtEXLkemous4JBAIEdjX498Jq6FWo/NW7untxJa3sP3CsUvmEIaWsiym9DlEuHg
IwWXhHMrOzm4UeZrTrMgaRGkwUK9SJ2qgKmVP53ev6/ed7MKGpfFVBKQ2NIEk1S3
KaguFRYbi6WEaCN0UHpWFxD1tYc4IO15RCYeWupGaCO9a4wWYh6RMfTAbNZetCXZ
TaxmJIlr8l0Sm9v2E0T8Jt+Wr6ni5tr9YnKBOxnjscYas359aUPGSccMZFGi4X6j
Rtqc4M3lfcVPu4c+agw4HlGso3c6gjpzTbXQJ7tUw1kCsjTVMkrYZM8TInWD42qs
23Nur880fVd/T7abK13oSX+izXu+FV8asjlJkNiQkONFO/zucarWNc9+ZDGopJ35
OKTdz6JY+ByXWGH0MuYFHLqC/32U71w1zOgKjKQglK+mWLWx9RkwURuKehUHe2B1
Sp3wEW3uvostUFaOdAWLH8YtU+YwMWQTHumE3lDcuKSXyk23+IW7r4+BSYZK5V+8
T+FZfGXIz2lPliYzmBt6IKC3QBE6Dep9yyQWVFu5jRQw68SjcY4owueW6DLYvNKa
0slqUg631BODit7Oihs9OlTfXJBcjIuHJsqy3XLMjX9fhN4gJfduZXMtNKfjIUkN
kBJPvfjW3c04MUFQxlgwl53zQyyg3DXb1bFv5frn5GOtc7+u3noVcvga7QkZx51h
ZpkNx+I9e5U+CJfY9f/iFu4x+uKJwerzXWpCYqvWqfA8CQ877yP01iJgA7vcwWNN
86lQqQWTSVxumy+AA5LV5ZXy0RnEaNeS3X8m60l9nk5WZk2T61R3FBMp9hZRvGI1
rj5EDKse4hThy/UgwHM+JJLu/dYI++DEfjn16mYIhSMf4uYzWMKPECcYF8ghPxOc
4GRJFqcRxWmNAXRbVC7CvpC5KXvedPDTOhgdrgS2bfAdvqBPFe66NsynVTCR7VrE
lVth/LXeU7ZEDxU2hMFCCdcp9EbQhAjJagZLs72oWRBDBtYKX9TxXs/hUBlcZy6y
7fG7gOMdmDyVwzXuuk2tHH0YqzaklUzKPp5YTaraOdoH3n02v6mvSLaU6JkM7mEN
VLkEU19w0Ky6q47dWyluQlRiLdyweOfZaLydal9MSQyFBBajN1uCt22OXJzgANcm
D/74fyBjwhVPGUnERREuNm1IeYC6pGvVAU9UUBupCYrzO2tXw2ajVb7XAcgYcQ8X
6TEopawq+2EsoL+EaDWUzKT6/3ff12yS9ZDyXzwaqp9+EfC+lLL3hNdtOzInR6mR
uYFfkJT963pLY3XW/3CX6DhTDl3ktwS2BoMH/oxrTp1hPrcFXjg/lV3x+kNW01TZ
EkHpk6ko5w9SEiL3QwNB0bQgKhmz93pJHStKCttRgqd8Ix4DPYC+YOLgJ0lbg8EV
s961pB3vtplQogmql0+EQWlnDWtN+bPNcvaZc/+KNtnudH2Fho2DUXEDWxvNf9l5
UVhCeuM7TrMp5AAaybwt+rPZVQ0pUhl9EaBDznv5DHz+LZavujN9skw46OSjj9eC
S+Ozia2iN5572i24+i1icVvPp0jPsRYPtnioLSq0I4Z9oASJFMHvDbbqQhyuN/PH
gKNm3g5SKZxHGDtk7PYThzZkwbgPi3OCQ5KCMkeYUW4py+5MWfMjULHkCtZDKuv6
m6UfGbRKz0caDyAMTdTw8AqjhYLUstjY9dIpkhvB4K3KqDi6zPS1LTGW0BaGL1PW
PDi6QgjK3x/eb7Q4U0wlzD/mVzF/XCwbJSG/slJ8PhfxaqIPNgeXDegM1qMbYF2h
eQHqUBTJOurkOa3/SoQbs8Gv/SfI56D8zbC8qaoEUFwaXMDOexMgc5ZZo4TgHm2P
qjeplk3y3nhLoDINRK7b+T/idq5t5odq5te3pVYTmUyoCoDAGugzbC/MJ10ubOwV
7mToVS0M+cLmrMBL/HF6khYRpedHY4LHpjsNz8c4HNnSk0egfNQHFwnX6kAfAgmV
2gB/05vXv7aPM/Xbnz3IEj1pm5K3u/8LA/FWHKhd6zg59ElDC17UDmLesUxarZTl
REsYJM9xplB7k9x5SMdiX/iv5nZdybGTAsrP84p0UQVteXF8Yv3hMGY7oKMJH2Ur
yhj7GPHvGapxlqp/5G5doJUypRXEiWtM7rdNX3L0uTqC7uxsj6Nu8MymuQvvky+J
n6oyKagFU7ioMQDUXH+pVaV+UKafAKkgNCeVS05bNq2B24yYbRH0Q1vDnTPweipK
cWIZPMH/eWY/GpfvCbWQ68vFx5FGe4/H5XdnDg7yBEZNKRazEvvIYAOC8pxAS1aS
8YqeifTgmBasxqaOGeSoO5zNZJSqlnf7MSs9GdOU4r8dcEZ875OHbk7STwGg6jf3
SWQ8NXWFifXP+v5Nw7wzFq04YgpHiYMJx8aXg/CBcHOgbODsPc5gUxdGKNV57wkR
H3QpK6b68slDctOwYI57SeVw/nYN5C2i5oxHil/gVCKVYTMdVX3OeVS5//4BjyFf
YOIdNjrgZxWvnsLa8YgVVd13By6Xq1JoFhxQ5OOcnCWAWtoqcN61sTj/28qvcq0u
TDF9rbXdxKXMZfCBn0lG9nzJmYrUJj+wFgh0J3yiJgE0yZD38z8LHRBLn7g5Y2HA
+tO2DFix1TcP2KU4QIHKpgoJt3WdBAKVUyiJakgv6mtrzokGeMwhYIQLn2ArqP/1
ROWRCWVn0WoQXcHX1TG7xAWJkaWtpkyyYC/oUj/Kkt6tz9V1aFa+D028y+mcJUjV
Wo+TDv+SQme4NFzXWBw85GVRqwhjwPmWrtQDW9VGp+94JuOZDV6S/gF+dT47RjK/
L8AZz7CrQmcoYYktKbDpmNKJNc9xBdpciT7PiMJGmyRmZXKp7i4WuJxvb915tszd
vk/5RTuST8eKvK3DYGg6xzJDZ16C0lwWbojS7US4qp7bQ/mWNwXgesiyZGpEhYJE
n/DP9wQE02dFFKleW0hUG0B3QLhAk+fQgZNWAGlrYtZjb2lowQAIWrdgGOnnGlnc
e6aG7i7akyoH5EPXSmz/hkencbqyEFpnxCqh3D8cETa8/lEwUK4mr1heTwzY/Jfy
QrI1DwlkXjoRdJZZR5NFC5HadCzSLmJEaLXteNXjz/1WHVyxIbmOZ0fkP5ifAPFJ
iUawz8JgdJW7Sfb8fmIpsphssmMHP2uFWC4bVFSTW+81L94BQtdu2ft3WdCmLOui
2w3hY9eFYBxr23UjarzRdUebKRbBbRc6TVBopqBFI+lPvjO6hnhHs6tYyGcEteyG
fzmyulSVwf1MPBr8IguJvo6IgWub86LAYHOnvfTOuR3mTBsQj+XmFC9SkLkTrtsU
kveM69uN1ZpH4mv66253Lng50X2VqMOe458vnew2N+Tl53wJa9rQ7/4iwlnFkPOL
7vwXAIZiPmJWj1ol2rTbe7ckLG61WlF5+vY0G5zeREyrsc7pbWsGBROvqDukCPw1
doki2IwPFDT+tK5MtjYts0PQZR36sfeKZIU2r9+DDuwhlgbKMfZ1+SJ7Ptc61ZhR
M0epp30qFP0oi2oTgUAw/Ugv67QbtUapquMUIOLFq+tDqS3t1JakvUKrBOmHI2nk
OhDa76OvKTgwkRtu1fbxbN/NlsTi3ZL6NKKwksSk1Lv16HOHJBSrie2ARgZIXJ34
q5tW8G2oI2xpuDje8X/XQ9grWuUpBhaiyEsKPua9BwEJLYE2m2DScnF+7FrtmqQ4
i0jpLnasEKcbz9EC85nK8sPIx4Cmn8053V/l8DcCrYi4iniOwQ0YnoUqmwnNteUd
VKJuhA5tLhJf0RID6tvexHpFobJ36JYkN5ivXv7T/7DlmSAKBciXQsnuea2u3VTz
ndLV9EV99EsN6KE4mq/m97FI2mx2BAzX6DnR3D266dQerKdm6OzE567bs9KodW03
jL5eAnQ/eJkVgakRe3zmjzRnA9p9+qamTkw8qroUDxZgHbRaaMuyXqBnBjgBbl/Y
9RVTeCKLkx5c1Cf6S6heoqwt6ZjbrsGQ64BDUY8aT4SkAQFgv5iEk3csg/vN6aCC
PpqLXdBVidLv4buWDtIlliIkPuetIiK3RCJ9kcx923MYJU5F3ASX82NGwj0+7dBI
brNLkKOrUTWOWKlkIKwztlehavRdQGD6VKoLdlZaglQCyEi9/0CeOlZsUYpB3jKb
UWOEzqefwZNFv5bKoBPwpmaWZFF75RXlNLfL/mPHQvX6hOWyS6Hi725Ik21NBeT/
DMmTTEked0b0sH9MMlOZjMAtQlwKcMSaFNEi6kd6GFGHkKg0VEXH0BZRAEZsB9Ve
McWAGGnX5KZ2d3hRq9L5fGJAUsZXWaF0cEiZnHHFrwW47GMI5PRJzTyQguw4cUJF
rMgfXZN5/Mt3jc6h5t1Mpju/UOaQxJL/4ChiiYdlSe6Cx88V1Kxq38CR+XrDFOlo
BeYGJ5uKgLeeA9ypVIB9G7pZDXxj2S9LvIuWn1T1stNsp2O4fwkRXfHj9HCLIfr+
kXp/Z3qcrxGRpaCeAixs5KB5KsHjvtDZgJJZL7HkcWCO4G91/pW/J6pYAUkh4ZBH
OGTXSae0BtNJwi3HREAqhUnNTF58monDE9m6wsy4ykZy7zG4ovYoE77+QPashCC/
VpTXRtAwKI7e0laPF3+iRMnT1kKXZL21L889PDqPRmJNs/Cx7U2CujdQzMbk0ARe
teF/ez4W7X0LTqDBpz4jcDXNcsIfO4UOzxE0EVZA/r7/bKHn+/6ph8JuPVCJmTHJ
OOcr2KIlgPyY/f23hVj75m+cJEYUZHRsfgjcrbzfpxk9ybFvJ0i1Mk4naOUFUACe
qVoQxWf55Rd9Cv9WohNPVcJHoR6Iqs7I+KX1zyRxNa2EtfYO7bYXylqJfgSUki9X
zSCy2g5BPPI1HQ/uVCQRkPZSW8UmxFjds0ch83LG/ta7U2yFoCpxNGheq7xSyPUq
axHgeykMyq5USWFZY6xdSROv+4ca+6ZHr7VJgHzaBNjxm9pA+IRyZ7FCTcQGS4TM
YGwgSkJm/Tgw/mkjlbSd63fFMayI3mcy3ivBBt3r/MTWxUfRZchheLvHFu73SugC
DS3wsmfqNSt7XFWi3MNCC4IhVR2k0XhbqcV0gm7SO64f8pVhqXoWvl6Q2nCjAtTd
cgS03vdTyKBjj0db0KoAzZhtbSuHNAyFhWksVGCgXPwP0rXwWt/YkXHSv87srRYi
tPFRqANxWV0B53oLj0lscjwij9OliUhupwQXZ4ytnO0vUCT9nlr/Jpzmak/voQ/i
aRNhGcP3aTdNTAF9pQaPC5Wn8bJ6fCz8kmyHtBt6Vnw+4GS1JBl/u42m2b8XUzvt
gHAc5SAmBFzq8BBFrbdFaW/oUg4Y7oJKdHdVqgPuXmA1bs+jv1QzTOixMgefvT4X
nCjcRuX3v/LvmnumLy2Kxk/YbYzXTpOHU3P4F1DxUnVYSGSu/Ibww/eEvnBen6fM
da6FJVH/0VK2qfR6ygS8R2J634TN7ERCrQr35tMa2MnjEPPr7uo8OVr6RGEgxE1Q
npeRUtETNYdBsnZk9Jm3NkLSzie0yWLMY7PDWO86CyuVMRjFNI9adOTdFb8wYC68
wJe/sDLokOyPVvL8tJrm4MSpLDLeeEeFsojsk+db3h/HMltP5L7MtuT2DS12o+Kf
w5KJcOxayMW1PteudRx3n5yt/I4KdlxyAQ0ycTzQPtDNhhObwUHBKWkxcl0SByD3
6SCRUxGrqlZ1Tqvl3OvTMtM1+9DhJaJTcM9JCyd1WshyGc+QcDJ7tsJVSpM3bvoc
geXTBXiuaEcGVXQNAcwTqjNFBlFbGqbNBELMQdH+EElc+f2nLxgv/Ev3gtDWjBWh
Qlv8iizOocidnihRkwX0lkxGMZahtKBOREiY0TT2rjwjZl2N3zEhmDByWk35cfCT
SY4E3T5tQQ8d8i/qwOo82xZvbKrZRaB5eyQM+YFmXe8sce74QQwfvOqIX5yYsu2t
1FwtjrVmeTHDYXr1dbeGe/dx6X9cvY9Wl1O3FZJ1nspI26eZPATZBSaXqAuKL/cK
izVjmGAO1kftu+TTrwSiUG7jvD5owsL14Tk9wLumXiVtMh507DBIWvi8SYXVgA9k
9a7wNOHxNqC0bfoUC2JkYTeqUv41zuKn5Z0MsneEnRGKb15g29tkokD3rR8w6cTn
RNaxywgyYyJAG0X/Jku8uSHNMQo8A6F4VNS9QO0Jes4gAOe6lmc2HswOW1fiohH4
WIDEm13C6kCDAzEb08QgI0rLLmNGDFYszwoW1MxaseCmWPGwSCGIdNcaBueiMIkW
TyoiBmCjHxkXBA4Bgop7ZM2RYqmQ3K+TEkx0Cnr/mvveJ+HLAjU7LpVgybeEuXTC
gAdTnygJjHQSytOV3mvILEWdDExDWqDB1QLpVKxnNwuHHTOnmKqaFNuuybmjLVul
koKlXD9H01p4/C1DQ8SAiuMEdI/MS0NB5CCeky8IbpireIxWPu36kxAw74o9w0J0
ao0CNELhRLw23TTg2CGSyEtAtrlZYm86n+gkLa/3mUGwxNrYfvP08R9a0baE/NIt
StIh2t4WVvDDzE5eaGTBfV/NTqv7wKVf63j4Rk/v4YoPbRr4LL4lg+8gQE6HGg4L
QKYEd/5FHHWV0lppx/U/BePF4mKvoBCYswi/hgwYgH2Oxeg0CdwVQz0iaHWDHrg6
5603MFrhXSVR/B1AlqlEj2j/1zO/9523ol2X46go2yvECjq0mkXlzRMT12dAGkAa
sTZluz5oF/W0Iq0uqtCkjzNI65v0r2mA+huUPCsUJz05uRLe+bp6IuEJJWoBZQoJ
c9afvfIsf2WKYSIb0XnaJn9JV4OOfCmzRp2VFFbxGHfFB5o/xJ0b5iwjwuPhShPZ
9Lw8drkEAawJedhvi2cq7YhGc/76Z/zA6IgpptNZI4g5e/LFgF0fHJqWwF0ugVbM
xZrzLEI9d6D0Pm5Mws3npzb+cflgNlNK5r1ZX0UL32cmaGmnbx4nhdi1avpfZVbP
5OsPny1VFMZqTnQD+NXHDD/i0srez8lzt4mMc58TZPFTtm6Y6D92iQAVlkiuHF5p
r9YOtzX+p3darVehYwXQ8ZxpYIpv2TAgkZlbaEqlb5kvG2rp9ExY+PbBFRWphYer
6mPFbaEPsurtebfAul2AvbOrpOlM1blRBj/HpEZyNzRVfxehA9vw96V+7BcidSpc
wA36lCT5fXM0apVI0DQEEVWlExgF0RydwDwkfaJpE+pI0oUniS0BNNdp2S/icwLv
vmkH2GQrQ3+E1JNy9HYlsPd6n9myDWqPPn+WHJC0DNxrTXD3VKhjd0oJRnLi4vFQ
Oy0W8n6E9WDAvTbraDpCrY/jPVklgPYIglz9ubsIGyzVpI5WC8nSjGU4+cjwBoXl
FcqEA2bnVhqsLv9UKUDRAkPTsPh1YGASQ8GAnBvVrUCpW7WvAgja+symdfuSYgpg
i5u0Wb01uTLED7HsLfv9TIO53U8gUq0BYwtHRAhfehowxC4ZSdrHrRK9RpOoOHlm
v879kxCIXLaR7C7J+enkiotr7iR6f/K5+nBV6PvRj3UiqNEAjw22o1lDhuEFlerY
Cq6EX9Vy1XxHvVRWWpXoV1m78zvVAO20JrU35/QpMfr19X9lXyvhoCoCP6RAl9OO
JJr0VBf0vY4JDAKCq341vFAaFy/w5OOme7ns3AyyPCDYgCKH3oOj8rN9Ht53u5Qz
CJLWZoFBl6chRN3E6K5kCWa66Bskp+q5OopORbSCf4gUAY8UFLz+WwHZ6tauxBMp
h2dzaCmxs5KaGQdLnVkddpdCMB7vEjtJ5xnfCDRCHD+KDmsFWVHJFGV5lFtRZdYn
DtF1gVpYX5igimhlZX/Y/iaFuO6TiX+VUnJ5fDH9rIMmbV+4Re2BTtwxIhODcGgr
GxPFHbmMy5pUF8KxUbJ70z3cWw3fD1dXFKppKadUj7jhLY5njbEcZROVEmmFifjh
zq4T6p0X3Chub4AZEqckrM1hFmPSEcf1h1Ba0TndKu3qy8LmDm9osqct0ECqYCX+
/wceLzD4T2FCZc992Phb5s5vRMA4v0kqL8Lx/2Z0+/KOS3WOU3LJ2PTImEsaMOhE
ac8VDnxiZa2ITXmY5yHYfccvZw89GvBT0o2h0LtkY/BxO/uneDjtaXTCvNRgDPPJ
Ubi6HT2AmsJ5RphMV591llXqaxMhlMiwYd/fIb66EtZEyCUTI3UMcUr5aub4Ed7U
BZZVpgJU8LopIPSH0Q2f/QDAC1GEsRivMJRCaULS8xMdVIfGnrn6RqbOIxKCilJL
d3T+vJ/fWr8KbmwNrv55tUqtoJAoW3dKfX8baaqi88tLwiqDtTdaxIgP+Pyp+s3+
6kUuo4O4FyYsDhnXc8y95wDy0Rnw4yxo6tu29hq2+Y4Xe7rUscFmZtND70Yoeu7A
0AyFSUIOyTn/LPg7EiEKpvDgRedJmKPMwKTsOk0pnb2XPT808oh+gOMc3ztM/q18
d3JasabouygI7mvF9wKznrc+YATYunhfLICpFrwfK4ZzRRo/zfQtghMO4Ff/sANF
cpRH1ZF/WqHpal1JZu+gIPAj+V+FWZCWU88S7/3IKDgxcSQBdwUFx/Dv+u9mKbWE
bgq4AtXfLzke1vU0egC++BPjUfqAacK9EUtfSTSktCprB3O2YikVxZPGAmdrUg+7
i0JQfHBPZFiQsM1+JqMg5iGSYUYV4NgX/+H6K+aaPhNfAfPbmA6Otxgpnyzfysy8
S8vJR5vUF+HUZHJetsN44hNMJvEBPNP5PGptj0YVpkHbYW6/BAUIp0Pi8wI2BT/B
Gwp0NoTVVge+nKnAgaZIE9SZ7iucDMeW+LlgN7i2n6W8YZ50dXvMkiqgiMzxBgqs
y4gvSvDLMxUzjPoLZEQXeY8K732sochk9zDzQ+wJhCwLXbzpoYiTteOTpec/2Qzj
IYBWE7j8z7efgALwsxibHIFX2afiAKh/cJ+oiKeTRXRY7a7aiduslAiQkbOT4apv
dLkT0yA2GO53uuAGChFh8ZwSO1NWIxgLxQKr59JYoELsD7vstpCBZ0aJiK/lGdUf
sW5g0CJz1GMV68aVHczRQnlvAjmBtlMbCu58+gvz4Dt20mj5+v0B4yebj4610Nix
nOp2HAC3jPOIvuBovFX7HjC2OEyFPc2zr4m1v/NtprpOZN/foRzxBJ+9FXOCSukG
yn6dLL9xqhfVtjX8w+YGIjZQt3RTtQs+ZJlXOC1P/2ETDCVmm73IJagHpEVmGEFJ
276jwDnpIitlVVJ9VhBgu7ZKPno/ibGgZ4DbifYYpTwAFa4875+kSkqkb6Gb5OSc
wUxS3G3No+6i0hHesy0M5GeAJrDuC4OJ3ayrnrdX1ilgGg6epil7vDL2dsbgEBOZ
joMAoOvheeJLuuptdbdTxKYYpYIQgy/IhtL4h1XHrNLASsULEZDvFp7pczDpoiln
frox/m1rMogItyrwNam4yqrbgoONjxoh/2jUWZQZdv1BptLLyDbjxguo+Z+gAb7Z
aqAg2RbLJJvIXlc1sq0ecarQSw0/G941l0/hxvcXCNJbi8cGvaJY8jm25ieCgtZx
DRM8wJTavSmTAegNlN8diILqT2t6UYXQTlXGZZSS4LrhgB9Nv4M7XfgIQFT5Cq8p
KLZ2D1wUQdKC2EEk6Ne5cU0oARA0TxqOavzu0luiQsri2x4zTqcNov4EfkUcMGBC
0BtOAbiemxRlU+/YbIP47ByVKmycnZAsj6LCKiES+fYkt5CCBmeOYCLf0bmlcRYs
vsZ+4mrRJHdo21sBjkCYPjeFOe/w/yw6tRiCXEJ5iy8xylJjkzYnT97DML2jdDOY
ooxVbu7fynE0VvQxN8kP/8h2SaALh2YCVRyjo507YP6N26aHiM4pxtg138mi91Ix
97qlh1c142b7hQ80J8ItULHopT4dpVCenkKKmgO/1UUh1oX8AsMff3kzEN1Hs3Dx
2Wj0RFPKbqaTGuS9NifvOjNS/aPsxgrqxjvgcWWaL/tZPBM1dYl0oAQqjSci3Hqm
BFrb415dusU5VmyV0qrnLUtbz+tzmw4MV2ehzQAOaF0nFJSrdQBUuDgc9tgTreYT
KPQpTkJ6mwcrkPiksIEeR9ryoNRGlUvWzs/9HbmgN1Si2fyHEpj/nOO6Y5+l8wGb
nLQ90rXPEm5odkKWMYAjdSB5XQJ3DxXZ5x9TKJ11zM7OPujfe3YN3k7VCQ8oGkdb
FwqRL328H8xGrGNvXVlvWmo3rGv+jPQwM07aCvrRtoJbpPzOR6MSwGTaAk+xeGru
p90XMTIiiwGUt/pfoG0j+naE0TBiZ+r4nyVsNXk+f3SGfzqrZOhsq4QnFJQ4er9j
ag4RTUTdfZ7Fj1g7nuGbkPrMogBvV6tVMR3UHf3c0Y55yyk2AZuf4xd0VY0raRd3
Nv4u7+Q4bi7+6s2V2MnkZRAVzSqKBo1MngT2ftIM9bHHZhcgfV1ySLUTLuMN4BdE
Tqj+s0XNr8OIrDi+gIrW/NZWbfFp6kw88k+kK591OZyK8ojgABQoam0bjkl45UAi
J5vsCSFfbu+YjHvq4NUVEAT/FemvXGMsLCxdUju9vGG6Vr2dhgyaM8GdOaVmJ/EW
7ovdei3aCxWyN2NSehva61/ni8wqlwluShjzEg8iyvUPMQzi5wvJDv3DgpC8SPQD
49qcBHpQGV/1HNxID3oNms7Glsjd04h/OSw8H0tvHN4Z2bMR6ZMl2NGRM9r4RUa8
Xx8wSBynm3HGw00Wlr9wajbNtEaTAbraZEHk3EgAGKzlT7+gaL9LyDtM3qzXGZXZ
UuJgt+8idImDp3ue9wL7w29YpPctM/fLjFQBlw1TSosey7Pko1UJRCdK8lOjL+Cu
4GnxVyzVF6CmFH8eF4wuBVXicogbIg77W4QzskCo+4+FlC/T3cp8QPn861GXlBNq
3043FFfQ+3bFlyEgHn9P5K5rCBodQ0LIIaPax04OUNblOOv8suiF+8G2kyzrO1qH
33+96pceccpVRd1z0nZ/vHGpxccxxMo4kTbicRLcQDIeVzT5hW22kEPzIBHOaW2E
Q8+BwJSPzkfjwYwUKicGNW1b15eldXIFsfJyL8xqKFC+8PZnezzPf69hGiTgk0T2
9FvmYP6k22GeNud8BH5DNUWdeV1PadHGcPoVzsA7rKBsXOOHdEXVuZWxFjsJKGh+
zY/1luw8xbx9iUEghU+xgqgvAWg8aZDeaSN5vCMU782uL22qTye3yudrrQLWftFE
AkYtRHOaHyHtwlvoa9GNuAW66FD0bjihIx1CGh2HM/SASEPhHU92FAKZtAY3CrZK
uMKyoJgKQSGdMRE1so7pS9K9shHqi2ph8vD4KdNJW+o73aQZgvf37nYN94kN764W
daKH7tpD7yw2UYr742PJnQ/6E6WDnQJ0kFcCfONXQjO41XkvQdQrI8HollqLmbNN
1agNwc1DoLsVy+b8bXYQ6mHGStt29r96QoBED9/CZBd8EWtpYiNtAs1frzrqRoji
DPt5KQQ3yhO5GXVu+BjXxjzLWZZPBXCt7aeG0wK3cmx1RxpDFqObyxxtEqdi3j5e
oGlPSUlmf/+3c/IEKoFMopHiv7qmCyVCBRrOjRUZdvyKpA9ImCm2bGO/LRp58Cmi
SkXF1SAvVCzjvgi75j4mWNl3hiltNLhdj9FCy2DLnsM7+NNw9JKK9OUfSI5kQwDi
y0xRBGTk2STt35aFuycKjmR8DhkPwSgoViZMg0gbzoIVu7MMxypWTKPBt00C11/x
rgNE1kwLwo5hZ7jjoDtx601ziR0L+UrdziDGhDvrBxseoqcDPOF0EBfUWvD+X1f7
CyH7W++0He/6zk0HItjMhxIW+uGC+jWK6FZ0MTCucaG5Bz9NIwz48NHHiymcGEKe
VAak7FlB2kXNWEuTsGjR1Scp6/4uLmI2VHadil7DO9eDRre1CZQhregrdy3kFSjQ
L5lqcnYJk2DBTsf4Fz8zdV9E0VEe+AvebPAtyXLaYqXAwy0ExjbyHh1ZAEt2xEJX
REoQzdZeXSGYo2KzzDNZNcIHKOcN43lR3V0y68DRNQW2JNIXYDkeABzK/md6Dox5
uxgV1ZaIo3QSyU7EDXW6eeE+Q47JtNS6p2QJoclfOIqbWTPIt2IGIDcroUB6CDxd
QwBi7ux1PjflFPs106XWTm2vsNcbfR2f/1y2qplvadb9+6EtmSxx7bF/WxQppkuc
prAVxBvMBkjsLfo7fYgG90WTGGoweFLPVKeWDqqayDKAXi+qxtEikWlUT1PRH/Uy
dwOOoBu3deKMO2WsxfhHGYxKu5rlHxF87bCTWkC5JYeIHEkQeFijQoqOoUlV5W8l
vHLczTh/b3dmHFDX6rZ4PRFE2Ps7+2rIIhtftrNRLxRXHtqbFW2zBLU0uRHoWC+P
8xBQVual+jQNwaulXiF9NBqMgQfsd2fZ0uwovagKCKa+ELfmdHjrS+tHDc/MAz8f
xCsxzpGS72DhNnvtRS2dmF9nk/uf0wjQ5VLew13bYAM8nnfkiT9BtG/1B9IZuPRf
5I1D3Q3rmU6X47QT/eSJRevdA/inc8edgiKVFBjHoD5dJ5uYIFSSAFZS2mOfNN5j
vhe45E20U4aPylIFHDYLDVkg2bcJdkBDipMgpq+NOlDai3xT+TqD3QRfQ0fv6kAy
coNftHf9c61BBUJ29UWhUKHe/k1MaD+RSZrouEkHPjXK46L9xgD+JStDurMk8G6F
Y+zE5OWPyjYjebO71o2mQTUHI81zwkw2QXc9ay+UrR9wrAk3ujePcW0pho0gJuH8
rrg/MSNkAczC4tQP/M9llGQseM3OsYC5O7kB4BlkKWkCWdzQMow7EA//H+rdzCxZ
P05LjPTM2qDKVpsNefBf/nPoyok1sARGxGLnMcOIMQaG+T93tc4uFZ8qRgHFf9/g
wNHf/8nkKBQWmqbg5jQSuNuqkj6PIsNHPft+qLqeG3QzU3PqwNW+GuqZIgFz9noz
3F1rYOOS9llqT3Gxi9uWIEvozOdwnBKwIf/1nJHOZoZJ2fbNF9PAq86OTlCPKqcU
HBjy9TqzZkVnN1lHDGUc3tsA/bthb1hnEbM2E+5wN7Wnaq/QZNf9h9hy2/ZwTw27
PvYtVyX15kHwyKCMNj8pxIUyfaDTp4CUJXVKWr7fJKc2s1XaWJuuNDgeHvy7U/om
X1Bwd1T0LT3GxX40dz5PIkjGYJKfL8zOw3dwSlKmssflIkeB8eRZJqdcCM3QuKpO
4JYWNNXarkik7qeYdeBSuopOJx5G9mmoD6jjDxGmWAHdsCaLMLFIm9PIOjbpJTn3
XCKdlUIkx5pYOy60sbYET/DrTohwofcdmDV/GFjKxTZuaOWpdDV0Czq3iyQTiHEk
YlrwD6lc2CarE/HUGl+qVzW/qg4Zn0sjtkHZWELhEMSoo69vRA82CVu17A4y0s4v
sLoptwAuL0YYUT7otGSoOCxHeLf6H2btROrrauJ/FqvAc7+WwqClnSE2gHZurebW
wXeUGsPEmjMra+ZQg1H+qQxcXcQLKBggYuZCeAzugDOOeKCJLvSkHX/fhR7zSIbU
8dE8qtdXlTWqUiLgld4pWMn0EPSkL6XFHYOuJzbaHXfYjIfA+B8XPDqf5i6hUZOR
Px+gG52Z201gubFN7OeW0ZyXff5aHS7kHK3CaGi/f/AWUaTHdPlfrj4s/pzyq/Na
kDs0n1q9aK0yKioQLpKHOuL8G34bnVAnVTjR6QWp7Z6BzncyTi/LHC6W3yFi8BEk
CavxiKDWmLsHaGX9vrNHejXtLP44Y01hzq4zHtg5VFGYR9+p2YDcwLQT8b6zrBVm
PIeRHJm5CUcHjSZZlLZmZ+fF91eZHGpfDzmccJihAGrZS2/UVS+fD7+jLQW6UAV8
Kd5abCDsBTypafjbPjQ0ufmBZzcad0vbYmY0ZbB35FtdJBEi7HBl057ktMMN4U/r
kVC7BvXB8BIj+pIlng0ELjXDchdeXqkabqglDYGq9ZDqijxxhgW7KaHLEkIX6/qi
F8cKXd+4XIDj0HEr14EK7bGOVzqCRsd3aeKv78XQ0LM2q2JA2C+/tW23kiVJFGLv
YDGWZspfafzoiBsxY8u26p4qTz4gPeoE/bkqwtFJJ1hmSye7nJod+AoIvufmsRML
vyLGAkM5gAj9ZUdSJ143RNkqkblpLfI83yPUrrPmh+U6U65DrptiOQ29iWRpN4Wi
TlNjEXAYajJyJ6uzFZ8bCRwHH5hfxIT0f7N00cdDjsHACFNWEmm5Ge9NGyo+kuxM
Hl3ij5745bnGEZh0LHxUgbs2KRm8ZlHyzV+gFaloTS/2KQuAoIZ0r1yMLrwjZwzt
Z6euC0gp89M/KUHXMXSp6z+hrHrA2CnGe9+1e+Zn4moQouJCvGpNjcMvKutEwncD
jS0/Qvlui7lHx13eZvMxsB/FdPu3l3CQV0vb5DXmaZWA9CEG7Vy/7bO2TYFFTcTd
WB+5xLvImpXlF04Lr5S/H4yGK4sdkaM9QGprAFft+/nfWYRQRYKZN9o1bOb/MOtz
ZfRFBWKKGOb4UxlRqwhJTVKejWT2o494CoXuvL+DLe6omZ1Jfv32QzLEQSlmFZN9
q6sh7xC0lfNV4JW+NTtWNZHN/M2gqJ/P2AZDmgt+EHK6TcVL4ua8ugI0hnJ1ZvL+
LFDukZYxqrBGQrGdcld0Y6Ebb94IrlLbEZ/gSyFztkWp6kK46CPkyjl37dcyHIW6
HGuXLGp3QOC974/h1yw9oIbfDnYH2fUnY+Y2K4cQpvA5ocGomIUfKchTa0XObuCD
7+KqmqQxXtw8sC73kc3e1KZmFjpq/z+CmHXfNtt+SBaTfeUnvIwP0HC6f4XYbs1d
5/9FlAA9/0F5Af/VPyP/Pp4UogWdowPEPpzI3ERX71EBiOFZ4KiVQmD7Ld6U7/eH
8+JTMW2EdwT/6ArG6YCaTOdZavBA27h0coe9rG2vX5nxHCD+BQ17n/1auFC6UYTE
xEKHPQrjbJ4MH/TSOKSk8WqMApSk2W54YOXvxCcyE2wwiHgGJg1gAKfB9rPqY6GS
wiJkx5vqIpr3QIRin0lHN3Of99VrMyP3BSzyvwBKEfFgSMCGF+S1Nxk6czLRcXK6
LhsnL7dQW6gHVWy2o4HjPy0aVsFZTu9map7CtCbN/zswrUkIe1lN8sH42CoVwPCR
ZngScVRLgWaL0W1Yv+6gSEAmPBMLQWI/AhANNPEuIFC6Znet4CVoBguXwokH2aMm
H+KaMcns3WojvKp+L60ph50iX4vEjdud+cEKpZfyUcXj0XCAk6yX0IyN9c+W8X6+
T2zQb01gXcOPyH8P3wZ0XsdgzfglL0qq4rUUTYl8JZkiGYFlSsxEBz3GMaWwjppD
/ixMlwdVwmgVapKuCfKQHQTrpDo6ISJNQMiszWCP0+wVZIOJ0mBDZFtBwJFcw1Oq
NAEmPUXBRLATL4qdmfgYdUAz+T/elofdYhGwyzDzEIKOGd9ykHz0tfbEiEQAmzy0
2rWjDLr78Ri14mH/vAowelTA+D1SJQ06hfaP3wuQkItl1uuafANic5NsQl3Ewwpa
oGeBdiwAb3ergRSVY/6LAisFMkcYBYIIUkB5PACCRxJWgUjSnZSrTp8jzPDdz8cs
MjcRQ75o3WbOFNnoxBBJGpmn+FuWZSNsvwQl5qq0CrQ0nAG1H8LTM5nu1HbkO4sp
Pg2adbZzH/4CNS8DaGTfIisB3ivhC+pFwPXHoAfsA/zA+mD7l8Y4FIn9TSUvGqWU
vxsj0aWHghlkULFeyrV6cc3KFGmKoc0C17zhdK9MkZTZXf6DgfFlrLVJcbouoyDA
LD44dA8mBTeqoR8XlCheHDI/aVQU6kaOVr9glbqMhoISDVl233SojAdD7Y5dasgi
2T5LyZENhPGIGop27+34G4kVmeiafK9tto2o1d/Bmhz8A2+M1X7j4Z7IvlNl+92B
lYDuTxBoTBLoQRkaupRTtDFW25MDazXng97sbbf1TbH2dIm1a9ARTgs4fUvsLwHj
HrIeq4Q3lpEG/k+4yz0odgucDuiGey4cjrCEedKDksfxlTUda2NVQK746/PT8shW
5m3u5+mAxx3wqUAtF9Y9NDwa5s3ZclW0cjXHBgBn9Nm4WHSGhweP9YVe4cAZDNlq
liRvKruNoiw/2ewEknAOaGI8XojFB0FZgmey+xtll0u0aS+MXPtTySw7tlsOOkXt
MMTLUQkz/VE8XzTBKuDI/tdGsMZiCJz+J/bW92DcPHjJy8xrBTzbQSPaXoOh9bMX
VvnxMKI5myKVRri0XUqoWTSI8/a6Zgqg9r+7w7tTkVU1SIQdbio96xY2XBzYqnh/
E99suwcsBsJ8Bopkoou6VPAxFk45rKSBtneX3txsA0n0B64x7UR4Zd78Ap3NzIm+
gYVxhx3ToxC5BacWPwlsK5uv+APKyVuZSajkTostPGJTkXGzwlghxJvVEpttHeWu
CvxUjq6wQjG21aVze0fPhuWVKU6NQxMpHcEmciS/90BOk2w3pTqKGwxwkyb+aspR
Ae+5Iv248Xa/60zIT6Qq23pWpogr31FTzNw3f1uOGEi/wdoj/22+0gEw09zZzBZK
NZd4kZBp+Sm+yI1z6gs2R7xFjX40vZ1hMnugtBtkIZ+DnhgKEdmKFySM3FsqBxlg
ZZwLE+mAigx2FNWisdxboUGXJbqOHPuf0Mqme/2bucFpTy/RXVTm/BJtgNsHIWx9
vz+ocm/AO4UwNYPE3yttIYrQpLmYe3JAMyiZ2lHHmszay7h5VcmiTmu7PIdUrlj8
D1XNntGo9dC2FTaYYnXWxkCrWDVXynHtOARoccap13UeZ1kBuIHLUqaaEtkX4rGV
ktk/BnxbHHxnq04O0MiisMSgfji2e/SjkvfM6z2bso4hh8wf0NMXFbNw7uZrHMzY
RDYI3P0lJEfO9FIYBUY+xNFU6fS96e5F/6m00iCfoxNJPs0Ti/Gj0O+8KysqEsjA
ib2FdsL6bowmgJKy3NW8H/eBL2kljM9Ac4fjtl6iq1HyXNQ3SiIzKNlCNJQ6wCbh
oOFBNMbEOX/96FxQ/mky8F8akNp/PCqTvqrkRzgtp9O5Xg/tKUFD0V5y7Q/Jm03B
LrXsNRZHfLEekQC+pQQ4gp+tVg7S1ImC7gHhXxVQXSeJVrIEU/vBzBBSTj4LP4Ob
zXMtYc6Iw4CyHm5fbdHXFfe8/mwrE0MH7M+DqMrFGPgZXxYusaYFg9YKvXOlvlqk
mXiVHgeZE8SU2s+yY2mrhgZBo8VobEEz4mL68QuHU6LB5eU86upja62uPivgg0/b
jV/5EqBPxlieTfMECqJJy+YTD1xkI1Scn5FSW4x395pq23gHdWM5Cxfm+e6RJSf7
S9ylNdyqLMnjJslNFcKatOkXpTebd1VzrukJ6NehMMIyzfCBJVXGC4ZNrc6oTHGG
4s79V3wsGUXD9uQ0wyrUTCddlhmxHz5/AxydocEfuH2fw/Lnmo1Jl3q9A8mL71NL
bN4XmqVtvXe76iOdBbfKUEmy0TKx1/YzfwzfjDpoYd/d83BtlTj7q9uHJCsH4lU4
WVRhpN7XqONeF+7jecTM+KzzxjmefR6YsmBOwSP9pAFBEVS1mnNP7MHHe8VD8XWc
RNBhTsRYimF8WSl2Wg15MaUCXT37FqRjUdcSkpY4b308eVOtBX4FiKTSEV9Lq0Vn
g8/kH8ZDUbjjotLmLqIeinwCctDdAMNn90MIReQ7Pmg05sthyLF3vNaIZlTgiQZI
8+yl//X5knp6eq37ARJ0oDEIP4MPzEgTPKfdgMqx0ngeKAE3lO08AzbSKw5YgJoD
25Y9+QcR5hJNo925lf9CYryixKdLLF70/zpyEiiDaNNr5iiEwiQ+f4zh75COAJMy
Hgno2YDQClvaHpcZGP8f9iY5N9Vq8UCmBbQMUsWCfNZQdeUJcukZdCauJSeL5Jdp
Kvqa+/CQSOpzOKMcPOmROoTNtztZJvHPTP8Q/pz7wN3ncUjB9e1HaJ5d2pGNg0yE
dQRGQFtrWdf4xVCbPzalLa9SgoCxHjx6jGmbVJTQyAnqf2yVEfHJWHKoG091W0oC
mcvqaG+Nn6rWO1B3ARvBHsOoy72LUq0QaJhKPlO2rjzk6ZICypceAW5O8lOam7IU
nVTn0G4livSLzV3hd1pbCviokHCkoQBeuxZGqYVCPkDu/fXm7fDfYVqGeR+VT2Xb
HaClfDjll6CFzRecBPSqVQxCBkxAxsdd3zrhT1h1aLRE9f87gKnjQIuA+hVfORJK
xapkDNCLINi+g2NZyJDN+11FHxOM7sGllLcL2Zrx1wGcjHceV3/mV1AWDvjJHVHT
aWQzUiUldAhv/BGJXJM8Vp4gnEAknSYKzzvB6x2nGF5YQceAXDkghuS/DLJKVyOJ
+K79ZGwkX3bT1545/UQ8HKaiK3G1Y+zmb13nNuVxKzvmdtryScg8f7K6KPKqLObU
jWe+eAbygri//bJnewEHJKwLCRGuqR2CQJWL11BHzoqmB8yVv8P+v+Te5E+bM1YD
lJIvc40KZswccYnwNTy6KVcBlcn4Zza5vadPwFHFwunHeCmJDiOgaZTwxkPEjUbc
Aq3QiT5PTFSk7cgaJpnIH/jOK1EdsFBjTCT2tMcySKzY5rl+fl5K4U7cPDvmmK9T
n9BcyMl33aa4b/rLN2tirFQuj4m7yxzPjcTom2ogu6TO/l2ivKVn9zNDSDAn17YZ
24x3kXUO1HVKyTVNYTYMgahJ+UX364BoikQ5njs0AwugZd3kEfkwnmQaK17MAUiZ
YfvWlmC1TqTDrHzbe2g4uWomtOlM4JK7jeZxs76fmF3eKCyMCKzgzebDE4eVTOR+
flkhpOt8t86GhIL48+ndKpijlsy2yOORybizeIqJjgrACos6U2F0bsYOwud3/nkd
rCxm0HPMcNGI1bZYkizbXi7YGndW15E09nCrl1LzEasVS9Jves87uNBBMhF5LU1y
dM7EtxcpUtRs+fAtrxNufVpyhqqOcdEmT28Gdq5DfaORjzsaB1AhSdn9vVuWrOSm
yQHI+C5Iq6rZkhuH6FHRyxs02C+gULGLgW6n4J9d8QiBIrO78jS4/CNSgCZSLhjZ
oY2LSWAJD58gWm/CqK2l+PF0ZLugR9GMUj39JoKFbyEbJ7eUX0Q/uuDuvWe6gb4h
F9R8MxXl6wFMtoR0kdgdOOSfzgC6GyDDTu+yI5PsPBG4Go1/cAo5ySQouPQdHFit
LM8UASEFhg2slCiutjNbPeY4FDdEr3LC8w6iQ7Ugvev9Sn8rrFqVYYu5lJM4IGJB
13M7XZOPVA6GfnTnV6MgzzCvP0QvUAqOJlH2DFo3WH85XsDkT4/iBUCgjrICqBko
4iX619sazWslkeucaeoE5WLMbZMTczxrnRXGsZPhL3T5t+uyPChYgMQ+6tjNqkYH
lvA6WqF/x2kX1MkJppuc3+/Xzk1dcLSKsFszow+cw7uWRvtVXXWgNYx6EzbIeXlf
CoOoy9YUbOncgFse1AUXlWMZSj9z+9T1LgSK5pDsdhRUcfZyMmtPxYpBMeTivOiQ
k5anxlnn0403N0LAf8I5I33gPSLE8ZmaAi/M+j39wdet25SrTVB8pBKhouWfm7Oy
EPIdalIc6ySDqQ7d0uqEe2ZdYgzjMusNtbx8xK2LOorj7lmkO60QQWzXFL1WPdcF
W2Lrj4nVCWD6AnSp44kX/cGlfp461Q8Ez11y+PQQVuN2vS85nrDOkp0e9KbN7x89
r6H2mqqf9jhWuvwfvRQ/Ggp2YBHOOS1TbBzBbmjmGpez8sObL9d/lcPAFXGT8Ya7
MVnfuDJfSe7IrfTCrnZ6bCN2BxHJePfH8hxKyY+y9m6fxLYJfCmdTUHfY75P2Nls
S7wMmIvQPirTY0Z+Tmm1LWckSukWzzSp4zmvvov9gt2ic4al7jhvPmwZskeqeIPr
Pp/E77WWyS24i+9SQPQIq6RVRv6tdiDFfwouJG/5XbWkW6iyOXUDy0bR00IexvXx
5iC8tdgKt7oUhvzDcmfALtnwNen11dpELHoDfRN63gfGGpaKtXwuL6yLtACFDrjH
oHIyARTIXNErSwQcJHeCTe7orNAxOEbEgHoI7G32p1wtH+YS10eIIeYCdRf20VUp
w8UCz74QBnMRAON6sf5Yv4QlLrQ4aoEYt/B2seynToyo71+FtJQ6RTBf5sYpp7Op
01GDrR5tsJRs/pCR6SRToS6WF6AkOJ4M4VIfbCP8DW/f4Gq+QQc0OrCmrByoSzkS
0WEXmZjlxMP2041ozwdW41AL4lCa1VGKQtBo3pvgAZq/v8RLLwHikISwybzm9ZX6
OqKKTztL1L9i+nfjMAlGAqx75sqdIN4VhJJLohG5PL+j1+dpCb2u8/2jrKETm64a
w7FCiPfp/MP20/9ssHMKCAYKfd9AnkMuv0/E+0CRcR2UnXnZrFCbysjYE9ke2KqZ
6/mIF9uH8MeZLEydvIPXgJF7EgKDbiuXOXzQPd827f3Ni+O86e7jhcKEYIQ1vvPK
D9yQ3bBpgloAuuyp52Rx7xIEtFNFE+e/3PQCFiAoVS6fTHgLI1kT+7NhCZxI/crx
Ht5gM7h1+87NzraD/gx7F4LMANTPMZYAnwDgfmPV22kywVN5Uu8b9KsxlPu4JFV1
vpFEm8nowo4t0avWLCH+l1ucVUqTDPns/+Ldf67DqrEgvGGT44foLKHwK7RLSG8u
U19VBrBOF0fxuKOHo+8VZ69tLw4HzaWcJgNPvZUjBYZmTd9apv+gvg6x22ILuQJg
ZZsofkBY4xDOGYArGe11VpByZigWZqnKpSbRMHwIreSzbdXAxZAZol2yeGIyiB5l
YsYH99gBwEswJALDI57Tx3PNt+kePrlPlPhNs5swVGDtFqB59T973v3Q93nxsCJh
aIxWFQp33PU6rV5PHN21fPaoY/j2JqxoExHvLVztVYLClt7DSoe+dLUWlpCH/8Lo
5o6Zq52kTnxKsAUbkrmuIoC6mFLX1MNeGkGdoUV9RcVuKLipUnMFQ7gdTsrSFK8N
MnnNRBsG+EUVmn5T6RtyvMVYAjNr+tfS64pLaRFSQJV96oQDbDXrOO3Ssgne1bTJ
E4bILNJQ7rKMYMHhbwcd/apa8PFJ2B9rjnpJL2VPJGWYeLU//TumQq0Aen1jUOQW
sbd0B7IqL2WrtF7FrUUOmZXY346deVCs1U9SNhEis91KC0K7zeFRU1jfphUkzoZl
FmjbsAG1Y94SAznfrrZiOl/SrCPvOM04A/kgOvuivnLqNKN8hjmvJIikIlKYDDM0
lbBu/DFkCSV9BXKTMoYoG16970lkeL9F4yC5ZaBWW/IjUSJxD+7rh2/IqX49o/Hb
fcg1ylXVtq8xoHh0Dr7t8kS7l9T+QPSLKoN5os6CSObh2DjJXNKaGLS1Md6YS3JI
JRyXIqfSf6G+Ky1DTAyzbCUkmg6bbOw6E7W5Py5cq/FpdKCBhb8qUismIl/VBhxy
3RlJ5pwSmIaf7Ah4Xnkf72RvEROaEQIrGtNH2iVCLPNsZoMDui4qBNdGNgpNnPC8
dmPgquDp9iSmivCFIR5I862hPr9+wyRPAH+yHS6BIG79S/fjqdr7+bFxIlW4wmSz
wVouOeP0KPH+AuRjcfmXWg1e96zhk2oDRf4x3LQG3/QXcm+5iD1IBY7RF1tslG4b
EG3W7dFKtKAIM9lvzW11MYPi3rKxdV0ZX0x9Qdal2o8c7vnCSqIyOq6YVMLQ7b/T
MaBBGQYWsCqwfKuGMicnSapIgKPqzYxlHJRtzq4+4xmxjdCOPb419OzmPOunwpOb
o5hg8N20M2YakRwO1RIen9N/6qGIN/Jb1Cj6ESc8GxrehPzc/e0wzXkOUcqGjtBP
cTS173OeGET641yKArXoffAsqoLk1psQuJWbSrkXxM3IGPHPpEmW9RVDeWUWvm1e
eGwkojgnD3Q2v0dCcWVpixO0ElWBNxcbh0mUo+CNOg+wVuTi5r/uSx1bbiUmUY8Y
kYZPgpMjGaFfU/1vlabpgqbQhRODbhyW7XpXYDL0+m2jkpWlz4A5QFxFKR/OwT/P
6KLw/LoTFyc5LGtBfwMMV/vVLqErXRq/gf2t/40X8jpNVh+5lzEVYgp+zaYAvts5
iIbDCTv4Nb+jMU3m3dGNxA8WSBnAurKaG9pH4rxpI8fCl43qkoxbYctutLVeDkMa
ZqukdX1a3gRvpJrgbDxJMn1rWOQJKxEIbn5htOpE/gGu1XyqMj6x/1qiDSjdpBUe
U7j/LLmC0Wd1uz+j8R+pa2tbvoNNb1CDny2M0M8UpOL/s1ufd2UME1F5aHkRS+DX
Vlefobh4/vWxoMtyNF80I0vgNzZzLepWLcih+XHbaM+rVvf5SuY9TzkBeFCtJ6rE
kF7Q3zkWrLtZ6cpmcEMW2TtT9nynG/6VL27qtnSOM5SIwEfrbndUNs98h5D3mTQb
FI3bfMwjs9MNIKV2rErqc9EBveENI37roZR1xGZWjmuj7hidnSfy6EMlJDGPtkAr
wTcJ9ASqCE1F/rPLNxwcFXrMRM0Vwin2BRh/lq+jDj9qHyXM+4pGF0Q/PgFKHzi8
AJLArQBRE/ZnaHb2aVnHKG9AlX0WX2Lu7smN3iRO8hTQQEp2+68zjmK8quZnIrW4
qiAsInpfn/sd+fAMzoaFchax5zUIzhDl9HUHuLZ3vmL1Ug3rfQZ6K4N+X683a0uN
iQ5JnaYXzhwjcbHit1NlRax7WbYutMyKvU9iymGs/5J90HEPP1cUAOz1q8Pbm/xu
gMS8cPHCC42iZqX1Eg7pR40hYbGTSyhmqLbzG2NKKCwjMkEYM26xkUmFBe1RrWnc
NKrr6XHMA8UAGhwwQ+Flug+PfExT+mr1+qegET7NYOLSiBLYlb+uaGE3416n+Mcz
PMv3I+M0E9syf8Uaum1oDYppSCopYHuFX32OCdxlmE0sUYoHxWydnaZMzIQsiQ/i
4xCpizQf6Ats1UBFkU5IGRTW+4sbgKe6mhOxxbbtNlBj8uM5xul1d6sYE4QRMzx2
x+KDzJKH1zR9Nwb4PR7nuQhNhTLT88UreSGKVxFN0vQ0YyBgeAPtuPfiTblr4Zr3
WcPK6yDmFj1Tho9PAGXpyOwKBy6WYn7NNOlzQrTdJC8Fxu8fMZN1iKrLNf6vk8Uo
TSvbLkxGNBfvAo2JDkVlBNuSJGfnJNeBdELWKuEn+P+YNBTAtabVeAtJMZJnrHsR
PXzNduXDGw0Hsuub33Fq2BfNjguLzNMs6UHLbmUamUvj1nwHnC9GDPGk2pat/jsu
mXFg4pAMsqyf5EqDFgS8UY7nKj0kVbQ+BdI74bKqmXCL1M47F+gN8WdIJMpvnWQ1
nO55wCvXIERKp2xsux+Qi8cLBUQf8e//MXEcNJ6uIekuTzpPrC/lK47xy9MgLS6l
cfbaKoyQux4aizbzcTfwyVPcC0hvCatoZBMRCa4SHOSmMArptj06X5X0bqSKkUYM
xZlmFdTn581zq9a+kE0FyZH1okZO/e7DZzBlGslyip1bySuid7IpJDLvGB7Z3arp
4zhGnWC9XNBdNzjQTnRZozK7opsvBnq4qpaYodHWBT13a1HVs9MyNn1ayS3n7Dyb
bov7JiYEaaw0Wa/WIrTNA0NP1UcEFj1MY2gnmlXhgeDfSLReABUjBER4oWwg6g0h
c+so4EbpAXWF4OMXGiiNt32Z0eUmBLCIXx3zUdGw2Adjn8t083GvtPiYIXj3xbpx
lN+NDqF7FBKn3/iY4js03y1ITqjJtQj7P3cm+MBCh21ZDEqfFtnyEBldedzVSH8w
T8R13cP+Mcp6xIoPKmpGiziPN0dldBCt+D0NP6+lv1A7t7X3xvQgdw77dBt2lkuc
o4D0OpaqFPtzpJOzMf7cCX0nvbsHt5QRi6YRn/FW0lDQuvi6bx5fsBIDB3n3pGtv
kGujjMmMY9YZp0q+4LyOQVjavxia86YZbKQRCN+DlVpwGs0vEaMcSja1crMFJirx
hj94Ccvtau3s5N0TxIvrcebGW44wRWP5wOfXyCB8rn8Ux/yyVqdC0YzvoT2s6x0b
4+3gcSQMbcG8usw6ooQP/1sjGp41N0fLg1t2sJFS3P6zF+xkdrYzcXUjNYozy45/
yBJzBg/wUcntv3S+V2gKCknCVE+9hsdO9+s94mXdksTD2E0IYjgZzCRzLW/LX6Dj
Y6tpR33TAkZUpC3Y3zYyiZildkBh5ZXBT+zR1g9PuKVwyBMtTPbpqniYdgRSBumK
2tBHi9LDHlmXdJoZecvpnLFyCiep/vkstx0ky0BLtjYSjDqGzFMiEf1/lhKPbirh
1rn+uIHq/vvSfCzkRAwP5bY+qEuN+7nR/8PzGXYf6Pb4AiCxaTlvAPUm7s9Rb368
hueYYuvaCoQKQfnsuYgRkUw9C0BaMOS1q8OCkYIpGGsdd9cp6w/cnITI9od0i+Xx
f/Zt1MY83+rx3ZiZXjx+tVocLw7QJq+JnI+h6A0pBZynpt34SQvXDBI6BpykRTGT
ttU0Sj1tvcZ0swahW2D+8ypL6YtE2r9EOMKqj9PRmBikAaiOFuHOaUPfJxTAaXwM
0t4QNwYLFfFacPf4l7ZdWdjRACUhl7E4tAwuQlA/tlz62frKloKLMA/oPom1NFfZ
1fRNDpJwLCkmOobhtMJWEXnFrNAE5h2g8WA3RB79Pv2oA3G4tUjTZp+fusLa+Dy8
Lsq9I9RP9yTU4v8JTIX6y//0JDo/ws6pCMWzvETbT9w/StLCGXlt2vw75Sakv9Yi
Q3Xq+7EomJ/e9ojcJPEgUhxcNpQaZaFC0IYoGqeBIe+2DKQ2JNO5v7YVFHX7o71t
CfczVY61whpBfedaca61ib+6mCzCzf0cNlznUWZpcjlwVgL5evAFFMT0Ud5fKcEh
QoJQwbDOmBb4Rg+EZg0N0LrRGNjiwrzLywjYG3UZRQjX6rLaIrITOeXPIwWlJcXB
ZgYSZ2AeLT6YVqCerkV4/mr9/mmTEP3oeGiSIek7+i2sF8CdddZ8McMvuatdQXrm
70rbM1ZvzNS7Y0UTnk22MmC2an0F8lgcz775DBMXncMXoskbIYJl6uqf+sx4NGns
tz7m2NRUiMDVLl7uajRFUILvEPtFrm09yDNacO11VX86ga8Fjh+wVF+U4541szO3
WqcbwkmoqMyxKSsMCuAob/xzfzFuO6JYlfwZ2Gwqit/wmTKXA7upnVw2G8RqnpRs
eUw5LgOZ17K4+O9XyfA2xkn/vGwz04qVhCQpDheYNJpRD+jQXSwxo/VAMWctyAF4
jomzRY8o95kMoC1i1wFA8uqcM9308NcAaVXM1RkBqnyhVH7Euud1xKXD0fuxJoW6
ZsG8i1hjIpnVuSi2W0sjaaeSFb72dnUP2MBmDOWnyU7cBEavVEHZhvMEskolupML
X+tOTj57xMiCQvvPNy2oPQn+hTLRc1x23RSg1R+ikdiMLkOakxzHycderkz62Lz/
ngGISJ7Lo6ZXe84K1X587TOo3p+/NVWzxaylfCgkR6YOoWcAdfHfQmtpW1xvm7ri
kx0UA90rpIm+h86cHbf99b0No4Zz80att5A10xr2WtdkDlwizdzyNfrLwkMT4Nk9
DWP/nDwU6zlHVorsb0HrNmAsY4ha691skLw7jjM4CI4++M3x1TDAtVFVpo7GMAHj
tDmMrTs0aANpctlxfsyXKXAIMP5+3P3/xcvIhrhcvh5q8NXaDwlY5ODu1UtUEx3a
tlsRxkitLhMl6mNm+NETsoTJoSUeNIrP+2XxzFF1nkk+aiWVWtGy1CzKw8QDLpHy
0hb9zV3pltiLpqe9Tavck/EnbtG2SqdosbOKp9sJVRRljvPbtQHntxKH866VPNtw
7zEsqvTSU5VCJxiRjwvf8O7DgQazLIfNCtCRVZyKwsjia+Nj6sTrWFJk7kSBQdPQ
W/k783dgaECzMaIzDyWJotwmsQCrG9KD9eSz7DTSQOHTATKteyzITpHwx/MrWoLA
M23pFgPMz1jTr4ny1Bx44CMkUtZGzID9Eg5HqXGpk5obdI49Fs+oYQL2JEy4lua9
fiE+RhrLUQJNpGy396RP0zoTmlrY0AhSG0Wg6njcqZj9d9jKa7ZEW3w4zp2zaFEQ
O9reeQ0GbTTBECpwfHm3vdGqnhO0MK2tMoNMKBsoaHJ0ZvZIrPKbC0TPDUe0viK/
tOx34BnOgbLwM6OkPSbQnikP2peVCRcWQraP+VoGAG5iRqpPL4cZdV8PlwmRaMZ8
DkpMn7MrRCksobwoGhVHKQVU180LFuq+Sefra1p3Vpg38WoyUNjoThMJB1IwpBBI
D/44Zs2VUhXHitGYsvbL40HHNQ5c//dU3J7KtoOjMVDvUoDBhhQrPPZWrLIpft+6
ApmnibuMQg5uzpgfLWydYRlfXuWMPVRC74hA48hyGTOPeZZZ0jRe9+AO42k2LFWn
QN1ssrHVB6G862ExxMpn10WpSRWr+FII4TgwVI0QmibF3UKjdhmACirMUWHfJZ84
2hii1MELbkCIMMtAxmN5ir4VwYGQcDOc9imUSUhiKK3ZjIWD0Yktsj0OrXntKb/6
fY/+S70LuI8O+Djch2HwR3ywT0suZktFC26RFpRH2C7XyxyOuJ6v1JpodWxYpmkh
CVADbmRuKDcF8H2KlJvE9VkNZsDE5/zxNYRE7ROjbzaMArnOp0OYm6Fyc5HVtOVV
1YW4SZYfiWRqqMLgMiCJIZ4PvGbF0Z8Q7MkywRvSaE8AAJ1Jof0yPx/M4+1G1XAX
6EV3FHwAF9Ns8i6prueI64FPD1+KZgmNpoc//fRsLHGGTvH3MqUM/0DrHiTEeO1y
MEX6kH+YF48IwoIMrKxP8XsCNlvBqQpH2a7+NbXq4FdjuzmR0wc7Hpm5+Ug22p1s
//FqG4n+2UXX6zR4ss1K3QhCajEyEQon1StcsozSl2x9wmB+QJoqXi9Go0XEb7rz
NbLBIf7+QjpowtF2sVfF2L+WM/mOeFnNYuGo10aI1dhQy51F15Hf6TZvvdhS7UAD
2u+Xi5sYRx+cjWHGAMplKZgFOtN6+BgvEF1WaAxecVEReYgFzs5kkKxUC/b/Ib2T
ceNOMjT96w502tmpkNgeKfll/6EaRuCOcFYzzEntM+RtZVPtaZOkd1cLxp5tpr5c
oDhZRwO2Jt9WLIiyN/qw37Y5Vtb/yIZIJc01u5pQjR3xpkCb4xCsv+o37H8nGA80
DKQAexPumfq6vsezLQiSXxUWWCDNA8minwLZU4XWu5UK1PS5C+BDw8Fz40dgv2ni
UCdb5z4Fba+imolDkLy46kNp4ZdcqJWTOr8tdjEdg4XzQfxOSOFvi0UbWYUhC/wy
bOFhaR1w8TrAzB+X+q2PBv4SxN7hdlDIHZccI08eUufedPSnyiywXsPODzDU1uOc
UyMMokvCom5ioC//nabftgRNGXh//qBybPzyMt97l5gQPCHq59C1Zd3kTsdrn2/5
PGUFMPiVgGyU8mT92NDPeIU4/nozmdRpyoXXxCTRDSQkaMVE1+3EmomDuXfQsjEt
WMTLKfYZsetLs0id3IY6wQllxrSXFkwX9hWllYgJZCV8uY8bVtK0TNjpT2w4CSjb
vjkQkWLbYIg5i23GV2y91KDWFgzmVVHuyfiuwp6H+yGlNtO2bFWZeEVoVdDtUcSs
e3G7RX87+r46p8ZyedV0TM5t0GB4Z6Pu5D+/tll9HyKbMtp8VsdGAur2sWo8D6En
Bfeyw3JHQHgDIvanzjLJnmkUHsF14DGecG3Rrt+bya2lBqmYRWMfURAOzeCXb0Wh
q1TQo6oPlAK9H9V5cX8miKS4DN2wJqtncr47aiRRe8Wu4lmRGXRyG5bNO1iQESFN
1qTfyNDnJQvpWak2sbpHFuccMA7YmN6u3SiYLdUMYqpKbh165d5NnVK13yD96jO6
8ALFmB40NYvmuIuNyjkj/C9Uiv9ehjs2efvWLEluz5nshMe2m8eA8qiYn+64ZtGK
iEy3Wc3tWKfnjU0HpU6+a6QkBM05Rmne9eSKpZ+WIClWi5InObBUd59/vf+pjHm2
5OHkCG6NRfIDM1P31eGNlUmiEiDSGA9iBe0UEpZo8+gELmSVNLqq/2KGkxNrSWhi
rIrcGnwNJdh29cdy0EeuCkATdjnMezA2ErYDeDfVbFiy79YWUYyFL58y32Vd4aTR
K1w7feiEeOFE0KvvcO/biW46iwsaD8Kj5Fodb0T3ClruisduqpbaMmy+E4wKmCLW
Sqh3Oxb5kIVRw9Z0/Gawy8ZvtiJYm8mANUGSn08nBwK0OEXzB19F0/wYBXAMxBbj
DIvIp5wj5LEjWn6290dMxDYCSO8tUdpRV6DeLzeBiKvUk6CT0lO9Ps4eB94kvNX2
6TIbAs+m4lds31VToGuHMtYzQnO6ZLzFkJrROBLw9gMIKSLn0I9gwGySNLExTb/L
hDWKMX/0Ae+v7pOMXgiuCgaaLifHduAyRS8L19zJBzZAhjTDFpKsJh3a+Thcl6FK
gDLPgIWK68Qq7/5Pp8lYY7BEsDT+VGyrOER7j5SZKYUGQOKEp8X6oGPmD8UFIhaY
kAL6nxmvMIpeZ6ofoNim0Ru751FmyqdBYPCV2Jy57VSGOdAZLWqpkqFqLzDpszHN
J9xT7dVCxXNvD14FiKC0haqTWU6eszlSqxZcRPOD4ANJ9bv1Lxojdog4C0IKmkou
UOpz/ZX9ZT+epBTrWmrj8UdSqkX+ri2fLEUT1q/WxgluXFOg2RS6g0nRKnH75TAx
WlM6fij+PsrTaHb93hmdHNdmVJJY3h5LxUDf8D0BIsbzNVubvdVAA5B5UBgXUvvP
iZC0HJQTw+n0ChOgEp6SdtlRSaiZ3VhCbPq24K7f6ZYQFMf/Gc5tdYos5abhQ0Tn
UnBXELnx/+rtJH8+Vp3FcCcHavOqgTr0V5ZLceqkBFCFeFlLa6iTVe3xuSXQQUy4
zlCuAd/FzHmIh79mnCnEDfFM/zI1ker6YbSJQkpz4U8okocSTb0H35xflMuyPgil
j3SmwieN2yhMAshY2zUbrS5spfwYRp5MfgCeEGatOq8sHS4eAD6ApJnXWJhKiQEO
bQekAm+oXYXW4CkCbVVX+YLJFeUNnod+3lltVz08lJ5EszTHl2pE9oS3hj/LXSbF
pkajHj2FSTYBVmFWY+8zzCtYwY3lU5gQs2WvdnqvISIo4vnKu9Q2VXhAB3vyOqTu
eQd1w9LXrqG2apGTcT9I/sdnRIOWdkHzMbu9GO+UtQH5RHI+b3jCi49rXLtZv5Jf
iOgFP9mpx5Oo+Kb3jDmmZ6ZMXOXBl/2ZY02BybyhmfC2bzR7WJhQ0jeQUkxRgGuF
XbupGEAt0abBWrrXpnNdoUNNokBDLTenS8p60JrO51Nr0vDJYKSZLE8HytdzcVdt
JREi82Z+cQq+UASRrL4zghzzwZfwwzRSFWEcP+TbWGhWURBBptwp2ovuQUW8Jvf8
T6IEOBadxLWhG5foKZx7qyXGZz8xJv34/4bxg61T1VlQoXPMPuPfMWs81qnn9k2q
aHkuIvm2jbCLpZzoiOIf7me+MNTGQrLvt9JoAEFZ+62qAKfXmOkdm+mBn4vqP3/Q
G9NMoO4yZKHyOnp80dWuaKDtY7/la1ycq/kbunw8/7Sq/MGaAZeeHsxbbbByT4kB
bvTTWKE2Nv62qz9wF4XSUZ1/I4Qecd6tdPhp0b0nk2Tp/VFj96PkmHlU+P2u9z7A
8j1FCBhFeDTV0ayg75UrYDqdmDZGXawpMhN1lFg+1ICeHveV5D3o4xDhVo2o9CeM
KClnFLWxo5in4G+D11rq/t45q9v8RGD68T2uaiTReCuy8CesazUqyCUNEFkFfOYp
O36wwL2lUJDRP7kM4EfKW4lP/l4JwM+9sJXeK0+CvJjWVivJqpv3FJTWPD5spWoS
WHkl/KWkkdwJvkUWxbKPepO6bhzvQOfGzrcHs8p2w05gfKRob42iuVSV7+W24Gnp
/h1p1e5aqrmX3bjMDvae0KbokkPRPv8B4qL8SfaMDJAUzchVy+voR1tYl8/C8/ZH
YyNbgQY0rJ3Ov7p/ySDOLD15m382Tm+n9TfIafqNioy7J1b7FWEl6knHgOVdlj8O
dn+Cy27L9VYK6eMLWRu8c645zs+kn3+eSJc1mRok44n2rvhO6XvTFMtLAYAHJiSz
Jao7IJ7XI/9//eZK9Ll+isxaGIFaDp1tRrW6/4mHkhHDFoQAGlgIkpjcO9l00bvr
sHKfm807d0VBZlu5ROdw04tUZxWkZxynljMF7gtXylpZDLljYbWqxxjUY7Vmlclz
GNxS4wu68jU1UI477MpLhswn+Njkhj91mOvQqobxL5co+utBx8FYx6KNOcjBl75F
lFRZvDxijQ//8uQrP1kIJIyqx1U3yFpGXybZba+RkTko61BJxVkg/890pdNpYxt5
cOnmvjoFQMD5sFOS4zlQHkqRaHEOKioPp2x7BtaUjZrALEucXmktso8OQ/eo8BdN
qZ7DMoHRyND49qs6+E7yQgOs/mEzA1SheiBaRrN+ZcVZnMNcUH8lPjnJy/EbGQYt
AIUgGhZl8EpIPW+bVtIcnKMXPNy/UgctFQC/aj/2xHfuYv9dViqTf8kbhkR5/C7p
CZn8m+o+g8QBHtdeqPDTSciSMyMscxp97uK2CzwtJJ+xkCWJrFGcM+RenUPRYlJX
VloV+1o8VGZtCdTXl72lcUep8wZXCG01CXSR8LVyuxKKIhXVeMKJHYUFYWxRHEPz
JoWCqDR4U8LRlSprctNm7PqpxdCmhh8ZmMhQV7yYmrB8fRL8iSNkhalEb0vbExec
lMcjDa2CY2yix09gfE7Kx9NyD0dNwtnr5VzAf2FuXNM/mFKzdi6MPw/WkUijBBWl
JnXXMzWUuCCWUrsd+PEvdxbUeCzCmkDu6Sz/9gnuN6FRk2OnpHSz9qxUiPqV+GT0
wFpCN4LiBBaFDJO5R2XD+8/Bqlzx9ggbsPshiJvQHDax5fjqsjA6wyKPoFZ5CuNt
UyVCoJ4sI2Sg/aPyot9jLZV3+MKEm5cgRXxzJauhj25gs/SJi8INMhY4+qJfqM2e
OIl1KSgvMqsVal6CJM2pfRSJdXdIGzUHaWEEbDuZ0Gk//7wFCeFUBeQzjrV3OzMc
oTuIp+gHusN5d9lkwMwfwyLqORjTlTUIuiL1mOZKwAmimAICcHaEu30Leuw+rPWa
VPoNzCe3slZM8Plf39ozQH00v4X4nz/LtweozYomB7VCduyOhsBEAZNUknmRoq05
9MhwgLiykLarGdfWOGFLwg2AupDNGHCPAKjL+xyFrDyU27Flm7e7Q/z30kR8sbd9
IZSn4OF9zE1bLqYBA08a20U7xsj56F/JnlR3h0J6rdtpdMvmBJ14iDZoDXr3IZ8Y
C/h8mg453OKlOIvf+GwgLwyYVHJWfAXgu3TcGP4d+IZMluTmgqIl/GzmwU+Wbhyv
/f4NatyUIEH6LamDEktIgLOeh8pVSXigLZbOBFdBfb7x0ekxhw35N1mtQNdJtzu3
vr6fTdR6ZqdQ6v5AmnQl4X8saXf/sy2fOey+8594l+7AwUMcwDCO82/qGEFvB7Wj
ilUeDQAJ6njYksspM1cUQn1tpkkT4zxTFZm61Tga937b6VqGdpVo+j5qButKUnMl
NZIekijU0J9ghmexuAZMnZGjfCIRi+QAgrxxKTmUQqNOfp1sVR9K94bl+r5s11FK
n2jdgNQOVtqNtxsVefls0McNW24w0kSkD2+sujdVZhKoYlkoo1FQCAjHK8DN5By1
2oa4AWvjgqsHpRiLWhEF2P/RNao8dm1bzaVK/YPRf5+0hSUSzrzcfvi2SVJfeBTk
AafaSuLvp9BxV5gKBceiOz379xES2TqVd0frqedHtplMgWzvZ1cHfKFm4bA6TjC9
BzYQ/4fEhmGU2j3kbtD/NVLiLm5DQDyy27zN+DLbxPZcFTNgbQjLlTprksI5mAj+
aPnnKsG6Ug/e3PzlZPPJdrUKIzNzZg1tGB4qSIb15Vn0QsUqnwllw+EBIbN6LtyO
0FA2GfTVCcU7OQGx1Q7n6tmuS2fWiTIlJph47c8F7hDGBJrCx2WEVd+e+7XrqL3R
EVjsfqaB8O8vjLa6uKvcNcVqYsUHQh1d/drK3GB3i4UqLdB9JIAlpPk0dj5viL/T
TOHONTTB3OC0+7f2fiGKSIh3lXmK+y9GPy4GMgUIJ05tH9B1MnA3JrDXeIr/Y6r8
ov3ra947AfaLAiQff8nVU7pLkPBu99fDX2RT1sbo8/EeukPg9OUiOd+jOceR2CMq
enDWtnCouKzJ2D2Tpu8ry9yuddhlPqo8ILN2b1wf4YnzJlzhkIpNgknjI2hEk1KA
TMWhdZdf9BT4DZaBHTVV6tk+kX/SSLfXvdn9eNlcRwK8GiNtLbe3fHQCI7WY8/YL
MRsn2ZoKwa8YKwExf/c/HzdWPMmuKu1jpmeUzJmefar7jbHQTo80GXWtpcAENS7J
eln7EXjmUZ6037TPI5xVPSDsvFDyWLxv87XP8CPzzqJxHtz63n0tfjPuF9tvNrxA
2aG8FUW6yrg9PYkxTx7EEwhYQ2lRjLoXi2T7miHt1VUh6b17FGkTCGyKlDP0iHQw
YPSqZm/5Bvv4JdnmF6/ChbrZQ8JhTe1dgKnJSfQyZ2Kuxv4coUP/3ye/wR6QAoBA
l6lVN0FZGlIfsjck5B32SW5yoYjn6DQC1R/DFKTq9x8N/K+CUQx4WrDNXU8tAIqp
Ey43yVelSB8Lx+yQ+wA6ZW9hbvE6XNm2I2wpUmnS2Izkeu8BeeKMW/xVmTfZ+eGV
OfBzY3zGwy0PDIck7uf8my0n/bjAR/iDk3lzoG3tV7WQqV8kqMD9crDVjjXGEUqV
MjDEjD6yl1PdhBUySOJyBLINlKQTJaOCFvMyy8F//19gdGxJzHFDmVZyFU0W4HyR
ZwzNlX2Fi+Dfja86/7sWRyhAgaelv7m0L+BawYQHHBzP7bplkF5hv3JS9Ht8qR+3
x8KZASpoRfI8wVlxPQo4VTVDQ6eSJncZS9N1Otkwca+tbOybgTPraP1fCYqC28e9
WMo6d6LD+EFImtLRjwAG8FzJM4+gJM4I4y8uPjy4Z8Xbh7YQiG9in4kKgzLbUo93
Jg1FgbuaaHAKa1ouRhR5kOnVHbCJUIT4CZ3Qs+P6z9HtffvydcC+fkzK5iQF+tZW
qLOJ5178xdE6gn6J+XmersJI/bE3XyZ42ZDGkqn0Ehn77yCMks7vdpPyaFPeShz3
O8ZEm7Elo0vcWEvgwl+YZdtDv/Vp2nsy/ogP05RKpqfQBzQ1pphn/cYMmLXVGxYe
LHFTM6RPlaAdLYWVG7CtCg2bcSMM1Tr2HQ4f5+xbtdkgnippohiwkNkVr4uQQCOI
YiEPExoSSWS11txa4mBokHZgOCDDHoD6HGE+OeoxoUv67xZ01wpI1rm2DDtSwdos
Ampb/OLczFBbYzXu4LBdiLiJanrUnp/lgZlgK+ro6TY9vDxJGWzlMEzoHAQzsgeV
rj7XlIEtDsAP6fLIA5toVOi66EhAjBXIaZATEbFr6iUZlpY9EEA1zziI+c3rYw/Y
KF7EARRcHZiIRsmWaPPEgebfg+zbwnxc+bPxYOl8wbvE12+oTjjh+DdUgif3HAZu
zGb2U7xhCclZ68aB4aJ6b4MJVEOXT8wbpkoCMzUWP22ISepM8QC6Om7EHUqkfA13
yyWq5O0RJSHgQXwuxr005CiQAskvJcU/COMYm/Wxlq59IYT3mfCcMNQaTv+Es0Ff
QTdO5PGm0HDMFVveeSEOumTrn9SNy9eGv0mCbOva99bKtDjbLSygp/3FqUiph4iH
4ei3ZR7LMVxufBYS8XWJZh68EbSI8z6kaHHoeKgeQbRZ3EjVHDSvulOMsRYVWCmG
5gWLk6tB0W1bthCHVRIMQnJsciRPHeA38YhG7pw6HInms5QmbifcLlv4Ungx+6PO
5Rs9wbrOuVmy2edCrEKOK0JI5sQkMMDH9dJoVACGm9ubEmM6AXzmIAyVjq+m/MxC
otlvsvadWmjMz5RjjTLOb9hHsBslKipAXFT8+muwOmHYjfKmpPdXT81bq6pnZKnA
i0rsYfxZShrk2VryZY8HwnCi5DjT61SXv8I2AY8Us5YpoGAp2+2iUL1uBk5PPGl7
qi5H3Tia3/a43tvTyPYVIzJru1hDTWmIUNW5SMGbEGNjVRodI3D33HMeW16nPQj9
sJm6r56CwNxTFCaz6blxRKggE+sfax3x1QGu48XftB7w4H3qUnDcjZMjRL/dXfY4
AXFzfjTpGof5loCZ1hBn/9v0ekEoZpTCAoBJP4pcFmsuADnO4+EUTbY14bNZqC3+
fM9PAESfl/f2toxCi/1TDWkYIWQTf/MxOPk8+7fbbsSEOAeDTcSlGScXO3dro+Bv
dAr4j+I6ad+E2tP5KfCaEdMSpt4yvAbxgBYir+YHuo+sIzHrE48Kfc6LCPoiT4/u
42odJZ5OfB/yPsum7SBAouZnWhfIJXRdzl85U7oucR7uSq3bUtq0Soe2TKQz0sf5
tUamCeYK+jdzJC5Jal4jLeh+tiH7GjRFOR6AV+r1zDbX528tip99s+NDGCjfiHOT
AqTqN3vOlV6HStZhz7CI5wHucFql24T2Pht5dHoT/tinAFEoEBbP0Aujo8Iz3Vou
w/yhZxDZ6bkiBlVQE/5K6o/r1SegLNgzcGj6Q7iWg2/SVs9zP/QVmWh3wIhuAHAl
0zEQ9MqONYB8eDxOMQkVUHzjskf+B1sMiZIib1Cx2mShZYDbqy53sCZMa0NcV2ZP
hAkN2hkTzAKimZp4S5/N97mEcPa4AfSqZzXsi8JwZnMObitm+TF20oadNVoAkVpv
6EB7uRT60GgFsY+Myf/yAQEM9CP6nN97VrihXdV1f6Hd79CjmLxwvktCZOH6hbLe
Rc/76LhyzYCric1r6MHdBbBqJruefRpvt4uTbrcJXnlKDLEvf8K9CCbALdc/B8sP
KWTMjVed8F+pvFnRZTKOH4Q25kqHyMgrll2Tm7F21Ht1H1KWu4mUayyWF0MIzIua
e71XcPog3PAXDBb6O6AY9O9C9M1x1t+yhoWfvhekbG/R2fD0GHeKcUJt+qi3Xbz6
ZM+KER0w0pX2BNjUmudfZv6t2db+WVZdNmOSG/qHWbgAxEjZgFNWLmh87cKRxL2p
3zUDpgWq3Dd/gojjjAqhW23+Nkruw59yKL6+rB5VYz5iiP5qmXIbW+s9NcFOrY/7
0391guFCkjDBFO0CGw7FgBcoRjsfFJ0kF8MAn8f+g5Y9374S8wQWDswVngU3E9Ig
Su9v5OTXEMZOnYhnpY0+gkdwdT1KZop/gG/2k+LT5va75r+rDK1hQTGmJe9wCMZc
XwtXG7/apz0RaBxCHD9eowpyqIHpVAcgI9zAllwx+rKTO+hGzzzJ9IAAUpH1sgg4
IoOZlUOSi61tIzRyosmdHlQeMIeWisTbQOUCMlDg/hh+zAZx6h7/Ejq1rCW1+qFg
kNfkyLqPCm8YGeJClyyT76cqtsWvAU6fATA9dPsjqa8Pw2dLfTq+4QPUCSYRAQGR
In4/LeNGq7xFsKuJqH6cLmzy/ylQ01axnzRU5eYHcZMtY4kKXycbk9Kms5cLpd2r
pQto1mvtoiLJ/u1Bgaq4EjC4Ohm4Z5v/MFXyD42UcfuRF4WoeeR4FqWF5VfXNXys
54N7/DGiEMVYBO8Ejxw1SiHcvp2WkAzFDafy+RMHMk5o8ubxeu2GCKkcLNFQAOtv
gdTkz+o3ywOPbPeS3gqnmLtQvNq204el4wm9coQvakELgSm8lGdfigTnNpHG883n
GiZ75SHzFmqUr6ubAtbD7lG84qwP74Di55eOgtdIu099e92Z1Lfe+YfQzpaLDd0z
m3HiOPtUkkGhlIrYuYn4U8J85M75IaJZ92mO0mUMK9wMnKnHOCYh1XsxXJ6sYRig
0Q+wVWXWiD89A+/aT/yG1Pujq5N2iepneoqlJnhZ/nPkZYIiuDxuhS8yDeHiiRHw
XnqnGNsuoUTGELQ9qos8fha72NzrWAS5N05GgaEYREF3EyYGyS00VkxkX3Jy2JPw
vONsZM2Gp2OABSfMhyzStieOFt/pMdiYqoFEcaMceMieDZRkcRL5a/oiJTCL+a6j
G5Be92WIGUHpNxTjvtFyzF/CYeA5qi6Op75IFb+Ee+Vf0R5+8/ZyYlRhwKe2Xj2e
YtsA395ErtjPGpdPQmrBgCEVX7MG68aTL/xvWDahWLpxVKnmfV216RTnULyRiNnf
RKao/KUf5v29iYM4S6aGqv21vaEznv2LAEghgSjEJtETQgxAgIEYGzJ9dD7hZ62M
XnuNTGkKaIKVnCozezXlf8JDtXOsHV62bY1a7QWCjboPAgkhIUZi6CZXY7hPas1b
T+Fe/VT6nAqPy+d9Lpzt1Il7F7BXNHZbKbAtLzqM+MRH00Hwp1exP0t6SQxeGh7a
/2W12pedHsiaQZ71le0m16XoRsB1nHBbMseiaXqmibiIsBJSKVJ2t784vY4R+ALZ
oTL06yXq/scbyoGh3d+Y2TArmkYpIQxexubV1sG546+oIlVDh3iZ91PcOZYpmFM6
DkbaYcvuoFrkBs5Jvye1/RIzcpaX/bl5aE7Rp2SCMfzgM+IWHfZI7gdP5BrVe3LW
ORwfzfWeqvNYoHtw3gaLiqL3z12hK4BTNI5h8h225I7eg7WHTSeGmnos3IG8jOze
wCKpNurqCiQ0AJ6d1jd7Cw2VXJMr62mLIX15syKkD+ZSRUblxhdLXJtfqCDExrdX
NIL4lykN+AWVENXNVEZXw2gON4AQ9ZLkF3jzf1bPLOv95Mt6LTEYl6R1AGgdveML
nxk0jYT+FTiPAQfjJDjiGvXV3WYTzYAjSsrid3ivYatR71x4sTZYleR7gKFgpK6e
voDvJU0/UwQr1Us0MgR52+pcrVt3epWsYDh8Su6ozJuTRVoZ4j9xdvhY22XTrK2J
ooxKglqEieFajyl0ho7ebyVDMntfpkfP56PCyOJZMfXMXa9L/RT8mirCcXlLaFsB
Dd8Q6HaxsaJI3dJJ+ZXogKfEu2UTyjua2M8d7MvvL3qiWKqPpZEX5qjMLeIS+yhO
zSHvO9FNT7e7hyISfPHqB69Wj3nflVKJ1sfvsUumYrQvmoQLyzEW8r92ccCfhyea
Qm2NdkpBVDXpQVPUhSLK0MYmuH2+YjhwcmHEHMfA01LA7+p6kEbtA6NUDxHKncrO
+i5BrkUyiClykuOlzmH/zphTDfShPIlrJFKa0VjPm6E9eOKJA3Ubz9cyWnYZz2Kh
1H7/F34ZGEfBwaWhNLyt7CxM4KDTATX+uSdwZy1TVjuzokdji3I2VFb6oUvDWyoK
U9JkWTPZ+2NPZAfbncEQIWFzNZzSacHkSADj4Hu7J7A9wbDX3pCt4x3Q/AqcU9K4
b//56VyEkWMr25CowmfQZ1anTbzPJEnehd54EJ5xpNuNOIhdUk5m3BJf9oBvIRpo
uj/G/Wsw6mpaVg8p1l2nmoHcqDYjeraQVGGw4NGVMRrtAD2DxLq4QU4+8010RPjH
SEYxh/KouMRGhh+vTOz+w6d6m8FaBai11cv0NZ0ZCxDmPdGKmII7Fp5IXCYCRc6p
gCn9MhFd6pt5S/HyxINfNlM4b/9C6N3z0f0DTgwUaQ4TuPHF5uKz+zd42Y/tag7c
p1jkyNGfs77utskBNht0ZO7GGy+AySLObMUYq1YYjYykjRV1aqgSUe6AHvATjSoo
JTCYgaLZJHWoh+fnrtJ/wnBcp+rPOLeZ4gGcuG2XY+EI4uyRub7c8cmNbNeKARGO
FNLB73l1tD5zpnQdW7Cef8GpUC7BDxbQHpg3ZadMy2qwOBN5wPgVR6kX9Z/WUZyE
xgMel27FrXxY5Co303Nru5djklU148R/Xm4hGJzrmhO9ZCOjUo0hLCMwdMy2F+hl
kfniBguTDg1ZuwE6Pt9HIrX1d7/qAKEti9WKtrQxUPusAmZ9N+xDiDD3ODjC4hb1
9BhsDokWlzvDYP9QY04gcLPhOBvxC+ty5a5elpyPwALbUTwrNTTOGG/4j+C1a7AH
fCHBYZNMGI0eCKpVH3Z4ZsBefTjVKhVNHUppKGI9HD+MPB7UimgIQdTtqsshwh61
f4yiUOy1EyEFQTCnJOzphA2t7Lcpyzyl83L6xIn2gVIQSuj6vgrO4PW0vsHnBC+e
4nW2q80xpE7lhbYiRIE5pWyjsimzrVjcCRABUFKuW2W8XhoxguRzCTKfUkFC/wWU
nhTdJTiCMQEseH1va/T5oVoM8MZBdtH3WY0YlomJ+8yXDfgoJrTAXd660wIV7Hli
RKn2YLuvYr8pkBxh/wrOVzfLULUwcNumy2DRxReO4TeAiNNluIF4CwNosAGTFYyR
PZ7ci7HBRBWGK0lkAzFKAftOLF1bxtLj6eoMRpJPD7qUWKCEPGYLtAh+f4GIHeTB
0jU6+3WTB9RLDb5ZboYFot3p+ZD5pdzhoHc56aHWIB3niadIn76r88t4BeB4pDQv
g72CY/C0H55j0CQQ27ckLyWzNEFy1eIDFy6IcMOtB6nbhQad+sXwBABkq1IfAZ6y
7RL5kB4bW89Jjtbc2DE4IYuVcXLZbgXlmuvClv64eVwPcO7JSdR6SwT95zgV1ag0
B+gZZ+3Eb1SiXIntPY1RNrDM/d8/9dHYD/KnhrYGq2VMViGbDxHzJM/We4r0nnLu
cHsfCG3OFlMSF6cZb+6ZbE82Mh3yA3MT2CvXUTMJhY6b1wjRWo+ipyq4wiRp+OeO
25Jmy8zspj1Bve0Xz6RcuqdI9RLsygiK523PMpEHF39f0mqONVqQ/ZwLZec+R3Jo
ix6L+IDaY6opR638Crc26p/naOwjWSv3JTLbzJm6fkghJWsNR4Uf6cSu7ktfgKdi
Zcj3DysiAotQ6a6nefELlIRjuU6ng5bxMNWcUZ8hS7jDSfpfDdwdlwBjnEFQKXTO
sUofVjxAVmdGsSTr3n7Nr6tRfsNnw1eT6vlxobXX/VzvD2R62SJwKoeU3cxexlwZ
2qXAW6OuuL6KgKjFOvcLQGKBeGnyIz1h7s1XAJCApdM9jjgfp5rZCedoTufFL429
6+WQSW/pxMJSstDGT7vrYQJ1r5fdiSwbGegMtRuI6MuRRh3WP93akL51VNluDtnQ
cjeY3COdxj29qgUnBigxeN/gIVjNrjVOBJckUlfXvOe39MBiJToVXA1ugCKwaHDW
1uOPoChe/XxJ6yl8tpadtgUfLobJva/snphjIeNjMjbORDODSR7ES3+acV+k6dbS
ihaOzmEoErKHn85WgEX40JoB4p6Jh26HGTW9SfTzJtQkk1k3eYwl9rTt5UqvDpFe
37XLtTMgYkUA8njPyc1KGYBkQP9I8ol9A8i8jLknbJGRBgsPuakOJRhd6JiBMFGc
frJLc26wLQxzWKrazuXhcvIpOWKQJ0JA0KfMXbmDJD3bDD1tbdwxlghg9deUbl+S
fYhMwJLXiAvQ8Dtsj56V1Kqf1E+UePo1OxPd/1V3Lb0m55U4trXHOFxLCPcxamS9
9X6Ej68/EoLy9N1hCaLChBDYDWgAruDWL+zGrjJrvkET5juRscTsEfnoi4wSLzpY
N+kYZOA0RbTN4ykZWvWFSFmW6tu+dvlxCvvdEhs4BjqLuSA4g4TFkgcxq71xPmAH
3MebHjNRQ64czJ/QH/Z/Xb8PAeHU9qtvE0AQ2vXFRbka0hT+6cPJROeX9ibWak6q
dATj5XITCoCD1ZlaN9hbmqvaTcG8ztZD60zj9li5CI2LmPL2z1T1O5H9zpZtkUvP
7W9QnxpR5/vEWN5Q1MVHXdxeOvsaUuktJ/WFTpntjTdMNeM55ZLG1/fZ9nUdDhQu
6O3D60uUYsXq3N27FVyRbm7zhi/yF2k17x5S3cUR1MMqgTBWn0Vua/fTncFUH+zg
Oeg+N35Y3Tknq09HnOs+ns7ttox/8EOd7wSZQ9qqCbgMWSD1bmWlgSBIXoK4NG2n
F6XKBUbPS57NEY4BeiGVIsuaOMbpE+wCWkwjQCR5qK079RlI/B4w7ntoJYCZupRL
NmtUIiixEYqd2j/5hKWA4zh0405yPTVIPSjY8k0Ov/E76/b8X2eDH5fFlNXRZscS
tEsc5fBIBki18SAvYhGEpRwL04qoouzQeZk6cS1AxBYQH+Teuod+SoWKwCd0gWE3
xMOHI1zBVLQ56SilFKIiKhrPQbNEdNGrWk0zOMX2mC15XKpil0UNXLJ2e7wVS2iO
KgfdcUS0/4EP959px3ndxxKpaGN3f9guZhb32CcdgogvQUukfdLyWA6SrwfoCjP6
VxJXdOhb7OSo294pZqkzx2X4Akouo+p41jyZf+uJo+e+yaa84gNT04oCNCLfEx5/
a5nfWdgs+EX8D2MtV1hdoFNIZFQ1np91vMpKk/pLyKMAecAmD/BqmXcCAIgBvV4c
3hW/8GxlbXSwj8asBkBrGx2964neba3NKXbajHP9pCjWc78P/w0JQMsij10rPhXf
xWuhlGUJDdCbs8Z9RssP6wXuZ1TtrsGfOeyVRGrHGNE/BjWnsofamPAyeAn1C/zd
bpTKFpTMFkbT1AxLPjaIFRpieuRNIl0CFf/u2PaAolHlQUwcbe9BFmVFNzlXW4fg
ohUv9WP/a0liTf1GJOSKv9pd7fGdlof6VNFF0kR3Cxtu+H5mT5WvMhWHB6yj9ibq
hxmWHCGj4VhsANZLOrmAeIdN/9USQh1rSkctfjAxifMxJVzdid6vgPFDXjyBl3mT
od+WacPMibzhoYNdJ0csoGKuCEcnvnomRw3VAiLYa1o6nVpq3uifU+ek8+in4mT3
TQDAFqU//f6+SpbSqzBaVDhAo8ssSvyMA+laZRtLvfaZbJNQCEbGQN2TaaDNi1Hh
2mR20tEjyV9bqYTPjgselHD5A9ZNlMAmoZ8rVNdjqypbikpc5lQZ1G9AK9yHMz+J
zH1hmCGvuNbluvlGx+GUCYtTO/4NLbf36QLWcnrSCcmebkyFpHXVOie2wi5NbZ/1
9Df9Jj69H8cWjxyilzU1Rp9h0Xm96DcVXhu7XtNGLISK7KcPXUpgSUuiFa0NSAb7
Ob8mAp+2s724tzqR5rYZgYRwTgFKDkSdiPJeiAbRaHrccTh6jMSHRqXM+qJlc0v1
5QbNxr8iXO6PoUCybT+M09rYZ2bB6xo7iv/y4VPGQjxzgETgZDdzHNCNe4pm7qof
mTd8KQK1QDXpdLL4u6rnApyIDRuVR1ublFAqB4iHqhC2yTWKBKqS9uQ1kNPPExL/
vpN3NnEixLXOn+1tLk1E30Ncf4O7bEFCtwvnpEDbKLlIu3hq8ZNHt5/RYwCeLUcm
UOzbw6I4mt75QFC6ISbbWIGUxnvIUA49iBgG5XBdZeTJiMYakAxuP4S24yzuA4N4
SZYnYALVOdsaLaaVVMEzTViISnNfPJ/oCYRrLRZOPuAdemukIC0+7f1ABeB3ZF9U
COlGupZzVu6jv26mf04c+k0zhH/ze00GHyaJeStakMRs8u+LG0fUcfoZykm+8OC5
7yxyFDNdvajH/ssVcPy38O0qPRyIRqCoTfC+ayXsusMHlGEzYnZFF8FOlUw2jM+z
mwsNYR9RYUhE3oJsV/mTgJ7CeHVqnYDp8oOwY99Chu2RLO47KfblhpSWefCRhyq3
9A9nC0+ofibY3YIFjR1BfGn0HvmYla6whFCTlrijRVfC9iE6SD2F/kFpdfSkykco
CXkLiyUYZPSESzUWCxd5e8dYSOjbme0E/02bvgzNnFBd8K6JFd0qzGlt87gAKTNc
8X85U0GfPdaj0cDr+XZqaKoI+X5BCAVRPkDHhfpO44ZyjSsXDlDuYeFZxIIxzEol
SGATpLA0L0dbstNdixbvP85H3K++5Pjc+YdyLXVoUrxJh/b1fSjNMZ6ziOFjiTIH
+fmgtiEcWxtwphjwvhKl6D7nPyCV30wLvkwxZ4oW/KoEa8LajRkVE3NVpqKeucxH
0wgLH5ypeBFnWVLpusv53m18nC6zVIBb09xDffy5jK5xtPBpyAcIQkYpo/IXXLQN
I/MuR21FBVH3F4/gLwyS+e6UwaDN3iHgcEW5OJ3KluLxpE8ilAbjK6MZJ7S6hTTk
7M9kPaS3Uvd5ahDy7R7OlycnszZd44D4uMsZGIqsomz74aUABCEBG9nmTaa+0E3d
pdu7MjUhTCUjpKPeZflC9WYP7cTqF6jmsnIhUbJhwByct7GOwliBkykYbr1v2LcR
T/nHnVDmRtAYirodgGpUTFko11gLXotWjSfpl8SxVEN+isOmMaV3bSWHy1nNhncG
eAnhJnjhoMlsGBuMuWQYqbt9Elg05X4vF61FpptZA1hTv2kD1OQOEdrldCMDcuBR
8Er2u5ZKN/b06zZJIuGI4LXd3wRkugb6zHYQnpzslDKaNrYdd9PDq9DGlgLGJUst
16cpdNs5XV0X0+p5AqxlnhXwnkUW4dUOwqk7/ooPQbNx6VBqkKCXa/4oGmA3FAxk
podYbokYfCW/IPH0LgY3e6XJeFSwVIwLkmHWm/Hhf0k42QWKECkXnJ45BjTGZN4y
ROD6KiC+W5VzBAipkk56/JogbxziJkwrtpqqnpYIj13py5VC43bqixHriN0Vbgid
Shsj1msv/fJK9h/AUFZaqmEf2Ce2OJ9aRmMqG+n4HOp5VIULJeM6na8fYwCL4fYM
ilEJwsB/qyu1aNT515/+vVEpj1EJUaXZBN3VHER8bQxGpwFpNKHQL3g3bVB4Nz5O
bW58ujLea+NmQnQlWJ0FAxlLyE3cUFOMK58EF8aRAmTWS+5v6TPLbaMWO++evt9e
uVg2dp5+dtndhLMeRZEsaAaoZDA7otxFdiTBKka6nH/Bz0559H6LI52bLE4HTxMw
COpyofSR1oro6k7sC5v0yzLRLlwTmnPevqU6AdkrHtOYt72dGBYAcp4Qxx2Nnm6/
uBHiesKpN2wq7H3H/vc/GxzGpvUGq2svyw0iT/3nBfkuNMzr0D4U4Um+XkyJL42/
IbjJtPbxAL2Y12qCfUvEbTJaApJojmVI87lpdRvsiU3uUkaTQ6SF2j8wt5LPaUT6
+KZIP790wOBHW95FnHOqoJvp++7qxp/3q3YYnolTN779xTNZ69zx1F+aUlZK8J9g
NXH2FV0jBRTcdjs/9KS1DcIPUXVMvpU1rxeGgVxW0KSd553WtBWQFmwarHhLGRvV
jjCxtT9pdWIaVCHt49EwEP9GGWCtlqLBeHrJNNMUMFSFtlpRMF+5KlKexh+oMmh5
GhWEQLM7yCpM05cAHLaX2r4o7s8Ik05v2Gl10RWxuHJp23B7Z87GlkMPGSd45UDL
LFCtLSPVnZUPZkHC6GjtcynaYqmXzrbnukIMaJeorKLL5FranriOyZcdwhzGLW9Q
eVGgAOvaDp6n+7A2Irrefyes6Qsh5n3pu/iYXq4/+wZo6K5PK4LfuKY8S4aPGTPQ
sTxYGTOWq+VxM4h9NaxrHBrQh8o1/odQrAa4jnXTeuvK4N/tu7I+OkKYZTImpksy
aNsmxtC8ZsvaZuxvvHHFHyRSHlcNzg/iB3GJjs43PrCNceet82gQJESY1tq8J47s
ga/aZzkWA0d2dP57OoYORgkOXFDKkf28dKrJv4EKp7rZnHnpxWoL7zibaqm+5ZCt
GM9HT42VhA7L8p1TrW5B84Xv55CRgyL5Y4Kv1suuKyzEZnL+ct/Mrr7L3BThT199
ZAltJXfwj2pUqPOD2e5A0+Hbdxx3+QzEWmGP2rkwvMvUF7FxeVxeT2lsBK/C+RWO
YcLHgnKxMoKJw7GeabgKZKMXKSH/kQJRJrm6Tv53aVWVwviZlx9XEFfzIdxsHH75
6NjgDA+9aPYp/EqjIhJ4B+cxDCFyxjA+KexbnCHGFJUZelYgRBvnCMS/FBZUBLej
woGcE+Vfai3iD5zt3oawOQbItEaG5dtsdvno3WSedBXh/tog54vgpmYmkzGjxJgQ
GCNXvsbkLMiDHYBJ/etdiW3ToyyRcyF8JklGN4Ig9s0BzwjMUam9YZqlbJl7XMpu
n9WxbA+T7Zds7E8HQxKDAHK2RSV2fmUAwnYymSYvHOE7i4ZhD8C6cTXsDXGQvoGW
RMGGZgF4Ic/lA4TYG4/nsl20WML7PgUWvYcBI8pU9U88g7V4dh9Gicpbo9j+VLDs
TkFODst9/w0jPNQo8JGizEj2ZbGJONzN6hiD6rjw22XL/DwGw7DCRET4mSzWHUwf
7o80jTO0cEUsegagyr3EU1H6rMR/gq4PUQWH6uS+qr+q0tDrLtmnV9kPS58VJEL2
OGXlB5vGHdcK0idDzdPfDmtGJRqsWkzMPXXo0m/h4LSHlnH9sMcwPiWRF2QW0X+H
KuR56hCuJ7fNfQr6y315b/D1OWIEl2r1Z5ilm2u1I3pZzOGbUp312R1WXI4s70LS
0+qavhFX7+grWF/wVN5Atk6BAVbZKd4R2ZM5uOHQrRMcDthpiesU4waMD033/+JH
OcY6oXinPfdWglBEfml89LnJKk+/syA3F+zDsjZF4Qc6W43yDgcfJTsNyyBOtGSg
+4gKWuZe0Szvmr2pygA+deQMBaFq4PWUNnvYE4XdxG1w/itYn/AiOTMX6x0ZvuHn
kOagG/DGGeibt7bjXOM6uhaKE/icx2FdJwytND3BSuSM310DOnu88TUGoSbLbwlV
8I+dYiq6hlNKnV5mQJp0+F6RBTJQP7VAV+FfBeVDaaWPjGZwW9Zob2EHi/beMhTh
1JFN0fq+GubuqqGJkBAHE8W/sbvrKaHkZVtDH6bUFsi5dXehxmxtTYoTQ9Xz1VJ6
m2D2a6ApFQa14gIxIwqNCCn00DS45Kc2qXobp+dFs3GT7rJWosE2iZoNYlqE2fsE
hwtgMpKejdY50R2IVeokcm0HdMNAKSdfl9Tl80axJ/ImDYGGmLK/jJELlOfaq7Am
yuW2P9kpvecaRsPdcPYWXIfR7bORQAdbgPTsbdrXhniBNKNLFXyzlMI9RdkLyO1H
3AjIXa/6j9FgNVgyTBXf/KiKVLo6QwYvAUdy7M2o6KeS9gcuEp90IMPLOrQHhgYO
8rw72X0UwNg/H69vA/U4emoMkTzdBg0buWxUtnj80Pm7M3AQFRKoJAO1MP9d168B
0HBo5+2de5axbhrwD1XxpKIBawOlRCJGC3ZiYtgeaPHoxK5PHgJsZVxN2DIpdwdf
mERk/PuIILa1qpPdbclM47N8m+buvKSwqSX0ijKE10DqFjr0JYghlraLH1qKlM72
MVeA5Q2MoP8JV0M8R0DVItrl9NZEzcyJJFb84HOLGUA8juN9wuG7NZagwS+W9MYZ
KmcY6dr/hdyPrnt641nJeY/+iArQd5KMU9J6mgfCcUp3lkMfv/t6grLqXscmHNd9
OBJSGKCvKpOU7hzUszqzdrxKKgD0UmpF13GgUGG6Z7tCUqIamg6BhqD5NvMZ/uvS
fmCoE0zWSYYvxTlIuy6K1t10UInqWcAS8/RMrkraKl1ILU83jJT0P3KpGoAUxRR9
FnXNLdsncxQvO943VK8Y6XviqiyqHnDX7d49bB6dbbRWmhT7Er6munaHC23q8cIB
xkujLqg0xdRyHSnCTWgTGd9oE1q/1zuJv7kOAaQdbpix6xr3q6ZjHG7LIguYmBsB
JgjsjXnhvilEbgHg99A6Ix8wnKG8mHBfjqlyvimtMgq3QXQBdOEUoas+esBK499i
M9R1fKk0r12NYrU93hB+M4yVLhV11txwd5yb7RkmH4s0t/P0G7cUEsgm8wylI2f/
ftbnz/23JfXCw5elCcg804fYv+vDEqio6ZHvVi9hviO0vZScuTu5tHhwamdr8NbF
pU50Gqdr4nuUuizDpNawto4t/mQeX6nSZdpqjEKa16pS+8Va4NgIl1ce6VT/dHFT
fUZ1UwQPECn72BHSkuCDErXqtlc9z5O1Y7JOiZkPUDQF5ePl9nUtbmehOAdlCyvd
XLF3xcKRmMqNJgx7hKeAe+Uw8h/cAqlvV9GxhwbKZWLWcqruMMl2MpibZrStAISe
LmV7tLjwGaDe0Us3WGYtCBCzMEGVpW2PVPtzUafIkPK4TE4iOUevyPtCAU+RrMhf
9JaFI5ycdo2hvqAj8kb5WfIa0KMWLx2hjgK9Mh0mpoEH8kpaC6Chx7ps9YBua3wy
7OcvTrpU1GwnYL2ztxoAhPAbD6SqGMjwVp0fiOpMIa3fPlc78ZG4XK9lIJoVeba9
mMr7q2KHWVO6PUM6m8RKeqdu7+hRx+xw6BCLypsD7T62o7xApEHFMIwgl41NYrss
Upu+Tq8PEj8MFAW4TQUjYXqQ5P5aPHnP8/wt8J7rKK9cEK6oJL+/jn+6ovx3BBxd
WMe9Z99l7Ij2CbJbVUAAcUvOcXBW76aa6nmI4fSzlRF2W7A8en2MJUh6NQMMaAH1
H9D8javmorg/giHIttzKkakpvLCXL6aCFcScy127xi9CTCMfh79Gbdpoybkial8w
`pragma protect end_protected
