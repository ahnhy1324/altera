// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
HHVQORpS/K1MGWhGYZFDJ6+AQvNRReKdB7szo3EqxVGcDeGpbna4cgbTLL7FxmrnF6xhlb3BCHJ3
AAzVbjxrtSvDkSdAUMbl1hMGuRgkeVHhUJzmztUM2UXlh6RsdEMTpD0yWeYfuQB0dKXIjtAUIkLo
H/nGer9tcbyNRef3Jl3Zk/C8zBgWQXDJNWZPnq/KF/Fm8envXEdAWbkLVuz0Jgl5pOnUu0aOXEG/
VzKPUteS+a8l1ONlsdcfHnSDWuqARJtZS810kyDzqmq+F6xbGQzkfhh0JVZ+R3QNxw+antNJrJpM
/2wnT3yhH4x5r1ENWQkAqaIn/+yJYuWh7sGHZQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
DHC/RayFXMXGByxNQGHbnn96nDUiw/9RtEFDZedaUXo0DDxJnkJrI3HiB5pNGe08D5nY28w/FmQH
SnQUhKGjFxIAZBDxtgirDWY5LBFTG5gLzwmW17AJvDNF8jOjrNkFTujnZWqCbx5WnKvdmZpDV521
MHSgX6Lv374RnTVg3AjulVE9MkYJiUBdN1XH4/Nhwn38CFvuaSnT054fBDgk1DL3+6i4rn0Fb2Cb
sJVGKS3aIY41vlxzt+OTwHU50Bgr86TZMBVWBqrdjiIKRdUeSYfkZlpdrSeLWVrU9A2GMdvGw3Gb
lIt9zMF31J3oJiD+pYAAwjMxXgwvFiov3jHityOX2AwgXBQCBxycUxUjPHeKKQXYEH1NihZdu9hK
4lX1TzmPolOaGIHDKNPbKErvhDaIL0Ngu2PHlihFqZZ/gEfatc3y0mXwJKqmZj7tEzehGtADAv3p
4AWLb+ieswHXfT+77CtF6AostWqNYJqS6tHqIcjGpKD08H9jEzJdv9IxhCiK33QHlbk8aH8vGagU
AW5i71GPfrvvpRBKqlhqAYwl3rdhvsLG2lNPd2cbdAlJDGga6rq+asg31V5b3Mx3rXK0auj7hro/
07lqmhzcOIvZGFVv7i1qOK1LnOyxGdnFu05ntz8FY5+dvOPD/MSTb4H5wRr4GJ1AXVfnzpjCXyRK
pu1R2upw3XRbgO0O4Y+pb+B4QsPJp+kHRzC/KAclyxIwMavSz8zNbme1PVV0NcUEci5KNlQ5YDbh
G635X0RiWPvuHZDoUBeBM8Ounr9jr/ARvKBIuSjfzsoVhNeRX5aSRJVvUrQV4iBKWvT2Cd9b+Rxr
QpBwm1SyUSxx8TmWxnCnThzjyt6oRYQAKrI6UXJO/wdmUf7wwFkXz3hhLasDccFJH8eu4BMnvLlb
1geXic5zQA4ELeSiR7X3A2+QE9A970I+1cR4N1fnmiv11T5Au4MoNwVcV61UifDq13RHEbpDwGAt
dg+DrrV1AEtFPn7jqiD8t8o6YuPDU9q0y8FBu6QXP2ogdGt6HkUy0T4Ka6ZtS8MVFFtWk5uZyESO
ez0hdOxVYOC7UwGVfdVBkT9ZhbxglnrdHKA/qAdC21kHlmd9N9Ycw0dJkc6vQM8xY5lSJvo2aPoX
wgCzH2CVNJkDgbIpF/yGN0TFXXLrbJ7CGtwD/9sB7pBuYuOjSdLi6Bmjw/7Y3KB3nYBL8BIh1Ogb
uo7jbjRhFujDvcfvbiUYpZ+VXbJz/+p8o3WKFzZVHnBjgeMTB1LmCGfz/atj/0uH9uw4UFiCsNE4
ur29rg+1Wt/vNrhhd1XamgiQv9REzCULnxkDGifWt4JkMDSwhzFjnQXAMDeZZUFw5Fd78p4rLjq8
fU43WuC/tv183Z5gWEbNazywfylbNir772oXAO8Jo7sSu6y5D8GXriEZnbXCKMytUzLOp1YRxMpn
+hnqzRp1JLNtAVlZgJlIMKvx01xkkZiiVftByuP8BYGWaOsPx7WbyrEad6tCplWGlgfIkfZXHSbE
CJJfLEvisMmbwE/wNKZx9IY8/1FutcdaUdO12j2U8t8iy/fcBMggRKeAaoyqwmLHeu5NQXd7Iss5
UcjN+xxno/DzZFBEJ9TwBvjn9RcZ53/wTC4Mxk4220VPB5djMI9OquYOiOkolKflmt0YvNdGQxZM
Te+scdB9wu/VT/IBJiy6llMMUUG26glAzvQRpxTHo5RZSfKKgs/AGpE/BVhB0kTMqtV0w7OQiL5S
40N57urI1NMAcToWbudcnMOeQwRmw9P3tlhCh2lcZovbcdh98I505okC/9DBVCqLV5H2e/96s6c5
THMqfh+PM6b/d9B65O0troak06i3LtOeDSN9ksBC5f9mIqi7b12bhyzx455uxJejGSiO10+Ce+4D
t4BtuiM2NUeeql8kXOqZhJi0fhL0YeaXJOJ/Qlem8ZSsE6yysoPrEnYmKjm3HDpylHX5Xavh+HqW
uC0VK3EVYypx0ExEXmfEg51zoAoxwkOhpnIGruQd/jAd8Obn08tdW0/BtunSIR+9bj8oAAF3AktE
BkXbWns61Php3p+8WNhsBf+dfOs6ht7Qo8YbGOUXBIZ0vROm76cY+va8frV9cXJm+VlZCS5Z0sCS
C3z8MH7pj+i7NA8ehiqfahVD6tvmLVbUI6KiGGtAFug/AePbPm+j0pHU0jU0S7AIVYa518GGIuJU
gCrZqWccd/0+Fe5YbWgNobIAW7FegjihEAO58eN9ftQb/4Ade7hgvB4pCpI6HSIzw5aWuQXLr6i0
sqZsJNmwphXUNlYejsn5EbEGyJ766l1VuLfACsN8QyoZBY0vKYrivqNuKX+/AVIBwCEYSTr87RC8
kqh6MMDxN03H2j7wRxlalNeUPCOn5gaXERWzrmngB5VwCgXrGSKCh09h4R1Je6QPzXYB4lbAjyZd
kqcVPfuj0uW0aYbrqhhbWLjR8EUwjMmA4OPsul50tblhInlP8zQ+z+WHsDHYNNWcLjV65R2MNIkp
urFfRb8c6qfAHeE4E1B954CvKUHzzPwNKkO23IatiRnYHKv5J3b7ZGpx7qpL0kq/BVudpslDgrlS
khwfqGLn+pviUFP88yyP7f+4XXZrknKwtkQXJoHtwzGTNMz4ljIXOq81c2wocMeWi6tf8sCyy7pS
vGhJJjpfwM9YuKmqMziS9rT2UXTd1iqIHIMMjGUCJWzsSnQWCag3/xtq3qyy+Qc7ujrigIL9pf/W
7ubrXp1jvKrIHo0Z+7O4mmm1Dx6lckeRObltpZDDcXdDBYqDvtIrV9KoMKFoxv4NlEFsQfLgsaNo
RapZ8mzs+jjEvMcD1Lg/WtqgavifKeuoer2Xt4jnPbmx9nZArqcktkQRKWyFWfJRUDyhrsPBRZ/W
6XCokWXGXYrk+XUTsCnGBHtmhFP9QAk5fWCU2ZO5rFT3111GFxsEeAbRT9W+JO+DSXAAC8XTa5Nm
XKPEsTur1Kvfabad92BGNv+Ds7fmx7DVF8eLQ90JiZi1vaoo4OvYzRC11893Zo5aQwKRwQgOyA1c
bQ/J6KMr+fNfQWJVW/epAJ+PtUzsPU1yngDiluzD8O/QfTmUEcswghIF3e2O4cM/c/0jJYSmDeR+
lb5rhOvpo7/i0xmMLgELtsJl3B6RYGc2sPLts4ZPY4QctWmWINV7sX7gogX+Uh6U/eRqURO12DtB
xBSbnC4z+5UxODR3YkWpRxbjCT6NiGFhMs7tBi73bboU12iJNeuMu1ckgNVo5ufmscRW/DX5JS5H
0bsbEurVVhKHObgX9O0sZEDjq9ydp6WvspiydK88i1NwqYV3euY1JzJXaFENyvNQAASCQmseHKIz
wtMXzLXXe3xa40d35xZfdICBYWibhnW+CjTXiWZfpIadtKIf7Wwx6nW+8kIZs3+ASwrWB7YG196Y
kxmhujvQvD3giTFo/3it0xAGr4Hu6QqwdBMLFbpVupziNmFFih6BA8UKygh+qwplJ7UT1KtDV7cs
wIgOq9SqxE3pyQ0Vr9J74ZN9bGDM9erapMuF8fPow0KmMZgk9UtGv/bV2SaXH2ZhzsRzeACM/uSZ
wBMh/aSUdPSpuzpbqfrCi4aiaVTbD7C3j+bzETJ4/yYJ6vVyq4temQhY0Xom99t/z+SUgcgiRYEL
GpyfLu2vmf4YGP9UED2iYGwbpx2uHiaQyn6BuxvFZL8ZmEVFzMh4pzPzFbs5zthz4cOpU6iY+Sbt
uJNYLIEaRK2dABHPjUCe7b0/Oqq+v4raA1XNWAcRxM2naKnudZSKZgC3VYO5JrxzWLZLGWqIwWdk
Do8+nXwNAc4fpy2iMQPTZ94y/P3+fSl7LyzYblMhAtjbKggw/FdwIbsbgB6SRmxDlfh1mhNrk/4m
dzXBXugoyKPBSH1sl9j3EtikZ5fAWBA9g2XJP8MrrNDD1ga4naqra+gBKsv2AxU39V1YPmgeS8wl
UjVUuSJ2YZyIX1IBh52wyvHES0YqTsmqtCW//KTHyKDTv63ahJHAEduZYAfEetH55xsAahoTthEX
F3Ocg15UuWPe4ak4+6q6CRAmodjErWTziWY18dBRIEHAlvSox9rJacdrCidkixnHGI2C+QQydwaF
OELebVIYYyRvjf6U///WEu/W3tmWIUKo5wJjFS8eC7hsYRadddhnW5BNKNY/kolfNmqpcp8EfyN6
w9uDHQSGboIvDQS8/ui0hS26zMwKoNvcleUSJ6HYY9dKV8eY54kvnCzoE4Nw7kyTdZFHlLeGDasZ
wiV5kM5W/FgxNfsWJFNMB4MPf9Z4NEcozgCzXJaof01BzEYRbIZUOFYKouSNIactYE2ZsVdXxtxb
G/phpQ4ls8FGr5LT2mCycDogRoAgvPYCUVKaxRjFKeYsl4SOw99kBPvpKEBaitrqVU786WMCzUxb
2uV1I3Yy1CzIizC+CIO5Yw/I5e7frwU0pEKLsRFB3e461ZO9lrNkHDKM4C+TEPSLCDWT10jC3zLL
XMGS0V11nM8a1VLkPz/Q4vz5tsX8MLoVJVQsRShpw97DjMEUf7e+gQ3FErO+2PWHBsLl78LnOU4M
WSNTpqNm/q0pPoP4OOe8ipOwT3umBjIpkUUU0uS/6H08rHGLpOLILTNArY53ZpYExEEwhrqqo7Nd
5f9UbwKSozK3eZ6EEjpBkk1y3U7CfiGpgf9z9DUHdHNz/98+Fg+fXtuQFqSZxi4p4gVy2YN6sjHs
Tv1Gl/MYjHRdJRGWCrGCkUV/s3ipiDqaD/olN3v8SyJZw0bkABIyOK+Ypx73kjB0mKqeHAxJRUP2
vOTrl3wZw/7oD5WUOMDu1gY/gtfEKaOhxB6Af2YNeuTYo0v5iuE361IK8LGS9dcSpwTxWL2Ovees
pHJtxiylf+qUG0JDulnXzAcMlJoaW5j3Ps3QJjgpNBPBMMDS8OB57fI8epIckEdSiShG6MqT72s6
bGpKM06+lruFCD43SvmEv5fc84bl/fWIzMcecAj69PBAFsYl6OcZevc+8msBBsgUJmilcyouOUtS
MjeMD4j/SjmTh5sNI9l+vM1GnlBMwWnkY5edUSULntOIcjJbZOTAGlG+eeGwipoHK1DlzQy53olX
izjnCpYQ/ztDd2RhISFni7eZk7ZC+ISCgMuObtKWGgzX7IDgTZlaaS3u5EgEBOI1oqvBu2eefl1T
hmkonIVrquzSDvc+cRUR9EUWr0CniKmaRANXX+OeF9/52QCTT9ph0FNmGo59gRFlX/3oev9mSb7k
r70fZJZE7OtAlmecP/n/VC4wgt7PWLsAHkLIMtEfcYhaCo2uhk+AQ+VJ0+OmBBEcJypMuSV7DMZB
7wVX2rGY3LWpibJedFczAlAnwdroizj/OSs3620lmtTQu6otWHTAWVjr2IAZ+dMinfVe0fRrqgY6
6pGwWmM4uFdMSQVn6FQeXwc420gssiymI3auwp/YBYFCoT20feO222xhxA9+rZ++F1VAqtcHQCyZ
uk9OdFfonxd84NYg2+oRI/84pOve1Mx/bzKL11pczYbXA9ShFvitUiRnz6e5BLfCqeDU4WpN8ag3
Neuc+DPlIRMAjC0QVC3XsPMGAK9WAUCX1MHu+pQKltUSjFNNqmqfkOtmHV9Vzfw0OUfegrhBuxH2
0HHf5iVlbF+FjWqt+TjtLX1JofBjG1kOhhCiYZU3koir9gfhmkhCPM/TZ7CB3DKOYlRJ85N2ZfSa
RuQ9/GteOAbyvv92dqAcVU/p8+H/pNtUPByO3RrB853AX6KCPDCLwOjjlv2jFpP7XMQWlluquvI0
1+1lBQp5PybQY4vkCS6fWbrNf1iKqCZSowXJEEG3APocOVfNTSSzid9xwsZemqyCmYczB+c7NV5T
kSg9wCa9llI0VSyQxm8Yzly96jltlLyE6v0UVE7KeuKafOr+L6kvYnKgs85iFutIIS2ywnGS5Vu+
xW5qxMWt6qXkjfTn8d+vG52qhIXkuQN6ehBYjEo6WcCT6w==
`pragma protect end_protected
