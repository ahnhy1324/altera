// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pTc+3qGyF+rxAGLzw4koCYmoLQPEfNnjMv5eGN1rI2QQWMXjat9dATcXBGYsRZv2
i+XS5K3HJg9XZSmpV6mnXGPPl8g2yX0EMuHT9BsgB0nbvp5SQo5oNhj+QKrfF5YW
ovdAsXnu/MEHRL0Q6c9hnXZ92DNzxPCZDriTM6zYIhs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 61984)
y7/JCfSZXTw0IYEjLVJhsJdqBbJmrUX6NxWGe6TEjuYmMNQFG4/MUF1uCvxPcD/K
N0FbXWjzUWEOD5GmQTeqverVI2H9jD43Y1wt01AvEeg1WKFlNaK05AIWcnLj2tSe
eQlozuKekW73OMs79j0grM5HOCLJzMqHdvU29LzPxofaEZQbC3mNh0sbNLctgidM
1HsVloG0OZCrEE4FqbNoHXKIg4ayaG2rPqrEzU2kAdmj+SjuW9H56QiUa1eZEpIn
2CQA3ApU1HJAUc+rg+zDIZksqUzoAkFb3CQgjeh/dklCSZTEvkV/ex/K1ifXemAM
kpH42zcybrdPND23NqJ2K8NpTWMMGRa8FO1wwO9H68xSyfFY5Sgncta5GNJU4+pM
McfXYPDObS2QYJehfYBgFkTtoC1Tn1KWZBLPAJo0VyLItB9EGiQClWJffZVLAB65
/y+x9M82eTnp9BcDPhHANW42qfVF2iPhPvu0PO+5jPNXHbgmjtCY8/+FGQXaBTGT
U1osOgvQTYLKFhJgqAyGC0MAe24hUGUpfDVPbI7MFKAahxJrZTg2LsO+SB7j9/1i
0eAYU/aKr2h5qzVxWnJMVaRug68GyGUWaQ5LFMF1EJh6Pyxq4SD6Ggh8hNtxTlYh
OrbLYjdWBwEh8cyzCOYyAziJ6SlritMsuB5Tbj42yk3a+xYF4KoSUvtUlOko0PdD
tlHNZwBclBELegDgaqY2TJi1JfFLo41uYqNQ01MjD40M/eWHj6pbY2qenk23URhd
vV+zPR7iNWgZmWoWQFV7KaQKUDg2MQTC9erR5tDXI7i0k69GyOsUPWsEXXw22Eeb
zS2haK5LlWqhwyEnfWlDzz+khPE7GBryc/IoJO0nOokUXxA8ukD628OALWQfwWJ/
tfYQIp6DIat1ALwuFsl+cFX3hZ9FdsVoThD/KsBsjuHWlrclndySt+WauGja3uu1
jxWYtodIdTTQUfVHMswpVpokpVTCDxOjM0ont82ggCO6ONg/5qUuapIT5QajSsQX
BV70dARjfey4cww9UwgN3KJ3g7w6gR2jKB+qbF4A32E1hQ53el5bqoHV4qM8GKhn
zUawYNcbxynUaTeI1Fc91GP7fY4CTrKa2djwpf0M/8UHjPKACZU68Kk77RUZGbBi
morKfk3ndScT3E+sEqp6kbKuzRbMz8kNvEK9MaP/GekRAqRFHn5KbPTrSTDZVRkj
A4EuZQcfRgtgxSdyAqNR+RmIrk7+5Yaq+FynqbdnkQvyYGyweAymCFjrS+81YXN9
zwhRtBWULiVre7hoWu82Tutj87GXtuE8Nz32mpHzLJ8tdJuf3Y2kBGoN1Ig0GrSA
XS3+/Qc5B9cO8FWI+HbdSwaTTh1pVoTqX2X9NKIzCUqHm+gGIClsxJ42JV6zMSZt
EyeGuDCs5rsC0gx8tO0Sh4b8KY4waT/gLvvgLmImv+H1byMg/cVoq3IqvO2dq8wX
Mhe+hJ0k1bkuK2hEL4NatyCkAZqXQqRAOoMKWjzL66oJMkTQ+YSMOqtIv4xB+BC8
Y5uzOxWOEkzWlH5h89TVbIulV8uH/7ij+oqs0LkTP8uDrzzIUr9WHAt3l93Gta5x
T0TO1aKBZy4uN77jVuxr7LGr986fXm8sa0KzjBOwgsvNENYzSVl25Qwfk5f6rkdc
ogtuEyPE6pVYuiAfeSxA8dReyIYPjNpHf6PehkvOjkIitH1PxioOQjLFiRxJbGY9
SWKqfdMmMtQgNKNZOlcemvjXm+IUK5URcDVz1J4ZdonfIHN8SDur4ny2QLPoCKgf
EoPAqVlJQWjAj2+RDgAb4gsToh/DmrblL9tLv0kEAobGT6QraBZ8ufIDPyTVaIHp
zz/uFxzZPsxpd7Oek8LyZ2HZrtdBE3MapC8V1vPqfhzYtXaSZpKhvj6jvNhkq/AN
ZCnCTsdxgm6WQydu2BhbAH/8NM1d7B/50D3z6Fdqm6jOuPRUn/R8Sd2U+lPCa3lP
oIEJm8ZPyj5uEolXmk5Lq2swaVuRng+8TBMtH0qF/akXB9/Y9Olglmy6XNuEFxV3
CkCXd6QCDAyM7FN3PsQfF6awIzdLYi/mqR/tMTseHICgMpTIwl/aW2eJHzpfavHq
tLQLaRsYnf2Ghn4Jswz00VzOWVkHuu+8YYc3KmFAXakNRfv14rn+ZNyaP3aMNPlw
Zv5dUtwxJqf+g+0Yhj8itnVDqk4/RqTKMaa6k3OWN12wpd8sHddOPFIf6NnI+754
Ywa/3PlOn1frcDBZixjQtGQmh8mY56te5esUYAF5Lvyo5k7sh2C6xdnZjbrf1mNM
sxj1OYon5WLs/Urm4Flr48G7Ie7ZPyBeVlA80eSJtfQT61fAOzjG+H5FIIRw1eWL
6PPUY8/ncWkPKt39d81No4zDUT+UUKey6/Hp9Cp0cWAgtxg+XTtRg3z4iScsyF1W
aIjNKcSnxPq2xdwNM3Xjb7Fj2s38T0bc5qlQX9Ybhv7fZH32j4ow5OS2XjQzGtno
NLWLQ7qcWwLULsfhCdB2qNe+nxwra3tjYRETZF5okYolljygYZ78PYH+COI2oOPP
fCRH5LRjC0J07bwifTV0Xfuxw+Zif6gtDBgBhaODjbO0U4fRiZJo3DaoAneXcc6k
hlcQKrWO9qxolOjZ/BL/utEn+MaHoVpaEQNzHbv2ymBQ3UhU7e3vDMrwp/5Q9QH8
f2h0V+KFdzwIudqS2OQ15kYuNLQXfpqnvkCK09u1vmSUgmOKC/PV2vwQOUuloGf7
X/aPPfcUmZYN9pzSm1p1oJ6LWFNuXAZVfOqdRh7yDBNvnszD8BEKf9gwzx7chSwA
8gabuKms+q812kLlrisZdLm0+lOkKo3DFXJe9kIo99XGNuaeFiGZcYdcZ+SEKXYq
qkTxj/pMM+s/VFNK8OzwnU+NI7jDjJU4tzcqNnbrecbf+gX61OQ6LFQ1JnHWYHDP
x4JUlyuseorls5ceDowRZgIWz1BtGo3KGi9N0/wUTivIedRhfpwuuZKpiWFSMsNN
DowYEQlZi8frkotZM6GbSAW/LJvz7Y1l8Z5MUaDKIWSDNLihHK5rcWKJTbyJMOtz
3A9Er6ZOc6DQQb0TeTfkkCZsUAYtUAFIDp7pqLmw6ASvj0Ez1MeQOheZZnpsr+QQ
iHkQUYxVE14n9Nv5Zu8o0jQ/TALQhVnsSMbcOE0qNY5LK3+0efUZVYTe0YEbntCK
93HXkDNcDARkqdL8B69OIjXgA1tRz2NKzLDADqw2k5AN+ewUsxZ/fyRBvPuF8vnu
cZyMJ/lj2WaMbUXq9qzTKNRJK6FwCMjptPLc4HJ6nmX4U8N8/OKLj0d1+AAjgjRC
bMD5MtXSxgY5AA1eUGezBlgFia+K2FCQqmk+Xj/GWs8WRFev8Y6m2tlCbg5liFHT
Y+lJyleDRkrj87nzCUEi6fNmpH2imIqZcB4LoYjwHQeF5qEpKp5aCVlhBxeMNBY4
JMhi9g/YsqHF67ZgCAEffwlCZasstXli74sX74Kg4UGTGj+/kX9IuPGVq5a91+Pw
JRAhyaBReciAmdQ+Nk43Ly3J/nJOvhvjPzQjm7j/xdufrDZc+zLi8AdXBNE0ZZjy
Xplopc5rTO0Pzguo8tG+gQGFk+2POU55FrU8yFsgFRRlbT1f9X0f55vJZPRceq53
SoQ7o9SWEs+ISm3lgydNkb4H6oB/PuBcwv99ito8LC0rAljHxCstsVN8dGQoCJ5B
8LkI9LnMZHaHjBYMptElHTGzXY/ItkF39d3YaUB4QS2xs2le/bdFtFZxqOIOlZYg
C0bI96wa5aP1+zGNPaoC1oSjyBTKW6pUmZXLfIJbGVpxPqOB7ihGYG9y/OK6FNVz
QtxzzFQtPSdDaCxpej7aI2f7pxTABbWLCz5IjykZdrdLowGuAWVTU0a9pG48y8zg
0AFMHg9tsL37DAwAKAZhjvZhzyOFwlPXoNCjlKuEMSpNv70QdWvEdFi5lumX3L/U
QRQADgaqdoEYEwjqBwbJmeElFcsQit4e+e59yizZ8uRQd1QMOfWEwHvJMli8sSNd
ykYGg0cW0PVCPs2zFN+G0BGu0wj5DmdCWzODQogJBNVb4QniuPeIk5n08RjqjkZa
Vr5vesVTnTtJJ6r/srreeZHcgGjl6pCOggeX+RfKfzembunXcnos03HqJ7udEcTO
rHJm9HvcvbFHjyfZDaFAesydRiv/NHvGavPl0kPXE5FegZAmOIz1q/yhvnkieFDA
Ubbx6QunntS59IAUM4OAFUm55ozR61w//c320IhkTj4sDyBjcPmLAkiJSq/0j11z
ZGQ2vBO1jbveBf7nE9RY+/NTXfseiOPX8MkTrATE7kP2eY/9KvgwASRMw6MqlPWH
5w5dCs8MQ2B9WQlZZ2Wf5ImZYddfjBoiEUDqlFRn5pXGqB/Gvjr28qqh2F0DNFzK
v8gmY13k3Ytd5fY65mtE8ClfUhZ7zDHHlB8g3JcOzrjpQq+js9JAh5TRGTX+XLaA
oeW+GdZBpiWkXkr8jzaXVz31arpy0P3sSD8D6OOqffjxG+Xng6NgFDdRKmFir/CJ
7LYk1rqqnGthUImGuWuqzW+1UjVawzxXdEuNcKSbT9gY8cXgxIlDyktpb/VR8xeb
h61sH+hSspsJohfyhorgS4RFw2BLQZK7fedEnNmjrU+GETU8APd+fjaC5+QsUqHt
iHICXpKI1YcqKdooNc1mbbFfMaQwh+H4YjgjxGdFiLvEeRxGB5R3SUQoEJIT7xHR
+uCz1O77TIrGUxvHwgaRr1wTAeFA0GMT1WlOA65622kkiC+ETcPwfAzGBR3htlkX
xpdHYi7Nk/TD+sWoamTVUvgpW16NhVDyObshFYm9Iuh0qUy9FW9vmNVNxHXSsz3m
IUvaCUdWqt/5fMDjcMbTWtbnL3WOedeew4wBYB/d5pnCd1EZJIGSw4ymFgcuw2eo
3xaMVHhwarJ9/RQgudH9U3UEm3ODL9E1ccx520fq/ptj+38qBR7xtsa051SFohGj
N7SPbx2wRdGm6oM6YUf5RzBEO0Ef6zDLg5oANZdI82db74h4G0tLKVioOxfipu8U
7G96MfwbHKzPqCWGNt6uc/9ZUc1Src5Be1ODlySWWS24Q7CzLVMlFihDAlaNpS77
4sIujnBjoMz/BorSD7vfNVOSnpgGuKOSUgVN82Umrf0u3AnE0OW+YuUaI8h0oZRC
GBVwCqnJ2GLLgBR3aNl6la1da9hVliSiXI0i6tpT8qf0Ax5Ce2dXvfvsjtQozLUh
BaAZ/IiQNBtazwG/Eai2RKXV4A0wYyRXm+O9tzUQWipKgbOXE5vlHnde5b28j5j8
ds2oN/+vrWKScF48YQuIjOMHzklPvZc+XsOneYSMSy+094jUjNpRSJ98Fv/ghlPA
8JK6I3/RXAG1l7b6bfMJhPovwUm/RCOTc8LGNCPbIP+7+1exR/7R5Sv9Mu13geNx
NqiQsLGe2z09tPGmv7l9VtTGnC9gbJlQhPzorPdLlC3ni5igXQcktFH5vu1oy/99
QTkn2D3uZUuMjWYw/MjQ5IDD7iySoBKcxK1wL3Z2H7HN7DVwrLygeMHm12Flctel
QFjqt7gFW+MTf2J+xTIrQimAPSel+n00LBdN/kRyllXdAU6s71VhYwq1lvt2UQr3
Tk2QFnoOICtXccn0v/KeHPEIyMN/VEdvqdII8S7GYCdfa4UleKsVlkt091Z+3Wbh
runTEsT/NVNKoe3YS4FaykcusfnF4XRyLkxVsvA8l0TL1Su2Y2jrGHM74VN6MdNW
HZMHmaGhxlZI7O8r8kawTkfp+S85n+R+1i0SbWo5gpt3KbMUtTf7FS289KlGc2jx
G0wlWv9m+nttU6e59J2TeWsejMPVgFD/7wZqWk7e8VUCMijuWSLyAvXMVovPa0YM
2BW4M2IpfgRBAHzVD772N9n94vB9jAFKaLyQm7+m1sCE4+nRTccwrjIIO4o6+ePf
PFvTSac7b8XA5kw4Ww2scNHqWdzZ/xWEBnK8XtjykW8MJCNIHA05FwiJyriCGEx4
yxZwGCjTCx2DJZmZfxfslT+XFr4NXCWr4TzadZYJI+UPGZzk/KNKLVI0UtMe7s6w
EVBEB0Y/92aocTCn6BgPmlW3+TYWEUK2Nasc3omHrsaDAlud1vfSt0vnAU3iUjmK
DPkKsq8Mw29K6xBQRhvZ5+Dd0FOu/3OUEdBarv4uFaXBYM7RWQRRmoHsm07VgKtZ
LmUsfHq3MzaGSOgrqH6mGpFm9tbU2utJarc09nitUukLsl6UcWR3Y1n5PFqCy7Jk
o+cuN7bPkC7J0bpDmf6QsL5DfBXVIZX+uR9JKM3RTWhbXVaEDT8VQU0i0HAGbYNh
ySXqWo7aTCKe2gOMoLtnbRkur3dmOnBVYbKzzP9KW05sxXZYTKG40AgHVaODljBa
/0x3Wrciwg+3WJ6dZqKYqwT+LgyNsE7Q7rQdW2KgA2WfxUcVR5290cPP1tSqGVjX
xBz/sxtg8eiRzAIqWqTymNrLec81+NOW7sLeUnJeu99lcrWRbqDXu4I5IjJ9A9Ek
VTByLE7QS921Yh6aAphCc9DQ1oPXRn41zDxYqH5xANgHVTKXBwtMh5o7hvNLhsa0
sD4wGJmS0NnQ+/faGHd8RZhY0BYxRRXqporAUoPDl8TVnF70rc2h52qJLY+aK2Uo
DxqYZD+z7i5xBHL1tL50WMSW8uAs5kWp417OcdW3CPRoLPkGl+80dLxser9qEpMo
O5U+8R5CwyMg4fcZq8wKXNGVl2CaK0ztlLT8TJfzo/ryh4hltkVx1BO+wlXdHnSz
rnZ0/h4558g7eb4iwl7z4S9jVuN+9PuLzzDfkEBdSlWwxR8sWMd9RV1pBJa4Q6/n
eqeKxrpelVguHzQhZXrYn3RGPexPDCrRdF2n2hN2rwOVlZKw4n8VgSn440DkafB0
UkxfTENJ48/0TvHBbYsg7VDN3JGi9F67XNuZXvPl1upPsj1XwvJH8Kk5lwu5Kv1C
2Unz/2U7/i/tVKPFX6MVcILDNp3r7RKxpt1gDTN5bUq82DkwiSJcHIP34Ihj95T7
MhtvjyuKB9BgJKDEWzvjLo2TYcQ0QCcmrmBguqc4bV+JuW9XKURz+9ls1vGES8c2
JlMFs5fqbbfFaa9frf3hLjwlkW7rOy8WLFxFAnarcwzIrbsE4rmqWQgezWSsxmoa
vJ/E+cnIGI5zlaDZVCKKkHwOznbWmlOQmzhTzgxPtIy5huRJm7MdJGb8EfbLS1/3
hHUkbDB4QPEFrsDh3ax9u/tW4SKLAwr9vU09G/DnFFQFmO4EI2hI6kBTiyMFoizh
T6iZzB8VGlkqZSLtF7rrDbmzFBYjD7Q/f8vryjjccEpXFNxKYgff6Tt+fdYdjGpO
NmQy+5wm/f9v3BTswOTe7JoDvZj24/3DgcNpjfk0LDXHKOIP1EAX37EQVpt9W2kr
ijk4zmeglvz1xLaYjwkmdLiiahP4/qfqJHHoYL42w5W34a8uA9b+IDTxO3C286VB
r9EV2lGp4waTa68L/JLc/notvjVBsx8CZi+i3OEs80ij6j1dBl3niV7yYPFrzAvc
mTLRrt67NctE6Icdu/mrO7K6PSNTUL3ZqOzlqUDbh4MHnQatZXiwCbcDSoclzvUm
o4SLdl7OKzhTzB8UEdc9gzTE7ug68MaKfnpN9VKaqZbOypdDFYz3XA5/u/1Z7RV/
gutEDrVProfEVFEHkIivHAgeQIA4vUw+6ehSypjontq8gMhcOzqfFWjEcBktj/os
u7QyFd/YVA0N7/MrdO0vwh7H3JvGWQ4e1I+RvFIuxPBFgLA8wLDBegKcjRuYaSHe
C39mh+BKVXl9FFzsToljexm98vmSeAZ0MuV4BzDF0d4h+J1jUE3zq5vGJR6qwBY6
eLTyq54e+FV6r6SP6Fc+KOte9jhk1pCx3JBxHe5P52+b8Gna59EJJE8gkCjGicNx
1VOz5TrHMd3dUxKbuZM61eRnSrFk8uAwBsO2fTM3lPrLbjUOecf9+tVGbxAFRCOl
dOHM5EnJRFB6F2EWdxnooRXW50279IA6CmYXIuN34kaeBZ6dQRaH02kcoxVCzBI0
jUAgsQl8cWpYfOwxewzg9xC9j+2usDJBeKCOfbdKpYkGkO9hkx+zn7CqoLGy4JC+
aWPPJHUgFIX3HP+ME5bFFHFA80P3+ZATl4SNiV90DLX6S/l93bAtBQ++5FXw/Wzs
yS7tbH5f5X3KtihvtP3bL7Mmib7usdObdSoXKsnGykrsW9xyxPZ4j+ODdYZMpTzS
n/24US0jcg20JEvq9MpT5xv50ZpeVfPfYYH87BrWSATHKcibwfPx92Q9gJtzecFW
vhWMl45i+dRg2iVJPPr6pAIaeMSzQtZ3GVSU9RVCe6eeGptl+4Z6eB3yG44Bz+3v
VIIlohKlFYSqD5xzyXBl7duei1RYQgetNsqm1OBwW22oY+u+5khisWmeZzu8lbfk
yqNbyBThtp3Kls4qYUSCHhfKT//bMCXn7dy5jfqP6wcjqJUgzRCiC1V/uiaKHN/K
86pu9drw/nnHe+pPKp/3qPYkgZ+aQ/tjM7SJjQZNEfXsGECPSlAP10DQopbIOixB
QWSDp45nweZL6hu/VtXeVbgSICxfNBuaQBB7s56CtFoYsRwO4OGq/kjiLOc09b85
IpEvXhzuEK4IVK8SlJOWZKyxLAOLw9L7wS6Uc3x/8K0WzszSpf8VGZzV59OfqKOU
/wDXJDNWyRuz6f3KYOCM4j75KZUy9ncOdEafzc0SC+38S4il/pD8xK4oTfzpEGl1
OQYd8Lcb04/4p0Up9eFyVVr8QQik4aoAAVpt308nRnP8pQvK8hTBqmAZ1z94c3z/
bzuB+W6XqDWjgQ9PVZgnwpUJf0iHfqIi5zRBJDsVIOdeatbw445MRxLLN4r87Xak
NGf5qHAkiItGoOJmFwDgpgsb0rzdm9A3eDnEjZezwQIH5NqI9mg3DoG7FyooTn5+
WWuPfxpeAnmhiOVl7M6xilIdkf1nT9xwdCtDcanhI+VL0VSDGll5lj9m+PfM91rk
39N+7T/tAFU790HpGOaRLIQyYWW3Zh9M/Tg9NB5NgDX3CBhcH4mlNcjTQA8Ol9EX
Wr+V6LefSgqxGmVZKHTYuqE9WXzeEm644lSZRfFvWR/2IHdIpCoLB7dFpCsI4ZEb
Ah+G0OaN1pQte9+iHRD/VFZACUZ8ucEcAOcKTcgpGKG2cPQmSyAdkdAcyvnHTNOe
jHd5T3l8WOEfexVefzkodmegZe9XnTDNzcjiE4KlGFt9BmPw/uxtSZo+KRc9796t
mcgHJHVZu6pbEx5yUOxmMUboEkPgzCNZaH5aQv5ekKcPBzghhpovERrxmvDnp4ft
mYKrSIEN/rnTeJAF7gFhjHd3ixpsrMpEKwkbNV8OSuNsGfIiQShx2XwKlyYLWbqw
FNv4LL9Lp4Jx+Am2Em+qBEGxj/Acfe67kIYwE7VtHIdC9CACGipv7Nt/df2ibMjG
rkshK57dodM9fGvJ1uiqKvkCNik938J/3IMHDd5MmczEg0D6kFeNIFOXy/4S5/L4
VVlz93+6a4eXgxz3fFLldnZVZDclJ8vFQSHW6LJob48I022rJY1D2cpznIZPAzvJ
+uzvFncDC8nkIRajvs0WpLk7e3jcmZsKPnbI1DE2BBXUF3pG2Qp8lZbDhThn9zeD
iVCo7vmq5d+2K351iodCYgejGRy/St3pI1QlHx3SGs2WtPnxZkDQ8tgd5s9QKFx/
iEiUsf22HjfR9e8D+Opn6yyjRQVOiVBn/6QNzesxjDxY1a5mFPuaIXSLSOHar65s
10N3pj5oK1oCPuwesw4urcH2cTIzSQD43IDvZjzvcmR8Z5svwPrcvZV+Md4oopvD
Xf/sy3/faOL+Iwawa8zzPUGN1labSemRWRSA3qvLe/KbPeV58XN/VEe/jp1+F6H7
LPmGaCv00ciP1v/dJkh6JkSTJKDx8amNZFb+L6oVjoxxwleGBTL/g55W6C7nwD0D
gC5OoPm5KUM7fs84+SD4GpoO4Jw2tm0iguY4QXbRw06X+SbNbjPvCz3NaVGKr0ja
QSeUkPWrFOeujqDk7Yls7zY93+FGdAXW5Sp64QnR38kT4xlsLrVU6RkmxtHmW9kW
wPghlTI9RA6EWZvsO8y8mG2PzTMClTLIKuo2BCZwcwFZZCW/AYfgXV38BgOA5a+0
yoy/i3Yiz0rMR/ls9Zy3SYlLmuGJ8vMLyypMJb5hxK/LZ1gX6FbqdyiYFFVH7ESL
yH8FVnHe5Fj0UhTm2yct7Y01Makt/mJdqrwCoxyUGzc51t5ZozAigr6fiUiEU3yd
rE3YhGTzM4ld8qCqEpLxGjJz+VChc/1TpnRAXroQBRR06dZ+NefKZDKHH90OnfFN
KGnu7hDdDYjZEIn2kTqXByNEd0cZ1hKJL4SFYlSMZKjua8Ua+Xq0BkCng5pDb2hP
OPXiy4kmUF9QCW0OY4zA4L0872GY8+r1JUqgTDyy5iWZ1AyJJpKzjvrxXuXGNX9b
uMqIHZttRHWdDX3KhCd4KKeZ1lETfD9v4kuWQ7m3wy9FLNMRHRxc2y/g7j8Pv0iv
Tnuo2jQorgmysPFQ8dRxC89gZ5aLTVA0pOLs0Sg18ShIt2EybvXrQIgP52igGv+U
hpovIVg6k114sGTT8q8fil0lORsw8bOWS//SGllAF4Vh7a0zyPhNJqHawzJsbi8W
70poACYRrI6RmP7mMEARSKhMEBDTVnLRoFKDPaXBfo4TNxgd8TKZ+ENCctJtorsm
cu8gVOV0N6BAhempiQC/z7L7c8/1q6zm9OEq2xKJq2ltZ8hAihdWdrXtHaQ+wa/Y
Hl+p9Jv3eQpqvUtINblJ59JN8GNGXpA8a/euK/r9CKr78mVtD7NranpTzuIu7GCy
lh2ub3Ln4oBB8+iprzMgtRjTbhv/1Zq9Qrc70MfEmwb+20PYwFFTjzwcLTJ7i4+K
pFILKBekygxRrHFtlW+8Hgrnlifb+4M0o5apyoHi6sMGKZ/bqYWvVSoIdZXYoRf2
qUq4P7Mt7UTnCmf+A0r1ukNHQIa+lrbo+fy63LYM5muWWd3dFNL1jnjStHsWU7cL
dCszcdC6IbtZAvmhpdhLtw90YbkHgZlIwzyMMbTgvVK/hfmDR2AY1CijNFOLVuga
WgGFR0H1KWjl+gZg0ePSR6xQ2ASWs4UOXnRrBYAmsEPtgT/dyCr0rabB2kwWbJSr
A/2J1v2hFiwwJ1C4zGj4lC0qcHqscB1LHcic+33ODriv2coSOu/8E7GDfFGpNSxn
f9oT4k0tma68ij6YM9BJy3pcX7CNOmMjRs4LgU6Z58dOb/llk2QazAwYdfD+f6ur
CExg16QI1+d0yR4jZAV7M5AE/SulLQ5NQ8JmLKE9wfJmiBi8K2LwIN6j3hOaekF7
Ko5J3ChEVYM6JqumQsHHBM5m2NQGLAepAA0w0BNlg2rp9c74v5wuxjJ9Re4XLerY
x4NXuWQAW9FcZD3wjtiQFdg805xXjS6EpW6ydbVrIYhie1aU6bQd+rlhMFIskvfn
syQ+VQRofWe0hPpwhEDORxG6hlMIM9+p056BmZXUaOAljlHKp7+61eO9dteLLoSZ
7Bp4aA0l+k4jpIRsmL5e6IHLZ1DxLW2bGmOKy5quk8Gp6+ZaaMI4tyC7DKommbc5
+nsdSUGXNsoRjQdbhintPJ0uzu8bkClAqQpkL/327G4DdZEYCi9toaGRPySiUlc9
rph4ntV9aInqWQtNJNqhVwak78ANizWcEshENkI2LK+j3a8lVnUY8Dttx2fqRuQ0
qYoSI+SePgMfqYiwJI3iMNjc0w65O7+W+hXf5yZGyFGGb91J+huGMGd2WEetacaz
IvrWG8r2Z5snA5yeCbIR5b4hcDeOD0jvlSOiaer9NWg4spWlVvJnkUJ2V6oPtxpg
ekGS8CHVza+B+YWYE4kawn2cT3BGfIIkZvCI2qZqF4XaertiXYDzq1xny1qmcbPd
nU0ce61EqREPdXBCrWGmlgPW5XjABxgCpqZmpUo3WkJ0YOWlmpGS3Z0AnMV4EI7r
4iqgV0/CO89pwpFURiwFVjMu7aqR3coDdeZ0/JaTd8hW9XKiJKG8AqT0T3YCsNiu
p6ILEwjaWBph8EdlPOK91UZhfN1YBPd7s7ZwubeIlHMEM5TysZXhxeH4i1dSc8Sk
WuKmAKWjWLX1ZLijZjFk99eyPO+8j6LdbQpjX6v5VOcYzwNz+TwKBZ8LMrRGSFZr
XIyHhQt2wJTP/PT5waEy3sFW6UYpOJkvBwQjYDEaLR3KU2FM1R4fr0NhIBylmd+x
7ry0/pcQc/8pwNecAmo/qb7zvihxDOFzrefOj4tEgrqku9Ny2ASr976regdWo+gE
A9almiergsac+YR/gdUxEmH0jo0nf8x7ginRYlk31G/5xs9zPszewrAMvuTKObWa
QGwNnFubzC+yIwsLU9Td8pgTyzYe8ZuyEQWK4gnfZvY5Jm89nOAW42I5BOvljuHk
TnBfN1zLfiAuHqAPwX/gm/lvoA2o8DWE3bIDZv1+gWB530q12wsuFsyhE0Iq0OUc
TgaSIeMhPTv8MG1+xFJEQniYewlv/XsCct1oUqGnF355dguXnHVKz2f0iOVYdrjv
1hvNTTojuS1Sn2k8DVhu6JiVLQdn1NgVKMlDfvvG1Fm+dQ5f9mAB44jas7hxI6hN
jhdE0hOk2jso1HClq+QUYJXguxjm3WytPbuFFMZ0e60xxtN+CjNbF4iZEB2Vmg1i
yypsgM5o7sjcppuWDC+zhAC9GKCBCI52veD459C7YCIGncgjs6XUNn5XqZgCk9En
xTFaqFbsZNXb32pJ98L+LCMLgJtnLJij7VWNJth088jvZP6FezezZIC1HTuFtIyT
As2kgLIAZaJGNzqRfHOFAnTmLfj7i1h8aM8D7PvGXchwZLSgUjBHSkjEEhgPbfam
ltl7xeQIOkswjLf/zPQigia5EnqIjcMN9kvktrWP3MTsaVRYWc7rA+xx5uW6jO3j
+9gYRALRC3jwSue6Hmu/bDTc4+V269VPMzsSPum8IdxiKLdo0Y0fPLnz9vdhgctx
D0PIv7fBxQBPX3X2QEkKSlxo5EqXQGCJ8A6hRffACTQNmv400klSNCm9ED+0yP2p
zunLNS3kI4lyFt9w4ubNlKi6BlQBLEwQscP5JbKR1UdJa1bHZyLLWmiu+oJ4/B+k
KRQenKJyWkPA5JPev5S3KJeJ8CAGqrvWV9EFw/qudWsmQvDzkIeIwYRFjYDgKk4O
DlkSDQdOagc7OhA5x/RnTt1hlMN3GamYVBCSYm0KPN3LhPULjrDhfenJPsXNkqHe
mgI+EFzUBRuokhYz8aQVjQH7+Gs5E/90NWx+WjwNJddtM2wnti/QW0V1EfSzebXf
QKjUGi3HaOqOc5vko8kTUGYzciUnV/MIHLaDSr0yTtA8NPhq9Oa8iw5dv/n7VEaD
ubBZsF+5oP/+pId0ts9wQ4wRL7aoAhltJk3N+0Rn7ysZyAOGO3PSSq8lzbaL7PLE
VQoOiUUyEPFCQoEGyFwqscU6LCquhGXsrNqXWDwPMqhjZ9T/aoHjfjh8sjScYdLm
xH+OkelFcL/aUSoKG92LB+BXO0F50yYwbZaH1lH9y6WzNhqWsU148TY8yLBAu4W3
XoJp5nJWppKs//W9xt8ym4jucA/c7yW4M/Zk4DJlSpIwl6KcEdtLG60bsHgHXZ1R
AY1UX8Ipzwrkv9LO/7o+eA9RKBZabyus9JI1daWeQTwBQyHffHyoktPCdJPDJ0rh
BOj0ilpofK1udhO6DLBZVByYm0uaoYLYNHGZx9/EXv52m2WnzO8sSlZ+sAMliinm
mR6DNr5u5jPZUn+OjcsV/qbT6W5VfPbK+M+E5lcDXh9MY11sxqzY9E9rjWFJKgBO
dT2naT8sFHH5i3i/856lSF7Ltq6jCNBm8TW/TOvSezHyaGHNNf/wiINc9GpD46ph
fUcWF/12rRA+D3DaMa1ungo51moSbzcg1xe0NnkePoC3oyBb3YlpOvOkY5DNHzMU
e9JeuuU6yG2zvBhV4xNyMr2WxAh2XMjHDHnG435uWd31VjqYIbxCIFGkTnDC5RlH
vIbXCbzKMmi/IIM2NX+XpBNwZNE0SUtPHw8dVVVZyhkKa2yBNx+x5hxRni0dULrV
xFbMVyx5teJDFHimwBaGe0Wdc5sSCDW91n034txPl+H5WCK086bAPSlZKrlFTJKg
wzC/VCyvlo8/ET2R1sWh6Ef0j57tskwB+iWwRuY0cy7sjXVU0UeBWM03Um5xqorv
q66eT8GoswRV6SCwdIQPzclsDBlxvABc88D26psoFvs/dfEWAN4Syu0pK81nv18w
v6C1itK+Xah8M4O30p/IUMk8qBmcvLy/b+Lp31gDZYBDYfRxvOeXaFnP7vzJFQcf
hoBn+4GFwrSOwrzev38e0NcigvI0lDFEKO/fm/1eh8PCb2Rg5FlpixJjenah8XPr
kdjdw2ou8Xe+sgaUjDVpy7eWTZrbV0se+fQCT37jmevTBoOyrKrRUMv8jOpCzIXt
eyeP5SOKt8gJLwek8Si6iQu+JTVvRj8zakdhYHhJjH9CNAXK81IjTDU5kJJfzcPn
wKyDmqn3AMsO04NWL0vRckY5YehgM4/3u9iBlNYbnwJfEM+lG/JTaZ0JPI+vPd0V
W63lz3nWAjK7z3tYMJ64G916I/jIjAtcLPKf6XHlwZfRmn8vPwpXGzTcVW6aJ1ve
XDYDl7TKWBouAW1cGVq1iNO7BBomLSi3stGSerxibT7ATkv6dhHhWdzUrX16BmyZ
MlyaOKUbgOmLTVpebJ9lc5JsfxOp/f5dC3xdeTpfEL/KIS0GgHGLp8yUnXE8waaE
qvYUBJ4nbW7kmjLRrFoWHVB3RvioMWiPpa0Vk7o4GF0FTBTyzvcZpUSxEcjYXs3l
He+MzLQ0KL+Y5wopwvq2ecw9OdVvSaVdQ9VIiEUKEQBigvtIQEPI19aWlwDPmb8j
Fv9nKiqtsSVxmylI6IZsLOTlykrAWLWtBofHWUiJJpcaStV60fzX/Ubu8v8zxyFP
HSht2Lh7gb8Ap21IWARx8vsMteS1DfPIwlb/eYCp5yjt6oy2sU7L7mrM2G5ww94e
at7IIjYc3i3+1kApxiRrALZ8S6bTgMOIGZFp0ozm+vNTYYmV3tOlYDcxV2rrmW/M
ISKyEK9RhP6HS6rodDJuzgJCy8zjjMeL1GFa0rdsDFkDquzzyTQCzy2FfIJa89MQ
RkQW2ukJnO8aV5+grq6Fs1Wh2YNdAb1Cb5vJxy6O9JqN/hl5U9JCwj7CupU/OtBY
snRawdw3/NsrVWwcRprkE3vaIvvtbebFpHRmo/XRL+igWH+SGqoX+ZKNE4Hg68Vq
TPw18E//HicHHxSbFj0cfoWlDJi0o4UhVY2OwjPdI0HPYwtvkiLRGPbTf4M6e0Rl
gS8v3qX3szlsRSIYYScHWBOfAMjDYtpkMsedtJsT92IkXbyZudQVCVkmIEHj6dBo
SVNOyuZd1Z8ZABSddp4/oDFZOCnw4QPpT+UhkCbEKJEnEnOQtAIL3cjTqFiCwzUV
cpsUu8D5AL5uQS6aSNkYv9zhO7EOYxKtqZNV+fEcSNTxfOCnxCToyrxp0kIbAsY8
b9mD40Ipks4wCYUNoXJPBugSFwmeh6LA4jMPaMDihU6JzN2bv+CHBz/+/c2jIdt6
FxmKl1VUh1LEkHgcLNYZQiunPAn0ohTFiQx50B/hl120/gJXJACZiiwXqhM32NsP
ZzbqZBVZL3P9Ek0W8EB3ZCtGfZiWguVYnZzQqcfjoCqkng1Q+7JHQI5Rmh+ewaQy
4YPCifHqRJkfbAfZrEFuGJsirp9S9q3WNXE07E1oQitGbS337BCupUZtEXvrDdS4
ncNyXB0gXSheQCMDShQJLadZD9xx06etq2BvzqSvp9mpQ9/vUJ/Z7ih/c3yL8TMm
2bMIgvNuNcY/MXHrmB1R8Dmkor9tol+epKMCHuYXLBVZQWGHR9fY5o4oTKb2PL+t
XcK+TrQLrmW9MR4QJ67lDe0dOl4uWK47yx8TbtzxzOpr5keO3lOkCWRRkydwvW0c
4wnK0P1GVhnAqL8lwIwls39cpgDzf1H8BDRV0LyW2pQszMf9DOlLiPctYwei/RtL
I74mEj2xLSOE8IbWtv0imkjZb16Bfz9Fds5Gax73jM3yME/Ljy/O7zd0IeZWoUnX
Hhx62PibBePrl0Bq8XJYlTGnOiHLzY3kaQbj82ebOpm5vxO+y9rOSJOuAWrz0Gje
iVpEfjSnpizSaYIT+h9zHIWRH4N1+et/pcV5kN/owRvUNyQtnsVUAZ494jTQDbMr
mTE82wSxwB5zYQ0ptkytvqAecv4ULvnFW+I3qUwM2jdrDh5IsDILofqS3Y82I3uG
Cg6XeJDvLVoDqYR4XdzEGyrjG4Ma4g2XNXkCYGSObevUsUaz5OtO5PY7X/BX2KLQ
0yDTpQBNqcwwrB2fJUMxF48hHU8UGn/LMPIdDqRNK29mtrZ8WT+93iG2rK5yRNX3
IWQu96fzUjbSjsJY8gxuFcDt16/ZB9lQAXeIQtS8SCxPNKFNz5ay8b/l0IG7waM6
8nRIOsOjYIL/cZ2MT4aPtcvqtXaeTNo9f8IZlIh0v+HopiZp/sXUJM7YLseY5Ynp
LXukJ/avk7P4pQ1mksf5XlsLHhEAWOhpet+yZH09uUEYn1jN0tgl9AKrsoyFv85W
RtzrPXpx0uBVJF6QYbU10AHOFOG3xSy/UEnN/YNTMMlLEyF0TeQiITLmCsPAQA/P
Gg/xPDOMSGloFC3zbFwhIxIoIknApFEvaENterXUbW9zUP/m7gQOf2d/0XFxP30j
HW1nX++TToIztQddGelE3y78zq0TPr9LlILF8JV01agfyS1T05V10lcaR3MudBpz
FiA5Et3KDI/pMzciEPCvidQLF8OZkUzmN8A6SQFC616xl9UO5Lv6xVCEXYnTB022
mdD55Q7l6sHbRuSnJKRkoo3YbJTRqR1RtExgHj5dgbu2Ez76FXNMarl3FLS7JPua
C+Ppc67UtGBDDPHSasaLHIjkkc9o064AF14BoaTEZi8uS74Xi1euu25pxPRSU9gj
dOuQwM/75lRTk33Vs4CK1qfozwuHwpKlhKIxNfT7LX8jnR9FRaWdQWX9QsZSoaSG
0CdYa6LcKGJpnQ2iIoKAE9jEYpo8EoT6eHeSVBZ0t8HLnipsnpQDfyTmOYm/4v5/
OsqVp3svAAu2s2JOjJ25ok7ZV80eTiBzgsM6UKsnIhxFweBVEciJtfEIJJACsLEr
Ov9kMjXaQGU42CM7HnwRELBcrw9/zUTYjevGCi871wAbRdkcQZtWEkep24IKvV6Z
3/+lrr0hP407Lkt+dvDwBE2oCVnrCAMjAuCXAt8/3cInFNfv7QBcCIU95GDwMOER
cWzmIRlNTXjeOxI8S+hb2033fdHgF60WvlllmKhvug7mwsv1bYpepPr9m5oeyrZE
GAzL/JHDdFk0Qw5oqpVcO+K02bjyIzdoqAvdSWo7UWyd0eYxb61sqZTfCDc3Dlhl
IX3I4tDJf8pmvoVWqiwEUvODPSsQ9AP58FCluSmpy+s9ST7dTa8IQ40Vsahf+xMe
jU6ah1vQRA2UGQrF2af5Hm0nUqtMI/1HEdR1956R2nY+7j9cE3pSjOHIj3dtnSUt
UJkoPYg/3JpxOu2C40siUoRFyiX6lmAXtaHxRHlC2oNw17TPPlNfRJbxBUU6IDtb
Leb6tqZqqQi6u2RpNDspCP3kmJ48ITM4AqpJ9P7DllRzR7H00CfW0yi34l0LMtNR
XQlWsOvmzepij1l3WbTIKN8Xi0iIGoYFB1+IO+1SyO+6ni4TR/cZKwX+wC+dGvGD
dDFSEeHgBkNfCokPpkz/eJGX+nwAYZciP8a1xkTFwfbssc6VRk3C8KlPtPsHFAAp
XItwZt5+NNInd8gsFWoSbg4Z3xtnO5/UJbf1+EFSZoFUv91N8V2wrJQPgGguh0Wv
QxMvju+k7s25NCWFpIl3hSF6B5AiSyDjERO4qkH5mxbY9qG8kenMM7jPtR6qFBjy
Bg+6T4A0xwao3KP4A2IZ7p2V/y7vHKG02iVXCFO+nV2mnPwYdim4GNeAIxqhD70M
l9U2RHVSwmXwY9GBj440sFcsEFB8vew2xJmXxsYQOPE7SURqgqKN9R76XauZpjXE
C8fc7vR4StkPtXxnOs1xf9bkdv0IXPsw9tWmZYtFVdI8O8QbQbFPO5mKGvKeWR7v
lF4RhI/uRaFOBUJY+BH0e/2IKTM/Ygita/XxdJJSMTO8GbxuqxWL67Uz8N0KVvpv
i8i6531TgrKudSLotZb16xfyfQtiIiMeL2wj3mRCM2HiBseT3e+qZqjb+vsGVkM1
se/SDZjOSWMu9/6GcOEtl8vZ3wnfUNEht2wPeptR2zWdLhf/myaaoWrRlXOiMG0G
+jrVFcjBknglB+RDNjKnL4KfOPJOb/+duyXoVfBCR120iGg+yPKarPOKzHbR7+Rk
D/fk1oPynnPYwHGCx0ezXWuao38PySr9tnqKMLz827Marxv4onyD3Nf6+xdVX4VX
syZswE59XpAcLCGk1R5rGBYyh7WryH3qS2LNg1RPs2IqduaZf5XVBUN5/UAK4cDs
IwZgNrWyrx17Svyc/AaPXpFb3QLAKUt7vunB0oUijL1BCw6VD/bEEm30f0jBF7Aa
fmJynDm76rJkPzJMC4/SyoZQQS3WhQ7dAo169cUHWaNXSrmPpxs0eZMpd698BdQo
KMG3LFcVLwctUwVtTRcjcU2fOV1V54XWsFL65cYzrAfEA3FdgPLtbHml/QPgFagw
e+8+qPTBLWtia/3jDC5mkMbXDzTg4q9C4HuADsh1wKl5C8cznnuNd8eLiMsQ6GJt
LpBznqCMWOApm2QGQqgWkKvXwg0WR77x00W4IdM6btjB0+WvbiElrORrErtkxBQO
wOsJCO8hw9aeFTkTkAuyeJnFpwVAX2I1z+jAaRvst9FmMu2vNmKq8yztlc2+w1dj
NkeIAp+TCEp7yAyGd0b/Ll4YA99eGFTZYYc9McYc+v3UltTGMaBwlNqomT7JTdmp
SKdB3YpRHrea1N5u8MltqRBv+d0ICv1+nzzk5eYwq//DJD66ejqDUb6DseekrZUP
dJl7uNcM4g33DDvH2O7Th1qRmZNJ49y3R5vHf45nxybzkKbSggj4uUfGcUfuG06A
9iOo6HEDLymMfLbM9ZDPO0VX3gUh8MLIGeKep0QGnxfBNvgOCOTW2sRQShG+S1Wn
YXsrnpJ1yj7hmijjDSR6EpsEzZLzPktX96SpU7kwiHTjL4FZ92Ez02Rnl1SM+TBO
KbFw4DJnmFR84MX5/LWhnDdZOif1Gdf6l0lIrlOzlq/Ccrlz/cbuhsSticlk7XI/
UenYYmhCTXMKdMBnPt3dZUgXxPK1IEH+xA4EnI9XzHzu8rWu+9xjL9sz724r/63a
aB+eelklOMsehmabFNt9OcGcMwJkYBVoUb0teBDAoJYfbw5v/HfW1D+k7I7yZEq6
eD8T+hPNE0SjmLcgiMkeccVhCU0HptMCfr2U84xBFmg5POjQM71N6yR3r2LBmdRz
8a7Q4gg27mvNY/pRJH8ZVqSwWk5c2VdjFBa/gDa442SdIhdkoV+WIA1YzTqBvAKw
nzebboh59dnMXGPzwNMtSsW2akrLUBrmecDehpD+8dQH2gv6VhkgTTJaEKQqh3OC
aPedYV5dbO+/53inAfa47h0axZMy0562v6IY9AoPDexeuSl55M2pGXPnI3hIeBK/
VwSdO8gRk9HCZKmnMkvIesN1E3V4wLlkk7TmcMNJdpT2lICcA6O0fGjhuLcmabYh
Rq4zk1CQO6wnRdgJCsKa/tfb95rDPdDBRwaeqtTgHO88lge1RDs9kTsgkRwuu246
EIfI1H/jasShtvLZpHd/k/Ic6JLN0iW7faat6SjzjR+Wmw/vJsumVlqbMAHO20hE
QgCGzwAuYIud2nXSJ8UQCj3d1ux0Z/yP1HZIOVwA0Bas6iAZ39ynhAdSW9xTTTkm
AkUbvZkPZBhYkhxx8ddz4X3zlSmwmLVxHKESyJMl4GBGzGvF9AOs8L4oFLgpEa9Y
uMajTCIm+M1/o05ChGLZ/2NWFdHRiXMz/imuyDrdxB58YJnnb52Kvjz4HxHCmCzL
AIUfDY9wuL5x771ebusAShMuuv7QXzmbhHoaAXf+zxh48aHMaVKjV5rKi1tQqLl8
L9cwMUtpYPLbROqrqx1o4ZJQ4Y8P3eU/0z3DAbA3m6XtlNzTxN4aGXgBY+wPRnXE
kWyyDLfnjgqLpNpiZo0Bmoc9O5Yfg0fsoIb8/L+kjjLOoeksBnVNIGcdqhw/NqBu
m6H+mXV4L2Im5Gq7xNLg/KtUen6iUMnEp6s4yp0x6Yxpsokv4Ift0q9meOKLwu0O
LA1HdSeuZVQPkq/cqqQ5mig4Zx5YVapU2Da2mwWttgUjRkrbT9yXXRajbDKK8D+r
vPUYDZpTLsTMunZf+7GIuKuqGq9diXyThyNSf9Xf6yIb+vecadQsTwEoJonyMy0c
lMgzpCNQetk3KWbYqUtOFqW5vb7NBPfv47ThXxIdLleCmX9buXnrmw6Uwm7k+e18
KWjsJ84Xo+dDgC8Ht4GYT43bt51CzNdrVbs0MtzvXc+IrSvfjeJierdIhsxkbAKk
4vsngQJcx3o4PIIKF+gJlw7CP/LuOLhYC1yZULLKZ/0NyF7tKlCcVuD5ogJIesVI
trbwFOMZiBePuDCEb2Z/+kP8hRBcpFi+mdyMpGvr4yF1W9goJa7blyhAGliTl8PQ
hxE0fn40o1hFdx18649XaqVSFflhAxKc0Is2fRlpCwnFvd1BGZz90SGBdNH/sQvh
zLg39s/+MCZaX71XSLiT9/+YMAHI58wU0MSlf5LW4tZisZxeCYNwduVcKd5qscK3
kXvEBI0QxZJbyF86srsz2K2v3/J6QcjFjybvXV7NJQWpKogyL1D9WQaA5DlIhYj1
xCravKoX8LtSkM7f/sAljpBuFaSKRVP0GTO20WqieLNTbZMjioz0FRxxhFY/zCb6
XGNgqsrwz8WtGvjPfVEkBO6jdThPzT2Iqfg4s793gAGFxC4UGk39ja6yiKdazqKC
tUkSzfyYvbxrLpyMLyYZMl+Uo78L1OZku9oDWalZU/dAo8SDwUpff3CxN491gO5V
DeZ46iIbNoqM6Ys0gWQ0jQ5six7eCFNXcaIr0/1JzVs8/vxG/kWuuraszQlD3sE4
vodxQ4F2D7BgoX3fbRfBl1/3WyM+UotnAv2aWJ9RdsWaKcxKWZCfPPCo3wJaL3lX
IvMsj5ZC7YwBS1clMxuXgk3GMYT+19gBOLlih/geSWq0LjaX6gqRpt1boqnZy+Fr
Gc4XPmUPdxq+IITSDU3/RopxYCf9lxrTZ3ObkNaRVhqW0QXm3UaieL4SD/z7Mged
icBht2NGU5ub11G8gnLCm+4evnuUU2CkVMJWgjU3STRUyOA0j5GlHVIsBYvWqx44
GzDpjCx8GfKrER7ZylxIU6EDWks3sDJg9YLLxPLquAsAif1fM83hR5oLs4zyKL8B
kxKp4uynfqo9pp6Ubv5S0Y6v+vSgkmoBzoySMd5wTew2FWTEq06+FV5kXo6f9c+M
SxHAoEl+ssp6dvJtUlvQAC2zASHT8AZokVnNpjWjoDkaMsHUPG4aAxffbmr/XVdm
dVqY/xLa3aGhkWQEXJK8W0wBVXylbQTtBn0n8gWP0v6dDBBoQXIw7k++k9H8m7hl
/cfxtIyOjwPp62iCzk8q5htHaAukk+oInzDtCjrXZC+L1HEiWd6RDAQ+7QtZw6gg
ytZBQvvR8JFrDCOF9A0h7K4z2HIBg9e9hUHezbnERyiXmvXE9uouJPQq1WVcF2k8
UrMsEcK2+Fl+UHMmdrzrgxMbYz9oz9KwbHz/xwi231gHbI96+NlRmTpOm+rSeoRJ
siS/4WgPYkDhRVNWNhqGtdEO5WA3TS5jVeIhPxvxpd6xWKQP/6NlaAHfEaooqc4J
5n/p1cQXGuEZa020DWA4x5CFeGI/3UCJiVn+eS1Z2yUymNMb+xGgpKluRwpYLfHp
qCp6NRC8X0qssx3KyCSjCSHEuZcsESFATSzcnRssu1McJ982UfJIFlygRZaQ9cX9
uMGaKVieJhhk8agYt63BBouy28tnYTiGB718CFM4KVj6kVd1qF+kyo3g0JW4VlBW
MUBJTDJkinG4GHKNhJ/bm44tarv3Vquk3bV5OTJ+VkzXjMDvDXMPZJ1xfpfHRVTh
IASdgN/iKJQ5AKem/fCAXv7CsVZXgQNv8Xtq4pq2wlQ0upzdtAVZVXHXBlgSQETw
0tIja4Hp6eCZUmy22bIc+KPc7J/Mzjxa0n/KPuRoFwJuBbMIErVy9+/JxiCQAJdX
/dz3OzS6GR/5VpPuiOOBSokPhs+F1BAL0nodqYpe5USPWcDO4wITd6j1mcxSWzdY
O60luLd6hp7o9nTgIhCmEJhUD4gwYVtN5fiC3/DYHhPXsnVEIZIAChIQJXEA4Ekq
XaeYW5udN6enlWnZql854zfjQy+xSBt3EpzPXeGN16/z8tcNQ0GEvmISKtMceng7
FPE22GbxNesyvQRc+fpHYQYqH95dvWjGfCZrAtoJTs0c9vJ2b0GWHQMv1AAufEp0
1yrDK6M+mdqVs6xax+TKInDFBb+F8Bnxd9MqiXN8LvP8jvw7SkvWoyDzSFbdbcVZ
3TD1AmZXdsH/89YcDwjpfjArejfjG1Og31OKvv6eWXC4LO5MQOQmNdVw9f6gBVjw
XpuNfyN2zbnH+n2bxXxo1qsvfar8IhraqZT3dBHHibp+W9qNAJB2ld6HxW7jZ0Gd
m18Qrwdyo5POP6FxlxeAufnTD/qSoGr/BTka84JQ3gC3wYgL+baMp9j+o8ZofzTM
igN2NnU2Go6hHX+2R7uaAlMB12iI+FLp/yV3wJUsIyPt7Z63vvIDax3hgwceG1vH
zQ27fso1dcm8OJOg5aoiQeDdVYOoiGV6FdFH5AKaFMjO1H0aSazBg+hwshItYxZJ
TSJHQAyrKS9xKF0+7B9aCtW3qHxgAtQg4467VbIC0phXk/3NbUuWk4grsIvBVlbp
cRtmes84AomvX7aCDXexonUn8cT/T3rskeTfau8fOmih4gD4OeKTY5ee3ruIcxcy
kzJ+fL2QFl1upXpvb0Nkf8RQkzB6+L2Gy5ryL6liS+7jA9IcPl7O3yfRVGEChsAN
7HMEI0lmDGGAsI8YjK8rVGZ2JegvYii82i6dbayZrdjRod+zyulaBWMYJyCZ1sn7
RdvZNWqYylP6mvMj39n3/AirEVzTmlKEsYp6vcIuqziIg2dWSXFuLHhQkXg4dM/0
6D7PwkVaIj+xrfDm97Bt1wcKlcIcxdbnPFPIMKkbrAWVQNs5aXCXtZTe4xonDhuJ
aXhUHMQj+lGEd7bt1XW6n1226DFpJbWU0k1a3pN/Q9Eh8RgYiJl4s2wR7Ve9T8VA
thCnWxkF95+1V4u9ZPtcY8Awdp/UPRUa5kGjqtvQEzhysrYYDg/t5/lSXgELIhUB
EjaaDl+zrQJ9UDbieNZhvf/z8gCrCTZ6bJrqjU6kkSLhkVpx2v1TPz1CfW20xX6L
bUwVTT7+eS1r9q5TOPFQLodBte3ty7mln3v3SDcR0bSde6Tm/Ae7RaqS/M7yezwh
jL7h6eLJKpvxaf/WMo2iln8xKV71MkY8zZbncBewp3CXRuw4Wl0AYzp1EUvnNKaS
S+rCoOdzQinxewTVe8D9EtrYWz+wXVuYzy9sAMNZK+viKH41IeVSK+atD1AAl8Ir
cqx1Ec1uay+UMhXjehTMVW6XmHBjdv50IsAOCMZZ35X4ahfh1Xj8dMkcWicK8JJQ
rvXM2xC7vONotwvuPBQHs4vRxAdovqjYTsE7HyZRAygZ7L1JhA5HsPCiSj6WIfZp
3C7FYQpXwvc2vR8bC3GP/ib5poshGvhD1GqWZczI82cBfqatzkNyZi95aPlTiMy4
FZSqKVebJgtdeGxtwXhVGJJ03FqHql4G0ObuUfCSq8y5bGzXnlTa2VSpQ6v4yLhr
0rhfoGx8PwNWuGWBoqXasQq3wozCxyjG28AwE0QuiGvhF14k/ZSEBZVTRgMh2z8N
B6XjVhKQ+mgIe57K7nx5mWtj7bm8fmUrcd9GxlBO8faFyrq7Ft38y73LqhFoVC5i
RfIN/3TDTweyHhvkie7SK+jSJlrABxgXUfsmlzTYhIJxZsJoshn3TG+Z7CG/j8M/
Dw4aQMBGVi0RgJmGy38tQP6x9OLBPjK05OqMX5STLnktSBgX56QVGWAeTVEoUgMQ
lQLwhlK16RepKjxDa4/AYIrIvLFCT+2QIMwiRjtQ39yQ7g9AakCXHjPCVE9ki6fv
kZYPQcH66vjg6c/Yy2qNTcl76kB3Z9qnviGQHBwfYFLdjmv1O4mQY9Ui5wDng2+i
KOMIMrtZowIjx0FqUY5cKs78kvds6a/lG4SYozIgBi5gXal0iK9zrhPzDxJwKgiE
KKWKFizog5tb6lkpnqt1/Vj84XYekhpUAWhfgrBjOKcdDt1vPZj3kbXAJmpCMCmi
WniWqastBELaFSU0eExOqPqgwTQlQWhMZZvSfqhaUaV0jUZfGPfckxRyXtuO/hy5
0oemNDHDbWQL+DB+e8BUu6SwLTIHP6TLeYGWkTDBn2ONy4iCh0b6HQaaz6uxfjdZ
tt4auF1JxS2eETIrDWO7dmNr5hAgKvFoYoN5hh80HOd51+zW49brGG73Z6xuBVix
EFSv9B4PqSoZR5QOC/nb27nQwTZoHtJE0tImcCD9Ym1fQdGmjYUbPNI1CRebdXIQ
+DRJ42SalIhBQGOHyGzxnpf/N5m/7U0Bc8Ce6w1SJ9poMYUdgztjwFvA0MXqJEt8
ZlcyNa5BBfCf79QeoTLVeddBE4jhlIrQcJ5kX7iEzrK1amGtnhpDkuX5xi1DSP/l
5YSQOv4G4ni8gwjAFT/yyeU/FoEsNvMatb2lW6F6sYFxjJghIirtUHYkHR8hZwrL
TMobTvUvWAwlGUj6yfluo70blppaggExq2u0xSP/qirkJj4NnezWC7r5lDC5eCt4
qG1htZEmWBB95Mv6Xh6O1H26+OA/YdzIJk/3aa25geuuhLemrw4d7opnzITCKVKi
TGRQseGkvcEnq+GLvsRSH+kJYjqyie0hUCfC5Mu8R3e9eYkEkdjLkBJ4IGR7MmpT
y4/y+c0R5KunlfdfHHRmul02L5NpAS/ME1gR33GmPOJbnPWw96IkK9gWYHfKDUjQ
LRkZXgKE5MCrrPeNLpikrGm07oq2U1RM6fc9r6x3+keyf9ajG5tTw0QX/jvWReRG
f9k5wl51Kl3iwWpPAG3W0ljg1KUIBw3bqHN0LC7DLgHSC1viep71YiQvx6UaJD50
lNyfFnT5pUH1N8YcUX1EgThQX/rTfHTqSFu1V5jqguXb9fVbvSV9nLkNvBnUXn2v
rSt0YZtK7kOVv+WNdO+4V85eZO9KB1DjzQd2bjFtodZ9jErF4Oh4TC8eGUcwMLvy
C1z0zmH8p8cCR936geVniZvV8G/5Y9SOVHZf05EjKDh5Zc3WLQUo6B0Nvet+jI5x
sbumrf99bV7zttfQt5OPq+pWMYD9P7yWeVVPIjPdS3+8VOhP01PL/VmGLFtT+vGy
7Y0plf2/ygqykQ4x7V2HUWG75SPouoZ//Ss5GAWnS2tnq0EpxWUjofFPcUPUQnn8
tZSr5dVCSeZiL5OircK4BwQfV+//VgBMVL503BnwiyMDRT8flK9zFBIVFqJ9fE6Q
aQ/Pl6oboLb+59A8k2EJBp/HsebHefoNGEEtSV0qsvyvQlKHuYPC4Pyh5gOGE0B9
GA9/wBf8Spktmy6eB4xEbRy1pfsyZBGNsSyA6w3A625CIvH018RX4OTq+HhDjl3D
JwAPd69stYPbPTTvmyvJB6y2lDfrADL5ye29XCQpsfhyaNIG3ss4o87S1F9FHlFd
s6zk8ZeqrVZQqkLY6QtpANCKUBYqKtV2CT9pzP6ZDsJKemF6Q/KLsQOrGJXxf160
3sEi7NGMAPxWkDYeSOvmcwS2GZeQy52Z4DEDsAjBg8fIFp3vAlBRhFsgyvdfL46U
3RX6TlOeawGrwM5wKBJzGGzgC04cX64S8J6zWMLCJA4AXkc4+iTP66TVUqe7X9V0
GJr2e4bt+gDy5iJjgLeuTJSsO2XxBsuFRBof3u3zp6P795z6eQA2eDEuQs9JXIfl
R2Vo+zwzD2UN6oO+g1ReSRrPIxuNe6ntJJyigASWOnobctCatTsgQgFXEDoxSiri
tQRgrcprfsXMBuIawHK7+DvOrjyDNy1MpnpTYKSzAzNtMk2yC42UNubVpAaaT2A8
U3TJggOO5kY+/2fbNVlPV0Ri+YFjCA/hVlQ54AH7ovpoHGe6H1ax/3tm/8cAYHHS
/ABYdP2LscmmZDG5moz5S8yesZCnj/CIkivq2mRBqpGxkcvPhSg4vDsx1un6+TKP
qsxk6aF7qxeDIxFgBonNzrVIbzziOudTcMRZQKTTpp+s9ls70OnhCp7Ou+buyWiU
K9ED/2TfK4WRAGoB/z2YjaejGZvnONwrQJOX7rJXaTE0Fq6oZqJbnqqMB6PXYaa+
h7D8Gaaw4X4l3Xd7a1NsioR8QSd+8yKt/1QEv5hgjB3o+38j1Pe+daXfIYqrSfQs
jj4bee5UV7KjH627aE++BgpxlIHzpCEddn8Hi5jSf6zTd0KIYXNmZRlIu7hhe5YQ
Z1oV/b6erwGgvah2utz9QghEWkzt/09/+UBp7ctwfmQBbRZZxndTy53oIT0DavAN
CrKg4EJ+z5hs+5AbC8lAAY0B5rA30Zzzm+XcHT+S6RcXvvExOWmaULZgoYz7WZ3u
dDlT7GMKJOWERMI/L6fqYZOrRytZSlAqWHaOi7SgpBKOdhaCWMMeENDbQGfG1c9S
QtzI8hGh0mzmqT6BpwRxo727sKL/jUVnmwiJDkfCBCE/0G0M0nfx9Rk2Djcs6UWO
uoegcjiys4dyvIC1gKr8mlLe/w5CPOJ4so3Ps4tf8yfG92MlJqakgCQ/6SJ6+LhM
zWnYx6MKEcovxmiN+ZqVNQAe3RtwAUjp0evFpYxETtQLK+hFevxyXffQsfmjSgL1
w/zl1B/AqzIJK/KShHKBdl/4zeTI4rszC9+K5LqLe5/B2oIpgUEaTkrQ9JiRXpWy
csnN0bIZYERFg8f//V8fmuXcqglrGrsdoPwhVQThKxF3guWdV/LiVrB2t8ofHdqC
N3ORGsLoso7RHRGGp1D/gWPY8r3q0wbvIv9yPoZxcEj6AGL9RR02QcG17Y9OgH4C
rhqXXTQOXNR7GKj1gipoAD+S/6KGRCAeZKLCSONu3dFhUN5XAp4ZXBI7774SJaUD
87oOFEYN1ARg/QOUVqRPKhBtWNVfV6cXCHG0bv9+IyILaAuX69wLvrqWqfJE5mog
10lMcmPZ7Wkv6a137kxGfKh1F7SvgX+7wf6B9rOJxmJ6GO+zJOn6/RZ+7+8nwJk7
iCiS6/fOi4n9a/QJ1xHX23C8qD0uH1EYg52H5dWpKRTvve7eY5LBFJR8E/FbPJWD
mrju8mGZfD7E1KfvsXes40XxAZkYS687s/208lv1dUsolNbDxjlMCxCpnKSDZPST
X4gwId0+iefbx9pMtYMnsCYBzDdM1F9UQRW8DuqtphPQl9MAsvNc1ZS4qCuxkCGf
f9Cj0L1TohwXxMJRYknz33MieX12UZKDZ6c4gLkvqIH/88mAlyTtRwDC03QOR1VK
cn+qSi9uymfYEKW8a9rXtvwkIpSPyhUuPpyg+Vl9/40AodcDYTM5dIEDLh/U13pm
xm0xiiK69HvACUM4VmXpn321MEfnHPLG7zu+j0h1NWeyu/77kN4eoD0Z6wMo0u3c
CVYwRiphftG7xb1xEsY2GJHumtjFTyZiWd5ti4OtaWIQV8GpVWkGKVZbJx1p7oW5
ZUg9VvbgnkfJ6q95OLwQde23jvoMmATJa4JojgT2nnwEEvZPCW9acFReOpWZlIgP
1gE3WJcAMRs5ht8UjMnuushGZlFIVeIzaSB89RlilYhlBlNdCDqtMeQefat6MI6i
/2VoAxe07iNog7jVViUbGViriU/UnsoxJxdwovpLqQdWZs9Pug0UkRlCTpWcy08d
hxWYTnS7XbT3NcdTBnhJHh849pd50AbhHO+J2dXIriviENPVAZxN7OD7DIpqQLw7
37OpFyX4UWpBzC14u/VUFN0eCGQr7rk4lxUCyi+vKWnPzv16hqNmqqHzgPAtkFAY
/tVFahCPIVl3RoV3fdmybcdDvntC13CZUuij07XDctMkDsdM4xS1a4v8Snwu61iZ
8iPC1DZlKOHbK9Uzh8nigscg4PvxnI0TppZeohGhm72x2/e0MVvN8cXhAsP1uURU
PCXHebf3m8YUrxanycRVItKnx3Ohxma3isiSuLUQKyPmh0Fg9HStrEiQeTDzZXEY
u2dw7OvGxgB4Y+7Gk+uqvNscTJ5V/yRWdKXgiqmdCJUHYj8DP952FnlpJeBxtukC
ySxEmHhwQGYUz4VYAC7pz8it2nO96H8/cfgWUGtMdOcqaOaKA6h8Z3e9zMP6ZmXS
WiXQRSzINt8vra0Rj2vsXskxH0l91JRaQmfXkIjMcTvg13zkUQfPyh0iElaAA+XQ
8WXEDGjJ6TfjquIvlKvRCTJhsvkAKvB/JrmL5PtAgJzieqNfT3pSnSR3n5+NtOnb
CoayRD/iHJ9F40df/NtkyGbiAKwRYxQ/c6dsw+LIupSoxKjQ/lgxsNODP4L95hXm
rrMNKXzmh3z4ogBmAcAOphRMepHrzRySpOiW+hX30Weu2O1/+N2BDUvJfQIypg5b
eavD+/h5CUa6rZPApciLLASFkTcdOVtWHJCNIpqV4Mwz8HoiyGGVi9kF3wt0jrCV
zwb/RjTSBkSYeYI3p4JkSMa7/4ae+F9kgkuY2nrff4F1zKLiOKGVQpsgyBNLDtoB
FH6jsHv0RPU1B7n1PVtq2Ls3NpBdfcZwWOMlak1/r8MJpoQyu1+CzQztqb90F/iD
ncVOxTYtnP2hQHAlbDSQGbjFRj1gx4flLLGi+WGSOibjKhCV8IXt52hG1rW3F/t8
YJYJ0I/WT19wAT8kzUEQvnwpo6YSDk69kbpa0gu3C557c39jYBzvbElAxzlz9r1y
9yEhtcOkyibJQ4dtvjFPvEaZ+KZPQisM9P165+Je7/zqz0pT3DNCkkns2A7Jbu4q
Iwc1YDYhhx6m5//sofkaCPp+N77CHcf6Jgld+PNfAf4cqz8u73uqgwcTevJlyl7m
e1LONesKiTBx5ATIy5QWREj47sv7UTBo1qQTj2Uepb2SZPvFMPO3FVGRErttis/Q
/PZZ+CCr1gs9p6tJrVZUiV9nC8f/DkRY8yhPBMte91jSXwI5z3k1NN9aesQEVneH
iwcc2xVSXWCNkMZV2mZmJoqDmmbV9MNxp86xVvjSxoYqMIAsWZ8Yd7wv5Y/EvUK1
ymbQav6MWXCPnhbj15MtV1WP9kT0O4XkxUHPffGpuvFlCNeb9CammvtGBB3G417I
BQtjsckhFqvWaK0EdgR0Rk2sCNRzw13zedwtIlr5nm+/qPGvRXmwvjZcXn2a/e1c
UAkAj2BdxdJC2KkWsV5Mq8fArNfp8Kdn30N4aQEq/zyHBjM62lVmqzmWXrrtsaf8
fi8a67qqkGcfX+drFVYgpwx47Aqofo1KgfptYO+jYuNMGknBVh214n9qWEDEG5al
Mqg7oiV50kcprBrw/KtIvS/EEE1vkhJUMetseyq2DWMNZ2061/P+eoGVcYp0FGr2
sDKBmsVJUPGVUbOkFjjRVqU1CkNNd9zKUGo79uO8/r1Xne9Ybj/JO0+j5VmEOWXl
/IlCOjy+tM6P1ktJFRDnc6JjNDLrG+PKx1vRq3Ktb9eoZq2mDzsmJII72n4UZRDo
kHE2a/GomKEgvSdGkeYZhwKVqgivUCbHsbYEg8Xyp9cmeWl+aI0l1Z6f29zKsYKW
TlDvG8FwB/rOjDtcsgj2vRPlrMbcpHDbgTearjRfzSf4FcHiAgepCJaYYku3fDfC
ebv07YqIOFpq1/R4xW5B1H4OVdIDIdiUfFnDs8U7jvfxgPsbfnLn5c9liBD2olhv
7HkKTxcFCcOrMkYD90CIomLLmdcuvwZfW1TWwUmEEx0vPm6TlbOZcMoBIwfsQc4X
eMdbjVQQHbw+RDzMiVXLUf0szC/bPIxZz5ts4+Eh+bE4UrbjGBoEliB6/5IKWFJS
wYp03omke2kE8Oq9lwLVn6kHbm/FSunEFvJhom17RZUFrJeOFJgdWX4dageS7htS
o8j/inLnkGWSNb9Xpe/VSkkRSY8kN99lE0rgwEQ+x+8UeNkLXdjEk3P/cQqc/hXm
B4hLmFd++ksuci09gXbES+CA/P9JdafyrgPkRH7zXVT2afX4NfD5PnDUZt1/Cnh3
2gfE+2uci5DA6StjWSkflFE8gSKcERZlwWed9lW3/kpFVwu+rYOffGY2YVg2kPN+
zqqVJ2aPxNQzmqzc3qPdIiAZaqYg4EckEGN4xP2SEv5KOK/yUHgycTQqR52ijjV4
1fFU9lgpVk6HZVRrSfu56T96jRMUUXexp657KOe1YUwyu7q5qWV1XuwmIEntQUU2
3NX37kDpgTscbI7xaEqZCY1exEt0Ain2s4XPcxhKRkaFX1Xev33K3xVz7EVieGOW
MeJkthaNO/9abGWfMqX0E9/lO4NsTerfg0Ki12EJfOhP2qsVzR56iHJfTGDHjwYs
oSOb0xOVQqt7KYwTYSbg/ESylWeSv8zoCToY3RBNjzAQVpCtCGOgMHTR+L2jEDXd
irrS0r7qMkDRzT8aKdf+Yvd3QWHov4kCgoPcvBhdXKtr93LcbiUZhcx+WWUFYC8S
ZRAlJBnj7jbotcfxLZJ3clQR3ooaEzdxHrQi6Nl1hOFnU/he763Zxrc++O5w2knD
RQJcm2uJVQW3DRiEQAR7eu/+tvi7EktyrUW/zzsy3ZdrT2uy4ZQCJ6T39POxT9ZR
DqgEpMSKktKmIYRbdOV9g90JZVwt8srZCIdmjrJ3iwPvgtlShmrMMnYr5VKpblUX
udjMk1JV6+IBgpx+MJuflLD40gx9gjd9pNO3i3gvTcG3CPYsJy9MuWbJu4X6N0yc
Uza1ElZRHKTHpXZ0Y2qbTJz8dMtAed7qDIT1FC2m4vfHcvTNTh188ex2rdowq/VH
7jKlfy4A9qbQAAwps4CJ544c9rLc5hDg34SC4qbSstUDlQTmy8IpEgrJhyh8oaWk
EQhAVtlTGUW2iHvb1AgVyYVaDp+XSVOGKSLlXNwzmzhj7YZhqSYOzGnuKzFe82vA
hEpYbofTibOnrY+gHWwpJYwYjq4F6KG0rbTxjwqupbaQRgk5P4K/1cVAt9vuTjhU
IT+kKa37BIHkvwoX2/n7P1sjqeO0lG+XLQ2VuSlehhZzQMVqOkIhZswguI5elrn6
BNiS1QwlLTuipWrEJbJORbVgURwRfTS2z1G4dFyccCcneujr+i7lXHDa+oVnEqjF
uBZt1BKt2lUoPLnCxtRdpAZRERz0E9c6m4sA1A9IcJ9ZeQWEnTf71LOs3A8A/25Z
6Z88+1rvrJ8qPshEPEMKBpmYraN+C1tfulPDWVGMesMx+i9duoyjHZf1S0nF4UsU
QEVI3cjziHNI2cAH0hMVXcXj92042S+eQm5cTaQZsrYhcdoLJfocvrcbx0EAGE1Y
gS3xUbEkoYtppQnVfOQHsmF8s1MUT2DKNgb9juSmxvS4STsRDgndN9pppB4e01tl
yjx3ii2IIsGguwYusk0ipNfuSzmRLEPYkxBkT2rNiuZdVgpRzNd9FRYD69TrAuuN
M10qXxDQhsSkKjk2WbqonRZSaqLl33fSTBaMxgi1Xsk88WhpJblev4EBpWKWKi0v
ZnrjT9tSIc/y7VrsRQ/W/0xKa+0cDcwgA7svbkigLdsj0W1Iglng94MsOVv69Wzk
Oxj7N8fLB+fRTjlPG/OBy8L8lg8UHfX+w8QEpGcClmEMq0v15jy4a829R6l9yDru
p3MbtnkCJDhOF4J0WvzdBIKNsOTefolcaiKPUkEufxjdrbT+rFT1yWI/a/FG4BKu
7HiqunAwfpLsAYqgVp16MUDn7Vx9qpGKXPTvda3MEKyxO8Ef4zH/IrUQSXTqWNSf
4Mtqm5s9VE1oa1RVNhN3133davDdp0mjMEnhzU2TD+j//TovO/RDDfrZ9RHgcHMW
7+eqx8gBIuGU4Y5ydHpI1TaDUhps3pdYwLNHgdTkd/un4WbFvnbr1Kj3smRB+tZ6
i92ngQFGwZ0k/AXAMTWGxFSYascCZmn5oFKcuft7JhPjzUyI8AhwrzRPeW5c4jsx
xxZCYdOePKDm13JfwJvFcMBuK32J4XTZt1lDLQhWsrzVH4jkzlG5ZjP1a6lMSCEu
5dMnr+/vooxFpLLsXB4wKodVwjMy+0z1fIgADWeZrRAJv60E8qd0roENm4nNIz85
opuxRs+TPOQUXKzbEbUbwPZhFdesC4bsnk7V0IKH63AWXotC2gJcjJGl/xAA4sqD
hdQfXd9pdnyH0MV+kVbXdteWdkdn8HvTsZlETwO1G5LNcHytP7S2YLAUYgi0HQQ9
+yATAFFfNIcE1u6ZfW6hYkA2NNZTtrLHnw4+tIcDNMo8IUycXIicqOZ4DZG0QuxH
DQBHGl+hjlhfrRYATJB5pmadoheYmHOy2Ttizw3cuZLlPGOCRvV5/MydsuyDLueA
ZUGJlW0NPGdfEQ+oGyViT2mn82nRE26ptoun2EDB4TPxJ7VakJOUbqrdJB47QsdR
GCaH8pipgFyMg2Obu6on6COi6CBG2khMcbqfTOxmi8gtF1Tg/dmwoaS5PcpcgoJ8
G22sdlaFLMrU38hB+IMkiYRq7k0sIJ+MqVmRu1BNe22oTB8OVffeIlifA0ye3Adq
CnTTjq0ngNo52VwaKrrq+0sP25moY+HcraASMS6eB0LVkRSP9efaT2wF7eoYIgul
O5/7fQAs9LRvGei5P1PD5ckxO+ZVfR+RJf/Leeo2sF7OwEWc7/9v8kThZwdU9b7g
+rLn8H6ZNZdJlq6R/h+Mi8ZuNkmRpvExciINQ/1Q8raOkQdJiiKtA0v9YDJb0Nmw
JA1zh8MbqydaDZxBgoylVNtGFt/fEwDKvCbqKe7y/6UFXExwKmqjZfs6lLbPR3By
mf2JNlG9vWeqpZhcj9wG5ud1ySHfU1cffWRJjrgJQcsP9ezq6igukx6Z3najxuhF
fRVmLvfSFfQ9S2MFdVM0jPwb1tQbFDwjHHOu9dX3dNr1UcWiz/fnTnA1Mz0ZNnvF
P7ETgos2RmiabH7uwZfBe226siL9zEXGIGP3B7D4blK9Bs0D39gCZGunIUVqyrqI
xv/gnUTlCqWtDVS8eImyvOnU6b9QqfDdDaLl/jMc/haWW20JqzbKRPTEJEjw2Oa+
+6ojN8Pb/W5HNvGlVf1gZdKmImYfBeEbEYaFZDBqfgcl5nAvwsLkV1cgZg0QaOEp
YegcpqwoEeiyJImkfpvyG1zvW+EE1cLRzJ8x4KXAE7G7Hc0M59FjFA8j9i3XzmrI
GEUtRZ2xQpV4Jrx24SFvQuf7yzz1EVGTU4WdCg6DIrIwngnmXBZhi3l1xmuwSrQR
B8pQiV3NobIPBxOJZB/OcURX36LnoYrxpwX6CvT+pD9780lTz2Si7KJ6jON7gVrs
46v3xShvn0tEImY0k6rWIMFDZ2bguacOamOb99wqNdNkiyFKxb3xC+NJ1ml+t1s3
xWAAW0OesIASBaSN7a+rGBnCG7U1598/+iVEKneNVpTwjjrlie5L/oZH7b7q8LWy
xVQePFzzCozNMXs2owIkaru7IE4oUwN92KoeD54rOj88gE4GC3teU46EUyjGBAf/
z8Fdr4lSH/flP7NzO36HBhPYuvxaDyAJ5BKc2b8vkXBXPBdbNqy+itX7JyPowfCU
bv4jljcSDamqMm6XCnBR+IMpT16J4X7xKl8IgsSilfVTX06EKZG5ou9EknTXhC7f
4zCeg/lDwXDuFfAhP/uUUBK2qifRmGBxpAGsc4q2NuRF1SOK8x/vx45Nhcuos6V8
eq+Tggq8lq/7wj6pvfwhgMqkFjJMsj5VraLJBSU/xGhdK9W+W16/f1CTiiItFjsl
AIL/rk04BXk8pGfiB8qGZENAJK7JYj5k+rgX5VOhqjgc0c3NYOUqyCJdJnyM6Qbr
qYTutZFbcLQOLSU0aOLgX/oisTF+ARPertkrUalt3F8o78aK7wjxRtKsHXmk3YwY
WQ+celKUJ4sL41r5Ak8tGMwRh0mq5uZ49lk/UAIXDZexwdgupMoNolMvPFyUgRQk
qly/UeJCtezyjMpC5H1AoBLRmyU928SRWZS4rtrQR9QceyfRPEyxZljoeoVgwOgH
UCYMbxWDA9nCDPu8ggvPE49AX7MGuLxsYUP7y+xWVjrW60keRjhSp/ioNJ30nD3J
ZgeQsU70hfdOapPhppMMXeCiRjFOKucPx4E+NphemAeOHzxweBg3KOvyIUWWj8bZ
IsIbnKNc4MKrWZKmRFNDl8hfQ+KrhSAhuJ7vyzFcUEv+tceKt4dnVRP6S1uAn8Ef
1pBmx3SD1XDmOUiHfiNDxhFzLJZ3o6vu5fUdcqyOkNdm/3CkDB2/GTWYsGFrsI15
D6OFsiY1ZOudlprqdzvMcoTXDGz5pcL4aCK6CeKL+PUtnEnQwJluFP7B8e7CIXS2
nF1orwA9LtQ4vdcGSWLQVltvFBuNLdbWbTeSRqhcx5QHYzezEMFc/UACwWGXVBNu
ftvpM+BvDJZJLAK8OOZcXC5P/eqCB7lA2sUsfhDTSDQGvU7R9HE7XP88d2tEbLeU
ip1XUlLNPa2nR7SK1QGEt02+YAaBG3KwyKp4jYAimErmnfwwfDOW3aHHaxW/Ycju
bmxXV7vCWAqnCJVXZz51ziGrkkNPrQHv1Bj//Q3A0NPzK2mMf+py9K/YRkE+Uzg9
WpuBbC/d0HS8Pc2pVT0+hrZNlAQWB4AdZLnT9TBIJ+2fiPwjgWuzZaGMCVpmz24A
wMKjDBAEoraqhGPIaq/FsfH/ri8OwD0N+heV8M+Mu3FveSr54wHsVgleNkcL4xYZ
0WFrujGjXLCMriWPYcq2/a3tVKdVJDSKZyP6R2gUHGiAbJDoNQ1ra+KuoQhXkxBy
MKhDU63gebtXF18WYxRdZf07YgI6yaD6/PZPnErPLjxtNN7xHY+WPxkmfBIPH80E
aF7gbK98n5uKT5jgeCyVaQxHPoHIVz+htetA/j3dQJ0bRU/7kVy51V6DFqHzK254
oeXLmMRnhmBxFBgTR/+FrtAHjIQsDfSXUJf64O4x4/z0wPeQf/0tr0I/QaRLevFt
O0r2VJfvZf7gh5M0w+RmPJBrJAU7ninISGLaMOQsXsYe3XoPLzQloT9cRSz0Hg/Z
EEPcOyYDh7UoUx5QEC5sJCPTs3mY/I/zsZRp94VAnZm3lc5km4zvADHPJCrx99Xf
G6u5N9TDpEzDhDLPbD8rK5DM6HUD7yE9hDwG4zRmmujM/eihHOBs5V2Ems5aoTqs
+9ipCNqf1bBRVby8FiojOUicDEfuANmiF42v4za8zPnmm/aBbrfdesU7g6SB59RA
Wk+K8Su/DJwSEIYn1unPSa4JLw/FtBxThXK+rOxnsYLAGHRDXSdYfDUc7PaBfj4m
Dl0d7/LxJXOtKJ4R/VVMxg68DbrP8hhUxErHkspAkHTsTJ9Szav0B+T956L1Qghq
ruPsEZhexHoG6d1jckUHUHQ56Xl5nup4mYxhbZOyTbPTBrx0Sm1DQQB337QtNt3u
e/lOrLuHS4Epw18YtARDMOK9Nc6dxPQn3uesucOYGq81Gyap5dz8ccBXjQvGZuZn
toAcuCMzBFrdt8RQZUxbnAE9xeL9FdZxbN3qZisKvmVBWOctxkAfbTlMumvL3vVf
zY4CmGIVPqXiTpr3o6WCgQPNcj6tmKp1vvGZne5tYK+BYbNUPXROPZ/dRadRsdIc
ugBusVCAqn5njbiFmhYo9qJ9FjeE11Ci+icaciX0U7uO6OjQ+0adll0crnoIjsgp
tviM49ozLp9V1F0EzTt4A4lrTUAEpuq1J87yG5odi3yaj4d1vTIN7iJ1vB83vT6Q
59m9PPQ+aq9VA6pMYNRkexQGIuYuu21eoFCN9EBZX5hZTADO6gxuMj0U8RAs2lyI
cJCOfPyduSpOhMmpo6Wh85OOHQL2Sc+QTc0oYEamTn2457rJFFYf3YQWOwh8h4+H
UoOBkCEtaD4x1hgus1Kcd90ifzPYd/7MyuxigFPTxcdhjXioz4V+1Gt3bc1U52km
rb/Slwe9uHFDuW9f35JeIM4aqSjkX5UVh/JhCIz0bdnrIFQ2qbQuBuS5nIcQ6rKP
iLy5NxF+q8I+ongq9yeAvXJtD6YhRr6in6LLQG8QXDo9r3eGQ1ym4p6MifUeINoB
f0G5ieZzFa4JFP0kg/GFvdjss7yzlHZh41JK5LMegMNCQPej9jk5Js4XtzJn7ArJ
CUkl2h6RrBQMuhX69ZnUBGtXO8G8Jede4Cp2hnWHLV5QjtSw+uUSRY8s4Gl7X6nz
iZJQ5464Lftd0RAzP0oY2+whwZRfAus3+A+Sn5mgJuCKzOxBuKWkx2+b7WCKTVjn
TuKoQ9Lrlnz+LDxZ8BMdrFU3HFUKIyzEaekoB2zmFfJ35UrFissae7KuICWqwJnh
OGGeOSIBfrMbv2m8tR3kXIaPPiNgwL1HLmulP5nYoxpTg2762WHWOEp0GUWkjdL3
Xihn8lamuV0+3VZSJ7FGBupi139k0dlSHy8hFPJjAcRIpttwzm79/hfivxIq1sxw
KEx+RrS8LDxyrCtwVCKou3WiH4LJAv62ykDrlTkqdnmt6+42ZF1s61YKybHDQ4JY
pwvIwOhIP1DLQMp49PKRY0u4lCXBzqemU7OxtOnYX9bIdwl44pjbkOKmmOwxIGLP
FJtdDd/sCV+TnNd1LwlLdlZZJKovLK37HjUSm4cQJcL2QIRp510BqtzMzYoqOTyS
cvqFWApmlmQmI5pfLQckraYIkyPMd6zdhKL2tf2XXYjoySe2jXQuz+M7U7lcDCle
+akyPi7Fs20Ve+LMr0hKpo0tcWThfUXtDwOqjFUdw+7EUQvucIgaXLc3o6R53lnE
0U5rHO71TNN066diK0t0JkfaKGLIa5U3KsUYYCmh0rBzyzfOYAfLWilEnmTZoUAr
IVWhkN12uLSVzoHYNp5mkCU04ZIs33cWoHdgSDuKsgwtu7atPWvelSSPiZUYY0xG
GNR1FGFRCwAYXdatt70B9bghCd5bgSeXB19EtxfRkUD4bDFFxNM4zXcOwG4mfMhp
s3ZJSE8jB1JMRrebvISBbY5oCStQfYP44/pm2WdSEGRnFx1kTrxZgV4u9k0CU6Wi
GnFutxICaTqY894JgXwqMK9itkAE2CdCpOsExF1F4p9CjczXBCb/edX2vR4Zu2Nt
/bBZCAmjllowInyt9Y1dUYbIByrmkI+4RLv9zHsxLcfH9nzA2G/6LOEbIO7iELCS
XKsTBEM466/WHeuePg7ggtDj+Ni/Zt4ybKyZB5h/dgn1IBfFm2SIy+IaPdv2ASIY
BdA6j0N+p2h0skKGfnYDLusKpGAMG4Gsh06RZJGe/mjiaFiwlrLS+yF7iVxuMWGm
YUZXPJqYySRWXPdCBPL8JboiePtjygcWsSMKILedZYQuPE2OaFNCVIRnCs0XynVd
KdAJ0hz4AyvI1I0CHWXy/TApOuHCqeXmJm6yBQ6bnwoMvIxfwQNhKbsWFRjpqfql
CeC/vCNBQ7F3mtymMwsEcpZKrmloViNzm5DNIVYTWVto2lzheWeZGUa3Thzf6z1+
MPWkKNv6SRkJnsWNk5Y+1XmvO6HhibJW53arY5XRxpSNchvYOGCdPnnSydMmVEQz
kzazm9KfFHcL3Z9Qr82qZczOjPKk2doqydyGAinQl0i4TuH+FJOdQp9Sg6Dberu6
nVekAHujL/8ZDI6cvxG0/zhNCFXKHv/8h4wJK0zEX4/ZkSkkxWZOA1OhBk6YAIlJ
PbbHy2p21LJ3z14VpbrIsnMdD2ZCaZ4Qxo/r/uhe4K5WZL+HLmEKKSFIQwV/x0J2
Berk6BkcySLvoysGpnqTPCUtYGLSfMYczqW4+MLt1wrtD+jC9WiAAvOyhEroh0Vm
k3CKDqQEzC+5oBqGXwydtHbkb0Ee17h39r2LkAC1U2gZLl6yY/Uct+0ANhfw9GZ2
WSZaM1otYWIGcEnrMV61xT1vgovxRvXWu4MY2D55lUepIPa+PGUmv8i3Pr2HXPAv
cnGax7Reyh7vC/5534CBuR1Tud3cDHXrwDg3rW1MBpGDipe42Fdmp2QQlQzAkqCR
7CSvDfdDmQ6tt1lewfRIOojI0a/fQ3jjJ/D6KxjjTb86WkpRjZMPstT2XIHaeCma
cCojIgWsMdPnnJRt5LSfio9czMu1R+sTZvMfxo4LTGRf3snhbyGz41G3pjuPdwDL
mZ/CZunBiVt3gR/EyRPbXffmLyhzn0mvYtwluQs1Ys1uXXjwIUN7N2RyALzRK5eB
Dn0GCwIIbZYf1fC82A1BzN/HQGRNtcaK3n4sccAdqpaohz9hXvnJxogfqo8f93NP
sd2gMIc3vpzhfd1EGZoG3MEfzIMtJe6cVZJyTCYoT6s5KfwESy8KsCp//UGk5kaP
CgbQItxIydib0n1QXOKZLqygzQOFXN6wZsfkkt6XIUeJOdIa8+GhC0U2RMg8L9xY
fMr7sa/RrobvrF9dKERsBBmMf2pBrQNJJ3ORpapRmyNkU5eGIQ3p0Gmd0t5hjkv/
RHkrarjz8iXhybpCi5cqeDhh/gXMgI7K5rDLImEuvG02/EmPKTLd22rxVbNBwwcZ
baI5X8JbgxOIE9G6LiQAzwypxgz2FGuFntkVi24n68CEwlCO0S1wb6eaOAf76WQr
a6mjjdsbiKvB0x5ld8+q1UiX7a+foDhiAm1ieiHrAhbIixaazFPDzN0pff/v+8wk
xr0PD3dQTb/MSFrH2ttTwBbn3yhZ0IJ6yAk/b7sYRLI/G04JlBYlgqduQuTD2UFG
VHJ62zBU2BPjviXrQt15//9W8Z/yoIeCFf8XmUY9carIcPDLgg99VjSyNq1996Nd
QPOWXjHjLviX5Z18KDgUt8Igz4rj/E8crhlNnaxMWfJfC8zgdlcdkEdYNxInho5U
BYNNd70WzYQuqaRqRBIJES/IiPZLB8XcaplgoTfYh6lGIvJHCBYhdUaKBgVau1JZ
G35UhO6G8PIjKNme3i31ciyqR3AnR4e/jPq8KINurT7r4XJP2eY05ZZXuxrZFV6u
UsDW3IBjyr+2Ti+k7swT6pXG6NkDBf6wZ6DVRMtJEjckJZLdH3STY9JCPbVtEKar
i7XBCsl0940pgAN6qPNatNRFarPkpD6kX2QyIXbm484kaKy2P65Ei1Q8FfHA+ucg
+A7xyhIvUYKCl2JEuDkFdXfB45s+x96tNHOTS6A+XPVbXj5d/JB5HJGHEV8C/k8h
j0FQs+OuUr2w7IQFfI9IPzbO99C6O08gLVFaTWxq554SqgmyWbCDXsH8wn7co03T
3kTQ9W+ddmcx1cD0nyihSNO237ogDb+2qkovK8MSsE3I4R4X+6UZcJYRVLCxOdfg
iKJBAZYd8t/8uH7ZjzM855AurNRaaucVXTK+XnNgwUMDwH3Yo5tkoKmFEuWYjkUp
Fqw4uABjB8YoJogoEzHOmpZstLA03rJDLiRo9GWaxp3MsjGtzai3VywmUpk1XB+7
hRVvzIyGC/nE18M1UWAb45BCSpqJOALHndOMgJs9auHjCl9UAsNT1tBjngf/mJ2/
WyxRx/mgt8r4oMd+QJ2E1kjmAAzJn9LTlt3CNRE4FHA3RV83YbKpywrHPkSPlB+L
TiQsqFOReEu7uHHXzP1e7vUnYOw8vH9aOcYSygMqT3ZVCIFVtk7CbET9UAIQqAS+
TEiPgfX7yF70WGsvCeHR9uENc2dRl6YKBJEGMq2SPO98b/rXAsCbkVCBmT5zwZ3l
jeCODyg3KqECJjaOZBYLpGAinyoJjXDW6N1pXeArfSvo3JYYXCZwo6KDAAWuEnyT
qoQIrijQABKZ0nLjLgCXsDCmY4DjDyXPNqGJmv3V4GeB72jHKpMqilq/17+0VLIe
o3u5lCnCdpxsDBc6H/sjXfT4W+tQNQlYz0zMx91vZg3wAcfrJrGgol8VDE23pwnC
JvFGS2onM9OAhd1w/t+fY0FCp2UXXrBGg8nfUGnkqZRkEn6+FkqI4AZT+HgV7js5
aGlbTJ++1S3hyQT/UONa5r2/QlHYdq5cMC3djDEq+RrCTLxC9ygyw4NK28eWdf+G
eVLewGTfh+4wo8qe3ggRthUTeqZs0Z/y9t5qvkpksIL0dq6oGZQWKP1FgnzNWUcZ
u7X3D7U3NsGznxT9d4SEnew9h2nI7It3IGLnBV8AsTnYhyJDiqR6cB+OrdtwcMzl
M+Ic6EFDmptU5GpYJ7smq8BdKHqExt/3I/+tltWbyynwD4s5ccSCYVFvIaR2khka
BaJk47LNVSIilW3MnByntPBXKVk4YeOpgzKGJ8JpTMPvF5Vd4UiU5huNkMnJ/r1o
4S0t3dchEoi9KpdivzQFYE15y5CsuAJ0QF+rKDt11Pq2ScX21hUFYL1rUU3U+HSM
JYJrU9MVGbNvqIZAyi7QsbDdVQJc6wDKpb00o+75k+vi8DN5nZOzW110bM+D2qlD
Nz+S6vkKg1GSeJv9L2+51G4EuOxhMd5KcibXKUgWckWdq5Ej8FVhFr8ZXjt0X+KC
Ln5V05RE+njAfB/k1HDDjYDiT7Ldg4M2+mSZgAHxzMUoDw7PgN43JEgbcUvYxV8I
jEgZSRsLOnZI8A6ICZdKhO+/bo5Hg5h44w9ouzi4Npx6fUxV3Gh6SRLvy4BpDoYU
+H5egEcMWLaykRmBlCy1/L9cVYMkzvlRRQiYEcVOS1r5tJz8SAlLvbeFQiUULUs9
8PbWPu21xRkqA8LTWqEdLTlZe8gP6IUPjv6uiBDtDQ5uINyRaMPxSPhpziJyaOWF
0Tn/sl2ExJaAIzGtKXgC2LngEWqM4w5wgZ5KMSvflntc797ZA19RrODzPOO5Xifg
8wfmJWj9VVmMZc6M+2Q44Lj03FejRs7ovfsqYeeuGkQWfDCnl0V2s79emuOl/FrR
ymCMqTElKFfJHfQvG8imVX+3Wa4lr9jx043nwKdA+VQ1POYpQN9+MKxvlFcVtE3n
5KDFITtyPrijP8VzBGrna/xha77pR/xmjBJNIMsm3kfn2CiEqndA+QaiGawnpf1L
NgYxx7Iz71ltwpRDesV7qkdLedelQ1Y3K5Yirm0i/lUfpeecxOxAD/fGqugGFZAy
oCCGly/L61NGGg+lnwbOkZIxXIj1eMCdiq1EPm+0dGiLttlCCe72ut9tf1oUDjV5
+nMMlHI/IcLer+aDC7a3cxwkvm6Qa+oTKuH0DWg0H6bWnrKETEon+6oXbou1Krqr
pVdsUnApOOUmmWbDR6wOImbeRcUWihXLnYA1iOZIHp+Q8vic2Pl1JQhzJ53AYxhC
Bys+qOwtycvQTR8ekK9bBZTezpHp6X4eAHGjSdWi8zV+xZM2vUMoeId2Y/maBZ/3
XNr1J6pbXZU7jNYTlc2xAEo6Z/vOV9gwAqo097djHhCpnRKMjadSTNT2DvNDcsmS
ZPONaYKBXJG8RlNMqj9J50YrZWd1q4VkAcIgu0JDBn0ONbDsVathO4KVcu6tTXw2
zFsMTCAsD6x2lWZckY8+Zmfxvm3T9EMglOPDQ94SEBy9r+RJLxg1gNdQELLOKd8d
PdEmtbtQ02a3Owh5lEGCs3wwbJ3rJD7wV7aDMuQ0jI8o1FvHirT4YahTMOBzSmWH
dRcg9OE9GRvxsxF5Ml0wKlyS3FC9cLwEzqUyiJ9cr4fUjqmNw5Mz51AYym6dN+v1
GPIJqgH7Sz35dB53+qGNluX0pBxfjzYfMGNaDadD83hp0wG4oSwaZMAvmqdvfEB0
EcHf/2CLLAbnveexNoksh5hyGnVJEi1RVihpesLoaiL/sNhE4Wi93fPX8r8rysuM
ejcru2vwcuSSJkhWTspnci4jE276EgiMFByoCUs+WhRPqyHQ9MzjUufxBs337lx0
ck6uvHHIhI5Ll/SOB7LT2p6C0tD7lAb/v9THjhhcp2yWEAUNqct/XTLOnvxQbFhC
OK8pI7W1a6sB9mKIO/AZ2Xnl7UTQ/aEpDEawJ9gFvJFKJK6IUF0G/0qFW5Jqqj4j
hmAJEsYZCv0DyvkKU/ho+aSmXGbzBwUXGLWjxd9JLYrkMDiNeu+ovmBbgoAFCdFe
Yf+iIe/YtOlM0nUPea86XJx0aZp47qhQ+t+W8/B/ikrA1ZFp0blepKzEEYg6jr++
ZPeW9LUbH/ncaJ5QPYnntnA7j1LFKqJq3XXKTsgtHHqC7Mqq9jlhmLn2vJnjVIDX
QhWtbKefwGLa0f5KAQmHdQ0MH8Uu9AlBLlyNnjcPqbEe74y2YaUiPVfpuglqMn/e
3xKFJwMFHB5Cqso4XlOkP5UgJKFZSEMr59Q+89JgZ9frb6VTlcedgRuYFzFdZJ0k
ixXzwBJndJszH8hWvB67zSfu52CU05HU2NFQF3l89ho/GvMHkJ0zHOK6TA9GWrUT
rf6ywRSLZ9EpvzdF6rFhpjP7zbn1oaVGS55qRwmJ99KqraF/OS+s28AaFf8ldWSL
+XY8ilXrhA8bj/6eLeQHuRSTTh0LQHR+l4DjqDahMN7Xmd1yhbLHnLY0O30rTlzW
8JFNL6RlLu8JWLeL9X2Ga98tK7v3Ce7VkVQMdgeftTmcfzIRvkjmyZyOsfdy6VTq
b3ZcRcDX17z9hc0oSqpEh86Ua60YV2SnTioVURYvcZBpzDeWjQVWIRRvWZNG9wdf
WhH8OvZ5ebJV1CO/LR3f9779g1RZOVjQ/Rk84O0c4BWXNFqY/ogpehKj1Pu6qUza
DrHfpi11t94ovLd3RGkfW36H35/Eu9ZFir2GMG36a8uefONja4573F7C11BH+phq
vACbT4PwW6gr/A2vwH7LVGcD/kpFJE7yqGgtKrYespeLHUlT+uKuE6eZiKI2EH1n
i6Ec07+FjiVqWZQPTPcCJd9a/VAS+0VfZ8Rr0FvouvZWeDxwItUfcr3YPWQyNigr
9Q3qoVc23oPJQ4aYzjVOxQognqGOHfnFlwD6ovYVakyZZ5pdwb7foQE8kaygx+hC
PNBY+2+0E3riVJTEZq0u6bDOjHcfPsRYJRPpUEDzcYZJjJdx0xyCf4Sn25z+yYEM
jnBno1qixnqWBDPYQ3ckmcJL3m020gUE0LTVpQ3vi4cu0xo+4s3BUVTAcX4zZPMk
i9G7yaJ5fgX7cI9gXpOA7abKIOWRqSOxcrCQQNj3+dwu2RCPB1OIl0KTSH8/7Kju
W9x36zpTz1x0znFekl0uGENvGl4uTFroWDimygHVG1OfjmqrwcdZoecLRFc77PQ/
pP4ll07ECRLCGZ4+anJMtdRBfbDZWY7wQfTT4/ntstUYHpycwhOgpein7fUWfV+W
eJ9fwmdojM8ELk/rXbjVoaQ1ViaHo98H7JZoJ41urVEb/wN5aCSD++99LWNwOhqR
6Pr0gRq2Fcp/n7qGcITLcV+KXFda0i8PPc20KU1eOkNHa0YqcRNoUOncDn7eRLVx
zbkVofIC23YSyRINEnEtRoZhIKXgaDAiG7OfG3SESXdEFLBErsAmMqE9kHL3Uvga
x7109Sqrld6FEZDg4G/plxxzEdtA6eoSDgosJi2XgYaClcM/DidsDW+feMPUxQOT
GcdkuB6bbVRnakSxyPgMpaDVcXUDw0SaLEWlOD9V5q5PXZOcWKwcLPDIt4cm/cu/
A11ukmtSTjhKgZRob7woIgq/jKBPZMvorpkr8kXne09E8MUaSIPIObyN3ZG+ZMQ3
obQ+HxCzG88S/vKRAOzYxczwRvcN71cE4lAkKe9XaQ06/ueYjQtjA7gkI2ymWdrr
GKTFpbZaSS6p1zqDkno2WAnL4hjyxuntSsdwFQwjL5mXy70fcJ4qyOlhKq+b2n4m
tMXl/RuSub3VO0c2WvE/qclFxnmj01Egfg5g03HCT3CkztiAON71zfWr+8nizZiU
xWmDT7WBDpToFQsukq7zCaP8UoGwLqaEjVqycSmh+QTdraWEMG/IELMp9y/BszvD
Hm50JXpqSX8YegkXsKYkKag+mFWlAPGMy6GsTG0zLZPy8fsq9D20pd6NA4iNN/Wp
v26udZDNw5nUF/ynVppKZqVoHmkfp4uuYIVKe1o3zhAnaXq+T11VC3TtyUvy9LYN
1L2zM6+BfCJncoKZw2XKFAizi/DNUB5mBXTEXQDu0TtKWk0u/Cmap+zMt2agVTaY
SRv5ZARCUBQ8uwDBxDXdz+09aNO1mq/ZMD3sT1hE6awZQ0GRzXmCKAZbP79afOjB
+mN6G9p0bDZNJ7aUZ7rSpb0EvnoWHPp0sG2XwckmjscjbcIaFbJuDqzGQViC53Xc
LILzevZjwNAS6xtOOa0XuXcXoj4ZwJwP/IH/9H3clyU2TMdiXj9nYEVKr64R5d9N
GVbC90EdteqcVGmx6ly1SEfACNMK445J54kzfqeslMS33SnwY1hnWKHPeE22DzOz
/kJJIO8YCFotZiNhPp9aVH4wZFmwLQLeZ949bWkBy9I9qUrZvNTYLT0GPYDVq4Xq
1TodN+++aKQseYANqrT5uldEP+ZsUj8wPfOIMf7GuktQQcP2EPB8yk+2lDoLkQ/Y
Ybxijm9zU/Btei2jGmJw6SVadYiGkR/4Mvgc747FgjMVH0mK3q4jSYToWBeOQTS/
yKuoeHQiNgIkG3331bSkf4hYXbuiqCS/SKPoLyaGCijljjXIGX9YeFlfyFr+xxr4
3XImFSy8pwTEsic9oVF745svZK/moAu4e4BWZIgujI9lmIXaoGxzSkW+B7dt4MT3
9vjYob0Oaj/1F7WcQmgQPu38sMTrX7J1n2yiZ2z0U8+RxDkbQUF3NfggPIDhBmlg
I+xwXoPyRseOtVwFurATdOPAjyHcZWg5MNjUmZ4fY26FsEe17Fr+gZiGtorTeufy
RA/TFDC7vcGbZvArvz/TLIeC3tTXw133mBqAWIpFUtU89hLsU/kTNFAs36pO5Paj
7peBNOlQgEv9aKaE4uqBsxNnfN0YyA+iZ+MeLm+bJVOe6VtGV7qJkTwkxjBiNE9y
bdZ3bY6v+lkOJXTaDNebl2U6rDRR3kWDNNnXfpc+mokNVOl0dvzH76HrrTmKQFxi
yPwULz5rirS8oxJ2ozbsNzQFRSHWdX8KF7tYKljmKxRqDxtCPRSCnQouyLopxUW4
8Xu+y+lQvxEQUUAu6SACKygC3L8Vq+3Rk6tlfRuCreniR8SylDmuN7uudkfWuTv5
exCIqF0QalEny7TUt9rKPE5x1sHH25rXX8T+VvTGKcsD5h7iF63KXgAM9MLWbk8m
zZTcPRDQZAVnQVRQstex/QpNJM3dsyFtsnYXjYmPAZ0n0Z4p5ViHCl7yK7f4lVDI
Rwyp0fMRq0JY+egTQ6hb0H9oJD31pgkcA9DlINwTFOBUNQyherQHaEXqKd3OrV/C
mlLdbGQvhbeu6TciPe5asI2O60WRhJqnNkZDbop4wj5nKoR43F5rjktD0LsFbFjn
eSQq1N6ZLXoXpTcLdYCtInZRCrBEcyLhI4YA31PS5UpY7fMS8vu5fhFi5TGWi2QA
cRakMnVke8+bMok8rxZhOMsW4786wgp3hAR+jBCQmpAAA5m9T4RRkxtT9TT0Pk5V
460cgGHfNoyq2NWWh4Ou9RSqv93j7kReocxaFJJ7bK6F3IzJ4/uEouuHfJkcg/+t
W75T37IJJ7HFWpDiUazzkrmhRLYAsfXPfLq9/f6hZLfujlkbUHzoGzm9JKsUpYfs
VQheAoLkvbGH/41pRz1+ToxpIqe/RUUoBQMXOeQZMXWy8OVyBogCQB/zWlwnPmS+
SKdpSYD8owYnLA9EX0nBoj9WGZi6Dx5LuRYoL5aRZ3idS+M01d8JAz5XDbEOp7YV
mhLG0wOB/E5R1aoMEuLD7qisfjpBVtTaLw5Il46r8fhBMHMkROJG19Wf3PDUv0nX
uaPRipAf0g2HTyOaWRjQC92V1Hn/LOXhJcRbHo7QezdvQaNGIDmVPFhVULN2u0JP
kc94WMPyY/NZY2YMxyt9J/X0bRWX2AWgSep/naTYJt8sOMBBUsNpKFAT3WRgnjCt
Jwo6tYjTUnRhh8nS8e58qjlL3MdoCl9q0L1ac9zN+NepCPQcswgiL1z83ZYppKKF
GUQe6MhKYhlj4OLu9o0rRHbWt1g68qEroy1zuotGu8puIHOCWhaMZwehRsBug9Lj
FQ/vzBKA2Z/1scW8NDsPCEyL4imwJFGiybmROVYwxKXsGzLWindseTEFRAptEGib
RZfS1rE9zTP7VMKdDqWaCAP4qAF0+E40eIkOuDM0cN1+7yWl1cME9h91axeKa/tz
NqHY0HqQxHIc16aG3V62KazCn+y7wa5m6c1biC1LmzJVhEOZl5Q8MGbfHmR5QlMQ
inXAeCJTI3qSespBTl7nTyz5B0mXd86/uA0oKPe7UVhbjPvYsKk8zkRdYWd9FHbG
tpgspFDZ1BH6C0uIBzANIb65yPJdxpJBWTp/Tbvf+HfG1vNF6W8NDnHUKnAPoad0
nqpiejOe8O0RgbB4fTGxYbelsxnitKHdVBB2fhbpzvUYBHMrHwq90QIq4sttKdxu
gyZ6gvotyKxSrWXpUMitviLik0gjBJDyxIH1s1eyvL/+HnQBSY9Hws2NpNLlIGqA
dAeSRZUHqB0jVfhYMg6KXYZXzVEH9l4bvuULH6i7Qfj2nPKWKotI6z7GM6UB6T+V
O5p2/14tkfBnYxAok0pY7kFovvHRkOXRvL8N5fAJ7AO8iiwEV7HFl7JWe1GytZl2
nqZkVcdTIIUFWrKdFfA62wZjHz9WaVRMxD8rf3Ss/OC1jaWywcGH/8XIvZ6RUHcQ
Bv0fYcWNCmWQtnS8pBI8CosTTjmN6+iR7H+Q6u7k04R/vi5WCdANDhW8g2Ht2Usw
yijEBu/RKLEDvKpq3omoBp/sYCAXx38Tl9bGPGv0W0yj0GQCr3Hwj7Jw8FJZQ94N
PCXaiey4rDpw1is8smvDjrZnEB6cQ2I0kriKxFf3BeakuDFwGdLwEYKayUTpEPNz
OD80z08VgTF7tv0/BXxY5mWNO2QyNGviUK6IkRIIqLmoKpNuSILi4J+v6Kd9bxZ+
0ZBeGb0UWDl8dQRPTJ5TPfYlXfTOXb69iAXEk8Jq6s4IGk2Jue4CkyXTilJ3PrJF
1RFxAfPPE9ehTlRJU9cqEUqyGLSpU3EKO8gdpT2M955GXJmEMLBKjEQ7muP/RArm
agiaW6Z4KJF5qtOOG27fHcYG0MmfRxi3xdvTM/Og0CohwMUPPikJqxdATpZNqwm8
X16TBjhMeNkjUdZ3Gng1e1+qTDB7BtkaixIsHsl0X47Z0iI9ugt5Tp8yBXKbnJbZ
i273EDHqOL+9WqINxyteVVXxBm0vhmIu/CoVRqH5vr69+AIxaCK8Wd6rLlyGph8A
/u7EVeHfM8gLvYfy48V6pvPIMT6037hVZ3pAuyEwJnS9cscoAEagJFX+rT2TzMlJ
anJzjYb+Jm+Yewy97d/7PEMMJ0tvdFPOCxMwhRwS92Sccik8Gp3sW96uolABFU7K
gXySPge5++6y9ldDaS61BNueZtrB6OzkR8A181sKllQRPbcO6GUAXg2ubbJHRxpD
MBqIwqRzRJdfA4LJAhCRo2I2EESIh1PjSrN+Wk7ioZbxk3NHy0CYtheAt8LQQoi4
QZzm3zyi8uvUg6uq4agiLNeS1CzjjDSgFE7Qx2oDAjTL7gjmLx5d2+rBgx3Ws+lm
RI8d8L1xreEt1uTeOMI9CurybGXlEHGa7W3i0uyTSG74fzirfParIIcvkbzH5e2w
rvYJXqlmqzBTpndqO4XjsY/q0t50G9CAjba++t3ODlIwx10YQWIImaKPedn02ROz
kKhH9WWYDP3pZKj/9p49kWJNVNhEMGAM6W+E/DzOyeCb9LTQzAc+DreloHpA0Wxo
xZRPoJM16ZDgeJHpRCmpCYS794cVdTt6iyLJDPgMh2tKtnNUSHMTBO0DRS1UXpoF
gKpf0/Z0TKtPfwHrSOAcxd5varE/L24MXQHJF9QrJk9Rcs+qnyiUbYijrqN2zZji
b6BFAJ0VYYC3QO8sbrkGQpd5nnIGTp71sIGOVuOwTQbXoOzxc+ZIiT+3MJMZZ2P7
+mLzkUbJpobcKGY7WnMFp7/PJh52oszYkqTMI82IZpRsa74FZNTECvakvp+djXLA
/IUAlTD6ImGSmWqAignL5jBieNY/NgIGV8zfcrCP2fhJYV2M6vKoT3k0/Stnp2ge
ybvjwpydGG3HR+Cmk36TSw78AAe1oxU5Nv0WT8621FdeIRhqseaxttvntpzz0IvB
zdZxuNfj60YrzLGZ+ADz2kkYQdEvkEa8i0XIkbKVs6sj3kqMvs7SKG0a+kQhsNDt
ND3zNhsCyEn6JDduSlCYPYWepSAft15+WAy5MYGdIBifGhVFIBMg30nFqTo9GEYk
O2aYjMP4O+kcEUbZ8h+ZSu3gflPPSms7COeGVpTN4elVjqH9ZoqKnmWKxJr7AILe
ERYiBi+VtuHuckMf5tLtN8g7dFQqC0suWE8b1769mku6CmW1OQeuvwfcWv5zaiHA
PxwmfbBXwWtsiSgBFYTGZC+Na5NfqVlcE2nTF80mpPKj36T5A5ENpT7PShc7xKHG
FGrdBt8Jmg15Ncw+f/VY7UW1SlMgOQiNWwpsRtbJdKqj1akIdMrZC8SBo4T3duAx
dJjLmADhLnI1849FBce4+J+70DVwlFXH9CBQTTzl04AwXiZY27tvLoUn5iN9ehid
KufBWLc8PEi38BmbH+VHwdVxfK5Q3U1UF9ic5D/3xdx7c+9qxTHqtas9BKXkQ6VJ
9Z3SnfFw2gfZq0S1a0ZosGLXS13xqWvfIdDNqdEQrJrpePbkGDLwbQSNv4Mk7Xge
PoXFYQppJBuufR3ELUakFG90BeuzzjcnvBDXKlorjtNnZrhHr3/sojjPb9rbZNSU
l2tJxUssLIMVje3MQrtYxW09zOcq2V784xdpe6sZYGRqCRwfV4gRLNXd1oZcegrr
J/Iy/R+yoggiQrn1x9WmZGHieGp3vLHMFXNsL+YUEKe6Iy+eD+3ooiAzdj4cCcmI
W8dLExpntBtHFMmpal+WXyQ2Tdby5XuD8MthA/F0L0qBDFdgSTpxStEj25xkT14P
6d/sn5Gv0Dud9JnsXkA61BbRiUXEwDQ5ekJtPlMTHSK5Vb3n+G4yoajG+34rfWt3
t8T6AtQ5bftpCiC//o4MOnMy4QiNzzUz1yiPpbOppcrXEhCSlpL/yRTTlPqJ6v5L
we4VEjYbPfOxhhJwuN00WAeNwhRAKcMC/sTfZbFRr0l2kK8KsKiXn+6T3HTPkCgs
ZUAsvkYu+ZlzYnW2MUdpHnn9/cPl1QSrt3E4bqW+pW6ygBHaP05BVxUjBNr3C5rE
a5v9iN/h07Ui70o4/RL1rOjU3SPT9J+PDw8mL/o+Nqdv2a9fz+emK5DL0iTHN9fG
voEX4ONelhArnS8o8dF3vGJBPQzw+ITQPWmilNjhgg9/N+bMQTi4/XZRqfrUoD58
v18a8FE4oeFRpeunEU3F+hl4BRT4+p/SEd2NQOfHtelzjfnweveOtAW6T7gU6vog
F85/Xyg2NHHpaIEzMu6PfgiHEsnXF1RdE02kobVogBAoBvUHut+4BgXKqKgP2f6d
Dw7yMWtQTCPqzvOY2uPqCdVrTYW8XkjlYsPcyuqwdixfYYoaJ5oQm1Hw+5K2jTrT
3b36gNlzHJWSGGnMl19unhT0FOqq6kN80lT4IdTJsc5GBJwK+tngxa13TrBRKupF
5TaUPSKtyuiOe+J5rK7XcmJdeZLoc4YGebwcgc3fQUnHlbKwLekoRG3WsDnByqoi
oGbJnBCwkAhLIzMM2tlu5TOobj6W0RAjOHir67wcPhVM3XFAxrPtKJf/znVRwNn7
Bnd5KOpAARSxUUpfbDiF8sHPw+3KdjTj3V95jzmVBexerAhQpGScJRXowCoyx+b6
xwo4W+6GnJv2RLRlo4nJlUs0y4BhR+DQd47kxWr+hbeI9IXFO6voYImRFkYPpYPP
8F+B19wi6SFGySDAKmM2nt6NXnAcxPGA5kAha9pPqMR8523XB4O5n1dKzOGbvgHk
5U5OUATKgUPEMKxuBkTu9V3qOIXekZYhGt6AD9ZP2+HAjHyAE1dztTOkhHgHBzv0
l7+dc/SB8YMzQEU76RF9VxP5v6xc20sJZiaQ6ecKlsjNutTYfNFqQeUfKq/752Xr
McaJFhalGCvVIC8Jw1p56GPzRTvVnoooYRWLUdE7VGyHrTRz63jxDTjr7/IYEt/j
awMiF2D1yr3RqYnPhRAD2oXWKQOryGF+/lqOFImdw0iMvlVbkX9o7g2XYGGaL3xC
3l7gSh2uye1NSJ1ghTgkXWwm2pNbkDZrKpof40LP7K5okQn5oWBzPkgKxU3u65p+
ItIYNoKzK6sz+X0cipbizUxZ47OAt5BSmqObdURDtCG9PwRnz8zxtzeS16vuyMKJ
Q8c/OdUvhwDxxEW58aRSCsvVrswrCTZhu1UXVWTxnV58yJojKKcapCBv3r945Ov9
1vg5uzFBlkHYenwCDmHiXfV+TZmcPEhKpKDawWCcP66Jt0dXDy+DY/3FovvLtW4J
TRY6PgurgxZGIjcvL/Ru2++IJ+XyAOA4V79s8l9QwsicfeS049gVQul5xFA4rzRN
awc8tTOJDR45yeebnVsjxH4DZiTn1bLCYShPDyWv+ITAovsX50g0XiY89OnNcSCQ
8vsXgsUub9jVllWgwd6UjqOkMuKYKdQN6HFhkeSCeuZn6JF+3fuT3daK24Ft36ox
eg+/EffQ1PNkQOCIgg4G1qybwpYZP9rXnTFDWfxY//cLe7EihSQHsrcHDYDWamCS
Bf7dFgAMKULF2R9KiAVbd7EjmVpNW4SejREuMWd87PLhLzpke82MKBEyvOayIkPu
STbf69PyHOqO4GJ3kAAY+fIUzdzPiL5MSEUwE7q2+pp5KaymuhbT2tKplGu/X7Vc
oift+4tDotrpuAWQcZwUbQuo4PTE3SjzS5MblnKnhPOkPcwseJ5I1pTpn9K9pYXT
Z2jgaXlPjSpW96l/Ky7aNZlDfMksG54XAZ14pwccgiG3RX3+XsHgCLU1GGkktHmA
oHNUOabD/on7Z6bK+ot04x+k/D1APihbvesVzWWxZobp1SD3FL7jjm2rB9IxUetX
Vn6N/hZXPQgY2+/aJn/uk0xFCpUSL9oc/Nk3IyuyGae8WkKymfFCqBp8ldFUeOWw
KD37wY3sB7+QhSAYwCihwVLo/YMJjWJepYgZ+IOBL9Gbxf7/KTnCbotzShgbhmRj
XS5CnISf6qUXmcBQAukb+SB+U6g190bwFSHITANwlrWr/rh7kMFJnt34eHbINlMd
sSAoheNBFCFLNTtQ/WDe9mhs2O7UwMIFoceLkCWaCOCziBK48ZmK1pICKXLCZVSw
9qdJdaeC97Z5MaDuuOaStmfsnjH2/n8276wl8Nf64KykZ1TDcJSExDgHySi8/Sw6
UlfSnlOaebGE4CQ9LufCIj44kAb4gc76kH1v9e5nTKioG+7NU/NK57Yzx1NZ2uyn
v3R576Knk4iDiawgGZQ7Jfy5Swo2pTeo7je+oz9N7HFVDHQajifi6aa7mTxw9zll
6U2gGfjNc2YJlsMZC28FDsuJxH4k4S8aQoO2s/ePkWTMt0zfZAa4KtWp6303VUrN
x3QevJl+kCj4DoqZLYe8eUeBRXijxo/N+2rqx5tRreWyOejLdrWwHiFiKOf0+lka
6qvmoDRpqP4/omYQJRcDDzlkgSuN8JoYpbwTU44K6czihNmbSPYZXFoHAg2CJQdB
m+IOwtv03OXV8Y3uVLB8EmJUXE6vx4NDLWLTIlTP19WNxkgH/2lGJDpKju5x3Zhm
8KD82B+yH8g5ROjF3qNZBKi3UhKyX+nsysT9jR3wGpVEUZDlk6KwiILWdykpKldK
RhWYPzJgvZ9gKV5Mar77I5nLyDJfXGpxu3i1plODYkgDGJELpOtgirVsCRgK9SnH
AvnrflrEqIDxVZQcc4atOuWiOgecaomkvjvgxblNVwVeTjhG1Hyd45Ri5FExZPHn
R0t2I+OHtXBF8Tn2YLYiROgMzseWtapgTPnVPMUdkFNtHh2hgKX9/K/WTBi7OySD
C0k1hShyS1ez1pw3Z6Db6C8IVKed+vDx3rT96LIqxa9vy7+BfzaLDjCQNazxNUC3
7WGhmrsd3dGNVZh4K5jlqbKS+APMAWFdTJKzk1pPkGj4Trdv3Z5Jy1FXYKvxz12U
wLGR6Bwf4PoYuLBUIFiVrxUownYRPS5qMHrF1uu3hi+EL4FA0PrKF+ZKtjF34yxe
PDXfu/d3GOtIgxL5Z/pkaWSxPcO9slzymq6uERbmG2Ri2YhIWqGjf3m3Z1gP3kXN
EzJ75My1dQfFSHZmMEKxT36S8tS3+rxD5x6Bdp485Tpd/lOgs3ZBWDv1yZ4apP3I
xo2ef7uXjSPgCwqg3IBtcT9o13XLzXqNqsNo9Bv/EZ0ubF5DaW2ud8wz1XkZlWnt
ShNt+o1kMRutBjjnEL+mOKcygaEFwpD2UOEKl0YyoLgVh1NAueRUIl2umcp5x+OA
B21pJQ5hceZYBjpZF1N+TVKJTC8466pWsc2gnrOElGmZgkG2K84cLyVuISeifVFx
FLA0kf9A17UgYT/o01hUFLiPk2hOYuljqLxyKa3GLVwp3IacwfYKklP6W60DplQN
zDeFcnl889Bt9aWyf9WqercAzkluDWxEXenPP9m8QGdcvRwj119wPrtHL1rDSr0n
HTKGtUDOTs89Fj6zq+4Xpm98oRt+ftkkfr7VRHlZi0ASQnbRO33+Fhe1zg0v8slN
jd1Hd9yUsi9z1jLdKZpCasbNzZnchgpbyMVY2atmSbrrllGyMd+W+25skQD3JOVG
uRzG3py32MtuEUMoLPlPreIgI8dFweqixNFS/nrMu2IAva0rwd9voWl0o7u3a1XI
sGiEn6p6f5DEBez6wv/dD1qaNP+yw4BkCJU3gex3Al8C8ID+mRyJK1APhzVpOQDS
0ZZaL2CjV88QaiKdiuI7oZybdoMGX9y0WS1fsVa+ytoeVGYxp3GQAEj17/BaJCV6
m54tZBGH2/rzcBjF5vl6Omai5sl4wQdxZj5m7441paV9LapUq3MpHSwbvVpmKt8C
gV8/Uaozpv53owhMQJ/TvTF8JsdHZl0nw1lWkOXbZjuVR/Se+68J8+9bTO1lJvMJ
50Ce9im6yixeiU3eKlLg6iugXVWFFlhSaeZw26pQjEs6/5q85H55KhL5J0ViqLSf
1rPvPZpevLtv0ysAVk3AI8oYrLCJEj4LWCMszyJDfhC77z8NurgSaEDXEVUtFvBh
voI4TmlywBiI0oZ6+xs7fPFXYRZnvMX91Ji+D0kwh2WWmAL5pL+31pg1xcloAnQk
+7VrrTQTsAMTqoCFdi6731NA89zKyisljdiYvSi/Cn8wXRFq2OkhWHOoOiUumu9K
werdmJ6lWpwLpfUWVAh0gLpfcVG5SQPr8RfiTZvwtKfpjFbJg+0hewSVfu105/C+
DOTO287R0tKEYWEkIQRAsytNCyGSugy4O/Tg3+5dr2TA++ATVh27WMswCWgSaVMe
BkB/Or5XN0je0OZEwNLldMsYsjnz516lC2KNfEDWhaqyNpeNGsvOltg7VXkEk/Qh
Z8xUiOLi9hB9WeJbVfsSc3woa5IB+JrjET/r52Wc2Cr02UNWKB+YOCOk7Hqv2t3V
zn+wvI/aFer9V2/+epeHphzUPVQ89zWia8xyvmyNMXnZCfba1bhkYdJJMbVgTXRs
0kPXlgeozC1ejqn5duHLgxta8b7pd1b5eyi2Q8VdkeArWVRezF6x/I6jSgI2tfX1
aieBawHjim4fI9JrtodjxXxeE6C7Bahcob1dPqqb8Ri3u76DmjIBFSd8ge9IzPBD
cQD0ra/eY9NboT8W4GOwBAvBORg/3Dqn9EI/u97uu+x4F1KaatHHgLAz0ByfTukC
mSB1yN0DDXDpzaeeAQ/msOFsHzaIE9HFG/8bNJexbGm3M/8Brx43Q70DHcxcDfUh
lFNNGjRxdy2XWGEaj64jbXlT27uEdcCIQA88HbPb8tj12eftPjYhHLdKhAShW4DS
nMBUpB6/6kEzRU3Y/Op8Rj1ULzjRo8YGZpc6zoYRkiU4lZin0wrZT14bEIuX/Oys
DUt5YQx+59yd2lsc+LVyi70bvLsevkxN+k3kj8N75z4HyZ7BjQ1OWCwtu20FZasy
uejbqYFi5HNhzBDzM4jWLF2cmfT5rBd8ej+aey1sycnVeuGLM+9RPKjxaVzT+5pl
leHt9kNdy8c+XLe6BD4JVxAx6Ki0fw+OTYNjlQCFtJIGTJhS0wsApxm5/VFtRK81
xWnSoywgGm/87mCv6xauuAY8YReolQLkVW+vSqgk3ZvRDo3TXC5I9cG8envdgsB9
osQ8FtfjsRtntDNeqRmaPFif0QKNoL1PU4AlwFKObQ6NHMB4XVVFt7yMxy6FyGpo
OE+ECHDDWOfvN56X/ezIUXY2oVLSf/AGdeFfWqJH5qFX+c2SgbfS4io2GnNGiRVl
3QADl0nur5fi+YNJs5n3xBWh6G2ltUjwXzQEADuIswI5jnXHQ7eLfzjtlyUJ9+1g
EK9ntZxrkQqzh586ad0r+ROmCkGgwUCN04yydFUsJer72gUdfbwbQ0rqE6iDoGU0
NE5Bkt59xj/XyaixFKWwl2RmjZI42eBO86Zcuc0tgpeSXjDa00GVV/S+ZqaTAfbq
8QzZlmz+/bruOQO//5SlpIWAW8YaITS3lx1tj/xzEHywBh8ZOsiCaDvPA6MXAawC
3MHDw/YjvqzPBcbKwbhgRdIMa1ZrlPufvKDN1EbTR0wrT/Q7d4ACjrbmFKvUwGsT
idwrX8oIy0dM0dTagkDnthS4QMUXWOHFQK4pImqvIZbOPtAYG21z4l1+kSOnep2a
lgowFjB4DNM6+wtvSGelFc3ksBPgIkxwG/LzPXeGbs21OpLLLV2Xzi+wYqkC8OGx
HuGzo66opLzEvOVKM0GqAMzlaYOyHoCG0mIZV6jn7CnJxsM1RA1F+KMdiMb4fxr1
gg+JPeWQb3Q0otj+ykm03IG7c7E8+Ie8m5XPxrldr+q0oYYxDkVHOc94AfwuNQeo
Gq51gBhHTfILM10/UTo7k2BV8HDlF8jw0A9evoELqodcTkUup4hCwfH5XJWT9IUo
8jhMmozJS1TN2T9SWcYwQtHZJbYQQH4JND6mf31FrW8hgZHsaXawkNwmes6f1KEb
TSWf9uN/9r6DB3lKSEZuOTG1+9GN5ihSs8NSMiJr8yp7MGS8mh1ku0Y8YS+96che
j55tE6W/EOVvY5l7qQkHUwlR3arpRrW4SgN7SbkmhQI2/r5SV3V4BhCLiSBx7+Zd
s9F203rwq2EEaEg3Ozj8RhlZUe6ct9Af3Dn6+LJBZ9R1+XghuXXjd1dUsXz9xGQp
s5yv+YNCer1tyVXjTjxtwhSmjsQiUCPLYHukX5iClg3ezF3VNDjV37Jb1MvxQJqL
84czHehL2rczD1pIG/xTPrL5uU/JIAegUeWkcB4zEKnKIIHnJb/8ZxE7p3x9se5I
3kPEZAWWh5a5hct02MCXINy6H1Doh0lH7G96a8QmKt45q0q9hizWxyhSS4YPpD4p
iF7Y3mELEV5qDrRxySmHNilmjxZSrXTtMOnsn9AnBLPLfQEFyWOlczUY8Ns9USnF
3tucEQuhpdVBN7IKuRbTQ8pyXzXqe5Rk0RMcSMbDsdS1A8zWtzcD2pJXukZzqyFu
tDuL73T/3sOonTSdn2Ee/Ha+DWlw+ujMllk2SNI9W7XUAQgQgBTkTUfKmI3HT6Li
YX9I+3vrbCSwWkFoPspDrPGxHdhv7QUkCRBmlIQkRayeFhcTHuIxdTIBa7pYscn1
me47zLuXH3rnux/NcdJEEvHxflC/vrehkuG0xGHredqZZ+ohgeLtTBpmPsRDC3AJ
kbImUmqeYNsqh14YtVm3ooPm5yaaXBmNt6vPrpL3QvB+SUqoIhP3LMJmM7e/0k13
gYsO6EZarqREfFrmWctV7incyh4vakFrhobRNxzinVY3ksLHwFJQQWU+510b+0wT
sMtwrSyAMwqcNVfAdRK62fm1VikAXStmpIHkjBqdATIewG6jhao3NI5eY8zyrbPw
YuwQKc8mSum1TFQDUcuasi10wVvPYfSJ5ZUVq1FIZ1xO05JuB+sUk0wPptKkRsVi
MF1JfF2q6GWHyoE8MWPm2OK1yEbcQf+d0jAWVxvbzckJwnb7Fe1LUIep+5AKlRCY
c9cECWfUKSADmfnCx4R89dWHXoqUCB0MOEgb/bIx56QMPFzeaXuHdf7z5z5HpMAq
xHc/Bhd2BZ1L9/VRBwb/9Kobz7zkHmMV8lJ6E4YoVCsZWm3gg006WnWnRG0Xjah3
Qk/sO0CbrzHTWzwrTgL9ICmQM4nQYaPYHssHAy05ZwUxWPbkW3MwPw1X7+AeL67m
hSoXf5yUmlox0eriElD+99W2q8qtbcwIy31LB0U9lHF86Drr5lbh9Wqi/7nHAUfk
baCOWjbpsZbVaVXflU+TBBCOM3QDiTvte6M8QS5ZFbu+Sqm82iQWVMZPak2C8f8+
iPz0ISGmJ+MCPa/+CutGuD+3pg4z/PerwM+a4UEw4iKXUts/9w31xTgk9iBcywMj
+nNPlp8OU3rVni8HLLA50ghXtraMstm1S2u3yNPWB/gtBVPTZfclLpO3qadVxEqC
NO2GCCO1Z/JfL/QiNkfc5GwFPDum0dnwySPUb7aXaLT4oUWXCtv3Elq3z9bmob69
kr6J3QqzcFQN3U6/GT7kyObqdnWU1DK0v4HfFoDI65pd6k23YbCbNST0CUqhuVQb
Py6v9ash+PUg60TtyIPivGs8S9/vT4qAvMC3pIl+N1l8HNZJnBVPNuiYQoFU//O4
Es+Y1PZX0PeOQjEA0lUvRD/HBx2lqDsIFE48KD9QX7c8UYLfN/WJsjvRIWT947bi
8XZAOZtKtyYR5bqTf4H7TV2Vl9wXWHVLn9Gp/nYxCE3caQCtzX7iDN7Oko+2BUF0
BkBkihPGqt01B0MiGa9UCszqGfWEOJ9jEOa8+n4iYRkjV8xZ0pbA2kVqO8h1RT3V
55QvxqLLgyA8uNVyuQSMAYSuA4YN2t9LyIldYg+GBTwp41bexfBhIy4Vt0BRYP+5
5WZx91O3rs9pAkW+kizAJXdqD5G0JESXyJzfr45BULEtPoVLTukdJsJcnGY4oac/
21WTbhyb9AgLR7FTIxejDjb/Dmm1VeXQxNMbUFL7q/Oihh1dqcmh7fLMeNVDJZM+
xZ4yhS6GRJyQ9kwbu2WmrzdOPCi5HCcUOWIL7AEmaQKtLoLSl0d503ZuzR2DQyL3
gLaKlkK0CUUOk6dWOkI5wcRqXj8KPIXy83bMkqhL094KO5iq6SNNf7B2fZ06IRoo
3hUIhXAIJXgG9YvUyWeMaRegKpy2s4hBzJl+jFscJVYtXbnc0WsXMwZCDhFuWu00
OAhh7XuFsSCztyfx98dNKH/Qsvioz6/bGfPlRoBBlnTAE9sdLoqLLNFSBChewpKP
pFczndc+DratRVIS0be4Xa62PX8yttK1mY8wkmEXdqUEZSbxZ+esLTemPfQmJY0p
xaAi2dr+5/1JzKy9eTfGdQ4UO8ygpOxecWcA2ImOXM9q+l/ULCJnsZa9ObKCtk3J
l9leGM5Sh/YyorBixz+JonT8NQdraB+cY2otpPby+usTw+bearnAiHj3fbNH6dZp
SJWFHTRkWj3oEpOeW09s7/GPaPRvXkxd0ignzIKVjaOEw7emyg+ut1pjNL8mlfkR
LTqVOXg0xgCvCDbZEjFSKI3LVDiCNn2lOZ3HYNK/oX2xuAkFj+9cqumgn4F+dg1I
FLuFR4uGEQ6Clt0zmjXspGk/P5yXmI0qvrAvc1EcSvPt4Kd2xFD/2KTU9fhaOyrU
FvmGoSaeHj8Hev9Kooa5JTgxRtrYU8DaOnI9vJ69JYRlozRALIqod7P1wdboS5uy
tJKqvUT+aZUVgQpHdv0LeCIimwKAzsmwSXQvfFUn+/Dt8XOG8SBo/yCgUu1b3GZN
NxnermYwxlM5ktDo9ZwY/KTMqDB2bHkz7npw7EciCyTvNImJEmWDh9MtIhPMqIrV
mwpK7CVHOtNmU7VlKQOSRj5OLzij5baHtxfGKRPuLOBJsVUC9hn4BBg56rS1FLaL
Zml071DrKezizG/BABa27gIIFei2SaJYDqlIEl0Irrhnv+JTeL/W68IVKn2D/u/J
vqYZ5BcAbWWjmD8DcvsVBokpE8d9BxVaTXJd7WGi5DWh49HKQxngjHVNKk2q/Pm9
a67nANmNoRxzJxO5NU9WxwR3R9GcMNGk6uI5aEY0ADrDYEJQPq2KUaE0CROVCDdh
0skGUhrxqlRyEcEysOX7blS9NsuYJ0wcw91Ajaf6OiWzVPU2b0+bR5wSHPaC/AO2
j5DsqTMUbPTi402yw38ElhKo8+cvn/W8aeNhStsY0m7KHQ6L4SLGeIyjPNHKmfPm
Fc7kJ1zlER8mCupDJdwJD1gYGlxK/4S4ppCBJUGIBS+Ie6qkWYZT5VQmllKmpU2X
O0zckLiKlI7XkFF7n95n7bjjdu1rFyWtBKWQh4rPhDxYI8uDmHgW3IJqUSMB1OTp
jlSIEOPHpWVNnMfKdZ0kPo+Fgg9WQrqTOCb78td1ba64+cN9W5lVkWSIwVpYBVz9
YNAh8g/gRmevHVy86xVZ/fJueHEuFnABRVU5rHA23a0AqLE4Etn1Gc2CnVWW0qyt
eSgqwc0F7W8tdMNVykL3Q5lhCTRWTGu/ZCGxjcnXg5urD9aRHe60nZ4hDwJQpsuH
2uGqJPepxRus2aJA19ZrnxNd2sJcD2x4A/7ni2ZvdDZGo+6B4FujqInu3EGppp+J
UqXj8n8pWenk5H0GOKHk/1AU3bAqrBSMK2XmI58xDin9LobnruqzyUVAmTk+63zD
g5BGxXumhHjGb+SbHldcCzj1SF4m5e3vavBtniZec4y9yf51Gw0I7ldEWwr2XtbW
AZ+CIZl7ivCGG1cCR0ujlk7sIrfZQ9lWHcWfnw9WP8wlegBrrnFxxRIE85/iZ37u
cWIuvX0KRu+JHU6u9uSCMzjMnlwJ8bP48WMmXURtTL9ouhFFU1+kDeRcR9/WD/rQ
acuhxE/sWFQ517rfgsLhJ9p4KVNLtnLJcE/9plHdOtPoJ2m2hyV1UNDNYj4uz/Rq
ePV14UeKEb4rpnKkbyX+uEKLOvfG6EXo5p40tTT3q8hMMFFJZPya4rf/WKUpo+uO
6TteCpXkPpn7Rb2PWfvDCXnZzo330PXjUHR87pacHqI0Ys2wF6gZb7BiJX5QQOSc
LJvrQwDi1Idoo/lmxl+75Ke0gXtCDMX+C57p9StJkVFZ8u9rZ0B2gaK+qCGbBThW
FbvBoEflil1XfLPlxSwj59mGBZmdkOcPWGROaRzl5uFWZ7Gekff1X1ieNo5LqJOt
gquNdpC3EzB6r8qSi4U2JdE4Udzf0M7ckBMoe8mySwlhJnCfRMuStH7fnL42Svms
yGpdeidtCoKfkI47b1db+bBBFk+0JJ2RYJFJh8go8tLcKIco33tv77KFUKpIWWi6
+gUa0bzzJ9/Rm3K/mLzOGL4JQiuvUnxu40QtoI3QXaWWWUxO+sitz42+zjji+/3H
/5zYnsS1zgw5F731gPszVPcOoppt2bDi3/JvgzDtka+b8XfoUmQkzPzD1p4NhBbh
pSLZseVE+iA+M+5NJUEZupykFa9hxk4TuVd5I+1eNIU2qBz+yPw6yLyQnRrGlU9B
nIyRfh+87rLCF4BNT37V9/3jNeAlyx8SU6Nd/2S3d26Z0vI20s+Q8gfDevD47UJR
JouYxH2lhUArWcZU+WkKGHq9r53TvTlBtfhYhblUg+JkqAC2fKMT/K7ZjhZEw5Mq
45AqiktAgMMD/evFshUJS/qXnan0SY4+O8YEDioWzzqPsOjRb6fbm5mf8g6/PSC5
AoTutq7+dai4EZXXHeE2UKPAXKWIea+KGUFN9ek4LX2TFc1aJidVSUCi7dXubjYn
7VCcc+/LgBV9C1+yhdwC6xKxOtCNOOr9oolyXZgeK8qdo0KSz57bqIk4KT8xMoMR
Qzn7ufxfFFFlJHwkMwdCfDM1klD8/Ei0IOe7poSsUMubmVNHM+hSqxTRyjTl4ezB
wYaoGI5ftEN1wXGfUSBNuZJ/YOyoO2Dv8XnPdImrORQ4Z45KwWqb1hMExp59E8ae
PBEr3VeYhFTAwW7K/+cbGzzUXWwJUjK7EVj4ji/EbaPPdWe1mq1uJ3KpqVSlXItl
+YmE6bWRSqdr1XzPbtK7rXauD+Xc0v3FWpREwP0KgXyRdiWrvPg/UJwh6UMTpa4k
RJFhbJGXiKX2yLyW7iOzjBU83JiagXlhySSRkiFymzrX2PM1v81cDVVGTNA+SYI+
h9jdS6r0P7rh3jBDyTIp1UKosZixpwMSQifIBzxcZui1ipuZszByOD5ZKs4q/kHm
I+FRARuFXVBSmLaNrvRTEk4Q0KE8K9SoRc8fF2z0fQFw80NdGb0arfYIcqqdW456
MVcIU2qmYjI8ppwWNtzU5Jjho4/qPz3YEUr6u8KhVMMI6wnRaN0vVW/tRFKdNa+t
+haWLW0wWgLgkDLtfUc5SpLzIlJPGVuQNZctpznKS4dh65FB2Tu13DCbwDV/fnwO
IWKLetrjWrtgJd925FMgqlHQkObm1qvNbpPzmGICbhcdx6+/+4W4b+KShQqDUHIU
DpydbX68ZRWHH0KwwjpQMkjw4N94aRvTPosLu/+Q29MhcjfNG0O128MzpLuAvWtj
sxRE3PAJ/Elm247Uk9tZMDEl0LCWX2iQ49t6beEZrSqLkPcXyX8A5LIOCwdEkc/X
4dGmdwALcf06YBmEA3DPAdu1xBLdalFXjd3e+9JoMp6TgFtDHmKL8mII2plAIRle
XctHcFN4gBLWjHelU8CIUOwTr+10oY96gVaF30gqof2BEcRboVeWrSDKwmDB8c9X
J/mOm2twwYQQWSq1M+sjyQPhGwh12frywC6GMm9zacvn9xJc7qlHxWzcp5D47tiY
hnun93FG8C+jy6GzcTasMhf0qZC2I0zI8xdI71LhlzskKVA34bDjIuvCAh0k4gm2
mK0KkIZfg4mjz4HvCSlrptIQ5YpNNNCUj+4hs1xXIqFPPF0qCIT4Q1aFUc+ZT12j
rJao5TF5CEExxJLqyBKzxN9moxsEDf1/n2oM6kDJRleTBX14MiCz4CNNsBO+My9L
mAPGbxUl83uGkKMcXiXEse1JRHEMiAAOyTXxbndBTjtLb9/1jVJAxjBdgN4Bj+De
AFafLC1m3qitMaltyNU8vyP02Puy2nc6Bd+Wvfrg5iSn5lzbQ9eLniLOtU+y0FVf
4347yvA+v9dh+rkYpt/Wu3tbRxJghrkUIyTFr5dnNgDHBiRDKlBcTtDAdQHYiuJX
CXyw8R0p7vwEOY2LX+/Lb+ZI3F7K5zZN6qaOWWGYwPJ2PSu7by9Yn5xJt9Z/OHFW
5HzRYiaBrAJ+UWDKhDQPwO8YjUnwnGki37MNCt62uT02ZOg4t1E4Q+vUoofvlJw3
OgJk2lI0jK+a9NQPxLibC6pu8qi3076l+DKmRVUw34vtvyD9rVgDyznrNQZD4bIN
VC20+BGDkRwHFPIFqk4XQUqokFCoggRKKj7J+icqgSayNW0fXaWzcFduk0/+p8eB
jqmSXjrUf/b7koz2D2FAeXUN/DPRdNZPSSjNo+WeCwobDeDscYZOm+qHjf7hlstR
iv7tA1gtzJz78YtloHLznCq/p63ejRxMb28LzgxpJjbM0GJ1EuyxqvmajzzQUwce
hYnuJVr4weQbBxUtVoK5AfmETgb55hrzriv1faPLTsmCFx3qdlsJYY6N9nf0Nvgs
EoFx+jVOAJh+0kgRskWqIrIvid/ffnTANz9X76+0cDctglT471OfKVttFgwJcTWW
maBqLpfkcRzJewvpT0ezETfBG4CG5t1UTKIm5ZXBo3nipynA8Q9m2QLRc6Um+8kC
Js9nUWdFioMNyRxCh8PrHdf9QUy8c0jN3FxffQCx+ynjeeYzrLRRI6UG6g2cwE+X
WVxmVgT1e0g/bnVX0gplTXNOQCHAoIFKjrjS5GuD0Q4pXK8a8t0uoISGLh51/ywf
DnjxF+lqrgbh90dmaX67rnZAaV6gclenshbttNxXjnN8Caas+EU2GWCAt4igimGX
gKQPFjd5RHo3OQL+iRalOh1vDrD35TbdCtqhIn1+8cmOucSRFiEFwlvDFVU7KlMm
ZeSeOWyGsAycjYtWPdBe1gPjieg3WtOUIRnmvFTrd630l2aTTGM8gAG9xkGhxWI1
V1GFWgk0jN6PJUm1/219hUj52wU4CiYIeuAHVz1qzVEgvBsU4Rl2ex5afX7MoGq7
Jxq3z59NVBkB1hcajjMJM6s93KTmRm+Q1K1mIQVC68x5ngpAXwCAFwYRlrUUpx83
9umiZn+jRA1jiz8yHvtpk5dhU1BkXjbRmzp3rEOElQBqB/nuiHVWDWYqDi6dQzK9
ERPNGwyUUhvP/WiazimMPBmh5t2RdoBQSKtdV3hqGDojwHm1zYThW0w4SfUos9I/
j0yIyGp7dhj4couY+ZsjPy+5WyBVq4UekNYf7h3j2aIr1Kfn4z643JlikDjDvnTB
kiBhCfcP7sCBWeamFjPzmEGC2IVCVnNRBYdlm7f3NXHsr3ePiRGHgqfS2x4es7+M
Oi9ci9kRf1k+Yt94kf+jkDZH3QWM6yE/OrrrvMHg+5gNuchbdgHIGGdS+lPNvhpW
1f9x4Fw2DXeng4rLCAVxnt0n//u9Lz3IaQI2XeKJD8/ygCv0GGgGFXopx/tHuMqM
Lcw32Eo/J8TPeNnnezpj9Z13N5cnSBxE2nf9QTq/05J4dQ56KA2tqvzMp+Xf7tZW
HrqdLNQaBbAGAxOkhe6KsEghb0WCRzGoyYr/CaJ/BgvzTo2rNQIGTrCeeADtx5IR
4AOUa+uDnRHKaCLEHmKR5s16Vtj5MX9PPCv7RpQytrlVDywVhCSInGARDf3C5p9D
WJPKhabhITUDgqw/BQxRy94ODkDRkkXDnyEJhVVgCi23eTtkovnuqIX7oyqb/7o4
aNIYMl+Tx6FTNeBC03jefcZWLa4J4bmqCeUX+bPuKO/5daIo1QhOkG3LNcPLSFdv
auqICJjdZH9Jxfaq7q7EZ0Qeo+2X3jbIiI9eSJDSlAKHhn+w9TI7Rd5uYQcEXX7v
mjRMQF4Lj3I1yZD3cOss74rxdOxNGM+FAkSnrCGIxy51pIxl2FcDsEFGt5meUsUB
sSBvC+9kqYRpm8Pje46PhzBSWN3cwseDHi09AeSJO8lz4peZ/o/zWW2agqitRhcD
r891R3ObNQBg+onJHw0J/1vuriZcsY/G1p1VI+yX3UP3fLlclFx9HbSxhuG50oQ1
Y77zCAtZFqujYHvsiUVDVzf3mwIT99iHL6afa5czUxbVil859AqhMWUNDE7BxeZu
+G42JD4V7gbnvEKoy2amCxDGy6Pt/vcLiUF6Au+rtA9XPmUnR3l9EmbqTqN42gkX
RlSZdsYGS4FedoYHNEButl1tn+5UcTzd6U0PdbEBaaPUOe/bVy0dZ1KJUIDDw79r
cDP4m36+WoLbUaJ+XG43wceUaM9YELxP3gGvecCsFWjlv46uBlP0ZXdnPHdy2zXl
xvq9U85aX+wrFUirRd4L/0OZh7MAHfSITNqSNWZuk/7sLhaDFKQnskbEXpqcmk6s
E5uHm9aEBaZMLNhgcZGCSuhBHbgaeNOK1iT5y5Fq1PvvuKZBb/3OajeD4TuxxKX0
QAWUMUzUObVD/1I1m8CyzjfrAVQA3Td0S7NgSunD73pmkYsEpo1+ihm3fwBpouBX
mCCSoS0EM6l97LRbWhhfu96p/wZ5cOkDYDc4gsnEVY1h8e3HqOrb0Z5d6RxEiuKu
qVgOG+iS+Rpb3moxrMAB5AQRj1DajRIj3XllO4HITMwCxcjyX1Zn1zOGAMnUIjKy
mguUt+Eah2OtFOIKNhXSyY7PwRjFLU4CWycSgCLI+sp+1iNUSYgTssEsne0Hf03+
autLv1NoglSFs99w+UDMMq6SxdUlJXo39jPRymuletMUhBQgbBPtjcQOAY+Po1nu
GPFw4XcHGp4gepaJZgCzHy9+Cwog1+dSThHqO+1t+UUkB1KKBdn7EePAjymM6MNP
YuPpXzT7orF0Ha7laq2YijA/nJQ6mIUPYXXh89HsBmEvlPJ1aSZKLlcjElWn99mM
xkW+/v/KJW6IFK4ru96gUBzanAdK/Z4sHwApDbANvSDn24DjptvKR2L8TME1m354
wGwiKB0cX0/0fizzfEcNGni80AM1BS7+6mJuu91SF7SOB1ubznDC+brVaSr9vPxo
II0Yy6ewN2JDQwNzBWuPbqM8ofUiegNVAKspp0i/DvLoA55COZGmDXDJ5rBoD4mL
SHVuDAdC0rXETDCb3ISA6LZkXzSn/nm9P56OFZqqabfWd+ogJe9B3wYWw0jM/jRc
c+2zybbS0vv2bAUOST6H4y0n8xF+KmA4vdsxqgM1r6nX+bzvnSdMC0JXSBQvVDxJ
i8L0NMb8AronOULNpAH3ac50Rv3uR2oF1eOMhzPFwSrgdHw2oqa92JxV3L6YJuMQ
0PNFEdQuQg5ZWh26K5CjA1aP7PLqtQgCots8tzpvwmIpTUbCGkZxwq7erd98k8Eq
Cb9orournwHFbp1fw0+JrRkxOOZQWDCdFDRBYriXTPmnPiULyxkTpLt8c5ILdW4q
gxeV+PS0mjiMS3So9BXB85vAimHdLeZwPunYrYH2OGQe2pwsSQSYsuL4aYPRsjE3
h0AFH9HBk8BMRuGpLyguVq2NXOo03Ep2Vjq6p1ZasUZo1FR/ensKNclOXkwnklxz
P4fFExbcwr74XSyKhmMzwGXGn3Sy+mU/h/UhxDYnTbzsosfNFk5opbFkjMT72xnE
uaJLv6V012fWNkp89Bt7OmR7WtRj7MRcmwkh40AH+sDxGjQ3C/ehPKL5h7i/GJXA
/34QGi+DeiFo09wubRYlm1Mp1gsVxf5/hQbOGmKATn/T4x/n0gyorsNsOhBUij+9
QrQaS6Y/Yic6/YiGcukOp2tkseCiq7ol4HOsVSf/dARHTVyWRftZuqtlbM5a+M+K
J/1Il/+GcAcBPtGwbvAifgpj3fu3gwROtO8cH91JW5KeOmo1aRqjE1tNqt497J0o
SiaftAw8k21Y1/Frvs8I0xNIyDD+fhNsIiHNLBzGLfS4TmUtHNQgnoC4d041/8je
IhkMRL2Jtu5cIeYRQMstdq7tNW2GBBruT0o1bu42OL4qje9TL48Ag/Y2gWmG439m
j1XIDxAfNkChoehITtxAOve1+J6FWDLxT6JV7RxExYQBPOT2L9ieX7HF3GrTGKSk
oysDaEH7QtJWx7z4CjG37fPmXsDH2G3RGTDy30mVqZu946ET8QElR+NFz1YwjgQT
pkqL5JBuFONGyfdsjdZjD469TUgzL4+J5LrX6tr1aQlrK0meVggoObOX+BTy1Tum
oWbJqnuWFL2Pdqc84wpm/EV4MbgomvIzOVS2urWwrUfDa8IuAprAxX2h+tmmGeFJ
uhzONgu0tjKDrYCwggDK5ljykQuw97F5+CLLM4EvpuXZctCasG8Gnc+iFixm2dK8
IX5FdxL+toZv/UyAeDmRwB7n1v0nABvB7QB+2vxMGjTwM74spOY0in/7w9624CM3
YgZyY15P8PgccZ5MbdNl45FMjJXaNMx7S+A+xYjbxBH0dUmtRnjJe/DXEfuFIayF
u0OcGV8lcEPpXy+MqWorv7cr924smawvqrhtlQay+Kpk3h5DU32Pj9LLl2pKKx0D
AoHVKeIQHwZ5IEoYJlrYTY0TkZEnr8ia1+v0qtMlHxmiTZjh6QVtblrpduReeicc
/CXlilzqJkdcxZZcT7LE7Dh1R+ius/YRjt7L/yrjBa08wVNGOOGrnwg5IaWV9ss4
TlsgqHwx+6EFp/rZQXb/RSIIBh8hbtqspnYiGkPl0ZrgH3Wn3OnTZnh6al4x55UR
fEeFNaYeYvuK3/HGisi2R/EmOQ2FW0HLR5J6Y28WN+nSh4G72fIZK92MRlxkf6tv
2aAvrHtHK6pzX17GaWLDrETlcXXMwzRqEkaoWEXYz81HI1iP0AXrA1I8f05QpIZn
XEsEnUmXdS+q1RLeWyq/keeX2AIercztMqOrgZRchXNFs+jA6aQ8IfZqJyFT2JEH
npizrwGxpgfuTLe62m/Abpw6UB2ElkdTj+uY97auDqvfihbsihEv94DnzfV7kzAH
pYIfRVAatQwOWpID8/3iVmMRWS3quWfbMT/+8x5D0wMxm45JoGVr4zl3y6n+VhIV
/gWTHg4mgAjYwCQ1IMnq1gDXN1XMX1PY4SnPjdkGeCA6Fo9K2R+CM9FeYGDmzKKU
XehWSMuPkjw1cBtj22WEiOEt19nL/00IRrXKVFGLwJuuYEvu+L43BG6/xfUvmjsf
TLLRQbERiKoPWgUFhbHPDUIdCLrMpb93tUeWc0opEkt3KIxNtNSSqYuUsukAe/xB
vkN1tVF5sH9tKonJhqbZWNlLAtbs07hmMMEfMHAL3bL8WKq/EGs6hHQzXA6D9X+Q
G8eo1Rq+xe2GaSlv1H3LNsnjlCSKLV9U2kJz21/Q1P1DjJu093PjReuNERjFLx0h
RtEHhXBBnL6LNRCi0/yG4+xp1PIrbJwbdwml6LuHQw9ZFfeEol8LQA+NJtaXIrXU
A1URjcwqzc4gZBGqXnadXYB6tsfCRE9qnjjqkgh9XJnoYfC6VnDZqnWh0O8XOdSl
oA1LtLOAEk4S+vtfFH9UCsd2F4YuMrZ30wN/tWMkY37jvO7nvUq2EgVllieAwrgh
Rwd4EkiysPB/4Muz/41xCDHv7mIB2VYDtUmyOVk0+UDKP7ygnBxEGNNChunXVLRj
QXMTAG392eIrK9SBzZtU3N//5rPxP//EIB7/cs0i7zC27lWjTfAZdYGy7LglSDYt
Bv5mEDYX5yZf/GPqAlGGrQLphZwVjXBEMemgq7KVhNX5eBpIzhGZYWLYERO030Ay
tXsxomcYWlnxnHWkfc9ac3CWFY0T6ocZ4bD9ae+QGa9FcrLOxG6ozlJ8ZfjTFmnV
ad1lP235eAsLUjs+7SdlhmyXxFudbMBYGhLUPbcmC8MNY/898MXdGBK4XUAIpQ7V
Xjksm1DU7G8ceRZ7Fo9ctvW3qrmV6PTQX3v+FSy3BBXSxV9ifpfi0zbCctIBIRVB
CpYNUiI3qWq49LLDD39KO44pFoZXZsdRvngrjDAAYw70QPbExfTOFkamMzIexrvy
TdQ3+7hUUOT2mIy7/10DPhStyzQKWGrWPKK2oTyX4A5OSMKTv4Ss5Y3pZHxFig4T
wltAbAVm3N3k1Uy6cczYCNHQwLdmg7MdcMDO/X9sKV5j12ilTwn1Ue6TOpReAohn
IE96lLPnraAVnUyxYEhst/z0rfxSfhfZLMT9yk49CMjdyqc/7bt2XNwt0KNTwiWv
SdoUXmuCk8+f5QALdlVUi1af/I+livt1rEZhkk03yUoSLGM65SNXZxPk/wodS0tT
BCDTPcE357MksrtTwSTlzSRzKBu1HuBOs2RAH9YzSYd9O5eYbwfPK8CYzG9qMjNx
b2WsrgL8Xaalf+9hweXHHZ5iRDmtHAinbWb0F3ZetCn9hhLyFq6IBSRG0ja8yHMn
3Z4P+IJvrwX5uZShyWy/Qs/3OFv45PoYs8vpVUq5kT4XAkJRrNPgAgZjuQMi3VEp
263ezFinOKw8xWyNKJfvmiOLIe2uFw+cFlRIioyz0SrkfSF2MGhuGAlNxYRb4iya
X0aTpDWRB0pKSCluFMge3IZ1tIxZEyHbkYiWt8de8ZHrBG7tWnZ0iLniapWedYGR
oEqhFpmQQUC6yJBPteKOi5RM08p8eEqnsekczBypFFLqQQTrP0I6eWv6tqXwTd0q
IjWOhZRxNJ/ngk/4A6tTouLRO2UKGP9gGaCPr+3XHCk+vjCdcHpEukjUJgCT/LNu
TwxZyE38B2Cagj+YBfJZVhLjS5qbvz6AJWHgGtlW3aw+Y5nGzuI1vbBX0/V65KBm
o/44C7WsKoXmEZEBSz5QXFOQBiSuyG7jHfIhezbdP3rD3G3nylGK4awpPO/mIMD+
Bi+s+cArFTjal+HtQwZhUMqzql+L33guQH5DzSJNV6rasvpP04Kd2e6H5TYXFXaR
lF2hjqpwQ99CvDUAf7iDKYidGgpWNII7ojp/f7k4lAUqKU+yyGST5DJc7G8azKSR
HJzMrsTJ0JFrQ9QH3kP6tKsjH8uqz9f0qp1e7iLbDPoRYvy25Zickyz/NNjkXPnL
TPTANsn+tM/okyLVJXd2Dl3Pk5v6/ynnw8HA5leQFZjoH1bFySovHqkJ/pUlh0bt
6svrBYIo2vEuS+jXomJ5FH7WGJGx+YuOJnxjEDjnOmWQzqqt+cNj1J3ysg0R4XLQ
NNqp9Rso/gMTg8z95vrgxVgWcTn31+QQOXU7nmZIM9rbGQAd4cR0xWnJZal2rhFX
NcaVJJgPYnTtz08nkxQRvuA619ozslTYaeuyI1D/0EnltgVvaqZAoBUWVN5k0W9+
thTWyAIFqWerU5SAfQmJYwFfIvYfn0Z2bMyTbykpO6xGpofyuLup8y5tCuCwtvyn
dWurpWM4iVHoL8L+nPd63RfTDyQ4cUl1pN7fO0StNwUbaR/5OyvPOxPmExTYlSJ6
QWnpVGT/v+HoOJyxGWxSpsYQSfYhJDYHs8D/kHD79mFKevACx78JL10QhUw1VIJE
opoYLbUEoh7h3WOYt+LqzhGiC8DCNeyVEi9uzw50ZYWdqhe7cMK6wGD1wnuisyKR
U+B01C/iEnDy3i0VInar2bdx+3MOyoIymY+lfpC8DNA0Rct8besKfbcF5Fo+YinF
YkQpxoIBS9pk+IAAqwSvESlv5++3ObNbviOH/IdwfRK2/4T1QpVuBbdt93twhAxr
A3nQwPwybm+8zKnZQp6MnDBY9Kc30tIpYFP38KPNkelHUxnoG3NkXw3tQ84H69y/
wEqviPsLkm5DQK0JXb6iPtAqOldeU8P8lxUG90+gZlWApo13dZnpO7jNi0fgL/mt
jL+XMFYDT9JRz5mVFYawc+BHZPiKtFrIY+7fD5+tnthzTUgzu4SXSwNUVrCGMcij
lysb0jgUHxfSmKKssjW+CBGMSSxqM9PRUVA7NYj/zqz/0qdH+10j7d0ynM0g9l+O
48/OytfU+CRSAqGLJ63L1hjyws/ucQ/78YD9GWH8d45Z4/PBTrRc0UrIge/De0/U
rkPdkFXYPajgEWUBtjo5rYz/8ofjqvbgMFdKM105Q2Fots7/vpGnfiHbDEG6Lfpj
8AvfWOMC5olAci6MmEP1/o8xx3bgXs7S92p7ozcvzWrRsaESWYRrJXHRlIHVCTrI
t0rKOfzJMzhoRLHNhoQol7OQkKtn9BILA2ALstD9uvjcG+VH7xrkzoz4DBUFClHI
1Rc7Tppo7SgEtkPRuBbePBhurCkT1ptg51pR93C7XaACwmhxpV9WKoreXcnDm0QD
OYyL/pOwxcg8DhYmJO3F3+L9R9MzSLkLXsqJ629Dow8KSwD0EhJAj81pwWS5WyhM
bZMmcnA+yOewzQkN5bL8jJB+PUo7XjiJtl3XX2GTxwg9d4Fqr/CXtNP6s/ojcsI1
+xSsX7QvVzB5KLyvKGksWt5n5LsUMe5DeE4BPiSZ8h7t0696bY/AYTB4+IVWCOUl
wX5EU4OYeTgHxdWSJ+Cz4vL2NNuKNW81JqMqLf07xK6UfGmLrJYqxXafGRHJWrAv
coWx6l1+zNQBcARKZPrnFffSdapU3UXnDdwzauzzcOF48v+TuxJS/JhFLslaoRqJ
PQZIYrhoXlgaj5r+2qkbLW+1kKIYKI2bwblWREtrcEl0nXp6U11rXtumL4pBOeL7
05ceXcAGaNzc52Ma8+G0tPZkwMGfxzJJGi8b8mm0S85/QC9vlMk5C99ePRQN1pAU
64+FLgzD4NI1eFIUThH8FMwgdxGf+/M5BtXtgs67bAWmKemnYGkH1LBmp/gOj7rb
F/a7Iu38ETQ3iHDmwfl2yB+KUn3fMfFSmfI+kGOyFotWKBo/KLsBK3k0qXY6at4I
rqjIs9uPBXzGZ4Xgytdkorb+Ou8NoLg24e6B4jX1fhfSeRD55M6cbzYc5BRJjU8W
RFUPkj++Ge4MD+QKrQ5/ehagjojDFzFmXNuHkw4N4EVIqOKtzojwyfXCMYjKPWuu
Y+OIgqna/pMfY7zzAzPaX1QsrfidL9bHqx/acceAKZG9xy5umlZiEhJEMyfaNXiG
M+zwg0GUXd+enfgabbtaYyWnG/cbmYmRXCzYm4poe5FofQYr122gT/WOAAzjwaCX
lOt7dQvkeNc8y6xOsl/BuUQZx/IE/4A8EGE7jm6B9/t0Te95BmrOuvdWLNfYfZIj
qfZuV5PA7aQnBfwneMTprDyIMejc8DKdVO0kueXMpgExvoS26JbQgYB8yQDKiiIf
XS/RUWWezzQI3C75f8pG8kBPS3/cg9PL9wHcm1pq6f7X61YYV/CV+Pj2oZVHDP1a
QT+lIlgC8kScNQJI/PziCdkscPWrrPU3yhNBtsdN0GYfvomk1J474swnT+kybocf
z4Vg5A1AmZtK3RI/+pxbViMc6VkVThZErsZha5W110fMi+9Z5mA7zw+OHHx1cFrP
pbUvHQMuO7r1lYpV/SPY+VJmDrMWHyAFddVNQyZmDOTXfUuYyrqw0a4N4TsiUCyN
UMffehI1SjH6X3/2YXK0rk8qOEdqDegIVHOEEvxfoqSQLidFdsc0UTMdBtNJDQf0
McnDv9V71XzASaA7nk4d+ZfdKctto/awS2oXC6kiWugKuQ+mC4a664y0lp7lvSgL
SUeSt9Zyu0FmeqqjiHLzJJWnwhrQTqHm3pz1kECK83qC3GTaxWDzSjal/iU63ZjI
+F5ztQFgdmZLGNR1mvBd5UX19OCwItZ/i78Q2UGA/jJ3w1e8/c2106f5PCEl+YkV
Ebb9eHn+zLNsQOWh8VC6aCUAZDjgXfNKm+QoMGBkfG5Q7X0jDFFh31+8BJqXdK1v
zdze9LCLbJcCRdt2tj5t86Fjn2wP9Q98gpsxfO3ojfKDTQqy2eFUWcIcwvIL2IvW
HwEw6s/Vn9wMRJ4XIlvAQDiVrJ9oN9KlkOFCHb1wbtibG5wnTKzlfhLqQYZaBgs3
dnHJn05qNKsM1DOBpeAXHS9EP9r4+2Q5zncBFjEvmApstVSMUnMsRHbf999nl10X
btv3XsIZTuEVaciFkMjQHO7Uu/d8EPCy0jyuakvYCy/Vz3+H36s6ZgiKoYLvxKPw
TZhOhwHozcuGAXPbxXM107GKemqyhGK17neS3REw2/xokqrcDi7Z0/v3N9tIOuox
yqtxUrzscDYRDMiaaSHjPcjPgyOnb528NBtxbT0XUq9/vDbMfNl6BCwAw2b464Rz
Y08RLo5c9/SKcdH4Z7y4FyiE1YdodswYDhs/p8EGvV6JEBPQRjOk17NjuIcV1PcG
B1/B5lngDtoCkVwi3J8MLcwRCPge1EoqJRLteZQMYxdADldXeLbJijo52mYHyuwy
fsGf2Kx4V49EN9OF0HZPBQXqN7VDU3N1jWQ6T5HCPjBS/HoMopoT0o9aWqyMEPcB
yXCJwahzZZ1hVmFrUKwMrkdCJ8wPnUEJDElL9YNnZs6EByBQHvAwBeLCrW4fa+jq
Wk+xjVNORz8NWpzF3OAWLgTmpngzrC7FgL4Q5BJr+tuQv654plalg/bM9XAtnspx
JoTk/qBTxvvY3OWBiq8Y5Er00ebDqBhStkDx0BKj9diKIwoaJuoYr/z6+kTs4vX7
7sgObqhrfMmIS7f0d//H/5st2Ub7R3igWV8qpPW8bRJmH08W4ZC5v9Lg1w0GYG8e
Cl/jNktetjvIuiGUAW9Ud5ulY/t2pZHZeppY2msDarDckEifap8WcwY9kgybD19/
u1iVw/8rINILnFtNlKlik7/ZvGkIu0gioAkXnH73fDABo4UfiMxf9LhRL0RLOqi5
0B5EEa5h0NQYJXhq9YV2N7in5x97RXFJdxVEfthblj+h7RKZp0/lSmdlvXPT+S/O
2X+/7wABk0Ru4M3Uy9wxWfKiRHiNMhERzSIk7Hjn1C9Vq0fysT8UyLcuCSNA+j/1
pDnFZCyeWgnPCm5f33/3cyjvehMWsX1o0P0UmdL0R1XUsyFF7KyvGix7JuwuDcY4
zrYntti3E66CDPy3NqegUxWKVVbTUj91PJQ/xh9qfJnll4W7NAKQnuRag3+DeBEx
08X2JcqiLGslqjOwcLyoBUSZDv9DXv5TOeQ3s+YUYtu8gH/CfpT7tatHxcWUlnil
GQf1FDjYVbO/8kjBap1GN8WV80X+MfApDaKZle49g3Po0u9RVA0jlkmRgBo8dEc0
4+YhjUKXMMLaLGkQVGJln9qWGCueoIb53Gb+Z2VseTOqfirZUjhFGr+TVMyL1cxL
uEmUemjn32kRliB0iXKjsvHElrSWu4g+bilA4JisWnDrF22ZYycTbi03O9ZOT2ME
DqzDtT8tD8FfHtpNDliHmeE9JwkjStajK4n4SZ3ZpJ4bdynyQwXkz6Iz92YvxVLT
ToD+N/z2PmxEFntbml5BGprQo9BJcHI0CwnW4zZTe9KdOZ1Lt52/qco9QwcbFb+u
FdO5EBw1nDCHn6+g1x19unLViqn/JfBw8X/xyru87I9kPzJVIkTNUvsLQC5hT32p
N10l2gAtlsCpGzjlVpZnrIWe6X3RH97vZRgovqk3y6ftv5KR/AZN1L1iVr1KMVh8
TN8tgHKjE0gFxsY8JyVC9I3tb1ekvHl5e9PYsT1iUbclmR2wUNxWaebY0Ut2gnng
1D4K18pMMcuMAWZAUIhXPhh+7TB2lSh/bZdp1j3kryUYQEzBVekE16jVjVe9GE/v
vqUoEOdzyCQpDcCc8RMKpd/jOo/yYwG7bKhNNzCXPo9RA3HGzgqlme0u/FRfbz4w
z8V/d89VrTrZbUuTt3wi3JBdlhqVuj8NIcsM1jz47LfYJ7JOWq/9lxJVbmPLtxab
aEIA+3Mc0Ny7V+N7ZePTXRNxmPz0w9HbrwDbSj9oxE56U9Daa/L9dUB34B9xaKXa
Z8rAJk1V5lRoP9l1uLQNoMD/NupC04M80b0i4XPbhdVDe2bHayJoD44gaKamIn/+
VveUaG47JRspbN6FrpyPjQhG0brA940N+SqtqC5nG/tcx6Suz3B40dwtL+SnPlwb
oMQyjodDEpYrWIZO5tsyVJ+U6U6sOtzmAw3UwynyWk+RNdsCtXShc31vADm/fVm2
fSDkpbMt6lkAT0feg7qNs9cfywcY3nZSeBCN3AEIioxVNtclfpIeC5BzM8ASqF6V
g+MtZVRBUQwxk1fKe+150dDfULoIGqo2qtaUb2CSNT40Y84pfoz5RwMr7VY9Uuz0
yUH2han9JG/qRbvuV6GN+hZAXWSAe5bevqX9w5vfZcOCbMYTzxQNb3xjU97fWF6B
M/6y3aAciVUWWKe2l4jl7QVnLL5L5Hw6S4xWq/kekHuxRe1ilKxLw4WQnn+QYpwG
+wDlr5sDA+BLGalsoGrzXDPBiGbqqg8gShVugWKmkor8UR9uFeJWCpJfPU3oLhhE
k0+LoWzz1CzmDNMeSCDKUOhNQ6SprRkzpINULy2o/w1GdMwp0JK8fsboYZ9re42e
kGhleWDYsjvY4fAmzyQyDd4i8jQweQtu1l1jv0sikwxd6ckkF4Qby1PRGOG+p7/3
nYJl5E5D8O1ZjzJi1GxWaJcAc62civwOOexdDJOaj/r42FfNd1KGowotk+l9yntY
H2H/E2LQaSiUDXTIfaLSEIvKxAFLM27IuEjlUzHGVlgrvphz9ZCG5DhVd+ZKZoZg
sVfDYwUSIRKGNc5tfFGSwpFyaZ3hNgYFtjUJ0y6l2Q6MzRnAyJ0dU+Qxh3x3Ka86
QCD6wGjyL/emugbhSJk/RxAL+uG8mERtjTItFX4JldbsGK5WwKcR8B5B2XiaoiTE
A5WNHa92Owe2WKR5szOxGWkfvPNShGkvhcFTYYH7IN4DwTwpNAkMPmQbgcsr33CA
CKwuI05bvjk4jh4d61DzgOjVPUw1xykz7qZPw5YYU5a/s5hSkj6mkzsUg9/dyM29
AEFbBCVHSc+Bi1CX1JCZs0sEgG8F45PThRtoQGIndqrF0op4hi4j5i+gePhzcduA
sCAfk5yZeuU2NYWrgnVjfJCoTQzXYOjSe3s2PK2ykY6PsueillgK5uioOhw8z1Dz
JZc4YODbsEhzzwQl4J1yHj6RCQoWWwQZDEIAAdFnPozOScTW7CxYNQCNzxMfeyjK
VuUD9Vb+eXcE8RrZuuaVk0uXQLm2opycpAe6CgcVWqdZD7WCsjD+eY33UuhT8H/d
m2e2wxb3vgIL1XfcTCORFezriPXbRgtH2b9ICraTrpTl/gMVDCFE441/4BFAThLr
oV0+i16kaVl/ilCuXkieexfEBFPVBK9t3iw2KbqtcxAeHgHIW0lKS0Cr4VCG8E7X
QwnMsyGfh3W7o3yQMcxtAV1P3CbDSCg8XC5mv6c1OkXC4qone0suQfbQ530gGWod
FJLHXOWhC/KFEh0cAkRW/sit2IFauB/T+FSQE95AfgjUVKYLzAYOboG9TUGIPUVD
2ICSiJZcbdDjDna1qj2PzzAbO10IlpJaoPqEd3oF2m7dyjsOFnqPEB92hFIbQxmw
p5dm920x3c0hJ0JZbjE5Jb+lzrkpYONR60/kv8YmwGawGyQJ1g0PcLovWJrGR+A+
GutDibp4V/bAnsriP9CQlhEAZXqL16a3xjZrucU8oPkgrXem3lVmy4Feem6Bx+W8
GDoJiVAvg5RMS/SUDXSnBB9dlyjweMgVS96knP3T5oH6DfI64U+PsJX/rutif0Si
vnd+KlIhZbxBmyzvZ+cRAW/5TtucO48Rxu5nmQXyvPpBIkIoZskpnPxnyrrr7Utn
YtGx6U2YeI3XucKoMYUf+PgLyfIzkm0iTcz94YyE+/JvKpw5NkBJwJ/mpjFDoEyn
t5UlahMjJ7WsaYuGwYaEilBtLTaqdowmI5kiKzgRoHePTt5VBaBPkNZ7OcRajpPk
vMYdlwsRwDFihJchS9w+lSDipVJCSAUU+1MOoR1L4byxQaKHwrBeyv8UTWNDgDwo
M2ht3jYduMFxETfGiFe8L7hiDmP2gn4HAeX3cTtGjl6hsnvJwF3Do87Fo6kHXntl
cSl4nOmJ+629QZWJDcrmK6AH/3M7gWY7Oc1k+1C0qLGXDA4A/ISed5xh5HufWGOx
XS/kKC7oyIaINN4INLCdrR6joaofBAlB399ps+XyR74RY2bQb27ozv4QLn8bDLTp
FvqFkBHu2ro1gbBs1xgKBCIfYwpfHbsWt9uG/A7i6gSMUIEhjco3gMUkEqgDu0WE
zEs+M5xa07zXF60lLYQgvzchaCdOl6bpTgPTDOydf1X5JUdUsuZcK0iynci4OE7o
JQhpegVithnjIfsezgp5bKGr9kCqirJEhnWOIMCzfTb7DlzvnTOVfceXU11rHfR1
8fdF5A7vkQG2bKUTPOAqN6j7buOx/kdQgTTiHVGVTnogMdsBqeyUhlY9Jy2hHyrz
tvJv+eVKInYVCgidIwNfhpEDcPrfQpL2hODPFUejRScAZBI5CWVePKJq5DHM8RGu
q1/75a5qBtr/HRC8Ax21cZpifTfC54NSNRNnij2gczBZhSzeCsS9ln0WsiwKcl5h
QXTQz5TL7n+3SnLVC55u3ct8axoA7XYiY3DujbKSrv84ZkShQUGmjx7UoBhgoUJf
e8lpP2Rryph5ug6/V44ZbAg6DrhzfnYHx5HTRZx9WHrOwp7xEWD4UW3cFHQDnkBR
Bw/AmgrewV5TB7Pz88lImxPUZJO7Hnheig6vF2m8ocldi0FFGkAp5cDe1X8HYaZ/
BA6pEJNWVKaqzjsoShbjYM7tpCYHe7Unwn6WnATOgj1Ey7C2w0Y/I3StcPe7Ja7F
ZgUaTqpRruxXW36W4Q0Gu5O49ozvgAYtQaDC8ssLKKqsR6O8BGh6HJ4j7SJ5bvvt
bw4yMIaiaKuaLLAT7zk6D+EzMLtjnfpIL5VmWsmCLoCdWls/eWmZF6+J+m5a6ilT
XICOvnKkwMii0LgefzltgEwOivhzoE81VqceiFtHvzedoovYl04fSmJlMC/8V6qu
qlHa7mf1hAx2YWWpXDEvHBlPaFFbhFLpZ8sKs66Hsbc0XTxWLSBIIFnJ88G5gEpt
wwTd7IKiiacPW77/3X2F9+Yvknsl7LxNnQ+8avoYm2cF6onGHOQhR5FVYVjjq4xH
fFz25AK7sI4qIFNKbp807/zBHG2yAwLRwxzgPjvkLGFWT8hNlt4DKwEjG2XkSEqR
EZGUunErr7MkJOEx8Z5J8ucgrOt/GlmZeW5VLmmI8wckGcKHEgwswr7ruh2Ns1AG
REGcn0lUl4u9JENONd2ja5ql7iMj4RrUFxRXEKfuEaC3/KglrhY/aWl0TwkHGJrD
Nl4eWropGPAIq1r80lofuyaIq42kDdtEd5aXGB5laeWC1G6wkXiRrJ6+qrHcz1mR
S/LRCFR2xgmizXPGytaM753OTK5SE5BT2Fy2dMLY+nyUJ85lGfgWtnRNFezKKnK9
LpHEo2zZVW1x9sIwb8Zq3Yg3i9xlffr8RuF+RS4U6VJTNBWzRQ7gRYHpFjfGXFL6
d2gWZxx9RHyQNP1vHar3rUI1tZA3jKQhGEgBVvkLylU2nAqj9/UP7gYZWFIT6OA8
g3oW5ESMheJqrLmVKMbdk60LKNGX6wmNtTvUQorCRT8GhRpNiqLMMDKm058ybq44
ikDz1vTP7kYNc9dZiwLS6yN2uiuPRy102D2V1lx4Rsr5kYFwL5uWaOLYLUXEuyuy
0J0ODHqjEBnOasr2LWgJLudMOfIboLAyZqz/ibXLDWLqFcTSU6CuoEy0zHcqePwY
16+1P+Eqvhg0YHZCYHkBji8oa1HkJbBwgd0UXyzeTixF5kcOYoMvmKOw7bafAxoK
Y3PgM6CsVm5MrAS04B1mFsF5jcPidNsBAjgNgLwoiLtk03QApquLIMsvI3mju2l8
vxdXsJuYrA5vYww6/+CHbG9DwcFtQoU5oYHFeXpca0SXiOOUYk2N7eassXhzDt18
UNX/ArDTnhT/NwIkAGlGW93Fi4RCPF/X1PNowTbH8gHh9jHCnPrYRAlb+XGJrKIJ
FkH1fh0xnBZphAxcF2v42Gr379np/+lCIiGI6x8zUyvpWhNcLuo5aLz0vYIaZcyC
ANBLmfMUoDldhHJIxk2zYwKc+xdc/mUL0Q0kfJ95uoravy+TUAMMRGMwa1L8bPrx
5pL2vr32sPavpwC73Z46FsJ6YuV+xhphinxNkEPE95/hNp3JdXDSqVy1N/ll4xFl
Xbhp2QqhnvnOKddV0NFJINnwEtQZQTnzkTavVcusMgbbJpIarNLyotvk5tfm9BAD
3DgIu9XXHKN0wTw2RjSukxgayG4mj6LHp0eKNGjKrVXHv35BMyFdblqmLn/c22+r
HuoxDKA0zcBfr24HYGjr/hLacYOp7pc6xVFswTfjb9Ydr6+IhSXV4pN4aTZnUZxY
90RmHPIHDU0MCU6ifR6NPr/VwD8LrcXJaIh14bV9vJYtiq8C9TBB1GTdBbZEQYQX
A23vqhx+CZypDNagC91gddxyBxg/jImk5QoAQnsyIZtH8D0ZbGIlPTlDvmtwsI7t
tZaqP8O4mt2K79qzu2X95AaEoJYi574oaAhwAc3Ktb10MT7ga5WFWM84kIohxRyi
qmPeBtGRWtJ0GeW7LEMfc7IQohyXD6fBi+iwZU3PBO7IwNpT4YANCzdHEK3jq9Um
cfy29Ybqa0ku8Bqwq6Oz+omPTON4M2g8b9qdZErRYWMXH/dNkijGgKjBtvNffX75
Ni+aFdNVxoqxzqnHCcwRR13kKLwPAzxQOStuQ6N0L6h28fOc0nWBdDJUlz2JdFec
qQ2Sq21iM4R9q00nhJDwyjHZRhF0yMltsO8QCq6UjqLFdoYkjTes3NjeZWrMB2e9
YwGcLtynIGmnBoQFnDGfDOrtwcTbiarDVd6Q2QEpdpzqsZKGj/w6+bH3J2LwMP7r
AWf2VFvONaUz3Wn6OsIBVRvnd3kauP+J+4tYo+mDbNJWM2BEDGTEXYSdKNfNrOFe
NNVTn7uKgl5q2LpJZgDR/N5c/0po8aoHBesVKrKTGqs3HSRZ35ghPcAsWYMgdz/k
1Xa1egTx41gu2tv+77bxjuM/hkPLBhTOmg4O8SIuyM+gzUWDe44/IiBmYvV5g9p5
yD6KSB/yXKp8e6inRmsiPI3JGx5a4ksKBCdGGkTtfWK61Sq/cM1zfR6//ZHx6QgH
fyeFig4I2AYPUF4Feav6n7jzSuRgjgrwrBQvTESmruu8wd7JieoIZcAv5uTK2pwA
g6LTwPpLC0O32nmFsPQ5opl5D1I1bT4rxqMGn1AU0Cn64O3DcfNXQGf6vYGpPvUc
MzRWELIS3KN9OiN0ojVsBA2U7dp97oECDM5I0dJ60cKvN7qAA0p2CqTUSOZi9y81
rdtBbe/4vtodZK510xRo4i3AokXnd1oNGA+I7To6vE+bZqz7iXVFGfBxZOwPxo39
CkrLZ6T8a69iHP89WJMctWqjldWrg//VvYr7n/rMEztp4mF3CgxCyDZWjwAH+o/3
AEaKiU3l37JotDPwYwHzFFQfpSqWcUrFBjgU07d5ji6363MXurvX0HVr/uxWrmet
RpRL5R75VxcMnIRoGYae6Zxw8ZZJK0F1P9ec3lRRSNYlz835gFjvRpnBQ+ptXrwO
sIpOPpl7guL82Tl3PoI/sppvhnjrv/RAHZqUcJXEp27Z91k6IDfYBdoAF2em2rp5
E83dMCJrl29A6z8QBS7ZAKW2Y2c17lpumLjueqdhK+Uj3sHe09Fr6Uy/P/UFYtdk
99+m2dImOS00UBYVWQdiR+a5kNt8KkVu8PofB7sdl4J3H5143wQjyOek5AJli0rL
1cDi9Q7JtcSkCpBwxfCAaofVU5Sn0dKVr0vj/wShzqDbEPqVYrVykdGha0aXjQLC
6krnxlq7KudamYpJXA7ZBFZC3VS73WKuJlV4oBtWpfI1wkHp6tN1W0xLnb2j4mEd
k6tfggKFW/LASk9DEgxmoCQMfB8oO5g1waNq2Ug0g2ND27JSPU68MbXxZPLj9044
76PXxJSmoP3i4pUh+DPqyMEGQ9b2hEmfpjaff9rKxCoLwzIcAkWufDokvO7vauvm
Tx+87uCBfYQObRNnYuEn2GP00MVPRny3DDc5+MGYUPABnzR7JwbEdhk1WBaYuJQ2
q6jN2Jgr6gOz9vlfI6fgZV9/A3MhZvjb+a6sBJdZqIF+OC69fHYbN3HC4L1tfFYE
XcpQetoDnCl8WT0KeB004a1AvTRWk0/mI7ix9La7u5zPEj8uACgFmwABOdLWn/3x
B0T81RHCwqYmNSz4pvMuWp+d6NPE5QtOI2JXwQtbSTKwUFYmmFCBnsTUkSnJjk9a
2Cx6sVxIWv8x0v3dqdsbV3TQu81ESMOKepU6LNacFrwJ6hP06EXkssx5mYhFkSVF
nxDmu5Q+j1xXm9ENDRVFK7keRVLC5u2HhkbhyhrgFOCT+Tj/7tbE7R33lCth/6G6
cpwjzGXMEpEH+RgUKVJNyR11HUOnDi8KCg5P8pHch686D7Me/xIX7IwufoHuwDZp
WvzKDoGGcaxToTrut/cCKusDuHbjW6OUdUws/mXw0zmVSnFYXDlfoDADJ4BanncF
IDGi+yutazHFk3MPU+i6DQQSI5mkxfLwejuSTCOybITQqwXn0g80Sjl3TfK7U9aF
h194yBLd9Wr7yJ1QIfrADn1JbMWPMgl1arjugfbWBb+ala03u1P0SVOUkNddtWCM
DU9pgwZuiVzvL+udNigO3xL/7pCTQsm8lfwQzodrUkLJZ3KoxJjwOmBL3hFiPEDm
wSECdqlF74HR7rZj5ACihJAU/neidYQjn444FelNYbtNQgl+/8gaO8CisQ1wF5Xu
aAvTI3i6oZVQn88z2E7u5l6E5bmSIgbkkXES4iBp1wZn1OsIBu5LtotTiLnt//wP
ofnO2L3aU3FgHpz8Won3vELvNpmmRrqcEBKDasyblQ+0COnKlDut+EmBfhZSdB+6
GxGrbW1cQ4/pqX6ZLylC6XPXm9hkWUK5mJZSMgfSp3Jl94SIKtvPMQXp8yNyIddD
Mjm/H2b2YwAvtIOMZN/6zeO6DClKiPE8QOGOSH7qYf2b4ZXKrVTgQoOTiv3KqEUy
EnWcZNL0uSgXIjAfo5aPXGwQHkj2A2/vcHsfxez/Aw0Uuk4rN5qNyR7ATOiXxMto
p09bh9ojYS+tSY6UqjX78VeZR6CMLttXrlBSOkBZSrf2AyiXsvVExflfXi8su1Px
8vFCpPjMvbtCXbGkdkbsjA1JqtueCIyDyAsaEQGSocl4qdIOHJ4ODBRdLEYVC4Xn
bAmdAsD4Vd+ENWC6r1KWc/2dkIVgihxC6oRavbPOF2cmNjTn1ckLvBo3WBtaFklK
0h4Myb2HsYcuyMltRYi1Xn8L7IAtIL2jh2J1eCUamwQ99q9ZLcpb0f261Dx8VCp6
zX5TbMeSxW0tpH9veMaCzl1Bf5jGdwhbLmuITQP5ZEHdnlKXuLUEFpz6BrwuBs8y
4TAqYjfQ00SKeCNXh079VEoB1ASY89I57PXxl2md4u78tF2WGYBWupUxx9P/v/jC
cw5m/pyUz8s0jvWUwEGKdriF55PgL+YwlM/4n2nPBD1KFo73uzbCEAGn3H19KOvI
bfu3YoAoe6M5FAYuMOLfEq/gL8cG2bmZIYXqV1jqteEcpj/IoFHIsHtcNuY8ZMK4
png2lWkWGG/YcqkVxxK1HXhq+MmXKJ31CMav5+tPfxX3LK9X0uFOqmUCAyuofOSf
h2hiWVNYlXpb+2ycqH5FrdeULnbSbLvN7GIhXfw042Roez/ELAcOC2gg4i+r5+AW
L0O8O8Ep7EVPoqxL5STFPdI8ruyYg3OY3F0PMFznRu9OJ6EgakOLaeV65qVnnl9a
YOLyoexXT2bs+9Y89lt2Eav24QOsq9f2WdLLDa+l4KpLwPh7WKLWzrKCSk25f7nd
U/cctf9krUgE9zA0MGoDLHGXA80d1B48g2fds+bgb8z/OCNaJH5QXgXzfWfj3N7y
6GFVA7RO2LDOhzWreqfVWE2gj6NvYcDIH0pirxs7rHbx15uCDKCmvlIxLtuahTF0
FruTaxKA7Zqp37u75ZSdy8YbxSfTky3LpeTKqnQiwW+N50PbPuAQlBkgobnlvMvL
4SgHK+XEdXa/O9DZRkZYFrEUnCiKDuFr8XxWhysbfS8ZCc5uwRBLGofT69d4990s
SnAzDCOxZAfFai2gKwwQLetm+0dr/17KP2erq4BU385vxSWGl1tvqOTH8PZ/WtX0
cHJ64dkBKKgOwuAvIYf4CEHNmHGWJLNbzhXt0a3D8Uom2AAOjEOUGuDQtAypiwse
R25vG0Mq9iL7l7I00yiGfnU66pL0q0FPN9sDa6hU/N5z3PWy21KrBFXbu1Fco4S0
LNd84KTJvhYLc/Vkpgxdu/jUhAVtpg9Zy/kh3v0X244gHS6sLHOY7vGlQ8wq3RNt
NG/O1BKeIG22p6o/B3akvgDj/AlTG4ZPALyI+03GKsmwKWi9pb5eYvLkiC85EhRv
G1Gu54k/asQXUrwR7CDH5lCz3/dKIeC4kOvNYMQFOLinXsiJxXJqsgII97ikUcrf
JhkYlfTaDrdthR3VJkDD+0WsNHeSKMRwANHtQldO+b1EYO1ZyycHoOEzKvYB/406
xjS88t1XrMnJrOyXD0BOTnsUMhoGcWOTM0E7oDOW4w16LySahc7O02VSJP9lo9P6
dspzz1ToRX75VtiW7uqTKRA0CP0+xhJT6Tnu9RK9xqAuWNwv9WZgjoq1k+A1ZQy+
/U8fuy7qZnrP5nsV+UuZ5NjhyW6lyO+6TM+RgNGKwFslfYajo52Tw4Ue87PHnKVA
Y/GWpNs1ws/N5Q5bBD4HImaC7K+1qoCbzsYZOzajHZAAp+qbSxOtj/WmsXFL5rok
1zDuU/6Zwd0oC+NRyy5c5WHWp2Bh0FmVo7L5UACbYCn+mSK1qjmT989CG0gvpYpN
SETerPzZAtv/1Sb/B9qRPq/wI0USD7QENoR4K/YsVSJRzz8th9iEm1MMienEBz0V
RadRpxuVO3vlsg6lvu6mXVWp0mrX/eMBd2b78rGHxU/1htRDWCkU7tVg/cL5Htjf
3TPR0Or5Ewuo/0GlaE/sJbHMmC2h9QLMJnDwLaGG+09fUB2hdZPLpEzkVheRuULk
Sp9EWJ4WIoFBp/314FO/Dg==
`pragma protect end_protected
