// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UBRGbbB86l2IEar4s03VwJb6ksToPpDEx3wyaOY7SFkEVVuAuJIfBl+Lg2QKQLEU
SuAmhvdjksMAk2r2LX2g/3Chs3UmanyybyL0hXZLKOAhYk4Kj6dxyMvIJdXfmL58
U63j0ixqmlvm1xU1PvA9znUO6MMuxql6BCo0SvEb6l8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9008)
VN9xcEPoYqW+Kb5psPHUfkgzw1nMskPvRQuqgOmslrubLOvse8zbOgUrfppPiEH5
XJ35eCFohpgK3YRKY/DBKrNmUTVs8YasgX2IQfVIMMOG7YYF0U8O+V/cOz9oYPwl
EhIKHc+yYsu8lhlQAJGYizHPIl7wNg/U2F/d1Qoa7DuM7V4MkfV++rnICjyWn/KN
PKSof7ICHQFoqVe+SL+bvd1NQAl1DFDTbY4L/A5NOL3w44mSL5Hm7Fxx1paX0pki
4y5l5q7Zq97ojwv22cEsWs2NQHUY/y8Fno9HAs86AGu1t1iHr3W2daCdN7+Aky6w
AH/vYxYGcxPmdXefrzp3TCV5igoi2WUcn8uxgPL5sbKguc5w1ZHoytdkX702O6Ua
1D4uGqYiQ+oSdBBkSDcT6LUZRBBZBqtHytrcL2y+M5WSWx/mBU9oFFQDbQ0bnqYk
lwCNpV7HmV3i4biDAeEsi2hLLQmDKZqNTAqZZ72d53LTYhn4BUHX8Fm1TchI2oXt
harjDOnToBADBM2jWCp8X6fKTjWYkPPRrzrRy5IxMQcyslG7KexCFiLednfijXqf
ttZpn1Ix4T1Lk/RwHE4bZDidu0pafq+F0LI29KnICE4r4qz329DpRKHKt2KvpLZm
Et6kjruFwxy7s7+Fm6wTW/mJVZhEYQZxPxSG+oF8378QbEK5MhLieOVTYJKARjRp
ez3n2u4xuPTzFL+v+HlNurv07Dp+G1x7P3oAOYcDB6Wh3QvBiHYCJnEgjULADZJS
k5Fyc6hTaiNm6zbacLZgIXF0X6OEUDe3blujFW7ZXyVWiW1K1iH8mMDZoDRGiQ/9
eGzTHlLuRJoz84Me/0f0zGwkdd8qs0XmNtzZowuf7vgo8bjC3TMCnAJEGis71XBb
ssCd5dQgDouCXj7J4s7HGkKpcA7keXjVoW1LQpPLAtK+DeCawH5sGY1RA3wa3Zsm
srEUvjChplgHZ8BenCWvF7saf1fle6BAPSfQdBDteLNMhAFWDXio6xcuyHCeqw/t
dGpoq1YMATid5qQ8GR6qAjr1EA1q+dSdf14fixtrPFfwjH6ohUkMzH4ugkFLa+Na
69TlIPHEAos1prMx26RTCfkbqb1qsPcrUbn7/vmOXeud2CC+SZXqdvTUeWJsXPDX
Zgb73V5Rygn+fvafVAatIOTkDC9rDmHEpQi8hzTdy3sfdx4abia/hDY9DZTi3d5K
3bdb7/t5VNP/b6seOH6c8yGnH6C3/yMr1LjLTf38ZIHE2IMCAUYNu5eidx/uKM0s
VTO50tEPYk/zQfj016rNrrGVyTzeaoIvcRTq/CrU9W0pPS9YVGpbzQWtt/d3MkzO
olVO1E+r0nUlvlMntn87dLZqPJL7aVoiBRR0kMsICs4hqNC5UqjwAvkWi1VuLEJS
Y89E+BU5RquPRsmBucjYg/5chjryoJYE24ljCYJw6PilfoP8lmvuW2Wqebb/B3Rk
vFH1n3AEsUvqlgXzUZqr1MIjbmGmoCFKhJavJK8ykWvKtjZhzdur3tzSGUqvZQ/d
irgia+nJG4NtQ4J/UIPC0j/dqjMbudWcv1i0i/R6UknnQdQ+A379eNo1wWcM2i7x
Wg/k8t+ZoXIbDCGJVypV0GkW616Q7WowX5DYIzxp8AWADg5qaEfkXDjgeq9tbRQN
eFY/tV6N7NG21lghsxIaXUC6SlkBi7OzW5cSi1nHUvgA/oX7SufjpMn31C4oRz9i
wWtEbp3ogAWcyy8itspx2kYy3E2KdxgjfUebYODajVjOl6JJftlv+IFDgU+iLAOD
YeuxBpwW9CoVD+8ZuapBXjsSRgzn/najhXzA3n8cW3KxNyVRzGq8m6LK0EnE8BqI
coQrwtZqrxzxomU3YJtDEk0bcycH5pSNwKucR8pZD77wuzaFAwU2qzQCQ8pIVpkN
vqa8+rl1IXdMFxoyaHHqCsZKQF9CEfvkI2qC7S+1zVQy5DmlqYRCJ/zVLEgOPjPk
250Q+vr8o7ZfbVKASL+5bbJ/jdSeWLkueR1fmzg48piwvQhNZ8S+taTMCfXwVTfX
ygl9RM5is5pbfzLKHViWEsecLorL8E7pn3FynyUXPMKmzWMIr3K2NVMxx1OfuyyR
arpQfU/Yo29Q59XLzeI5q/uWVy2fwbKRt/BQ7WkZ4c2i+WVTDRJeSJMn6vIdqkix
SYV7em80lSrSfvPPbVP5ZU68soksseWh4QUJq/i/hWVJUw17OiOwdgclznEPRkmX
d81p6rX21jzr+15qv687XL4DahSRboCtXKxCtO2LUPCrbgtBQBNIS6Pk/0A8P91M
3uJEh0Wn+A81w+lRvGXV5ew7TsvcVYiyxD8ccMIBpQepq4/FXEIVY06I4LafMYGa
VnxXKX9/RVxs1q9iRmZlNhBUw/+NXu+WPyNUOdvrZz14tl7+IgESX5z0H7mEBWH1
FXoechiJXkcTcvh2mDgJaH02rrpldrrst5S+0m+MBK1PWQLGP9Vtdtbdn8UwaTmR
bF5BdPKiYzyoojtnyR7QwnlKPBTNuv9hJjRadMXTMd7YMoHiRYU1RJIoSV3o0g4+
pXNSPGdioz3L5JkrvISdZefxdK5RySsry1bTFZbdm2ZWoWDQyfuknpSdNFVXqUfL
Hw/rImzDuD6tP6j5GOQWmWt5VsarMjwGBtViIfR/OZJvIchZ7Z4X48cm0d1V/fGV
w9TvS67Sf8FSAEHrqvYqt93I+NE9CGSjRZewnPNgtIojxN1MlxtGwjMmPgpezqpi
NM3Wa6PfUfialAw6bEZ2nFxDUd1YZOFDRl37QsTeJsB2XjAbyOICJsRBpFnaMcrm
XweuJ2acALwiPQX02YRq06NxTBA9OwEjMWTtdPAGCYA+QUvwxZwBSBna4C60Lfle
GH/ik+u316U7f2/I7j9Qq6zoU55bvr/l5W9QMfPOeKEtAWUjbzWrsTVFCcaxL4o5
hG16CKm7DZW6byBAkCJ0bqnc9gZe/UBWs8h4ZhEJ0St6lfnvdWfBTtLSo1FxNpcY
xbi5PQ8ZNlciEv8bJk8biLJleEhcm3jWbDlWmCm5Rh9HggKOqsfy55RIQHm9AInv
NbTUSr0CgDb27AMCoRZas2+rfXprBIlB4z7jI1gzTdefjSYvalkB/a2FqB1DEj3T
fGnkNQ3GSObpGHdb/lOLOXnBiD9xyzj7aCRR4q7JYwGZgIgY2+jNO0eQR0KQ+dOD
PezFVEpGTuonMk9xqa8WxeFebbhKvSJdwHB2rS6f+iFFkBzC5rg2vU2XkW7nBQhH
Huhd8tVvYQvU7C/ytkES6eq45z/fDBaQTObsIY7OWdNbc2dp1HyRfLUCk0rZxZOs
oZMEQhHF7M7o1KzibEzzKoagdrbmvmL6YB+teKuqPQRTokcWCnkTO8XWx6UKsYx7
UpxKhl/GmXL+U8A8DOVaTbRKk+pemLFFziebGEEKYMjx8AFIOwtF/IxkPazd2pRH
HXOp1Nhb2ZtLDtXowHdjl50wwwZoMueaYxsQSpkgtYIqEBf68FOhu3CSAIeU2il6
TmnRSOQxR5UBGZaxErlhDD7y1djnS6hDEyGHI+nBTSRnT2Phy/oPJSu5HlzizMdQ
HJfG/uTGuDRdN3D0nbi5fBmKbHNzKR+kebYmQeHLMYky8hGyR/QKw6+Uvg+yyxHE
XOUj8YXgEOHHWqP0mqO9LOpGB0nM0L8K9t/nXRYhaJvDLAVR19nTvwR5//DhVMVm
7KDFhMeYAawF8Ser5vBKGZ8B7j8CWuEx/MEVfX+PLVeebWI/IjC/3iDYsscUJDuN
Hzd+n19qcEA8MdVIhAGxKwckNckLPOfcqz7sUC6A28zYmlX4o2xJx46Q5yf8PfM/
D2FPagenaHWb5Avypug6qXFhm0D2uSqw1hjfyxPfvr7fiEjHd+OskCpAZNdG3l1D
/vb62LeSSBhVxV6nh8Q3TsCRu4N7N19TQbtXYZHN8WCfC8hNeEhA5h2JxBNdrUfe
htL+lldP9v6HhxrTsruySBcNtBgJeLzfdL2YNYmfZFVtF9VRx0/3FrlJwofx7Bsf
K+I79dB5hD2T0D52EPq19mkWGhsbo/TfO99QO0IfOxoU2t3QnviMCpWceeg050gI
NKIvjK7UQZubxkLF2kGn+HNp3exT/6cXK5rK3FTdjsEZljE6/iiT1uqrmaBH2lhS
USx9voGpPrXLvOZNOKLuT7j8cfKsV3YGczzloeswW+XvBzmBItaHrguP6ay4clgx
QPoJZcsVsKIyOdEsqO8AqQIakpefDsJNp0IS/oXVlHaB75DwdqUr/FttzojCxy1g
Kjwtr/NqMG25rgmLFXUUkfphcw6GPbNOZNxxPcm5j3nWdz//IZz4xL06f5RvAtgi
JnKCOJKiY381ZqOrQCDNRtoH03QZMNJ05qjfBHp2hZtOPRpZoFk/GLMqrFjoID4L
DiMfiQvoQy/V7E0JFHihyc8wstA7VL6echu/7pwOU6HZ61FjDiuTYPnOWa1NdzVz
3FYGyKTa01TYZZRGIrrAlNtfqV7HecqzkvpeVkI/2F9iNiPtFZvIt6njvSnYSMFO
0hWsTWwpGHpWjV/x0JYpLHUTt7kyIGJEDIiAhNOXiePKKitgC23mWvl0DLl8gBI+
jKHkfbEvwGS0aiVVHa6BqjiR/Cl50LhkjSzkfPtB3Bn82eOU6DNuQ3xNq8mSYHwR
NRtH0QPOD2Yer76oxaSw4LkPIDyUDYVThzooJK/TDEmOQPTWkIOG5DBQ8m05NVDX
0RYPJNw4Pa6TvWyVYPMmbWIfiyE9i05NCu5v1CWEB3ymADKkec15uQTpm42Xlyvs
OEt53rSSKI5riUV69Vc4UE9u7XTwzxu8RjvAoQ9kicKnqBrTsXwuWGReTFSSa9bN
51cdgKN35o12z02V/oiZa+k9Ov/2kHeia3d0OxgnFwXqGz1Bwkn2B8ZMv2AnZVj4
olYBUgAINLiZKuhpEHaPH+d1sG8GOALcc5ewch4Q762rjBN47iNBL69LrZHuug2c
2zGijReh2TNzM+P9peqLIki4X/O5zzDvBQ7+PyZqsIqFmi/9guQFsFX0x0Mf/b3w
sWuHgm0oHAemm90uzDMHR9vhdD0ZM5r1gRv51/t581WhNo6T3wfsOCtT/qsKFeZY
W3l0YE0PQQuyuzDY0vYM51VVfqbl/FqZRrvWmmkuTtxi2HBHfL+y+G/VdVCagX9/
bUiS+dEutn5hBeQ0oPJH2siX+qTx4O0d+WKqN4LDgydhXz2sXOr9B0y4L8GRgcSm
exXENCzBe8qBkWv3mCpSMPeuxlt7ki9zf+GNBXqfUtELjlNgYWgYpZpsAdFnzXrM
3Va5SYgvq42uhobQhnSSEvv/9+5Yan+gMHegf+OOZh9MNQztbziCHAk5PPCzSTwg
TsNqlNmarPUvzczqlDcCETuxQeMFi5zG9SYCR+5t6PGqJEUZAt1YDxzPzQwgWlta
1eZ2h+KZIlWqw3YPS1uLHdDYAy1K59OomNo9d0FmbogrsKevvic2FhHI8EoQUF08
KxC+hsMbt3QGGD8vlEtYARE+JWrI0jANlsgqbgi5wcFMW6jFVtj04vwatm3RVsiC
t3HafpKrkLI5nlSFqQO7X99uYWvbE43iwrKYwscSRTrkT9YpTVSDooppkYkIz5Ja
Q9ugPYvJ5k/akVBNdvfv1IBLfMemfpgpMMCEVYkrlJm3rFi42QmzB/IWa7byET0U
iCWyrXyhAr/QeGAHubWDrLd7MPdDSxNUKY5+AGiTVwYwnpypdRrMCoLC25GSlS39
bzBFjkxjVjLbS74S0/ADEGWqsUh+3yFYU65Ck3gIbe0ZSFE7j/Zmh42YXCWShhsZ
pYhtbap+MT4byiMfpHdHJ8m7rx8k5GVQHsu7ozwpB6/djLZvc337UBY1+K3r5UJD
Z4JSlu3YFPdDsRy/jA1MryCJkYxvfCsuzo9ksjPlDgHpn0bZFAuIcX6sWOtckilP
RT8eVn6tHEQT404xVKgomKuSBpSaiHaoJivKrX18QMJTVhUl6gE/U2HL6dMRT7gh
OdQBAQgdrc0H127tbM/UwpgyrzBoKNmxBExEHuDcoVwmLcbz0gmnnMVLokm4skyd
FtjRYC71h613Wg8z+exzvw09iM3g5iF3Hex5YgVxLYxKy6FLvphfvQDYZgL+IaFa
s2yqjYbhvGaMlDIkMedgf/lALj28cJoodVNiGzKCvkn6w5CHF9xVwvB01ePa9ccM
oCOLJc8GoJEVt0tJ9rv74wRRyLXOlm67NPxpDbb96p97g/Cuy3SnsRTD3OYZhSXw
3LKGgmWiMdwChoj7yr4vbF/WxP/E5iLhwzaqKKIgFcvkXgLcRLC+lx2yolSYVu3g
USZbcgd4od7EduHoLjhydpWWhraSMBNQxrvVOJ92FoL1B71JiD785/PMnBHp1JJi
6+IHziw7IJ+PrZb5Qa4UN5EEAODf6UzcYLDlKNaqLU9jW9gwERmqFp360UQwU0WQ
RdioCY+JB0cDn9uBIr/XjJDDVvtG1QmDRbNR4iEId1n3LTtqDU9RS5co2S/61Nb/
SJo4xoURPc9BgiQM9gNTxYzZUfnI9b5BbD6wckkTFm/AYZt+HC0r4Ie+i6+rv/ni
oidQXjrVKP79NpbH9xuxZX4YhJOgH9T5r+eW/evJ/lhHUteLO3Qo1PIg3zhIWsjf
VS8lu7L/z+SKfrwJ8o98HwrtOdXKtq6i1Zm0sln8amJceo30yKepjMApfbUBteMf
5KPJUrrxYCZxK8UeL9S2iaM7aq5smKdTMK2xWKAOyPjIR1sHarbPRaMtItySxtU1
8vVgB8elpdcLVLI/WUGjaRkFx9IkukhdglzlGSv6MRfH6NApvXM/56CikNODXjKo
iF8T+n4fNVfYFOZFMc4zwnCdHbEn5bMEOUsLEIQb1n2xiaCXkqShUTkCHqzNXGXW
FC7Xr95vGX6Rwba3h7J41vyg2ju4R1qTynBYJtN3j6bmgy9aB2Vy9Dx7Yk9TsfOL
2Nm4tuCJgmLuNP8lV0W5OMUlRP02zEX3P7/Sd9aUT0i6lVtlz1CjY3phprYH1n3l
Gg82Fp2HjyycioU+R0RIx7ru5vjqcHGkGItait5RRKn8oetRMZwDOkRNCU8MgRGB
F5Qi9cZ1mjL/B9PzKEiNgeD+PlbXr7lWr9YB4mkf3OZW0Ec5QLGvD536rHeYA2sv
6KUeeWemKTP9t7L2lqaPj96lcfUmjYmNFKmF+5MNc9SJMGSzf6O9OWi5sXkWihTv
cDNVQzPfX5HbF2bRvQx+or/o1+jmco5iFh6p+GjblWfzc8HtBxYRnCLKhTmkLx7I
G/HmHztHplcktKj+W7NN1DhDybBPnYeyEYgw66zQTf2pmOVpMUQKGZwQ1/2kf2B/
nU8c3R64wgaWHGHbqEM3Pr7GgWtSQv1r4nCVmevjuZgVPV/8IJ+p9Rpx6G9VWESq
KiYk56z2FhXZXr72pcdWjWWIyk6eI0Ed7/yP0e2XsvUNku00TM3JKynSO/RZk+YZ
5xYob1vnQ6MSD0wZ0GPKvp99IagrvL0kIK4E0wHheNVY0RTbK1fu4IWLXT+DVcb3
fpBbzSuNCUevO9hxCvujweIRspG2bfhJU90sa0HC1kPEcrMeMXhg+voHSxmoBKjB
U85n+3BnfbQmZBCXPwzx9CnOpkr6B7RsVZ1uDc4JowaKpPAXUzaKlXFri7SGgrSL
Bpt1IVKogbb1x3SbgtIT4Kohrgt5vE0RDxwQMsosEDLMYWEcEbdPHCPXAAQL+QkM
rmT2ooyYVM8gNQ/ydpRGJICHiHX+xfL4JQj7AebquRvnTHXAsr3LpNnNkjQShEAu
6nOksp0FLGYDiqFsDmWdzhbFH9lDUy+YryAek9jJsp+WaW2vZ1gAaeknlpUnXz6u
kMa9r8sMnsQmpHipILuqwlglHDocP/6VdNL4TH32LRY+fF6FCuI8swmnEaYlNYlY
AIbjfTONYjrDn3i1FEihqiJQhzQHNhoZCZbOZtsdxzoA5gFZTNp89bGnZc6VraWa
uwkitivKG/ESk8p/7HPCIxFyFA5j12DYHQlK6o+JzGF1JZBtzAN+G/DStenKWZnW
Olu7uO3uTv1JvGxVyvG0pKg/pHnNXnNS1kmLZw13wibW89lI78EbFiHF/zRRtrIy
2HOIemZfZnMoml26WzWqEDYCoVMTvbH8ajyU9iC1EgGxvgHK9lVpAHBdS43MZUMs
cHjY9lN4qIZa1POPhv0xEIIQjHovpNL+4hf525j5Ta4tHI0FPiEXdFbJNdrWhVo+
WRLOROkkfT64b5z8Jr3Vu87FhnHmHsMfqs3e8vFFuwI2p6Ko2bWbDYLDCnxwYmsn
nI2RWlQfiUoehREgneCFgk9zjGAquJJkMm1IvbTpSgWm69kVzq4k1cO6bYL6vWwK
wnyPRIoKvqD7UjsbrhCBtJOoZmMcoHfjHeY1lErrrK+6aWrnZXvW9NHyIdraChXF
aYd5Atop4+p6GIJspi8OFkiuw9H6KRJLq+v3L1altuY6H3J8k3hnyNa04dsZp02g
wNRP3HGYtKO00LwVjwdAUmX7nrhW/V/rBLKluKgOqNys3qNIXDDQxGajrsOGzsKO
axvqoyNsYAjTxyPz8jJD9AD2sIlxWtWfsmYZLQPHZtqLY9/9Rhsct8H1E1ltBJ09
WnegWuXzr8rJ3NdU5BrgsU5qsMgFKarKv5FQI71PwlTrASGmO1neFAbXrVOpkmGj
pIOiXrDzXHFjFV3uCuOj4GnWLro+ubsH/2KXCAkUTMiXHS0f+bBAsdlOxXjL/AFd
1zfAPeD3WZW9MJ85RLVwwBcNY9D58a9H7CEU+0knUsg6uyUjX+aekzHHfX1zxvkS
TOsvTrMR/miRCxL1BAzbBi5bL/Vb/R4cv2D2dq9kLN+JF8SgE3Hb/n0B4Tb/7Lw1
DNx4jfoFbizjPVIxahu/dwwfdUIk0scrqI8v7PwlZzZ0juX6C2/bLyuFScd7M6i8
4iRd1PpBT415QQOAtVJb5CIUuyLcN8qFZsc8LGIXXx1FM/EnUJaX1MxFhdVLXjTO
z07BxDfkvO3r1A32rIu7BO7BDkTFsCx0Ny4raXe16CDsM7D1q7fn1iD6yrGOO6St
70QwChbPRL/JGWyn5g7Ob6FUfIPbWG/E06SlGqHuQQvA6VRXl+Xre1wlSwg01bqS
vozpnaNoKeJua4B7MM/xkDQc4Jtmw5NIQYMuTjXH+DWRsteJVp4PrOaq1Zf7vFmu
DWCN8+qA2k1bN1iR3pZHk0SGFkywE0NAKaC4xgKKPdOTn1XiQ6EcAUiJ3WCIVmso
TWN+btrX9IGdpKlmIpTjF2eHJbs+AIy5k2eqnNgJ2xj2gp2fmNXDbOnrYs2fP6vj
+E02e/uGqUW24QOcq7Cpw1mv1HIvrHSYwCFIYpnkNy4FfvL+J7npu+V29g4hGrF6
RudC/0oJCH9TyJ++9zkIcPpxR4okiiODMG86nOK2yd9C38XSoMkxdCRsnzWR1yvT
eiJwEsrOzKX62POog7s8oaFxvbZmQyHS/JLEtiGgQkcI/4s9hzaj7dtd3tIYkwG7
7BsfFqLO+DUY7I2N0RoE18dOh8KfGeT2et1bL7AZc+H4PUJbUZqeSpJZawbk+iQC
91B1cAjq9i8UOIYrroNo2IhHKLEiEXc31VnmnVh/pI0C7kZlimZEEetuC2rXzuKK
QvdF6M2eXc2JcUqvRgKPhch7B4QTAH9ayBpwLQInV95yGqHT5rcBYLypaVtZDsx0
5/wPwu4EoaVhvUsCIOvJuE/1ju6EBmLESMkLYdlzvWZ32frkTIWrNtVNvm3E0Xcr
pLUCqXEOYDkuqXfkJAz0Dm4qkcqvqzoI0RUCqeSfeZZdRUpT9yiHF3S3eCzNuwQf
SW+DN2ra0A7d3k8QGuK87CZoKMJZ10xPv5vaMhmV1dmXdHDpKKE+g9QQnDG+ISUW
lszxEThsYgJwuzRb5Czh930DxmJcyazpuuxKf2w/KQlGHf7tV5qWedyGxLHJJj8r
MjjFpvtOcAvjpDhYl3gm+MQ88ZXNq5b14EXKk5AeuhmQUQsuVq1sNx+WO3YaIsNp
evHJl+j8Ti6kceBWhysj5U0p7yxYghntkCsi+u8V9hHRQfrM1sDs7aj2AGzn0PR6
tPLd3NFDrtgPpNIiwlSh2+acnTD7P6bivz0stGglTcm7xVVvtcdHt+qRMIhUDqOY
HChDaA1bKDbfgCMYya3C119438ZMO2NPoVS+4Vh4QAR4jNX7nnE161Cd8B4JQFfr
jnIWKgri1JtdCFOXdy8devebblQxGC7bJvd97zQFeAiYbSGvA0uAVvi2aVQftVDD
mHMC5XdNocghG2lpuf+dW9M+m8jCKdXfZa9YLRzZjMlvkoQQkm49R3BA9R+yPJl/
F2QnLssDLJf8p25f52ycvuJUJbvx3E6PsgslU+OdcdEifGwunpJVCnltMPNDTQPn
AYdgLqcMvlPcsQMxCPo0kx2RqZorJRAl81W1W1hlxR+63b14afSWHIulLHvTzsFl
/1j2TsaiYD0tIjBuBO8kVMGyFsjrRZR4vEp9UbTi+PP9mBz/XB7u6bFirjiL70oX
Lz2coi1Xv5+StYnAp3IA/pKwer/Ezj+SXswrGaeWhc1aYwbv4Ahe5s97TXUMWz6u
ZMZ049xd+Tq/Ge07PtMmdSfi99BzERNrtHgGZf1nxFL2MhRjXmmMbMFjNqi7SCQK
bozuRAXg6PvH4RgrvcN6K3AczwHmWRJuqrlLmKvpR7KHV4crGkgdXORGGx/hl+LN
1Di0H0egjDkh+S7QlgXvyg48MyBf41ttUNtYZPVb2ES6CRcEoUYt1lDH8/XEO09w
rsVnHUo+h7RammqL6yDP5HhGsjbgEWnsGDfxsOJoQFwx6TkicvsBXFZ1DnrVSj62
LsszfmrAGdn8AZrzPVSjuCAHM5P8Y04bcPT40xafp0U85Gjrcn07G2CtTg7K1/WM
OgtI8kukDw2O6/kVHKRmalM7XRjAPuyGdTUV7loX/RCxZapF1+a4dXB5aLJLyr9e
vn0/GITyNTD8wak+gzA+WPs+MDfVA8zYymzk+CbotOhTtGmCDs1eDiW3iZhfkvub
E8gF9jVY1OjP6cWm1C5RsL+pYFLyjjbZOQu+LMim08kmBWTuv6hKI8lynLqoa+Cd
7KZ2qUag1k/IBWgRjEeqbXBv0ayCVXSC20nRiXgu3Tc+CIRF/c7666i3FKk6Ifsf
/SbTUvxdi3tg7sIOcViPFEJCqutByahRgubcE+qDz1dqkT2r624eZTI8Kpcqkfvx
TbYw9EhhCY+8vvws6XJEV1GXboomOgnqaC71412JIKPGb1TO21+B6DY3UxD490wT
c+V32EGedmtUQw9v6mnGk8y98J2kOt8+6y6vOx6G87NGfRs0AVxGOghbwOvmSiYD
GuJlBpN7JOMAKETYTv1UEagn9C90KtIn0kkD/+Iwm5tV596XuZIeTbhMEzeOtxCW
QuRCNIM2AHjZFWqfGO6xVKI2DfPQhnzZpO+xs8NElR+pmDkKSeV7JzyvkayllmqI
vGcIT2LsclQl2gJJmyUh0n+eytWlX8K6/eD3Uuq+0tDQcE+1/WJ+g7ugxVsLeMPX
XfadzK6GbSMrdWXsE7yWS92VnfCKYki3H+ZMfvBGIAT4S+k8QKeNTOE0C2nOsSOh
lfQsLeT0pe1kdrlisagxpZjNIo7jO9veqjydIULTHn/4pr/I5e+EDXu0NLK/jzsh
ZWoVMJujG0CNQ7N1oW02+7KxaTJ3Ac2TLdynW4p4V6H8bZ2CRW2FpPDwv4V9ChZm
yvoehR/ziMPHP98oyvJ3z7fpT9nf+vK2LMb6HoTaceMmZnvga9T+Mi4u4ePjJZUa
pmaBZD4znimYFO9YXty7f2/wB/7wuSJoOfjgiD0/Icjl1fzDUlCOzPI6PZquOTqC
hDxIgRZuh5hzkEeVNwK6KPdUk9bthTgZSlMQd5gXR+i5GMTo/vi+NRbJ5WXhz2Ta
7zkJkv5925Sl62xh27ICn8YK6mla/aR5uAUiyIVbn2Q=
`pragma protect end_protected
