// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:45 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jPIKQVzwI266sq/CVVzqdRGvTV7g48z9GY16WsAu3HwrPgeyHVXRpzId83LB7xN7
xjwtsSY128a2bFa2n4P6qvsMQKvY6YUzT4jjx+fl0tE9QHzQ9mxX1pfsDl4W3zWA
qTVoE4N2FyFdh20NO9z6ocujpNkls2l4pgPu3ciwBxQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 53808)
FCdzQS6qMmI8YfOnwgY1BXDQ6k4KgG1c6BWijxIPnaZMyeTvLEaq98S2Ai8YeH6d
0kXaE1Gr9pYpVFTKC57Ob29AWQhLC6EQuu3+VYt5TheKM9vGesrUAjeay0tdOMeX
/kTzvV+GU8pog7WFTLKkfBhWoBjqmTHM5UkaZGYoKPJQQhlNkgYYI4bym/5HroGD
YQJJiD+6WAMtS50neMthfxvQyZcQGPZWLXD14tGmRZv8GPtQv7QbdJC6arjb6gkC
pMyZsWmujfbmupUtAMBuV1M7yKZJdtF4GJ7A/jW7n05mf7H07lWD174OWV0MRntO
fm2h/hFRK2dAA6CQ7kQpYcTq6UI1bOxlqd2Edk6sQr4zCvEV+4gNC8soNE2roG4A
JeG8HGFTJEBxoZqcLwK3Tqh1n+zGVoIdjaHi5ShdoyQ+6GBvVM8jXu15fG7EUQOV
SEjqt3kcVlA6yO+o/KGv8JMOaw4kjY5MP6sjE1ZUm6kwt1Q/66oEVq4shHo33Wvf
SGd3UYwiN9s6OsjGcJE117ookkKfd3LcNby7dPqbcSt+OtpuXBbmLEJiYI63W+LJ
V+0cib39A64tSPOH1b3JAq1LWj9A7ZkqaGnPecwxpQFRz4x25PvAVPOIHsCA9i9d
i/c4JFXkL/rQnOumnpnKZotMe3AmoAq/7UkiiwDz1wQn8ygvTTwJp6Qhd38MwOw8
nzyFVpnoIUia+3mKRhQQZa6UA/84bDweC9SmJ/GZcOkGRZNjf9/BHK7kojAIiS+O
KIZwTFq1byKW3kMZAELBr0JcZbtj7pOAEEXJ7FqlRDejhDtGVebCQ9EYqwVdwQha
j/mf7emBiyrWLyEeicBv/K+ury7TAATQoK5CBs3T4nbPjPYMS/xUp0dfVzxoHOsi
5E74J/WLnTFr02WI26G4TdqZWpHsxdrDQlRnRUcp4fDroOSWK9a5lyRrONpSWRE+
QHFc83K3dFtaigZd2t8LE+CWV9I2GxuZs3cDG5gcm0VjHpO2qekaBipJuE42oDk+
hUrvAZX//NEPNlM7gosH5TIQY8DtRcQsmvyEEmQOEbz4ldm6pIpRkL2WxB4RrCIs
l2Vp6ZJahhUj0aQn2h859dLMxRaS5TwpfulGa7CkvFwe7aj9mJ9A9DgdLTudmrq7
XPcbxIhjbp6aQYgs1E0HDQ63u/Ex7UXslTWkenVx7cjVlHuJt2OiOHPFgXxjh6Nl
Z9L8B5lJNXfse7rVHGPCopSaMlLU+O8G8zAR4HRaA/G+/GTrzCVffCs3IxVKyMpL
SSA+a1wRIJe5AWLdFC8G3Vy2jv8Rh4mXW/3H30dLzQWFZI0cNDwcwk2ZMngi+6s2
c76hfsfoiY7Ut20q22nC9OEZ1TLsJUMmHNPh/2KBfoxf4B8TteLR9dL6dxUirfSt
SY6p4esSebfPYdv64RfwdbTF9wYtEo1k9KK17CJj8+2iXcNjziDrva5KiZMQBK5n
9j5OW2TiXkwkUas9KGk48e+NGVFqHw7uMwoyfG4JsBxq+hzHHN5gSVe8tywMkk3z
61X7YhrX64HoD7bR/GxwdjzXnQUqc72v8RF60bfglAdSxe7QEEElXNXOlN0qHMGw
gtdKoIAhmET8aWCyO/xR7/IJsFssSCBOdkSjDUpPG5vK+IvEKPFPnTEILLkcFvsJ
xZPHNCYTyVbVNQI/QCM5HU6bIZvYD9dP0ocZmYpdvQ+6V1UURSnD4YLF1lAUPRVc
L/6kkR20I2o3RHhYiVmxm1MBdIC0iOGthdSa+v/rDcT4VfH0l2GqjUdeaYNhrvD+
c94qUewzkw/aoVNGhkWAe+sPd+2WHBjrEB9VYHXycrm2XbYNRDXDxxQ/8nFLvpez
XOLdYE++A+i7HG2ecaFijAenX3y5LAhhoD3xsY1uERA9+sSor1zO8G0gZ0WuwtkH
4xAFSIezFICJmhAPumNJ3rMFb6awCYCYMIpru327jlqeOm/yZ2OE67JNbbhF791/
oCVUzfz5zI8j7QZmluUeSiM1Q22TIIcrP6gkDuFC4i3llMUZLtDLvjbcHmuKZ0il
DRmUZw6MyRC1a7U0Xo4BPnPvNA8DWcXaSQfyhFtiT9F4voKXqA5dYC9CXeplk8hc
iaA0AnXlngo4DkvhNRbRjk/KFx6Ezitq7EKRIyomtJI78SEEqq/GxL9ncLVYiiPI
BOJlt75bSqtICEQXNt/3u+dxvet1SFnD/RF450fsVhByFuhTr6cj6FgHetyXvkZL
iOTcBXX+S79zTAVBnbwp4hMM8uYtl4fln612OztPgHjZL/VX8oo74xhhCW0h1iMb
QaIBu1XmUuwZ/UUmtLlay5z+xc98wea7BJdgoKAA+azAAm/Hy3GNDL8/3AeAVGAk
FGuRkz0LYkaUyF85j1kC15wq7oNnXnH60b4soh5S7uLfz5eNkyXlv27/vtLylsDh
aeoz3ADOk+phUPInj7iRAcXtenKkTGA4LlbwIoSJ8xZsK3CU/2ZbsuS3Xtx+u6Wh
PEn7a8cdrEHQZwmd8lvpHpZH1XyAMKSxiJvA9MFqgkBNfzFhwkscP47NPS4Ba17R
USHWStMWFCL34M+FeOwKB1zz3pOs61+DOI81UDC7POWWwMPw/AwyGSF/f1wPMrLc
she5QVBVEv67UUV240BSQs8OJAKPnw7YzInvdU1RV0BZlVDpozQ5boObeg99Hxjl
HQZkeQgoyG1x0VSfohDIYeZe+FlNMdaBsttdvUC65FzDO6AntzA8fwa8qSnFJFD2
vHUghl9WWcRcJekUBEVmZB41JkyLApWhLOQAyMsQuJFYx+VJqXbFlcCS1kgxoLj6
sQ2MBfLvV84avgqc4zS3I3Mlb87XDCRgHbyF5CijscdzMLxLuWRHuGnzKvFtjXlR
13iAgZlHR0jP9d7EaNEq1owoZ3ccjdzQyLElkB5HIbSsnufe3BVnkn76izPHdWhX
dTGRUzaAYuCBZQZPoZxD4yphj26FaifmGxrh3y2JtFAGJL4dDQ1QPSclbuSF+GDF
SEHfWIa5lXJDkplvMviBZUn/9FwVtStafvE+DWpTDi+16qegK+ix4uxgJqh8rRcA
ovoKa5C6ydg2+3BrulbaPD+N8m/oEVlyG4sePqn7cXcC4K3qkND8rZqA/MYqzO4H
asR1PziBUQ6a99Vl6sT1Moq4JeH/oHsOPLwnoBJUv/nCv38Sni38i7vxfaez5/MH
apf2ZBbjG6tZ/am2RjlRGU7B9n349Q/YIBLs8HRvoqYkEiTwDaYhL50+3lWmd/CZ
RZYZjcvjLMb6oz44UpIFFwytTHPyjtvJhyJkj3pJxlhvW2fD+LZs+UKKn4QFvSvQ
CrobiHZMPiosZ/0cMSkQHZmHyMhBTn0Wnbz/nmR8Qqw9sAI5FKp+Puwu3ptZ7UyR
M+UMqbjqRKysfRk6Ye7RJEDH7UuRqSt+vhOq+jjTaLAcqCos8PYr1ikTY2EhGdOL
kE4fKmgnWHxFBXSa5VSFnXA8W0l+iXXqtHtaY+2GbFnf3sLFk+7NQj1yhQhYxzie
osruTGV+9LoKiViUcFSalKph0Vd8gskk5oK23H5IITJkRG7pcaKykpZiji5ktZki
UIAz7Jyhhm3RnodRd9FQTwMJvYjGqHuFPtIKV0vY2OQCgrIwZtuDnqqnVwGLWINS
MVAEWNkOD9Uv3TiidZJKxBGdAlU16ixgK5qkXH+Yg5BCMkP0iTbnv5AbUM5kyzcY
epn99DmGkp5PHguGpc//tom2kk8Jb3/cQh5on4GyP6YqcRclhQNfvYpisIa2TE45
U45WhgYRXRmp6zo1EwFAFFRhSh4CrIXhYpz98WZrA+vf8/y0UY7VGbG4c/tY3VJ6
nTrXcZL1teeHceaKaVC4ZKs7TUUhBhPdNiP5J1ZuBHCeUUetpcngYiX/SkTU/eew
AsEHSxqpkdPheRBGNmel1/NlwtAVC901WcL69tE+lAjZ8os87JTZnjUwGUdsJXFV
k6aFGPxswqTDx0cdODDG/HFv1eRh2fIl9NBNAAm64c+swSxHB3+BZ2Sj9Swsoda+
fkGHpRrkAA79Fk17XUtkBJe6BEyWbiWhpW9kYDuewB44e/keIRCPsss/7elyo8ev
DhFzLcO8FXJ+nbpXpsJjLYGeTyV3HTQZ7mcQ+3CrZ00HTVc1NpPSea70Q1SfggN8
mjYg04IBA0dGHSYGr7M+0MuI/xQccRduRyW9AlbsAh4AkfF0IsOQdfeNMITQkwsT
ajVMxVrMZ8cWk4AzdQ0PaeMn8/ko0ioLAIsuP4J/fCVohrKzzoUNxCNxTiJxq3TN
x/rEa2xiqKr96XzkfroVfE9s3E8prSJjlvFuaNZIhZslQ3iukur5YGFuSFYgT+oW
mRxV/fhDJhSL6EsgsKHUAjhSDXbrnaoPqhihbkhTweq3kUlM/B1Ovj3kkR7HwWHT
owtFm2G1RG8oLb/C5q9t689YcM9j531+uZbuEnMVmeXiu5Jow9jn0VHGPcGJngQ8
2vSi5Wepx/iiAHka+WXOA3Fsp2CUiZ9oxCSBthyOmvEz7pnds2dscx7IDo/+IrOV
QojFZM5R1Nj8sLcdycOR+mg0VFNO4Lxx137ofmLjlXPqdjPuxe3w7S4fbH07hFDl
1MQNFhyn+y0YY0pvvRqBPS4vR+jKN4Kg2i/QjGWOX9hsTEi8y0ZXJ49waVydAeAs
rv8Gqnnm0umKU9wBdKkIk/pfZ80TJ7VsaJ/jWWfjST9Ec33ZIsj9Jod44AWJ9mjt
s1u+doIK5qbjK9p6OErhxwlzPyvIZCFotacSnnEPzjetZNjoZWwiSCZ5+v7UXx+i
fZMc7qcDKgPl9QPNfc8AjEiYvTcUUaMQJEhNLe+51xGt5L+HhLVscnB56t4YVVDN
Klw36cwDqV81Nq78+TIKmBUnn1iuo/m9ZuO0oU3fC/HTBaP0HDwTfmKxSr06Uflq
+6bAGD1V5qk5j90kY2qlqnIZg/017oXEopxYVcipe4oyifiJRA9L5aJ1jbYErwHF
aGic8UBpvv3yIZO8A+MipKFScOwuevhl7yvorvsMMQbGw+UkWbIOBLSL+SZt0lj/
rN41kBTybdZNayJ8qy8X2bX5mltr9tis8LI1li+JtsusBdthOZZ98PRoPYb9GeUm
VcLFjBjx1z4f9vugOR2S2dYTA03aKAlCgSXnJU8qViif2rcxC0w5gcKQzpBK7L0X
+s+HHdh7r9zHaW+/157RihvS1rjhrgcg2BZ37DAkcNuZRy1FY6DTcUPc2RX5mpZg
C5SoKwTS+2pDzKPeVASTyeaYLFv9VCmm6QsnpfB8PY77jF42Ea99CjFhdnSYnWtv
TwpROYpfdLNWRKNsCScjoorNYxBvAvyX72TdNU6MRDBYYF52Ms3lk7KLvviIAcSA
tubVwoSjmSEetdNvbFM+KzTzuz3B7AS8WH4Lftp7wPHzu8xedwgjcjtQ1hbrnLYm
UazqdEor+iJGrZxu2IFBlKEgQxcOiHKlcBH9vNM1FGW9kgHohwDEfPqG+AZ8XRn1
U00fhM0g2rgMl8NXC1oFZJg9/DATYANcy4pVZ/7mYaZ542GPJLQx4/HtJdaVkcCr
7SrpVTcD0NO0PGKLrMtY75MkuhL9lwzNNP5Cak8GjO5RMBE7Xh7/tkgmZpXTJ7Cw
u1SSqTshrQJjT6rf0bU2gPD3W2CLJKvZHB1/f0HC97f7XlOqJyfaJnmZp5mWXj/S
mA6fQTls85KbTrbqVN/lepEn40rT+J/1OkRvNs+3xjR88tYBxebb838th/f4xsDT
T+mT9jfOqIyvlcwhA/gssCW1GBjiHyKs3sJITh1CmnS0P4NG7VPn3/edIpMMqp0u
pyZgf2r1AOIciDYNHam+ZrVgYeVq38ag0phfBoWrHOnSm13kIC6HdxbOc5FSGSAk
vRWrGvIVR+r8+KhEqktbL82NkSDB4PCefhuHhuo9EWUriIu+yKQKbzzgz17/7p1P
eA3KMttIKpSwFwUnnd2uMLViZXTcy1n3CnTSk/CL2x/04BQDgL4xJHOxGWVgqc+z
0+mMxomX5S9x+WxBSmTPW6f+X5yoS5VIIUxz/qdKRrtE6amxtn6vO4nrstJVLEO6
UT9QB4PnFcK/5gHKRS5L8GHzJTyXCrpZuPAbHGdu+wLBwDLojVhjFBq4hu0qsmhe
rEUtJv7hEpMDEwk22meD6CW+2NVQcLijwytwxor7y8R+oCEAd+Ss1VHOA8vlEXMR
lhjVYmWi+XqlMhcOq3CuAdpQG4evAVekommm+9y6+key7FPlauZyznqelhgz0OO9
u4SGz4YMSPWqAaM1tMC0nk/RyuidI0ksTcuA00ysqPsfJUE+OGqMnbnRd8lh+I3A
U+6IiguOlWb5S+ewzUGUMS70ZpBz82fbXGX0pDJBr01NStC66FZ1StH1Dv8rntZe
aVErEHPfG8B8VSJT70vH1DnGJhm4jX9RK5JGuIj31spPfofr9J9/75UKERrmoTbw
1w6TloAMY+UwrT5fV2KWnyfYOBh9P5cwyysUpifVP6HeAcX3HHtGp/qEh9fc4n+q
0oh1NYPfgi5lrHL9Y30hHUNgoML7f3mHWY2QVRQ1Z7HiwyUoGWAGs4pPuZoGV7Yg
j+Yeeya5GHtoJpBYTggSYtMYQl9RmPl8ObEWW2wk3E9Wnx3zOGFq4m5KyflK7eUs
tWWlQQhU0ZY51e4SAGOZ6LLOu5Z2hq6l2c7g+tnI05BZwmAI6DkraMv1Mnsm6OWQ
ht/ZtBTHoSRFi/obzx3OaKksN7NknbmO13aEhBRJIbpkQXTSw8syPPQepTyQMzJO
VPGvoABKXu1GBloQbNDX6+muHC6dP51UVpGbbcF1Xy2ZBiqG8spaSTDe9FiNTtgW
m6s048y2WpHIbXaW4evPmf/robvSzedyRchamsTD97B4+s8VtU5YygzD3VEcRwNt
LHN+mS6TIgDpirP2zm47lIhJCjCiEEVwUs6djwvMePz0BBfLFKdBmNJhoftLlXZK
Wgc1PWRe3xtJ3YF56SJI+qRjoOdPVF7SU0kibhzJbNWlh7Eitp5AAkwEd6eGnuC8
QG6BzKO+WhtYerm93QwNjjlM2sfFPcf3i7kx0yHQB9vJI/sLM8rhmiqd/RfgOT9E
wCSSbZe3p8na/D4Q7Obfd68MV5oaV810RivrJBI96PN5cJQzUyYMESqIzY10828i
Y00FbHbgJEd5YQQimHzLv6QcJ8UEv7O4iZ9LOvwOi7cjHZDkthtOkgAezqDh4SNE
NM2+YZCIwaPiUBgaszKeuKxQCpQsATB2Tfh5XXijmTJO2Gayi/xn/gLxXM83bwKZ
dnoOG6oU5IK6pDJRQ32zQqrS3zj1gn7sulFHQM9AH7pNVzP92LMusvBwk3M2z1gL
1VwArURzLuBC1fsnWLjydAQTjiZVzwAIc+fwP+n5lM2LO7efXc7Dmxm73C1EiB9M
6HSFByfuc+B3XiFTMr6uTH/w+sSs8q4vt8gbEpeZqaoMcQzLeET5RviMgoUzyIz7
7ycYAd/i+kp0qHmxBrh32/D2AAJEsNeCvh9DVfHg8Z5BYk2nrv1RScU4AP4wkzQ5
v+WVXlHGsBtiP2kONMrsHKmUyh8sGtgdhb7fGauSQiaDPapUYviMw1Qtcgz37K6a
nPU+f8RxCTJ8fZmiTy/WC5zrqR4b4SG9naOMW/dnHwjR+coFDKXf406pfZQwpe+x
7+YCjkGygHbg4zO+RW92anqIKYUZ//9I4jUCVIOK8T8hxBLn8fB6Us/qFvXS2016
qNAd+PTUSjT6589OskqwJKZah4+EK4TYdjINo5uRGZtuprMuMscH/2v6DrdDHoHE
Ge5ekRkbREV3roktkRo28vb3bos8Hzi9ffz98WOhy2+Jh2qhuC6lYOR0Z79EpH7J
5HiU+lzJsrXloC+iHHwgb38rxi/4i9ZEVB+pW0/YMdpzvGopeNYdpcBTIYN0rfKa
CyaQtDpIWj01BhHlzhqPOMr6I9D8mvlabvUJXvV/xK87Plg32D0A1qWn26duIFtn
uxJufk8pRLdqoZT2/YAdHgvsbJsq0+LkRmTeedOPLPKlJM4RrdTbdpTXX8psBSs/
Yu9pcDYm0Zk46xPqj8hvYbQmvflPODiP4n+iYmiXD5Jt4msvBKaMIwBaP/Wv2/SR
lQu93QYVSVb1inskVJuSc3y1gsjByY27zr5oqfNOirYtfB7pVIy+kUjG01ank1tk
+Q5X/aZhRQRYOU1nUb7M8UWnrhehV7KtnSv4ys2WYB46tfCg2ZTnQemw+0BZEMMl
HSst0ks42E6PZcgdTcm9BxG3NkQTHirtI7CT68qT5w9OLHgj0Kfljhj3CeErQc9Z
i4DaEqD/7xHF8dK1VwwiaO/3woLwhhq57aNM375c6Bd40y9Xu2oBDLQMnFcLseTY
UakQuzxmADfcCSOlbysWEow3tmkDV9IbB+AjtieUGRw22E12UTEs5LgtoD+gT2qA
PDBM0WA572+8ZaSmU98njutK3Ql/NGB1RkaMkUvz/IAklk0TgECK/xt4dKLR9VIi
ktvuNAJRLT4okKz6nV833QkstUPDzg4niOACXEBkpyRJrKv8srkT2F+cEdj1pShU
2pNnpjufNAa55iSt/+yKqZYuS/DNm2p7aom3R4yXE9kC9D2RgRNjilh0b08FFhfo
5pmZGcTucn0sqJIrwISlRyMprCVTZFNxeC6y8sx/z1o4XEUIeaXPeiacmijEFPJi
3PsL/KkWiQ9ajAbUaKZEktfQpRhKoyd5kt1b4b55F48Ekj0XLGbDehEWAbU2J8yG
Mgj6Ucw+Eh/Lf08b/+cg792NoSlXLTmobHsOM/B45yV3kLgGp21/XMf2+F5ShHjr
jCh/SZttIvgOX5jCJb6ddPcPqcSFwDAi9cDexLggmwd5dNbeJ8dGwXVejDAUk+Om
jxHezNk4MRrRB8sa4On2iYbmc2q8qhBo7Koxn5L/yLMgNO+fR607zQ+BE+/Wg9pU
o5s1VX0o3VZ1W6uTHgqrz9XldwGLcy3fXud73XODienAyvZC7Ribzf464weKEQ4f
DTzkv98GWNnuLk369WlqJQJ9NRcB1eiMMC+s4xyVJ6j+IRSI7DiN7Fb6UT75jH7x
xr9Sq4P1lEp3ew7uIYnZIFKr9malN/CKiXrfwq4IfcYR8vgPUPluIENcqW/wSsvV
lPrN6qiIPJBZNCOQUt7IlErfi+28kTa9J4g0m0LU+zItGt96mMQ5AJEFIYEB4lxJ
FNe54pfOafgYmBGHYD7pvQI3YlfTs99Qo+MiewBHCLxzzCijRkes6eEiFGlWB6TG
f/CYJBh/vxt1iHl0qOIG2Z2qU0fnEaYbSRXGu4Gzb94n35epunTM3nIwtoqqkspI
aEWSDxfkYr1GGwj5E5KO/TCks0t78diHKW2Bq/zGpms4T9qtEikb1DDyHjfQEjEE
x5PB+fnWo6bgbDpDi4lw8r9wXWhW9YtADUW5q9iKqIbrxh7MaOf04NhgO5GtGqLZ
DYATyzqYvM06WneDS0bGXMghnUFxHQv/Twaq5t5mz9o0b8uInCxGZjSFFUJ+sOp+
Wk4bXzeixzvHs/eSgbMX2bFuFI6v3Y4iiLS6NEFfe+wzjsGewa0SFQZwKjH7ZzP4
AAf4G3C6F1LFfpl+OVxftdnDcdXWlwltScPY0/yJbbus5NGuWw6N03krMCBmm3+p
gWwog7Q2V0V2GLvVxBmWNUqcDLe1wEK0lNJqnYP1Oo6XOvHnozxOwsIHdcQ2QOqO
Xr1SlsAlNIPiXYcsPAMz55QCiFv1E+ilz/XB4t0zaPJPJKy4mqf0vrzcNMHPwqHj
n0Pnn3BGYLgz1f4893j1JvwvkkHVeWz415yylxrJjY2o/9DsBo6UvwGwh73ionLh
fkbXDA/SZLmwlf3R7gg5DdUUDEqgdLjgdBiZq1zatJXi0XRZUevCwei+t9C+c2F4
g8RXXQnWj28CiLCHlKwgydRIkx3u31z5xmQ5MvbCD3ixV1QArLbMokgCa8v/hEmO
9V4uBMzRjeR8RaXxM0LNNv3rhpWiSlQRBkfR+Ci95368CLLNYqAoPqkz+IrIR23M
HcxajKz6toyRxNznB0yRNKSIkSWBxIlCNSCjTOclE0z/Wt1vTmmm0jLuT2QODWDI
RbACnBFxEsGa4cT/v/iikCduJvplOhGT9N/B6WCI2hnXrccoR6ez6SO8RcLZmMXU
q/LusxzPCqZFhcqIFJl9Em2dMUkbVhaduVf8i4EK98ltE5GFCkd2ecy9vrMG//qp
dbT1N+3JXKQx8zIKfw46X0XUW0a23yIsi5xg42gP63TruZg8WveblB1ZXfrpSDLe
MniAata1ENB+mE5oW111RynFXrc1U3C1v412p5QapKokWqP0U3OjDq+3iPVhCHVM
gc9Bk2xOCISYd+9Hv+TZM8WK/vfMOJPv7YX3GSro6ztCsW5Tub1ShiPZzTrP05oU
9OAzgRMkmNSQdO3One/7/XWnyBS0UnyBzYrw+dTlIDI8kWaWOtNJtOcHSc1xnbqw
fs7/6PwCOplcZ7Gxv8Wbk9vF9cGILoueMXByROW+unDeOgD5nTJo1Bo/+dOveh1L
QUeD0jwAI2L8woE9Vg5asTYKhLuV2/YPCjMOTztnUTxwp6bPbFDtBJjasdMTsQrc
uGblCBUzyTFSgL7McLxkTxspHDYJ2Nh2sHNj2pKyBYzqPST30EQQF4JjSGxgb1g/
W32oibBX9j1n9XI1SxaaNCHiEMo8fr4B1lORcpUS3MIMVq1GOnXjgKGyuJNm0VFO
/a8gDza+bnpc/WagkFcxGv2EpTjRKOZOqfXEtOOlnz7fyYxrmBTt0wz986Ik3S5x
Bs50DhZPvFXUMnQNJrcnx0sbJFLAhnJ+jW4VBGJr5lDe4WJjnCE9DGARoEoN/cSF
KXgHNHktNGpz9TO0SZFmkhY7uNfAGudukJPnqz88NKllZbpi0Uk5nWB4wbhGAWNB
zvbPitZto8X8CIgxyQuahdCwk85ybz163H6JBHRekVEB3YZ/2qWMLnf+JuwPeExr
O9MfD7GowJ9cW3LWDYk7CMi1t3avoVOy1M76FWyzZneuHc/QseYgt+EctP/iJ6yK
Gj+qmupMutWwrCP0H1YWEN5Lj1cSqEH/joaB1PVJFr9znvwWpY6aI2dPCmF4FXQb
GHiXuFvKMwAA3gLKlAyUxq557Mt82lnH86SGMBfymrfNJHiwqyDGPtjT+4WP/ghG
FOfg+cImRP4CwEhBO4FDNb64ILzJVhrIgNUkhxC+sZ2beLnuH31/M7tPdraL/Yb/
OEBC5EdZ0VNG6u6cnmOmHtzzrUj7LODY/Du8Pa5e/XyZPg64Hcf+Y7bRZW0zB5IE
Kn03iWRcpVVM2359dyMCxE4RaYYp8w0d839atIpP5bzVPtLn69scv8NuKuddyOzM
GdVXHmlQwQAVRSzX0dL5BikB0LrG1CJCKM71lfMyVY88LfYYIwGRR3c7k2GpaLlq
DI1is8ECNPNrCZ53NukKhZ0XfJGRk+x/Zn9kZ9ysVw84DqhsuofT+kcWNIAEpXIZ
DoMVXHMnSafDoLRzRePCDqW/Zplj2dGVhB5HCWVEvISKR9EMKhfPVnqzgekVK0nj
YLyRYAGTv8NTi8xNDD9kBIFiLtAfUh4nobuDYMC5dEphqmdotCpa9uJUxtYyjEES
x0NjzelQeSzTM8ZJiR9kKuEGTADFowF+MyQmYLZUuJC+eQAklLzOo0odpjUlp/69
mOV0i1ea8bpEdWXUpWHt5xyUmkhqO18tcRwL8VuqOvAxnBWfAvaRxXbCMXFCVGzu
MJ6nC+M0N4uVQcv8SJ8Q2PsXJ0HchPg7rfkD+xNMVSVeDkbeZDfNU3a1JHUiLhTk
Mip9xSCuoZen0D4beVy61Du+E8LfGQjweQPJc+0YelBG/PlcbFLbppEEKP+kTcFJ
V8I/z3MkUlmKlmh0XQIPMC1bj30EIy07qzbBqrDXZRJ51N2wONyPE95GvR0SAGlC
E69P1GxjnCmTsVSo0gJQoDgV1hybLy7WqzxGi+TL0sk2moAp3MWVgro6tcMwNAlx
B4GrdBGyKRpzBTlZXJiipxyqpCrokO/aaDat1klKbEYhGLMLxXfYkhkNGv1W8pFC
ckg+bDJB2X0U5gDtnmOySRCSG6ilDwCXJLcLC3c5PcaMvnZazW3+3c3N5ltFc4K3
QD5LPO3y1w4yUR2wp0qhOKJHA9p+0Lft9WpMBwdD6SDUYE/YmBrN5hHkvFDrJgTU
gt4iwKUqtwubRODGOcs9qsgW9t63IqTHTSEqlrvfFM9rH7/pNpIuJLhmi2RqF2E+
ZDQAPexDyK3FSCrQLfJICCiqJqJ+wfIJCJ7dHQiRtA0queHe5phUB44mg5nDnUM9
txfPPpsUeNUoKDb4wNuV5KYzS+gFkOAUn62yAlm8EWfgAlXbb6XUebUeWvDIBDtq
nsiTmBt/3/03cLpQoLwDKWxTgEe7ph9jJtdq2IEx1T0G+Aw2Mjqyfci0qIZlvsTC
9bMYvQp6/y64SRqtoJfhhDCmiu8RGhccec/WSP8c7mMeC+FXECJ4QcDykQc/r26F
8WUt4FYzbgMlMbgxKYbSxV9UJaS8tmTdnPQyB6VMx2H0Xxzmg0Z+rEiJYVSS688P
NmlPIYFUrKisT1cNkKvAktMSSmVTec3gwlVqUVB+Qv0blUNAc9mkBd6VC5fkvyhj
wfHSiy/oZcIqNEdNQ9/1YNpIk6QparLBqlqbp+oo9qetcJLZftrauOGMuKpJ9bss
aQMzfV7QKW9OEqZMRlMXS3dpSIRg8nRubBbnsKN0rRe7tofkMKkIthVdi1QvWB0J
Cx2BuOcBcTTMRHPDN1rsIyAV9OJ3StEUISty0ESGvD3+IvwZn/G7GhFXqA+cIYBP
BURTylpr3yh5J4ppYy5PAs6CqieZ76YHr2Z7mX4bfp7z+80mcLUM7lBz5XKxyb3L
/jdvCNdgpdfX3S/yQLMX52F6kiCGl8+Por2viqZNbTIZFUY9Nk943mKXZD9F3hqV
48p3+zm7AQ2N7wUPjssiHlBT0mEeADpvTy+3Ki0/7yaA71EVJx5Jr0lMaFl55veG
uH9017Ij0vQEPcF3GSnBaZ5hlSqNJpMvRtqiLYx8DSvl+yxCB/+8fQm3xcISBZKM
j9IXS2uUEE96oZ2OzDO3FZHsZPkiSCO+/2m5z2pk1aoknUhQ1B8kxejx60565LSU
sUs9+9XVHs+8fWl6Le2rLaom5q74qyYaFsfW1zfEoInTtN/CcgxoeHkG+uFGsnxZ
SHDFyBRWh123fvenb70BHNApwZkPpNKXcgfdsQWVj34gF7hNtH2QLES77EZ+NUgL
qq/s7omFKkb6h4XvVFmMwq1kjI1aIhW0v23gWd+1/2dFDoqXI7ulN6rugEMs4Qm/
1tuVIh/GiYSf+WTaSBpG2hOBzR++pxW7KF4frieIb0+rdLK05SFLj/MjKbAHic8n
hlM4vDZyu40rwmOJ37/i1ovF6Rv+rbZ/GjHT2I1wqgUUV3vIRlS/OXv4YS/3BBv7
5HaA9GyJkHQV6ggnQDBsW/RuKQ0IoR0JJxjVglo8vGpmIpd8hVmYMPiMdwH6EKK7
Sf3JFP9TUBB4sibhJ9FUd9acAwLh7DN+XR1XSyEutmgI2EVr8w+qLJrmQFiEZx2H
dGVXO4MLbgyY8B/TQBsojDySg+kaqgkTiQ6jyQPjusO92AikpWTIKMq3u65Fo5X8
4LczaD1oeYif7DG7BhTKIfJx2Q1LPXHneDxy3PVY5FFi8rMiJg7G0QsQhqDqFjwp
a5m9YpeKEeqOdEyt4oNtu7p7ZqpNCIIhPa+5sZaJfXG7QVL6hmLv+YZ77FxytNDu
BRntFKV7RSX5/+IeGagrhVD7TClXnoJWZUSKX3bpAe8POzZiz6sAEAEKbI++UK+M
Lw7DQoQLAVKdc/B5tlzUM1LTrX2bXPpymqq8AFV9GPNLZj+frlPELrOgGq2oJpL8
uloPvDtD0WDTxlD0f1VGGb0aryf2A+Wzf444jy1+QTUVRJ33vtLeKNp8hXEyfqXt
42WSWGw9UyrL43yoB/YEeuUZlnLZi8ajdVDpbJcHqd0Vtv1E7ZldnXLlNU+UUqUl
nVBusLePHYpqHoNWvgTgzdt3NczSThvCyexgjsEKgVgb/pcvDQ4dCjx6uYnajEdG
tP68gaxg3zqa3UP7/2xdBFyy7nGsifNkIFf+GqITP18g20KIzDctn5rfFAdFFDnL
1S7IIM73CmXIjnrwPwCEUuiwQtDqAhwNUgND3PmDZMYnQsrHfza8ez12mfgtcQFz
Kj29QCOa18RbiGdzOFIiYfbHLnMjRPh7XCOHewfUmWk3TKH4PC3Ve+0he5RHcYpy
GYnmPNXhc22Jyb7f7gQGiWL3sGDMbT/zEv6VwiK6kn028B/zFaleOuV1YpZPt6M5
RTSX885geRbS/E2ysrEfnl6pD4u3aBlpO6pvx8MnZIN1pA+HdVL96S+P0MZQ6L3I
+BhHGI3SwXQWc9kwqF/4YH3VcrY1tiuXCDBf50sW+Pigyvt8pNPRCBH4rDm6f3LR
XyT7DH94vxdM/2XidK2J+PMqSyKulenU1M1Y5V8OUKNieNxHoR4YxcqMmzTnHSvl
eR/tflTsBaD/yEA1gLa6x54Lz9z+TjoDN8R44yqy62jfN2/TYYX5LRC4ZoDFFm1j
gh1tN1buov4gX5uf6rPtdp7Sd75QFszoCeNacc38EkGPL3GYmxIvn18368K+hhG+
Z11aVcOQncPdRUNPSruevQdhEj/5Mk410VVD3WRrWD07MSPJYGVSxdkImPsNux3e
0APPamAMIh21KwHWaaGqUyw99Qr/bf6wtmCIstP1a4RXhAMySmZc1HiPWZrvKmlT
p6u4gRdJpd/ctn1cek8Wa31nqrpB3UltbEDd+YE2aWAerWK10MujlddWjPVrOAxD
Lcj3DO7A2dZTWd7aGhWhj/41pGoY7MgOz4Skb/WmXO9r9uSr45UUWRfR6lRzmpPZ
ElAWv3gMeSKKPInf9ucoNpWVkmu1J7fHpeWs3SroqzlenN/LnDjPYyPfPn8Orbl3
YEglaOueQiglTOzbkB4htdE8jWTsy8J+B6EeB2DHU8si/lRyeCaGFnCYITjDk+6L
P2qOCWJ/0J1qX9e0bxy1EcfuBat+Y7xrBJryrEOeMy05apOZCeOGbtn526wNSIpB
XLnf7DefIAOgADE2V92XZ8uxIFVdDrvwZlbwPbCoIOXQ/Oxtznu+4K0QMeeUw5AA
af3oqwU8bPsG3c3O+BeuYgxE1yJzFK1p0LiG6EG6tkjtyR0Bw/YQNwPTxHgNUT/I
shCAGzua2qvzknEVW6jSa4XQuc0J+LSPqrFhYQm5N8gjwsLXPrc77vnZNBUQZAJc
sGFazfwePxAR0wnbW8c8JSE9y6cyxkdIPT4C7ly8tMyN6o2g2TH5Ri3YGElGu2A4
ooXbRz4nBJd/mHuCPaCbYOjB098LiQZdakS+mE4A6CSToKATf3J3IkdgEVqnmE/b
e+lCxqUZ7i9bQActcIBfRr9zmnO8i8/FUpeUeGrXjx/gGYm/RGu4MWLYjNCrp7KA
/1H2ignT7q3n/1a+0h3TJw+R6acMgY5UPkbzj3W03/VJYSMSaIMgCGimfKhGY3lT
LmlPYw+LkQ6+/kdb5Mfx1cE92L8njJMEibBp7zipZWmvWfxcGUp0Gv14KG8G86WH
r4ezYFOB338gY+msa87RaE3rZ5lfuai6GwLmsvwXGXGfE2ccLO8uN/3ITDfVVamz
JKHTXNc1fGub2siEQQymMDKd95Zsh3n4k+ljwCmOB/B8rgz5l/FZIpurCHJklZM3
5OEBbJvaUTUd9L0aqdtne/p6UjnjbmVwvX0vTCWsJ8fmcd4r9ejoJlycOtLWjsAE
LyWY6uZO9yxBAWBhtpMuhV5niQ/6E3AHZ/pGBbF/XTvg2uGCRACDXy58+eE0gYRE
B7Divc8WS+/A4bC+zOl85q+zp1G+9O+y2+FwxpUXrQ4ZQ1+DTsTC9gZrQdgYmPMd
LpdlVU5NQ/UDxzdbwhM+xYmpHcr5WcQ4XwSg0o/ayhWlMhFww4YAfQ5PKkTTib7K
aSde47ZuL0ENSyI7XpWYzyauY+wN9h/pzOtD1x/SjxaB+yXCIfvO29sG6Y+TVhI0
P7gXjfM6ofmbMryrvsHKfVl9vvX0d9aKJMRDUHtq+CPMz1rFmt0/TibO1nMLd2+B
lMEOM43vuWo3pfUKdbEV0lnZNM1X9w8QhS7BuB6J0+HgoG5CTkthTOm04DcJskBU
pKzyAs3sMXlt8LaVGpFHKSoc+Uaf4sHru6gOG4KvNjZncVXZVt0o4P+7ri+HqlBT
xC0ekXJNbQsagL1DXsvmbrAwE0Pusc21wANnOrb8BhhDrfWIQ7DPIRd6+yo+cAO9
5at85FcbABprolH1MrNJ4cNOEkjrI4QsyMvwME3A+lw3xU1GN4vfZSX+olgRjbrk
X1/x3jUkUyP0VZSOvcCYeo/4PYVsh3c4FQMwOybZRbYiShfJ0Rm0Q2IyEL0jN+DA
fR2Lw9HGMzW2hGEEorDTVZiNpNXNfulBoXqzr6Eo3LP9lUog279/uj0OUYl92zat
vaDgF20R/et7FeEw9KXG9mmCiqNsarIbKLeOz0tbqT5+YvNnbp1R0QkrQShu3Z1P
xmnd5L2m6yMSi7rpSYe8Ck3jn9DfwiDEYXv6DSGaHxE80yo12a0DEtPG2W0RGMmh
iqFXNQ4XcehVnYWTOuNv1E1bFAs6LaE8JTPjEa3xsG2iEcZiJM44h05ChVf9rJ4J
wDmZvZxG+usAQvU7YH5zXXZgQK8RBfY5tjO7RA30+ZUy4ogkyNAnRBN0AB8xvpso
Yp+YAtjnfRaKStd4o9pKEuhh9jy6AKoIYNDxwD/NuZAXZhVD0k8uYNpNwM5cEY93
6Ib7ZPmZF+2bleDBXQ4sDq2R0faLN2CCcwO50YuTKATRLaaVxo4yrfJB6oWyNAFo
fOXJ/5E1gRT528Aemctt6qGJ/WW0Lgcc2VToItKN7ghlGmgXaL9dtZ3MPTOmtVNm
RAspmya8nt3dqjlbQgN+CLaAvYM5HEZTNasmOOB3rCvZLsEMbzi9qsDkbYSgdpZ1
WH9z0osYSV5yEHEXMjkjeOpsA/Qa0RKpS3rIaSKmgdyyo9/CK4BVt5/IWM2wGAs5
ckknDAgL5H2rGmb/Gwo15jdx0t7Xl+n3CSY5jmcwUafBS50DIbKm01OYR9JkCg+v
LAIQ0Xa3FjtsC/3wyfYh9YxIVfcZWKjr41dGcNauuD79cRgufwTsKrhBUmACzO8G
ftbFFGftaEQ7FTSScGIQphCryiShDLhk79s2Xm+qy/GUSDusl3iMPmdm7Pl5b9iL
uuMAvRktQYUe53+dUgcLtDz1Rq8sP+jPYKUcIYhbdgeWqdhPf6j+hSe+vasj7N92
G1IkmeXtDeMO8gK6qXeQMYUgLTSnY/p1K4HlZJbcVv4d7Q8aDTLi8SJ3WaASiRLb
CcvcZvzwT+H9sMI2WG++HksyfshPLWWul8vxMFUKGm1rM1CQGwfB48QNR3HR7yUl
V/74TAq1O/Ojh0cp9rZTpn/PUCkT/UZuIJ7RFQ47dH/d/H9nfSqukTdXqaz7yZMO
9YJUj4JtslS+iwpH//+wAir+KaRNLfYdlmVUYEbuD063jhQuLGjELDrHWtXgTl75
wjPHVmMa++BY06bKXkgV9mdg5rCSd7xEBBl3Eh4zFowK24nO5HHKm50FjFHFgPeT
GSZ/9TFsCJoN6jfiajzlgos4g574WIZQquPUT9uJZzaNvZXOefkr1fMGPkxo2chh
pjpvgaHmpKhf6vFpAIntuy/Xi34OdPwWbBnlp+BF//pThzqF9Nsr2TAvJyhGBDhK
5fUgO+8rUzqI0qykjpPKIs39T+ILWLB90oHDx44pYz/l9b52u7IZ1MhkdAf3zWl1
iRZx1izDdOgd4KLxSQkRvuUJigLX7MgjXPnQf1PyVeqZqVqmfgnbeBStuqV6BXJ/
colwFZI570oEjCq/bOP2FHJCeMFAMV2ORCnPpvTh5JsadC4gCjhNoJGCuszIXH0F
9omC+c9i/21RzO7yZD8ieOSgwSttPrkkkhU6l6G/Q9+YEDxNAa1w/nseDu6xAlX/
y4r7Re9nJDk3qdDqqlCedyR36u1DCoeFp9qk3Ei3/NTyyANrO6dTYENzHzXOoL2K
Z+rXzIqo/qNiApQIA2iD+AO9v3Ji+tXjbYxEgDeWailZsYfupZF/rfkPdPa2t8Qt
lKRwgejSg+kp8vu/wKPhxT6MVBtrzIj4xQkuDXUYHQcss/1zAT/W7cko7TphPQEg
NKMR6WSHPky2Sg9xY/NgcKjEfpEFUQjHZE+tT7u3TikWQWZ2MB6z5PXt5z8Z6r3k
kYtZbd7CGG3tW3gshEDe0rRqEHzC9L7vOFoYLWNRmPfUiWtMuWxaj3clpjic+HOo
/ZnLCHhY5kedo/Cqt4BpPwtp7Ht2UM0Sj+SD4ZBFlLTyFVt6+kD5T+AVUMYRaX3y
dlWT56NTXp7uAggAu+xegVfFSB8I9YEvJHqkI1j02p2F4Y7rAgVcsgc576jgm5z1
ohrgar4mAVi0Mk4xLr7WPRzetvuI2sSq3jQVaJkQDIIPptR8C+fZuW816ywrRD+o
rznidu4qbUVa3zt4nQnYd+Sb/N04agSO0LQROtYzY4eTOWu51F/agionon6sLtSL
l3DodPiaj1ixUneQsnbrgdTsp3EZ+an9pIGnSxaEHPZqjOV5RTMe56G9kIjAdiVT
DwD0/RAaV1Su7RIZAnryKSykSvGglrivHmbs3p2UnI+DreyVrLYC2DZCdf0a5CZ2
TkKYkZ9p+SBBrbgYgDkXsOoxKc4eK/D4PjlCOlSuShSIgipVZK/QjxO2c5yalrCC
i7pCUZbij8EdYLruDwk+eFdtCoMsnl8A4JzQZrEy8hkzzYn/3+kakQoW4aEiyCvH
NPCaC2xfhqaeUexDZaYio3Mi83KFW6sgbT6K0baMJd7sVMh1WSLZfOC/Zi9YUdq4
/ZVFi+lasyuYe+LUqCDCNItrsrkzN8zGgQTGxFuqk40pxj7UhpK74Mpcg2Qhdqq8
ur0l5FWuf47sCsxSFCq/7oybnqr9usmtxJREpIQPMrQaA9xPSeBILr3AhgY/dzoL
PAnRShWrUR3vzGJRr7ytgYeM+Abo2kyoTRQXgl4heG18sRPWqvgjHiVQQSmbGe/R
Hehucy3JVs2ex3KIfzo/9s0w/Qz6O+6kILnhiwWtWsG5+LjSD4TZbQLz03vRaCnH
cFP9LakqetxvaKZ250J0JtqWUVtNk2K8bXcrFHimrjARFFYbqZsRYU4sIJLrFgh/
ymryUMPJVF++e+uTrx1usJBlrz1f86ykIaoEsIieetvGBPxiruFLEmj3lSXWZkiE
enrZ6TqlStNs5RjEijxpxjYnUcgfnp7Vz6TLx4oexfAd2EV9PymDsg7UlkonZ93E
s/UMsVzY7/1N2XlbUIHe8PteXrld2hfnbyvcYJsW6ulFMPnhzECaSLpU6CMDNXZQ
93hGpweRP0PcUQMFgOPmwmTAoFmp6lDZBrLFMgw9HskbZAeUJwphiflG0Nt/Xm2g
8WwjlnhWc1KyRBQPvojgDSxprTldB249xGejm80LZQKiSno9pCJ2EnlqMIYt9OyH
FWsMeaqdIomQJ4jGstZuhSwKM2tus4W2DKR2of4CM7E6VRL9D22YCT9xPPVRz14q
Bhzitw1UwqWq+AUizR+XK3+9Ef1ucZa/5WkjUTzlsNgk/U5fXzYVDhkC5/UQQDpt
AndkJtgPRux55kPR8Ym6RutX+gMFITMOCwSlKQm9MpW88c5yBozEGJXh0FCRUtbV
LPzzgJJWwcE/6Ie26KeLDuyuLVVVjCmbvtdG4486iNmOIFGNTWFjA8j/vGkIJCBw
Np74ruWm8tM+RsZ2TgcM0jiH/ff+9gNk5c5aLnfuhJlL5wyh9ScAwdU9RZgAe3Do
hrh/u8FLGppYRFLSQZoo7wYk7bawQ34VDFRoczuFGsHnwpYiRss6/XIOBXs3/kwZ
lWKPVXDt5a3l6cGlvLttGmK+6odHLqO1G/Xwr2I62QQGz05WxKPSqphAfpudk2jb
KlewYmGWuvSb9sFCwnC3C9jwW97kPU3wwhdTtYG9K8g3mzOVDd/b/msk6rADLgby
Hv1ykSdbHZnyTQnqt502bdoG3liGG79S7zI8zjCPPdMtOlXsBXsXfnrt249hq9HJ
MQRC2GmyjGJtQZzuQgskjoM7CNzGRI9ztvznoIltIxU6TiAFGGbljHIyfWb8EHFC
7rnIK6wRTQripzIuGc5Ra9hEm/HVMo1mW1SxRbuHXpiDJh+Bxmra6XkPL5S+vKYv
+nzKEgS1emly3f4LFrgbnnfwSUBRsng7i+aCkKLkCFKKl/aQOI+t6Xap+1sYbrlH
Q9KvYv3bz/qG73KGWlaK8cf1d5se6kKxmtK+m9WRAuulU+nJxXk6UpMWGRuhFRZS
3c/lloOQln+8VMIi+SaMe/tDAf3n+9wa68zeo7MMc5AMJykvqUy10TGhBlPCg7X1
nkKLdVbw2ZbXs0eqtpBqC0XFp5EskBfCypHCVHVys7iBchn4W1s+M4yO7tQcLFk2
vfOg0pBYWdFqwkrrw66vm63QTICRgglUQsvMt9V6b/xg7lquEZkGqOt1JITz1nbk
VKXd0+A2CBkq8dqNKAV5DgWHcSuK7KoxCq88+ECqePUTN/EYEWx839gOuDNKpvGh
3+2xjjrI8tlM6SUEE3hHew85zop+95IhpnANLVDZVS1HOI5Kfj5DSONC2FO3hY+1
q0MB57RuJVEJyF6P4wn5tTJm6L0sYdnF5xZoGTe63i3BJnZIJjK9pJqJZDm3EhW4
Gx1s9c8n8zd6zdXGdVDzeQZNQHW8QpofV1a7WUpFW0/MYzxtoRq3C9jFz6VtcbIa
AitbQmOBiZcVM4mibGc2hvCdtRqyUt9s8PQeHU3jFgA1jInDtmO4YfEqJIYK+EgT
S3XGiLnpnn4dIug1K1bNl4LkPuAbAfVJ54XDJMVFGWz/5/9j9lKLBr8oRBLYcVmB
VhrmbUAWywf0kStodeHiUmFa4/aMGfes8OIqnz2VIj/wVwFyqVqhqIzAYBVuVW4u
04qLlB84NbVWzse9IxuX0jxzptvSvYLWUP465oFJ4OB7jtgnXLCUow2t5NkOy2+4
2U3qpSEZyN78GDygZCxIOqOi3y7SspfpTignAcZmS891babqn90uVEKKxMSWCzAt
rUooed0kqfDqG4Kcg9bSdtKYVJH9K04fY8hMGRdrswaGNlMFj5NFOK3iz0OiOt5/
MXZMUu4x5dfSakvu41AcFNhlmZA/Y1VruK07Rm9SkDW/abRz08oHL6MuZ/x5Qzf7
So2kZ8/m8FkPvp1kNTy+9FDU3jyKoLIk5JZvmt9FrUwMK5Jnc+26Z3v53RfCXk1y
nqIEyhTzTEAa6ShmWoWymfLN8V5crUpv/MOSjHGInlN3I84pfO6nr9rg4U6wRDq4
KhOhMN60hw9SMkLaaiZ8Rw74Z/uF9y8ucexnBe7TlqwzARikTrUez0pbYGHVzRb/
OATe5FWFQchBg1KLQi2S7M0/rhzVmYkFD+AMJro7p1zIxiHh/R1DnfRbiSiFAy2p
B15T10/LAFup8PS6tcJFntWQsbd7rnJ3dTVyzkrcJ9AS/zJz6IvD9amnjqfJS9j5
QfTkG+etfyv0PKCvzv9VZh9P/8/zKqKQScPtuK/FpsYzsCoDoe8IkVNWreccP00P
nA9WfYM68L8aVLM3S64KHfVKx5BeucQjZyxJOjjvH3UesrtQzM7zsgCFv3D1RRlN
x2ochuS9XIWlDjd7yeR+UWiM+qq+vofbgb+Hg+YUaTZfFi+FQVSb6xoGuawlyxBA
4FVvRuTrUKpIfAlvL3pHRS+ceE5Q2z2nAEmQ0QCciZktY4nwue24E5LCnv9AZDpj
4TRIInCL44JM6gktC3a4GMf+tZGysNZeDrgIWkzheO9ejs8GJo3R2pg56RLlf0tn
Ds9/IwuSHTJkLvuaxxgXy1HgYIB1quSAfqO50wwDPYL2uT+0lcBVLsdXHPm3Wwm7
M3IUsExm/QBSwUu0jUXYAQo3Bnd19w1rudjEv0xUaKgjE2qXFHjwZsMuGwkOs+gf
MczpbJoDEQRrH4JPwilKYfZcJVBiQJw5rqDXSqcF23GR9KGc+fplqtG1oDlPMclg
hETIFKDPNLgGrdtR1h//lM6C4u4Tox9DnnKQ/mav5ME5Hhv4qnhXGmZVpMqmr7IB
T0aGdOtyD8Nn5mPovx/HzavsffexfGeMvCn3J7J/N/dCkGMEsQeZ6jGC8KSs9ctX
lNS0QDdM+Giws9XbZRq0BrFK/N39ZmKtCQNng5v+vUrYdXTUWQKN0cIk+xoT4wYl
JT8vlOzZb7eDUGpGFluZxX1thChqxIx7M2Im/mGWvoNsZLhJi3DQWk/AnxTIxaT5
JM1xqSzk4oH1yqKYWq0XILu0MpKU1FkXX9QvJMHPvvTGAAxhX31YiK9NPhr88ZdJ
U9T1br9GKxZU+BH3cunYqteK4gs61o9Q662i5k2P3FzpksirwHO8unw6Kv9b/aoG
uOC+iS/l7wBJzUnN+zG++DNFlcAr/ut1Tqi3Egtg+nSzHeasDll1SisMKBWxKvKc
mVpnHJXL/xgP4L46SFRAdkc5FPqKbnFGqF661dSf4LWLNlcDtkCbBFZqreGqK21J
ZlLgriIFRn1DIp/x3Z4aujny/VXV8RdkxPeQe+W19pw8Ue+dxNi8ofLPCEKvQwQc
AxS5BbdtoGnKNbzDfXHfPi3v8KMRbra+RGl/cJyoC61kzSb7oeCBxmEOlGp8wM9y
yTMrdTkGFulw7SBXX2VRhA1BW6/w2xsS01OOQgfrzp3wgn+A875Tfu28n7ToI3pf
RrWkuQEb9ZpzcvSvNi5L+C4RwsZU5VFgVi4CSqNmdrXHMQjgZmwHkd/5oqXBx6N+
XB3dmqqwSxHg+uT0LYFCVqDsE8CUI3xQ9jniBXZK8AN4YG2WDNMhe0U0EYhxHba2
I+M00UO4s2rtR2igPXMeXYMrxypeXpKIc+HIFNEpksBIawRX32aF72/s+2u8f6Ik
b6r3DQBddwVCpQJ1+M2YLuyHtD9bCanqDTNACG4ory8oLrkYK8mAWmN3WVoyX+AI
/Ls/rbQZFBvy9Ph8a04o3nAfNIuhX/58hbK5DmXo8TrxZdCRRpdF3H5LGkMeUlOJ
ZpUFm8wozPI4X5pNxeX7yKxDqq64TPMZIK+3T8qR+T1rvRpaL8DUH5RMd5oZGirh
rJeSjN4NJcFN5/6WuvOEwBmfpIVGNjxW0qwxzQxjjvCMiKBX9os8E7gFdSj/3q34
gPlWjXAW0Zhx0gG5kXJbCJgJEHz/I/1YUEyf96F9rrryr4w+DrhEThNva1zJtQsT
nQ3goISG1coV2dqhhyD95rJqXJY1M+nWMxH8RGB2uO+TFVkctQibTWS7w08Kok6f
Ft2sbWILqg9RCfnPbLcF8eYFc7cHdDL0BvwN6HprYSS+JXh+TKOYaZDVrVT6UocC
RzSCwJ63ks8pzZ+XipFqqXIWF1n7SdviO1ZZcKN/SF0YjvaiK6XZFsXyXV9t2mZD
eSj0kbjFg8TaLEvxG1yHdz7XFLwtsZy4jg7crryE8t+9IXjHuX2CRvI9hZkvEQuc
/UebERuEWYWF3nx2TEA13SFOh/YEwsidQLWeygpjJXSUgs1u3mnV7SelGEqiuWq2
CmpW4lUkvnaP+nsGqHqeRexr4Asp/5bPfhaEI3J+JjwLMAdWE1ClwzMkv99ex3Jh
uFRsjk/INN5zdhp89gSGrOdtrIV9KAT/p6CBO8qxnp+BiAmJYPKX95goGuxpMLjj
48ndwS3nMyTYfEKEcPQ4oAiq/L5EtP94BH3q6rYZBqX8NQuaYmx75eamrDBwqmD1
5H2oLQ2DYg90d88B3KwxiEtx7RxFXIpO4ZklTRA+sGir1FHSNIzRKeKfltXHa/Ka
n4XdwFZGDkUFmXMiLLYz4kCZacOBzJWH1bQgmKap9EOE6Qjx9Grr7PMy/GKqOaub
8jn0IXCb1xXw3Qv+8suQyFytCOabKU/NnV4+HJUx48hqKG69rzj0zRreMRtsMRR1
LFrhpC/SsD+7u+41nMdn1ADaLliI1bQ70H3Gh6D8qesD2YOvm5HsI06jaPwl10HU
yOnPcEtGl1l2U0ZGGNj3abSkoIXwVV25ZIPcyMPWoEEqS+RssaD38uLfyhlVNeqX
x9LsGGvgi37v33PONFTGMzyIxnwwzsqFhZthkEtXD+/OnOmbt4O3qpEXX5s630B1
cXPWbNd12kyeGZybyPVgcVKW8JreayZtqIhcGvEKk91I9WBN2fW5WLgYpJGsXVxz
Iq+cn+31/VBciQG4x6XlGbJiEMJmSTNscSuxW9lw5kaHvxArZaLeN3Ozsc1+gc7R
vFV+z3gyQ+FeaOaUt3EpdiSCwn44Msh8skJMQGIUPDNL1pG+f4G7jvZqJnljCf6r
4C5UCyvxRZoPIJjh4PSH9gjqmllDkYQfRtRcWYjsetjNYkJivqaGHiaajIhCV0Qm
jHBiDo3JBpkK5lHdmdlQUi747yVDB8cnwh57SIzAzhYZdFjn9gk7BORuisQ1Znm3
RrYY/wknu4hMaMs5iguTn7qiS8s5HW63L/pMP3DnYHrrkUARsQnuLqLDCqDWkUVT
irGM0upkDbCV/TjFKUldJHAWyafyc1pXPUbdSBTutdLfsXL1XnOs89fpnSfpW1vS
w52/n6DoGF1Aphqk54QCKTM5MJDs5vKIjuAp6uSkCxWcSPsYMMrBGPdk4CAUg2Vs
NUxn+YPiEEc8biUtLj01A+QbY8/Va563V7CSwlJPvEgO/AXjVK1PrjdL9RRhxiIF
Rb/Pq/W4o9FYAXdVfJRmY/OqVjN0duOuCzoh3k8c6Hjt8Zxs5vjCSLftsZQk+9a3
YMV6wSNOZxN86UG2INMQmm4pFCcANlNN7P9waCYG7mW7RS6f74o/1hec0vjZX0Yq
EwfFpC7hdihhUtR72o1xlFI7RgZNouLuZDbIc8Fa2yIfbDKLZ5mKf5NFUaiu+hwv
NZrr+T5uXOeINHg3zwqLIFNgi1pHRhqjx287SSntUbdVQuxEyzJLO1R0xx/jKuyi
WxzLy7C5Wnd+Ckh0jy89bhtwO/h3gZW4Z3L27Z58e46VemtSlSHTPsp45hgq/aya
SvWfPG9BxCvsgcjBvemBDr1gTmHakpuX9XVO7m/+hlpxHs57yQppS/zt6V50ly7m
YgD/kqo6EfxIZ8xnGpXXCf8YQULTBn6DRkRzfsGIojDUOedzGawydX/r0C1mJHWb
g2YMdSUKeV5D4cYD6x4l0bxb0M6haCvf33dClVdXExMAZnMc3062cY+TIA2mjga0
bW45TtWBpZNKyKgPrjzouNEOXynDYFxZ8PtFtr2u7O+pHrdAOsjDLvUBZVdKB12j
9p64PboAH5sX2QbM3O6CiKyjViw8H38Cowttb8thaNNtWE/hMECh3WT7tqgSc8kT
E6T7xNbXcEKdls3GfBOG/RXdeiTNNaTFfchzzgzt3Rsyfpg5UrwRwFS/d2X+RIam
GuW/q+ZZ+4ZFpqJ1QrbOI0GujvQRIK45bEyrsoMUD+GUYJFlVeIIqwtefqH5fmjN
8nxZvr+fkkhhgbie897gzp0WRkeIu7oFi09FWG5ZbLglN/kV8tSTPaNvDA8whWwr
N90794tmzAC8zcwxhf4yHd/2qgUJAw6PFM0NLBune6TyIs9Bb5jdTRqVNFI/Rk0G
CC3ox/ZuNcMZthA2Ut9CU40NX+HlXUUpm8Kom5MTnpSaXX99iF/CU0lvJhUNlnhJ
tm0H3rN96gH7O1ZD+bS4l/2sYIFp9+G44PqIP6CMOipW7FWIevR2gofctBQ43GMq
DaptBjXeDfzns9Fo+WdfN8ScI8czv9udVJth2Ouj34t4lmdJ2M02hvFxFsWbJKGl
pd9g31Cqx+Ba8Ci4mNlgI6XDeCcVI5OdMP3iBQp/SxNx1b/5tLPJADY7+xPAj58d
2C6HrpFnZIRHCZ+7VCJrq09Y4cKcTY3IwbezO3WzVm46jXviOB2Y6/t4q2EB07E7
/xlJ6leOAqT0u0aCPQGg8vdjylcB1GjOYVXiRqbbxprtYP4E+9MbqVBdPTFZ9ITp
w4daRPhVoRCNvjPEaVo6JmawRdohjbg8EpT9hYRp9GcH/6ZFzLk3CvAB+GMLa613
vxrqFxQ6KlfKQCI+96LKYAui89SMmsnEG6BKk4IEuXi2wFJxSHh+YLhT7RNMPxFG
ysqFFxJkOoZcL7VlB9H0GKvkaOcR4m7NuyRQc/24eaVM2vIpQxhPUDnT7F0h6/Uv
rA+o0Gq9a9V+dNh9qy2YM+1TufcXgm8mbCdHLGdj2dobR1uowYGvV8v2pHV2ar0B
pl4ktMSt/HKuHq8+V/NhSBtmEX4dK2jqXjYWahR47QBcz7p8tnRqGjIjRglC5CWy
1CXvqff1eVcgRqCQ1ugLz9ObgyrIGGEfg/tYVyA447nQiAVo1lT35lW8slcipZ7M
4y981u4YAmS5i4mOiO1/iKA8P3KCWcTIoMp1XVhLw9eoDQkkHgw6nicss99k27nq
hmymQhTmiuv//joRBHrJC6dnJcQ3ZNqXOvSpxrn3jatEi0+BMdLbuFdvNebmzewY
ooW05EgnngxyYfiFl2LMf6rh+hjMoPr8zaK2LTWtpdjr53GRSP1Ed0vVq/ZkFFRO
Yc4f3n1+7yqqkPIdBrha0n/sxq8rufeEKG62w4MQH4jq4Q417bYyy/9THXRTs7D3
gYaqAfR9Xm7LfOfVEvkcqhlMNuTXvQGoRbMJd4S37XqH3IrtH9VEwuyQCEue0+57
IN0B4090AHC8EBKv0beZ06G2EBq3OpXg6FdecRyBMt6XNueolpfVwXEhJK0enxov
ljWgCkTdY/Na4k227fWGUSduZvmLr51axNWQ/DDEh7d06cQ5UseP9emrUI468mIK
6AAZH6Yo7fqHDBnZy074gRkk/j62wZ/0xluWZZDWosHQ4pSjBul58PSMLrC86QZX
uYr0FWQHGYVYOJYx972t4Zjj9rB4OD7J7F8+9Pmvpd5eTNaGbW6V7SB7jRgnKZmw
tPH4/abfpivxtISWWJZkMQ++uUjazsom9Apl4oZ1GF1MKaSNk23pVwkk8egs/eiH
9FU1tQFWhPys/xO/ekAS3sO8Ye9wNz0b0JosKe1gySUfhBzNZ5Yqo6brN7dESpIt
nPLlTIzv/0O0XRx4rPRY5U/RiU1tCqNVP9b3XClSaJx057WOLxEkpsrHqZ7XjDrS
w4HVOUhBDkaAejhwnJDnJwpM1QNu7qo05jkWBMNky12znl+S4Z9Spa6XyxDSloyf
93IbmXfOeEc2Xg4zakQVTw7YIYCN36A5SFHSGsU2gieML43L2G0jw6pFmkQIyWAr
Vcho/hvFid46B/ZBSOeSx0vvF5Daf3dJW20zpCnIE08EJbb0S8fajrDvFsn6duqe
cig05lxGVuh/irg262JIFtlApvfyCym5j7vBU5oowPhhB+uBCFJeX4Kx9ELxQNwN
YCLYzcfOeN9kI+Xxz1oBavS8MqOonG7ynvz4X9xerAsVwbeOj8rb/46Xji8ZnTbC
l/VBGNjQyKKRNLwCzrkFTu/HijgNcm8da1qvhVqsCuBrddiaYVCtY+kNN8J1TKrM
1edXBWvwdI+KIHfunXim4fF0sk8DRdNYjsxf4Noj1gKTWK4/S8Yhm72sswk0XifH
QNbWm2MTt5mJFsrdEYEZ7KYuAu6cV7tIKfHEXomZOm8ImdYPZ+JjMcun5lP4h8J/
KS6Yqw+qR5+7ufVlNDSUr100+XYY5zYvezaVGJ4rqyjNWTZ2KOgVN7J7c374pJH4
hrSA5UhS3JiyydEVQK1PZ5+7yuV3twastiGsnbQbR18Q0EtjFkoxGdmhXU4rE8F4
dNf4KTcPodXpuXW05X51C0uP1gMDcslGr5/4Rs72PjcS1VHM8DcMbt77OUfoQhaS
SIbU/Jxtu66d2uOfLYbdmQPhX/fW1ZcE7XdgnlzCJWnd9zYspwYmlOBVtfp/T7gs
SNZAc9HoNd9NVbzDiw3NcZcY/5hZ9YDXT/fHSWy8dCRl/vs4gkfqFuncS5w5RaJ3
FxrH1jvErx+3e04SZSPXTllFwA7MU63tSvObEHUG1CbLIgTRHsOIF1WLOVgsgDAE
j8H6qoLKEJDwsiYNSRhxzSvbWdEVZBSPj815KUBylmaeZMZVT8EPnhwDgws0Vl05
dWUr82li+de87/PFQmslGloj5tZN/WI4vnEMA18co8yyxSjdtmxrpFhIQKit6DRP
3EzIXWUOn622ZxF4035OhPcVMFELaGGO6yoxhS/yGhpgtpi54hzrkytYqjNnGKhS
Y15J4hje9DucUWY4SN0SdNR0WuCVH6ogSrT8cnAqYEnTLxt6xc2Xgz/55Q3olMPl
HWtnTrKX9wHjPmt+ieC8sz/KsdyBBNVAOSal424Cc0IrewUeGlEhJYaLUgwrvPem
JhC67HN2Um7AU68eVCnkQQCIcXOahgCT0TQFL5VJInEJKQ8Y80WhzpF1HZyr5SBI
j+2DArCvqCyKdms3SxYAwkUU9luEXy0ST9BPiIJsnZ6xW7+vOvGFfZMB4mSBGce8
OWZb+3fdGc4hH59Hd+rVl0ee27Unrab53W6/pRziJb9/eCXmeZGZT9VtDX6x2w4+
Luv6FKrSjKp3A1wUr4znmltGsVtgs8jz5O3wTIFJiTLJ3aHQDB0aJUoyUh7NCo4M
F8CFZ8NGQKtrRdZKyTxIqkoQVw44kDkRaql9eQ+IaXsZs1voSe/fih/pzzb+M1aI
WYLjjjxhtqRHbrYqAcbcx+bWhHuTYEpUxwbKFSEYrXYbCyy8UE5/E7znrUiWNlQM
6RvYSu+4nZ+AFNju4dm/dcTl4d8dZE0lAEaAJloq9YO+2itCjzP+UTFpjhCKzfDd
t6LjYcUDJdm+CvVr8IlM41PQMb3aF5xpgGCxTyuRhcaQA7SKHHrTeoMC0cKLmcCT
SIQh8VV1FEIAw49/M9CJBQQlb1h+vbj0q5P1QzF5mTGG4caTS4G1AiYwc4YSqX+c
8LtW/2mMMnSMcm/f8Baokq3wjIkXtuCoQ6ExxqeeXsTGOSEYUCxFhWTpAhdMSd4m
5OfxMa6ylAhPQXcycvAbU6rMvg1vJmPecfQxIbW0Yi+6eGdcxSlVVKTADeUwbGZ/
7KuhiycNtBw+IxQIVhdo4/8eBhOt82ECwVacP7SeHaLJpW0fIMEHvy85EDSiuzLE
vsXZpRNY2rDA/C/riXeW8B9WpiDP3Vc09/GEWl2QBxB+twseq9ooZ3Tb0CSbSkrA
UodAVGZkAuiDfRDEV+FAHvgFrEUv/tKj4Bl5HzHdf84gpDJt0r3TH6yZGGiYyfci
hiMw2NSGrW1qqpM55q4YJWLrvBWoHCC6AqjeEQXAnK4PbI/lbVdLsx5kEeHRDJbW
yQS3X6/GnUJ7YZE9U2tQHK1Tx+jYPGAziARzEBHrEkiBfGUaPWu4Z75p4h3KTd0g
4w+Z1ReXACsHP4sGUJgQOlZzADm6tP707Zfbv69vnlc4WiENIqt66rec72vlF4XE
75LGxCgE6kvqW7FqnbDqVWkJ2ZVsJ5CRhBADt565IJGgmc4pWvxFgXkgQWk63Nqt
aTukLRXzJdCAD4CDrdjO4lu8w9Ioh/R6lk4RKhg5aRYmJbF41cc5yFcFzXFkS54k
V+lUkqIO06sQnDcfKSwQyDXgJy9Wy9L79lF/sLxBrKV66xq63IZAyJ/WrYDh7My+
8lAvxW7O5E+kIJgCF/Ye5P2Ynmyy9vktCpkqL2ZxsdkQ9Lt5AvUX5aqpZcjGrV+z
itihT1daHOqAlOZGpuKktc6w7HjjaH9AmntwKyfHV0rQF9Q7HeY10J+Y8fFgx4yD
IeBLpyGaziNTqgYYTK5bb2Q9x4DlEAHvHNA7ToEhpmG6USvPZzkjfST1BiIflWcL
6cNkQuwhwGYp34ZgLT+8ZuZpNZ1+rz0VTbCvSSbNZbC56cEWlaO5dnX6vFXDyY5U
BNTzIs5lEHvkMvZW2AZu9up5Bl7uLL8vnlO/7C186RDZznp8NE1sqRB12FTjkuqJ
zguUDKXcoPOwz4Zl5ogtTylDjA/lofuxTQ+fyIzcYOFqUNlvfhUXYr/8RVhoEkfM
IVeIAd9cEmiAj+vYs7Iw6dV6mGIz5Uu5mEhwk8ockQtjuEfEfeZu6vSQMxqzeBpw
VxmXewtm9ZdJCxXgUpdmWovVqEuv6ONJPOdUgK7GsaJCmPJf5NOtM7na6njomAzQ
GJBItCg8ELxsVH9Hq8gILFZ56h2zs5Opdt6II+X9j6lX4bUUld2s5SM2DC1BDULz
0rENPHavBm3/DVctOL/79tebHt8b6AM3yXBuCtGypc0xCJk0emA8wM2OoepgjOCx
5YmVJOD2o+PIVd4cIyYw20Kf0GPZvvB3gl3b7lWw2DCO8aEH9rZ7vfaBnZ0Yk865
pXRU/aNI4Iw2lV08OrNVBXgVa41foTp1uf+RKUqFIYrlOBwSIGaqrot3ZeUHFoQo
NFfzWS9AQ/UkbPjsm2ibEzitrDPxZ5RwqKLF/banmi1kblKc5MjrxDr0kfrdzEU1
Lu4L3R0ibNsudS9e6ynZsLb0Et/LY1nj0Q14n24hAXQIJRTxZbOZxXP5GcL+6sDb
SdO1FraQHBsffDp40xPuRAWI+zi/zOMuBcv1dc/0zV+abLUjIsiSdl2m7KQzbR8q
CHRuN8GkVKBWJqCzTPC0h+byAHtJ26YQhiyMJCw+v/HrY+yHMNhZnwolo6kLC0nP
rElzesXBnXNV02ptWJ5rxvWUE74g5zLinR/8f34mbOf5u6RvT2nBXY4XmxCeao4v
MxCh3TxzB2CFlP9Dkph89PmeuP3z7Z/69ZsESSZM7RU0xcMvnq6VgiOypFHqKlgb
b3S407R8+w5OIqRKJIe8jk0mqC0/S4G3kgb1cNNdwHvQdbaB3klJbxTVFDaMrJuX
TZOMJrugV8ROg5m2GBsZTdGfcu4m1D3z+Mggbpv54aAb8rc8+LsH6W4VE4LKh1AH
yrbBGe1pcTi+un+70khg8bh6+A7HSg0JBSfIl9IRdcjgHsEUHe67Lm4042BXZRLh
focFlv7O5JXsPY0ydMzH+veF30bmT8qKu0K3HeTBrutqxmrLGCBoEc2RkI4DhSVB
1eaGtI7Rlv4sn1gz5U3dr3l92EfhyqKWAiJ/VWurF9N0dpj90wMo2KJhBccqFtgA
m3xdFclx0OmF8eO8w6XsoWW2xj3hrmlTU2GflOhqbpxiFXxfysw/m/iIR7AMDxg7
CPWWpBclOZUbI8EbCEG+LqwlNgEJIwexPwF3o7EHDvqKbx0obUT9YdWoDRe0rs/O
bAv4+UjGIn2eMmrCgjoaqIrwLgmNgW8YC2Bka4qnGMvZM9fhaWa50YkFrLkhQZcq
dd08/gX+JYn2aqfw3sIugPb1qrbVJJS+Pd1347Vbm8cpnsnTcoRdCZJZLVQ+BpNa
gjQfZHf3uB0gvcMkresim8VtWSCdIauifsRTHxiowAKmgWWKc3fwGPr60miDAVnl
a1THxjC+U33avJd8S9w4OM06O0v69SEKf9VnOMelbFyRTQ5tdCEGk57bGSULjLeq
S6TXHSDR32qOVkbIaVWtyA9pTQ7e0evgeWU198fe2ALKudMZ0HdeiSqjFcw9LAbi
fa+K1wSBjIFHPU9ZzgyTPaalWuGtQikbDqtlojXZxYFvjWUdFLpgROjPb59owy/Y
g5GN/mr4mS2YJcMZTtjb9Rdc6uYMI2BDeevP18DttPyVbcRcZJzJkK1zyke5WFz1
0oB5ERxnUf9ozS8s+STlyincMUrtOLmXSURf0MfAQgCKQihIkNx3JI/CGwkvSKo4
JwI1OB4nvCWZXngIJE4yTLxBpOY4uMmX/eU2u6TasRS0WgyUd9AVW2jYLGHh6tLn
lOmrWBAMbuA4sfh6yOxpy3slT1kQ6R3b99YUhY8oiC5p+bOUHNsynzCHfsm0aq1w
8p45GkhwcynqXmGAz9kCX1IAnoQJh8XilIl7J/yKsmk7JIWahXvwe39Pbj0hwW15
7uyK7F3aXcQathuoGz2tfRrFfmCRG6m91cQt1S154s/o0QQzEXbvKHugsppHO0JW
rPdM2ahtF1rrlybqTWm892lxmGUNHLHKSIN6JrK2heHShBYNa363mWpJ0IXueejA
mJQPoh9Tz1VfrmNw8NDk/oEtjQ6gA+Yj3+oSu1eBaKbNsJ1OGX0QRH16zn5a615Q
nVyx35HX+CoUqFlyRAtKpDT8wHsPOmTjqAy9TA2rP8nRD2zrWCAIcqgHENgh9qet
ry6gx74+TQ5uJAcvBn3oYZBVbJtMdm2GyFqVfcfvWc/OQxUYkYIuZQWxFHVjyQ8O
y09chi3+d9ypglwVu6MldWY98UQDTnhDsnZGZNu4mrm0X6hfeXFk7EKlzljHmqNF
8OdGsv+UZbcKobggNVwGQdYzHu1R3lNKtF38gUnTviay0376XY7mn74Q5SbJCm5g
UU+BWua6ynL4MIzp0HUHk6rvyN1OliA4HWojLnsfwVKyK4azqHJijxXn0u8UDll/
J3JeICP31RCzUXT+YI4ssvcmvMH4a78IXZ4M0JR967+LKlP1INOkPZ3jPMyJILVW
N8/qRKzH1jbF3Jg92gh58uoRXRFW4Hc9SPb7pA1zmLzzqqcANivY4udt+NiqKQmK
faFkU02tt9zk50doJU7+guKWU/B1iCwO9pwsS6nJp+hKhqRemTNQ9xBJ92uzf5MP
pc81Eq0KWHNgiJVqYNoZhRUc3dV/AyNqVlhyidggh1kObK5nAaDhZWf/B1ACE2eE
RsXcqgMeRW1eMZe6/Vm9bYGGQiJ32vpejAqxXnCjPZfJWAnIC5ycG5cITiRuGLQ/
7Fll3vRLZxIgDdOCu828mVZs9AfZxVwWlogcyA/Dq47troojqmDQAxvKj1S13M1h
q2uw5T8CeLrqaUuKa3RJ20ohEb3zHHvu6phLz8t9sx0PCX3jHAR5tshjFffutWeG
a5J79NMjeZLaMjVixtWA71zESRHSRP1gDrmV1QgQckpnBqKWowpw2M60qTMwopFq
/PfuLVHGQBndcBfnb7BHAt9Ue1UUa8eywjoL3tx9jK2A0bBabPE+/8dANGfZ5n6V
Xzk5EkWfpV7wUQHyZH9T/Xfxqci59Y6sWWTWomFtgZ2VOW1x/EYoFj8w8LSi3teZ
exLHFe0xvfc+ge7An/Dg98p7dMHuVgvuQgg1AjIrDYVyySBSdnJrdMw7x6VL4k36
Lo4NP7VlRQUtKfvG46ADO6Kg9+2Giw/JY/hWSMl9xn1AQB8QysuOCiXAjArtVoaA
bBFJQuW3+KsGFIkH6q74y6i4lezp7Ou/2eFq/50Ta8LZRrG/M3HA/QvDJIIns2ri
x3ZcfgwFs5xy1F0k/2q7AcTy1a2qiUhGn4VVCpLo/6fTzjT922jykQFlOM2i0g16
vVA1GjrnK8EaRhSsOC9DzAUpb/1/zAn8oHDDEpCwcjqLIk8hyFvB/90hK5XYn3zz
3rVK4xDEqewV1wLsZvazzESZAkFsQATyiR8KtEDP8RZKHa6Kq1MDFZqL2mxHRLAK
QlLXTRxn9hGaLdV2sev342gUBam3WNAt8STT69kGwLm6vJGXt8ENg3eNkPZwOt21
l0tnfRzcmW8cWeDkyTCEnitNHL6wtA7w1AY6XYVYSWMR6mLzmh2CQM1Q7cKR96s/
zsGB6KusNK+dVH0UvviHRp8i63IdZvg3rjiwvQPv7OD4Stgpz+QLBhspEPG7kLJ+
q2SB/lVYXoGaDWw8HcfOpdXi7/+37g7pLmCJuK24l5j0RIg9LrEvjzkHB8WoppEb
Gs2Wx0gbW7dkPxTCp3ni8cmJIxOX0t6AIskcAc9oxIRxjiaQoweljk91ipxOfCr4
zGHfIPlm2USruBjdN6OI3x/YrTrhi+TwWI37AaeJji/RNRXAVuEFAk55BBPX0MB2
D3HG7O9H1l0yRVHbb9Nc5/29y+IByNEuQuK/gHwGLQNdhWDhEvgW91chTYZ7G+h2
fNXmidmn0gN3ubNyf+UyHtx0GNOXzcRiZd5TQ3yo72kb16zaS9yQ2WRF0stouFY5
t2LfW49NJs4sABwZ4jGfQ6FUMkrX0nwxpvsKlXbpAGNSoVxNxHU2glxiMQh3zvR9
ETOYh1LLQFnpjPpbzyYAHpj1vsX3B1Ba8CZUy6wtL5ompgVfod4Pd9ZNwTMp/rgc
8KfU6Wyg9CQo4vJOBy3OGPhCfIAkwFwiaR6/I0J8qbMXOjlMUf6C5HRVZtpa36E9
vJhpA448q/s26BlhTCEsXkEk6uI+cdwQ9764uvKCtfaEulXr2V8R3whWM8YxTeMT
ZxSlFxzHA/MQSoteLQlpiDT9DUssb2QsNPvLZA99bVZUPDjzwHqkBHPHY3mbBwsI
bhzAlr2+GtYpdH8zX6FOMaoo+SVb7LHZs3q8E9ecjIXEHjJRB6ouSRlZimCLfu1s
Zp9YVRjtCfVNlm+A+tjW0SVkwZHyXAHQEqrL9Ns3oFcAInk5EkLSprLKuBMYBXXf
enWJ9KjLqwzBwf6FUazcJwGjTgt5+pD/iR3RG8mg/bj5FOHdplfMCDrUit40BsuS
iw9FMNmEXsoY83cNX1D24OUm/jqLvM8nJulVeDATaZthb/LhoeBJQXxoiWsfB55J
rqnVFUi5Y2Wcr3MeEHeAt/AkLlehKavWDnqFMoBFMRtZ+t6AX0uuByW7hndCdjDb
XYC1FOcMGwLsWokgfV3DefZBiNUoGky9uiahzWsjU0ewlsKbGQlFHvy5BVN3gUl+
yUL9wxnMpVVnD2w/KOC/UdnUi4FllkZtU0Xxqvao7mgTHm22SKvoqyUCzxVKJbAe
stlmYy5XbydbgIVwqqRmsXVSEzPeHV4jwws3P4pole+HiUnyPxtbmgkazgzLXQYl
yXBn0zVzmfcT+rO+u3Mr481AXnbnEM1wbGhWI8EFxiJDRByTuBdj18yevjq49M3j
6mHA2mi7C25JkR0PlT/peeOliglwIYttEGIjIhPfmMOFrlp+QM8eA0FI/QqN0XTl
Mk2y23exKOgBMdV2KrCXm/ogc++OmQJ1tv+U7swHONrs5+2Xlyz6MAP6nIs62+WW
7zhFZOSz55pIBVe0X+xZN+Gt8daTOKDGH047d/XqR6qLq83IBuRqGwnUYQtHRlg2
OKQdhOzCOoaQkCC8Rx/GJtWo1Y30b4Rq6hyL7iDE1PFKNpO0KM9prkb3GPmYyGyO
4qV2QnFGaKcasUs9t2SEoB82xuVAZVYoHZYCzMk9lM0OMANdeVwsbzL+LpPs9GWp
wqiA7RIaoO3ZwKNmJ1ZOebbTQ3RluoIO0AkRMw6TdA1IreN+sLrKRwaH4lAmJkuD
lBB9BJ9Psdc0s9Gtfn4sPo1aSrInYqAOfAGZxCTdbm2IlyNNpRmiVFxKXb/YzLuz
AXTltYR3bMoNgL/cE975BPb13zlZs8w4kNnSpf8WYv3Y60RdHB1FRvMtfah0fhJv
IwIgQ3cGP5YDiTdM7UkUX2DjEuDEgCS+/9p25xXrWPBK3mlkhwUHEJo3Ltg+8Wbe
fLxxWHiFufCbugypgVegLYEDcdnz5cqpMG3V8otaV5DxHkhl4MFs7A0xt/SQLNNx
5jCiS/eN+Y/AjoRIaHhUxuBllmpTtZ3ks7PuYn0mqe9M2EO49/ZD4FmFRWWwuKzW
jEdePLHkoB4yXVOfMUrNegbs0V60b72Tas1pk711B28+Dc8L05Elr1lzg80NwOYN
lr7ZtNXhyUWu+Z0uW6zu2TEx6NxABX1erApk4ZHZvZhjSBZ+ydGdo3pwzvOKydjn
+OGzlvNkWwPjFTOBU2vyf3yvPaUcz1hk80CkMt9Nan375kUoVjf3EGufEL3GCjJ4
boe/hCHFnKnhS9MBAV7NAiND56BH0XopsJH/OITw4U92az1bePTF6AhacEDDkfmQ
hngFZFny1xlr8l6KkauH5q6vWGhTytGjYHdWLs09i2OjPCzaNpDLXFuYTqskVL/m
9x0pBIaOkDuIMgEGpYN2gZiCCK5FchXfhjyax9GjlG2E2AM78uVMEmzODN4W4XZb
BObrGxPMq2emKrzmp9S1A0hT2r1956wnnJC9eVyC+XJAMwepH5pB/aFFq7W6AhH2
JT6vCxAp3crx04Ch2USougVhMIlDk+F3/+fGYY/P+wYIbMxr16fYsv22+ieJsuXY
i/9BmpVLzOsGgejXmUVr2aCW7QCAnJrgr6q35NTPuR1Zbw5a57aIbKyEdX208eI5
MS3Uyrsmh4NK/KQrTTWTSPeOgfbAnSDFXeVMHDlHG6F8XX6QTJ9BnHJxL9XFMpW8
501hNI7RIKwHQQrtln8fJZeDMMk5usrGhtJZA7n3+vhW8Nwosto01GElBOIo8iYd
9hoMu+lzy8IJ8OaBHDDnA3SF7xOAnNHNmjnjuCe20ZuQkCvrI4s6rt4WCay/WOZL
uRi9uaCwgIjJJEE5TF/AwvNc4+l254cwZ85yN2OCDXqqyEkT2qbZpa5HaAgCJcDX
xmMxRnPU98P1JRigcBtMqhzVn+8rDxelw/M3d2tvKHBgqSbu3ijpGLYwqhQky6AU
MHe8NzWwQK957INva9m09XZjc0kI1PdC4HRtOOUD7YDxGXRNZzbH3jrd7qUfFsoC
exgHde6j/hXWus3qQR0og7yc2CskfeGzUkBMsEwhOM2vawP60X3SEj0RtA9IIScE
q9NSUcTSabGv0hpbnxCkpf37zdVFCXNPPx2q0sVmwmoinOaHmX50T1hui54GVpHC
q3GDGmIjBB3p4z1fwHuMiQ1I6XghOaQiPkJRAF9O3uVGjTpDImlXCrhNFpgWqeJ8
rNE+7crlLOO/eEbxPz12mLMNBHG3IZIJoZbpSKpg72CrGF6C8kvRW0yZ4PDa/bu4
UZxoap1WKMyuhGoWB+phcFpnUng5J6OBBzA61WTF2HLGBr+v5CPcq2G2ul9ygCHQ
diwtolhEK9wCdncmmNYpLzR4tWL2+bm1+U0/L45YPqxuGEpkHBasCf5PFbnJJg3V
elf9h4yRbhB6qhCJA6oiySHX1+7eAjvVN/PbQXwTtNgq/xmL+SuIORPXZUO+kVPo
6Cbixh8b9O3SD2ySMd+q3h+xtf/bjMcHxowBzMrdFop6OpwZaB8H5nGIf7Jm25kJ
Me2m5nPfacgNnjayYPX3YDfIyr+pbw76zwWMk9l8QA6fQhS8eXQBnT1c3vzzCyO/
PYFcNvsBwsHO/rjU2ac6W2saxASIGB/qOPGIdULastolMW5F/dql6F0LfV6xh6qB
dMNcw0hszOFyRH8WW6PQAD3r9e199jQQWhqwK6q+KJstyULdH6IveKX65ROS/Bmo
9WLGBGy3A+Z/vEDFy/UIENSArkaKfwOH1dVC3e/Opu7JP1hCO6roeBqr34JGKiX8
be8O3PFv9c+jAygBPDoXL6kM7sPngx2YyYuFLuUYkBgdE39KR4XHKKX11UUW2gdJ
1Ts01EZ6W7zELEOhr691lECHAsTuYYI+E4ceBHUD734yhDYDVQkj3YiujJN2SYNw
YtgEbFLtb0Tz/+n3K33qHiGzpyk8VrYEKzqsGYz6EHAyzQ3/sZDPuzBE77NijXBU
Wb0cFNcZ7Y24pjBzcvqrLmVZKjdRzrzOxXQXAtOsfebMP1/a3Uwy8Wvd65376zHT
KneSI0wKpfnHpoRr11yLVfQddtFirFDFugBMSm6iVy83jobyioIV0hcuKGHFZ2V1
B907KdI6cod9N7G5qBbsJaMkSbp4DixTF70YrJcZwtfaiJwdIhfs4ipZ4C2D//ui
I2HY6ppWockXMu6RwqhGpU0N2szQIgnS+ITpDYB9HHkJyAz87obxKhaAdGnw+EqH
X9naeDPFAs9VkiFCx3LpszLo4jN6HLuEDr4c8HcFBYH1W6fOrcnZJjq6y4NI3bCa
hdUX7f6sFFQd39cQJUa0KIFFu6HR+G7HauAOT0UMe8D021M3CnlTT28gS8CJ7bgq
EOoHlLPTUVllnAvd6yEX17KeQoB9IXN5StxGUKhr1LWxJ++PyuHSoJ9T/0ad97V0
tUhlPxndRdmiy496hUDsem3L/EN/0LLLW92snBFyC9Y7II71qRkSNndfuqVwxrAZ
wS3K+bAE5mRSG6qRXwNSK9QuxHaCbhr099VXNsHIGjSyHpuqwp+vHLFH/kCVnF/r
wRDy1nF7ZSHHCZKUboA+MPHIpgfQWFuCFz++i4makmZpaxyK3vglvT5BlgnIttbX
QSdlME1B0RIG4NwY/zyhlvpxy2xA8pjV5lgK1lKEmPuGa2K08HUctEFRcUzdcvqG
X5c6Z5ELWUbdcotCPzD5MufPChz41Y+DjShrnPskhMZNZ2IVzuu/fawmpiFZJyJg
BD0LUy4XWU/UKa2KEtwklPMgk49lKg+kJnN1baf5/IEZ+vdMR/rJP2nYG9h+OI7R
8DEh0ZY8TWv/D/zveU9439/v+42/cZIMyXaJLj/0WRIj1iJ+CHN8rC0PsdDcj7h4
5N/i8vLbIFA3rnQx7mOPZmsgP0URD+UsQ6N+Fh4qsHAHUGzHnqbnD5YfyOYdAWr5
/zhE5zeY09SB7k8xmZuBgP22dhUOFcPVc1gtoh6UwuRkseJ9jGC75HDKnMqb86wt
t0v3qQNzI0PTT1vHfHlijBaVdWGFMicJJ+RA+kXyRKa8VpOCWEkEz5kGVshGThZb
YHNAu+6waKRd8i7hMhPt0WVsZpxXyabKxF0qRC7K0p0cVY1SikuXoYxp9T3cNdHy
CS1t3LDzEcwFB4iiXRNHn2AYr4djviknKcNgA+x0V3IHtE2MLTBCgTxwT8pXgFZb
oaJ+hXkLjP/29hK8yZybEwU4Hfaf9jZLfX37zRTuQ6OwO99rCHp7KyeFqQ63VRmI
RF3hIe5v95QjkYUJ/7TPGtFh8QCr1orQsO7XpSKDSUY7LoOEDPAjOQWEaIu6TC/4
l4iOy68cCp2iqL8RB8OqXb64xRD1yQNdzhUSK/xDimpwX/eGugnv00hYeQnt2JOr
nPrF4qs1bwGp8zKGQfIGz9bKct45ywGBYGo3xMNsiTyvh5PoP8bgvds1ihtt1PTc
75Wa3MDzCRy5OYsZepb91np8IzYyeOix8MO63uvTDUXo1mx9MXpCt9331JuIsCaY
X2LZOz2YGr5SX28DxtVadFpZxF3OnidADySHxNJMV7rNQVXBKLLis6axFhTzzhpQ
d1cKFamXo2PV6PBWbEEW2CrKg/2RY0plTKQdHZn70DL0zFOqQkx+JqAlaIwWjKGv
74Ic9qqoNeDidI6Ihz7MIb+V3ht+CiTIPs+hnqqBrIeT4t3fctJUFBhgJCc0ibLo
e/YClfXqq+qK1+oWKjnnBzRqAAPwV6OGc7eLcxXn4uraFms2WLFrPBHEm3cT0dqk
YN0MWdpPCNdomYIymuaQdT/27f359eDcN6d0TdkBdqtHu1hnZNs3HK4qrBpTJI4y
4BSuDFXdwEi9PdG84WqBXbWFx/g/uj7spNlRBEv9nJtEok2LVdbeEOi5txZvUgM6
sTnVHiiBnCTNbOrnBgVUyh4renLhQLMS/398jg9/vAF5eeERs7NY/QIVxV2ro8gH
XxZEf+6r+ulOwnJvL+tTUr3MorY96pVOq1rt1tlSIvkT/xIBl1vpTPru4QhXiOtU
aUncb4+Z+nXOsruO2GzBSUWtZNZpNnXJWymNVanXThwjWrd2oJ+C1WEaqQtHQc3f
6x8wLoKllbyljH+XFbW++EzfaQyEIsnFDOyM4MhcOVNm/Gse6ZznmDo212kNvape
MFsGTpKHOBTtw67TAmNELqDcrZpMSC/8aN4sLlkIv7i/oLDHhlZQsbzbDFieMM9b
Jq8Pnt+gSTflfeCKUqTdq4hxXZ/Q1lBShV7UJbfwuj4Fl20/1D3EChnIYxzycbSD
pfcrZiKmE0XZjYZEejnhY5EAOGXUqNNRs4PCWarYEDkBtqHXmZgR2SY+QV7BmBO0
ucGJZB1guWJEaAIW8qB5qVGx72YMhE8DIrgL/ZYIHS6spuy1+RLD5euGhvu3KHKC
Bl/VrM9kxXIyfUddb6LY9m7atRge0OIX7bazBT2UxhGk6RLalUwN/DsUbe5QvZFg
RP9EcV+BpZlAPrVXNj0+Mrar/4ZUf8aYoGtEjAC+RNCmG9T9Mr+CPrkJJ6WKbZ7y
VvTOZMAicJNWM40ZP6OEBNIakpforuidG2bnZ+jxAR225IanwXE8+OQgXYGyBVye
8KrhH194+sc3jDMJlQwkW1i23AnVO+7n4735e/WJx7Z3apJdx5m7FabnuWNEcllH
AL1ApbIwdMwWo7HTo3Gr/ZQ8UBYNa7W3MMA5HXH0QGKyKSVxO0lVxfIAAPFfixsb
D+Tl5lVFkEat6gos1gKbq4vNQU8EQO+yXi1ItuddXfzttZpeQGFYUtoUQw/1cY/D
ZpD+P++N+untuYVJoYbn8sMrhbYWq7k7bTFUy6sM3UkfDgdN1HeWTifUKGA0uLQt
m6sAtZsUciAgjWTw/jjeryW9VqKHBPyJe4RjrawWNWfxTiurbMJ1H3q4GKnI0daw
qwgzPI7cJfeV7lR6M0dTGmq+uo2T0z6hPapy/eIsiJdRNxUPaSnwAFiDKOxdbYfw
GYeyqW5CCQHvov2qizlmRjA3iTRgyw2sC3GtfUoMYgv+ZjDvdAZvWyHH1+NWu6sB
/NZp+3Ix0QHkNDHlwGF4RFAz9OVsEY1QGhp9hXMMvGbmcyLQ/fa8weexmPj2y5b1
iJUu9q6M58k1UBuQiw7EbTPy/n9TCv8YpwTWbObIRQyn2Cbp3yqqjnhl34Pk9SJ8
Im625PioQwGbbLwwTo2LK+fTgX8BPLZLs+kMCu4gzEGQ8n1WN4sUhzh5kGmDbrOD
6CM7DXxz/yAzXKF1F4+hPxnXbEJu/cu2F3WKlJz0OXfT1/avlReWAoN1X+88322F
m/otqYRH9BurA0fPY7LfyIwYBPs7KWsYkLKJYqfJvKNCFzHSFq0OgQCktRz1sOAd
lx3q5qzrJ40Y7Ysw6h6c0fRmIjwQG4cl3mNPJU7NkzTchTNt6Kaj7AKRjyue//Dc
pCGx7w2sJM8yVhDGNIVa8JnrJDvesELuEJcRDBh/t2Pwehd+HmDlHkW63SLUcKj4
QM2PjMYhqwRwnBMjqus9ML1fM0MFeXG88aQCWurLxgIARPU91iDInM5+Wjjmi3wm
AyrHOso5iBHXQMqZvlezbgfslMhHnhgmDnx9l71fplmG+BwFXRmtXqq1CdgmIYEL
ZRIGMBdtXhmydJrEgclv+sTtLzG6i8Ykf0QEp5SaK4w5SvKQG40gAHP3UfMvDIdl
/iDw/vgHGi6yvOzxcj8qvl7gafDVkQs51bbO0IqqzPwZs+4/A5KKOWBBY7U8KROs
ePJH1Yz81l2na4GU7JZ8jVGLBhMc4m0pz50SgIQ/HDTOR/sFMq/UnCxHMK1pK0Ai
JeUvTTQnAyH8HUbdD4rhdlWWnkvUk1UOpvLD+ze3qahnmz0BkZy8FEm0Yy9wLTDh
cfK+d5LRmsgGLNSrSeDAzGkIgTgWrc/tD0Xe0q22jZIMKJT+PcBV0AwFGh24fdvy
htsipuys3IgAfFJ89UIx9N83/+DI9aZ0ytaM05Ws2e4/JGHLSJvpi3ep8sT/7WUP
gF0WHDWPAcM9lz+SWCXpHApk3vtQJ8cnQmUnH7CCcNbflj5ipym3gXnmNNtiaemh
wbVX4aVNQiSE/I3MpLH/yKQ3pO8KUeA3U4AiDzX4G8T30+I3h3kEkDpT+HoOxOHL
W/Yrpow3DbVmL64qa5voEvVFdclvTUNIA5g9KmDahxcilBoulK1Jjf7N3wlZ0RKE
uo524KOWqdb5HFPDNpG0TC8CsbEAzLOoFC/doL3StvEprU+kN8OfM4p/tNLJIR8A
nS5lz8RdBNWV6Vr49ROy+kwFDpVR3So2f1git9f0sG51TjIJvmSmhqqrUY9Q6dAT
zh5Ao5k66kF86L5awoUjnoDuQH5f5/rE+eO3MbFwhtmglelURLFBDqBnR6MMS4oB
zztotqcbLWuIpgAy0LTHAWuz+qRntXzzAVxv0ph66LI7D1UVQQr8qMJamjKvs/51
gdMFOhWQKCabWKld7dBiXMb/3QalMMQjEgu2FaC6ZRV7DE66UaCe8NLf/c+lBYO4
E7jD5jq6F01f4QH902Txy/Z/WuEsqU1b1coVhzLeSwZS/52sAJX9PXrpmZHPXaQ3
d+M8Vza8CP+i61aIPEQ9gEFlt4CJYaRGIQMX2hYOmFpcPQP++MV4sZY5JseZWCm/
l8a68VF6LgiGveJ7PGfmKg3anyaO1/463md9tQfIW/OL66gNNdVp0QEV3I84n63R
ubgTzBzKF/4vor/CTYTl3b4gyIscFNE0rNwp+KHxcW2zf0XG0DPmwN8uKGKmV6JW
q2vRQZEteNeel/jU8+tCFcI2/04ELBqcpfcLyKXcTuG9xXu7R30oFMCKHWcamFr0
UrzFDG/63I11qfWP5dL2zLchdtriqLYzwYU3CaFW+J5BaCChqfm9vn5et2ix2iOG
dUr2tPd49/aBd8vedpZehTnOvf9jRaTlaU20hkOko2b+CtzELSNReYv/mdWDbJ1s
BOiBx/8rvi//dEOzwXDQQrUF60pZno+lAnx1PpOibY9WEGWysFFGSz2HKxQcCQtl
BkEQKGmgacEOIzgDDJm+asGDNVPnxSOzvon9MV6brIR2wwJ+jqxXrL4P5A5mAhHs
9JxwH1GvbgrNTP1sYtCqqAPCa80Sln0oxQihaNNTfoyfFI/1ybdWfrpDFKCSSfid
tG0PC9x5EnGYRNedFlW3XJe0xcTnuRP9Ql9i3gKZCiLxI7t5mEbyNz5Zss8/Hvn4
a4BILXHcNs3Mg/hXLGj89ydIo8QS8B/X8LewOva0C63+UAsdzIVuG+QsVzAon92o
LBnLedbl+BtYmfDDYnaMfVQ3DwtXT7gcxNDr0EOUqdSVmdin92W3UoL4l7Sxp5J9
kODXOPWLzwUNiyLnJK5+qePb8ejkTBfd7/X1pYngM+cW0tV/qlYsNw1vGHJAFyWP
hOw0AxWjeG1cO0ASE+rxTjeMdyQSEQBqeQ5n7Z/WDDX7Z5fY2JKVGsd92ssPvXCr
mISm806l0YZi1Ru4dBjw/ns4EfOh2VQmrjCiQR0hIS6S1vHLtq09St+zEmrPmOKJ
fcc4b9sZQEb6pmTZhMtUCIx9YAUepKOwSguTDdy8bEIv2cbmn7ikPhmVwbqW1vIH
C76raC/7mqUUE3VTrMowTD9d33gMKX4qBbAl0yZpBZnExffdTolsBF12o36we+M+
UHalT8lEFtKSUbDcxOoc+RO9a0N85Tybdl2uLQpYBCte8Xhrqf50vRdy+kyG6SD7
DQQfxOgVxGUd+liQD9w0j56A7p31dPfmVcubOl7Bv8pSSCb9QgPws4MFl+KlzxtI
lDpbOid6noja6wxDr0p9IEQoNqvUYxfH7XLS7u3gBmhPDbaRVPu4IzfXYrPzsguw
jglb/Ddsl3TKIErH/0d4NBlYnhKXsG7C0Usruk4P/h6u9VxlhOXh9/grVGEVvGWR
aoDO/3dm3bPKceuXUVvVqhtzjug55miMx7tp9RW/c5yT6ZoYC62lFSRMbgrNGJWg
bRyRF75q/XgG1f/Ynv3LV5tLf/uUZmG05l4WV/fOLolwiwtcQfaCBoFUoTpuqMAO
PP8uy5REvYDdRcIqBD7NBe3LZFKuPA5G0lBgC7C2tvJZbXlbX5boK5daSm0bx8eI
U5M6Uvz7eEwBjxp0oAAZc4Kck+kaX5yBXpxfzWKVyb9DLZQZ01KC4ZgxCZJP7niS
QDfOmgl17UNh14Oe9EQMCLVSe8ibtPtsz2N0l4fUmlCN4yrI9tVKtprZhcYeVBfs
UaU+PJgUzlOBm1OoSpCaCVIOeVtClQdN/+Fms1/gnSnpOxNfCs1JTUqwe6lAFjmT
1rb20IeqAW6xJ1utKeHrE/bWXXIMe8LhejD1IOOaJpMzlpnrB//+Uz5S1JM0Gka7
5WcqSvyo6Cg2kqaUZEPtcqcsaZ9Pg9oA8/7XfnQrZlgWlnqj08QhIzL7A6GQpibw
55X2F89c0StzS3SBypcZ/CiIbBGDDlBGGGG0BkW4lmnzIYtcRukgpFIhPxcbI9fd
AbuphSs23DxsqJJp54eY97L/gPNO2Yd0X8hKz4gOsd3rI9XERCS+m6XwQyVWuKHU
tGa6hgsls38DijJfhnVjEjtvm2Zg+wEz0MOOAnxLufLOtf2l7MPTxU2qqlqbH3L8
4ecXqp+jZPf2VgMD6dfeeGevWmtFbdbp69zt+yRFfnBxL8rJ5jZyH7XqKRR/QTu+
vxvoQOY1t6Q+t0BLa+GcRwIyOOjyAGoQ+4TssXd0HK2M4UH0yQCFiOnVNZjhPybs
FjX7kuZabKp2860cAch3cxj5qfCfw1edo/Dk6LsJ13ifhrfivfBokBVmIje1LakU
20q9lQ2O83lupPnXC04+p15Hei7KslwEY+FGYKKu+SABu7t+oHcIBtv1Sa1bsRYA
ukgQzr+3ixjnzcv+ml4cFmcdTRz9WsOL6YRPeZz5s2wvcSzd/R/Cn75xnL+/YFTy
DModKeENZ6KmebhhcO6LjDSsZ0/8SvKTEnndBE58+MHKNA39TnziEsLYUTv0ohxy
ZcqLmHPm/CDMdQcrGi7jiwcHqxLr7GytGp4zZOIg3a3xP7MqRzg3RBQG13Px39Q7
H9B9v8YM8mdcY+Gw31DWyrkMxVerWN8Pou1qwezbGDtL1Oc4U6RFxXHGI6r45igp
4QfeTW+I4nWxaHZcPCX2E2wJ8+LgukNHbioYF2v3Pq3juulf1LhzCbjm8qehZVV0
k1+N4wwYFMh37N2vGafa3ZdhKf1eC4oEEwDeluKRh6RDTlFxuXHBFAguS/P9Rwp9
MJgv0U0miM4WCCarrFb94+b9RrdNCEk5CE1yn7qFJMy5r61KeByRpTY+4cbSODae
K9QyBXBJLHQVK7kJaK/d2RG+cyeCSYQEf8uPw27RpyRqHoaNv5Ca+7S9GsV8fxNK
tUKyIxEu5mHq5346oPSwiVf2IcPmj5qlH21GKW4XlK36ds4lxm79K2B/UVlu4nI/
ASiwufopeaivmiPPChpWNVPxtXYzMBYqlKTD0GSiqzkaNmM36G4d6Ojv9Ai65wb7
LtNJOUGBV7uMP0WPnEr5BfSwMPvxB0hEJ7PAGDHf5wSpllIX4i+rqKpyUkBh5LCA
k0sG4wTV2yCIrLjDsLWiPFulB+jCJ/2iDA0r8WT2JZPROprOzIDEqtx0R3y81Yd4
sKk3V7qANY9mdnH+VWAU1eywF4eeCjD95ogvADQzSCOXX7KRspO9IBrrB0gqJK2j
WbXuibRRCy/pVSWw4xoiyE79g5mNNwbwcVVWroYbrfXHWogxLzRjYc/eJSgqKqVV
f8t/4/wSOCC4goRt/B53biZNDoRNX0OUdfVgNi9ErVje5a3W2e3ki4C2hV1P3+GK
HPsZIn80Qj30PXiLufGE7Jk0RE2JPP5BazHtrobiSOfPdZrOL0sltp9WpF6gf8ms
MWLIx7T5jKE67g3BiOv+SUpyMlsiXBwimPYMybY5Zxu/qY2myYgsNKFrehiFvrJE
6HtO/pozHbOQdIaIgBvqXObdzpGIVwFLJjzP8gW23fX1f3p7KB9pId1gkoyS4BnN
5aUQAj2Fdd9fwVdMPwyeDW1vshVCZGlx2vtyLPma/tHkF0BXqxXAI8BsOdKA+i+K
1zgO5bnVfo7kRDRNXmhX0HcSKaaFq0FfNXKxzhpUqt22w8kdZkUWNss8FQDaThFa
wHPn/DmuCPjBnpWloIFgw0nn5oy5uT/HAsz8Z3+AObLXRuCSYqZdiHkAmT6QpqeM
x2s69AN1J6i5GW7HMhdk4lj4K/ZqkCRR8uybcOpy7rl7gui7DpyB+0z9gFG0rQ6o
aQfYnUYj1+4q98/pA+08rc1QBtwh0ruroa8PDvDCawriHQnvq+OSfRo5LJSTCCq7
wQWQ3N8X6gknlyTTeqvSYJSC5/WZfKXWqCikNEeX2eNrmB4dru5Xl9wIi8UJez+2
b4sNiObTnfRYmj1yqcGYThr3ns0tAzFDO/s7cItVQtEv/UVcuylxjRG74C8LLOt/
KnPdVrbEvsVnnoMY16XmHLPXdURK05INCIGk3d9FZDQKLxeHYhotG8/zIdR1LcNH
ss5hdf378j1Yxj3uFmMoIs/lXEOI2NES+yWsWsMous6bFNfdF89iWqaDpiglNGKh
UgY8f2g81i9BSPsjsFNnk+MCHpQXZlhBqSU/Idc87yEBXkkLF29XNvzvC9mtwIzx
KeL24+F/arirlOnAF3p7od8Xa3y9uw0x5jqjJPqKzJsaPsJgipN7Lii3BRAaVEYk
z7hAcJnAXDdpjgqVkcNA3Mzd9hP3Vuqn4Fva+jUIAxLL4k+j47/CN7yXtZMJ6pzy
z+ni/ExkMqSvJ3ErQguqn0c6VhyrCZLPuBP14H7s+QLm/4JTE93BdomaK/CUczAX
hbTS72NG2D32U9hA41nlwyEbmHR6K0yT/cO4/qrVaCoRX+jQ2npyddc3Qtyio7MI
17smB6HNDHukCoys+yOt+75a2dbajK4/w9cvvF/6mnbLepIHbcyz/TtghJwIS6YC
lXfQnBcpSqVlS69893bk5+iBav04/EOzNstxpgej53z+dsHYj+vjD/W5CdYQS9JV
d4bwVR2sY3IYl9P4ludKbn6xPN1ufGd4/bDRZzsdLkIO9r6Q3IOUMZ+MCka4btGi
TcPtOh03j1eq83Q2PjBv13pS+X3k2KElVd0XWr4OWivu3a5MZ7Xi+AZAtxtQwILw
l3BsjSQ2z3Y96tx0qdJN5DAi9z4jKpaTItYuhWiWwc9Y/CTNsjEoV98StK7x/+eo
cNIhYhREgSOGgg7Mq1tOCG8ylEWU6Q4IApeQZ07QSKOGDs/N6efHWQ3VBlrapYwH
JU8EjnddtyWCC52548yWkZ+WKy1tjg6oN++CgmXDlnzEG4lB/Ld/bOZlEmUuapaC
ofzDuT7jki5S2GLf9MtJfDwNRimxVff0X/M4I+KOn+pUT3o5vz6YP97yKclKToSj
QkS6zGGAwqV9GYQf+jBCsNkNYx95h3QOB/7DoZo89gm/TEE4EJqfQA2wjcMDpH31
yspkoiWp2hUD+i+PxMV7rVcfp/9mnv4wYlrJerhrXN6NQbZVYwfyNlOXKaBeIx3D
/0ozGrbe40+8u7QJTiRLItoxMOqfGKledRdbH31Fcr06xnTdmqeHLpmd2xwpuFpC
iYVMkh6Uh0tTqpUw/5lePD5NjcUv5qbncSn5w0xsT3H5s7An2jjteercJ8XQ04dK
9H3mF4fzu7O9c90SC38iOkN4TdvPX5DQJ/+9ofLVGwthwv3efU5CQNRCnFLfz33a
z0CdbcD4fR2A39rC+blrvF1fuPu1ZzSxyiyUFOZojf/w6LGR/W5j+PQqe1sgV0hT
bMJAObzB4R5soz9HUACZpqE5z8/JdHijmUwtl1/7S66Ba5OD9X+TEcnrOMdqGNfd
RVnTOXOA1SBY0eAvDxnYKcWHwvJnvBXHT9+I2MGXYsa0eO/DLkc6nCsFzU7iPyN1
R6mYYXlV06deHXVRGtBl+KlNdBKE2N0+ItgtEpNgWxnyYy86ih6xA5qkvpKPau2A
xnn0oV4Rv8A3ZGZO1aT6XDJ3fVtYueyoPer+HhopxYROmhH2SrxLs74pgNlXLNFV
QfdwzAzdVvIcaorxFiqsqgZrpqmmaw8P9038YP1xm7+5U0W6ZEk2YmbgEH1RBHSI
786DxzETqJxoAYWGTAoVT31ozNwPbCNCiTJlRXJVwyfb3zn2jMOShouDD16cXL2I
0Q5q1jD6NuIyYlW9hDzYf66IpgIfHXP28TU6GiMpFr1bAAq8LcVbo5zRyYElIDQE
tnmXtrnu1QIAFChpe1bVGcGG/8CUIygcqivl0kjY4URgHULCeTfOF3qtlLQt2nTN
oxv2jAcvy1HfT1fCb4vkpf9EZaYbBEwM/1pzRB7G93O+7zs1npCk4yGM0CtVBJr7
bB1vzwVLw6JnoQEUqY6deNkGhUaLw1ZUZi1hNRcAzp31ordDHtHDORvJLiDWYBXo
VHAW25kN8nmtUfzn1RqpLwmuJa/BsrcZEZ8JLS+VRdRqEIq2eGmUKLTg0WGz7WlB
GnBBL9ri3Znsxq8QcRNh+vez/VgRKD++mw9ea3auLcp8g5MzqHGoL+bVA+oWrHno
o6G5/6cCz/iUHzz29WHZEzOrxPgXCYnTOD6AEafHgm1JQRTAUZCe89FhdWqX/ZjK
ePlc/hdszL436HaN//Z9R6ZMi1X4uHYQyGpBOU4cCR2QSGkNhv22pzQVw7rURxgG
LgBqN83HUcnH4YTfsNdm3J33p0UjgUIvuR/ZZ0ibNJgaUFdsVIxpKGAtIbctazd/
d4RaSPYmGibKLI8MHaQiOkb0oCNI55KC/WBlxNS50rPurFLsmGwO8f9NvidBN3kp
YDSpHBS0zSYWgP65xsUgi6ri2MdVnTnFxc2bcynpyhLjiPoAO/leM60l9VUfCBbU
825gnaz228n30tABCvppaSLXEVSX3h6JX7yV+tPZNGpbzp9D2oUZtmY+jRZzaXon
hpkJ4xmgmtZllKV1gA9qwVzvulMdRMKdP0Ihp0l+nakF9pbm9MqLRXHSDGKoNdf8
Wj8yrUqfTZEAxxLi4TDSmo/lqRr8+92gBjUINuPfNe8tqE0d/WaNDQ1fmG37yqH6
kguqZtkeTCRvaqpeTHl22XdKWLgx0+5/KgBnYdhhX/4A5IiIdJ5eX2JeTHyc+9ws
ib8oR0j2WhRho4PAeu1IZxlaAjh7ih8eZWWdyBOPfDLskpZqJ6fu0nTgrISOK00R
fllGxyZ2pxRm42AZolTrkY4wG5umjkd5nGJIdaHzohQoodlXC2nFLNHWftahFlH9
516glZU/0Z7RdIgcMdelX6q/+MgKeGuVf7HrZppMxr6kkJF50zQy8h4N7sZxw4oL
qqixpS3F6q9EJPnHSnHQhtVIbs5LKs5LQ/ts93t/L8/gbDc+AEsbzsrp/dLQ6yHh
V1uTiyuS1QORB3mJreIpjRaOVm0rXh4/+7J3i4z9bgGp1a2AbQDlFVMpcz+X0sL8
WejMQJEq0YW9VaTDvEBiULW8yHPm4HHv5soYcWxb5ePQX6bSzBSx5H8sjMb7fRNp
7119X/NmsVhh5nHXkbYjkUgzlJfGFTEJJNFXl7fQBxHhgMPeyKwjDI3nyIclxdnM
rsIx53z2nPf2gnrbos/AHS6USAIqzq7qHZAullQ39SCZkbogXLMQoA2HMFcskQPf
NH7QKB7/e3rtucogZhre5oYJknyHgerqccYraNYlZ8nu2v5NGCZKsl42PGZ8ulpt
Wp/qMfE6yo01vhk6MbXgOtACBiYQGi/APNpEtwhdRo5s/7M9aGyzNv8chUFmHF4m
FfTNZFjFZ9ctHup/emoFlrBjKe6h8gsX1s0ALPBP6DwHNxeoOIW311GkXUrrpIkU
gUFqU8EqONqgO3KDhMqaVLG4wWrEY6cYeY0DwR2RYbeqWDRERYemjf96M3Ryt0/Q
ez14sq7LjjSjvtOrHkLJtrK0NvJzV0DKJzoPgsB6MFp3vEbmxPDw742GoID7DLD2
SOdLI5uAqy8uWkFpE1+gBBtMA5M92+WMOMoPUbQCTqinaGSNANQDm8/roAH8tgnl
pnQEAmqUhUm1rA8coe8XrLrb+foqnp+uVpU6fgvF2HqxmN5GcWLrvBggWDldo+IX
zWu8kLEgoC82WFMyoarmsYuuHrPVi2pr+UhFqgmIwAkjnaSSwgskpryCOyMT8AM4
vdKPVHkXy/NlhbmZivJyItCQPUx1TpUdwSURmXroqqJ+mxxfkBpuuzXCO6lpU0SU
QUQFg0AwWX86vlfekYq/ii0sQgEyoSuaI983wVZDbzdpCSqe/ZRGDK6LKXjHmzVe
LJBddTAOa/3xAtc2vWOmDZNBhH/eRnDoJftYm+Z/WFQiwegUtveQPvKMDRovmlLY
gfzEyX+HUp9qWGXWjRFPhQPyRI7G5ahPsUZgrzw7/6U5Fll+Gu3QtiyRiaQU4JyR
1ReORWVXOZKTUlKQ0Zcpj0BwC8AharZuBEN3e8NHjHGKsgCcgTRO34JfmD8jj6DW
As25SzX92vJO8nqeWXtCDHps0vpeliDyEE/FfZxcc2qH9uOFuKurKo2S/w2kz1y5
gzphq4ZFYvX3fB6ghhzg5/b4MNHjzwBa6GGV1b1p1VQ9aF9CSzwDVT7K2kutwFAq
cMiU8HdeYkbN3SGuM/jxT8wPQ9SMdB9LpXRrLqxOVmMIyemTV7s0uFOixGRIMbXF
WGZjvMHD6kwwCauCoBiRSYvwc3t20bANSNok/B5pvEvByF8ODWelYJIocvZvCqbI
AIscpuWnfVGtXd8WbR5suHkYSXcizl3m7igSK4LaBBa6XHN3d7eX7BTzN5NmVNCq
KnUjmsZX9ywnhBqM3/uqthNuyvcr4v+xVgyXrHl3oeHw9a2UBaatIbTuiAsEIKHn
z8TDHeZOjTWq/flL3SGOk4E8VP5wmMDPW3Qf/FqxmaXP4RRKGLQWOYbcGjD7eJ/x
LluVzNtUFPWmdTzOhWkjy6JgvdnunfXmW5WoRxWvphhvaVS3eP12hVayrvxg4RLd
vN3nHc7QS8MvRIveTBDUsyeJe4o2TZCmCejxB+EWQySrtCOH0DNSn8+sr+VNDHXS
gwrsqghFVkv+/TSEbWJFkBdPIhIUErFYeQRiek1oU3Hd1LfvZfb+uOdlPsfwDNml
8j3hRQGvFlG9tcRXUOz6CCeXCIaXojPrjCGsPQ0KMkaxc3QhezLKbj3gqbucHEgx
FINWlG5PM/kPxjqni3+5+7P0MD/xA7EUaNFpPchBw1X40G1TCfopg10TAeHc6yII
GCpkRatyM6B4C0VjMc0bK+8E/iu48BHobwSwV5gemlvkNgJiSZ/WhG0hCvTlDDPB
FxlhDafLcgl6Nisq+6+AkFPWq/m9ukCsuWxyNyz5L9a4NV1sy60t6knnlnNB5DWO
dqRuYh5uU09lLolndixoGJuzzBsWrfw4HkZX66nW9ivDF3mkyVnL9zsiUy9dBneI
1oDU4rrnYd7WIVnU0Ae7fG8Uh0XVGbcKn9v4HAz+uaTnZO3GdbXUScYsi9SJQ/ML
bdTRtNvu9GYmmy8K/cIyTRWRAvOGbIpPoSVkbrsNj3wv8KOQbe693VxYnr6XsAql
D2SoNRZOoVqx0y4BSFNHhW/7/ZM00z2Uxy5jxmCjjRcWcbPicoOWl2JdHK8+xjvF
buWfr3cnY1TiijQxc8iYk7hgWScf6QXx8XVE8r4SmRufKCxBIZW1+k39ooZJ1dCQ
8WRa4+uSrlwMI/wOq9aib0vlCF8ZUFS8lQgObXhE0Fqz5lMzCS9WXwmEC8d+7o+t
B/xYvTTSPAb2uY7jeapcsxwBaY56ultMIhNQaO+n4gXZwUm4iiYt/dtQd/CUFoqV
9wiYRzsqk0z6bTK6mjaRSNAiVCGXz6v+o7yi1V3bUlu2n6mEMNBwUVQtwOrjD3qT
icym6NXCXCU14YTh3SXrUdX8kwHUKm+bSHd9FU7iUHLMpiTIOYN/eMlWg7dGrzf0
FeSHzFxNfGkXoOK6Q9W3DzV8AcO88O26Mrrq3uHCGTlaD3NY7ryGLVDpl7K00ZLM
mcQPL/XJsIXNN/ymeJwT3VsReF4Ylk/TefcY3a/Nkxtwi7q5Sgp7nn+/EA9yHtph
Wac1izAMwSeL138q8aIm4mTNJRoZgZIiz/DiOZ4aN8f1zGbZ7J/nK8HqX+IjIM/4
nPdbd74vfYSayaxNjQK67wZUk+wfyUVNcj2sl9g6I8RhIphdrCErL20rODvWZVud
TSCqHs5uChVJwpUarCgoEUZfuwBp6YijydE29sAXzd0e72+ALkc1yei6u5bcSy2i
efIMo9R05R4xbsm7Hdj+UnTmB7rQpWdiNojV4YO/g58U4orskI5mH7zWs6bFRoO7
xwhDL75TAc5o05kK2/z79sb/ZITD5RP7KJWfijAJP7St/kd2w7eTolzUwm/bG4hF
Z4FmVNMIccVReoWg0RAmk5CuFoDSIQzl0EBxxbvxz6TGyk39P9zWTB5Kc0IBaGzB
7X5FCEDyZLiC0+Ence8+VduMsmbnrJoAv2qbbk79Jx+lRLNMZCp0TsHmX39JF5BA
PzKnam1Pt/Q8hBaTyqrWhLcmGXYeLzWx08ywDzAslcITt2pan2mFU6uWMdVIQwUQ
m7SmEh8lFvTfjYase59pZagui5UR+2QAj4VFICCuGuGv+yDF/YJ/IYHbYX0tPNkB
45NHkQyXqG/N1tZN2dWtBLki2STMarGdtEAPMJvB3Tjot2IlxAEQlNg0CtNcXqjE
DfJALj/BR7/nPkYfUdwjWjnPyoCzQ3nTTq8H6iJ2anM9xLm6TuJdmfQgmUYqQy+1
EtOpRFtlZmCSyYJWqEi8gaLc3363sANR5aCfzZeX8+w2Ta2sNGLaMbSC8WXxmVt8
ed7ZZGIjvK7NJ4ssRkJI907IOLJB0lMRLPSeUZTbrGcvfx9Ue46x1s+SuEBxTWQW
R96UWgCkg1Lujuxql9MNiZ2rHdpUNGKBKxf9uETGeSpmEydBtlL3dEoZKR/xTchZ
JmKA3r4uUiiP57KEYtY7hJauUXOlwXV4WgNrOl01E+Y8Rfj9yRQAP1dFNIuY5rAt
9AkN8Vh0gG8hR4/Gnstj4YgnxlKoY3MX3TlZVf5Yf4AtVmyd/GZ8TAj1X5ERIDfA
RIdOpCRw9oC32keJVGN/HhQZF/J5kv63ACz7mtxtISyQ8j7eveHhfzQQLUgiCS2K
jPDsI7ACoiQejAuOeLurUwrIekgKd7fyU7TEtbsqBWhehYotK7FDsj5q8XONx3LI
Ge/3tRQC22CagXEWmltUPA4/HWWS4uQHSkVgLvtdsGCVgTqF15aBJZdvsB1qXLAY
SOqRGb1LbR9QFwIyMsbMED/SDhur1VQzTfHg4AUyA2/KUTQimvwjH072tB/7unAW
g2Ec9BrF+SQqEhLmTWPep5I5vp1Hy/69pwS/GcncBn7pk0iXOZARo29fAI6jxd15
pMj7OXib/99wBcoQw9qH6dOqCGpdMNcK6AzzPChcoq4hKd9zTuGfGnxtM+fLQbQd
oT81/Z46spXcXLeF+U7bhtPYMr4kE2yS2rUOC5MmBvtKJUjQ2okTsIhed49beooS
VU4hyaaZ+IJ5/j0ZhLLa15NgtVGwM7tcup6OYU5WyIby4xVPKjbrq839jbAQGTvP
AW/l/7XpeYo0VD4PEE3vTw7C0TYjvTvLqLqU7Z8ykKAehaoq21q51vqO18LQ3tDS
JfvcmmYs+Y/3vyaNq/ZuAUFKa9lc38kCaonRsxGGarFq5iz2e3U34Tlgt0NUSS+A
RjvGSutS8p3hVKrcz3xunHaAlnewGz+epYVqTrkwT+N9JnjGl92SODtp00UANo3J
DTNS3tUVZ9VcMq8MzTtaVJ3bhZLSCj417A4Xg2uPIWNgaE61Cq2GNHHfEfjdnGxf
7i+lFa1ts9fN4+PWnH/Wtk76aLtPud8AcrNT+Pe7sb6vwi9MM/dRyWk3mivlvAxj
ufbm+kw5wcJxSj1BbGxrHJBG1zLMdG2as0XjLGgzqGaRlDci6al2p+3mB6OcelQl
thcY5OEvQcf0BfZEIhZArNtBHHw6Q8Vhj7ryl/C6ujVldRHJUkGuKw9hkzpEmeRN
0xAVX+vkguSW0qjEbf0nUv9N6ky2+s/JMOwTGBk0PbOJgaxKDEYALqzhNauFfgEt
+UYo+P3rpKlxW3Qq2NVejgN/OskG/+ECL/yB+sKQKQZ5hHOvxZakOKlOlz8B5yIj
iumrs2gKAkFXltGqJxYlFQSTefo1Zpm4Vxf8KrensmufKFDvqcBArXqbkXsgliXl
6CJpi2qCKJjCTxfU715B8fkKJtzPZAvs4FXauYemakx5r5H53jlU0JhlVhWLHlWM
1t2q8VDquSqYcSq6tNYxwyFBwJ390D7C57/F6NrJHiIMPChaEjh9TmF9DacagDxB
PukASVZQBAFFhhZL/j4obYTCAwmHHMzEfw6NozTlV/6T9ehui20NwZPgJQbtfCrM
Yhlffuk1zoHQjB3j1KUZvH3y9ZYNHh75l7ClAWDaXWuMHzZNr97185bf+8mPIgGf
7jiVDb/ZXhsKxhDTebpIUUDArvEcXFL2ir8/uyLbVrGLLQRziHkE4KBrsfUAh/Jt
K49m6y2McahCnnOw4Fcubjn+0A8XzaElJe8XWBFc/NmwbJmAwAh66A6Y8phorV10
4SznYK+Ciqwow6lGZoDXoIw5KJOd9kVIfBUVMvH0OQhn589e2q8O7cD7rlb5jCdO
oa7j7C5uUrnP+oBV7Btg0YoivYSmRBHvj13tTmInw/xydV7X3nHX1WKa/W9AI8yh
ZYc6SnJkwKH2+TVbly1sAMyUV0+wWnWO94UA6RC86v2JFBNSygiUaJFllHzPEU00
me7WlCmCc2ZkaPkgEJVCpOu/hFyCNBI9xg9PbVlYeYbdaqRcZYL114NWlSnnUXCn
qN+lUr5eUJTufd0NNfwqgFw3g4wNF1lT9IAOgPMV87hZevpnLREp0Qvq80U6WGVD
rU2yQ1yFG15hN+hFLP8a/K7DZkyBPF3ma/GMkUYgfsRzytuGUOBwiIkNgyNU2NPj
6B+0psY8bcnPLWz18I5QaRcyt++Utlq9xrTN+SbYlNH/bHIO+BHgxQgYZN7ARlC7
r/ycxmzMW6EQMSKpzdjsldIPYQgnfnIN7FYpbIw244VU/OzciD+9iKTFH2VyYqQ1
hs6IwV9KPrJzKR6aQlAWgiiCUcftRETwGqrP0ldQYV1/F+O/bU22eFyvkh8yMKMc
LQ1prkia9s2wMueeouAj8zn6ogtHHQWPcpc6G9LqLHmyVHcpgV8yoCkLB/f3O9DF
uTyAeFpDqytOX+Q6EIJrECUoFdrq7g/HZ1NpXOF+3bLqAVNosA8mJCamF8lgO5ye
VXcU/HhfKeDbNV2FSnsh6AkCw6NnbzhBYgs12wXGifnylwtOm+Itm09SjycLURRg
jf2Rm/nnclPxPLdnC5pyY0mwPeueiOSnzSCH4L1FbwCLPfO6igR5uCsFze5YXftY
3gr9mtlJTd7xdSiYC4FHB48YpdJ7lDyX9RHBQ7IgvnNSExjlJQAlqNJ1lNvz56Yt
KiLSRHWhV9b2kjgDQ4G+Nsg7tqB5+ACT/Xuezp6m8/hOWKtBrWOk0ZKct3I2YPN7
y27DfBuY+BWDBabzDleiwu+NuIL6L6U42hVZO4W4jKQspkBn6zeEKlHv3BrTnSBu
leRaDos4IiWFvtdhs79vWoyEAgLMkDj2P+bttrS1SzHG4E0vXmqitD/bAPWtOCKK
aDHrnL35RgnnX2aNc51RCsKspFobsuHwCzDi3U7dZpGXScCXreJQKEEaoByclwIX
1SDS41srp+5wO3wezT7T9bpFhN+HJCkxDMszUQYw7YrP57zJt/FfUlTpOsCUcz3J
+69a/H/aaAAuczxsA0XSL0sYDiE2wVOSsMzPujNs8v6QEq8CUH6QQmCqmlVKxT58
pT3VQu5t7+ByTunt97GmTdbPegcwNWDuWTRbATuoaCMf20xRU66kFGNydpRYH+ky
vB8eAW9y+XUTfHNFRuSjLWWb5YyWPMd7kBsHee3xFIB6ZkjJuFbX5joqBOSbEbNV
e5tCAauqWvJRHWTu2jHGB+7x2cxcDCvKF46JyVMjRMaqW9Fd3J/mwb227Ninvimz
vO1ZPQWPkyijzC6NWOgBI5ay152mD9OnCF8QGD6B6pRVOrryMBuHIm+TPKm+4R6/
4q29SfqK1AgfBMJ8wTg/WWXxIIhqy1nZpdu7G1J3m46/oXIf4B2Nrmbsvqw5kXOF
jBHpWLCb86KOz7W/VvuZJ4QNDeRtMR5MD5Iv+ZkKR4EtGOVKqO5T9bMW54OsyiMr
QdHSbgJKxJF+8Piqf1tqmjAWxQ4LBJuA7FpAicxeEyj6W9fpWMnkvuVe6K2BoYp7
PvHhD4EA1QpF2+b/ruvhSFrJ69PEpyN4DyyZyHo6PeUPEf+yUz/yP3j/tIrxLuA4
VNwV292Q/XG5TxN8lQHTDmBm185QXzVMovkdGNa/Ir7JJiZnIzkP0NdxjU12jEbD
+wE+k3VGNXlDe3jM+95Mlpfx4eZfAn2Sp1ePKPWDw/zvGQBGgVo5OIInlM2UySbj
cgUYCPW+XNzmLSGVTTt/zRIDDsgd8V7D9GkDlVePuioPbKLvdk78FUwaexeCvrPy
pP9dFGHR5RumeUGwSty+/qrSKzZnHl7gf5ldBdGACrSyuhodPIi24cAuMA+uZBTK
rXSCdrwRVT7fnuTIlhCANdAfaKkeHluP3Rqo9aKI7tq/+ZzOWg4XB2bH1PMFSYEt
nv2tVEaqFphLNxywuMLvqSouK0iY36Q9kGz2qTa0RvcUebGu0y+M15j4FjOX9HGb
Lov1UwIfAlNO2Qq8xIkw4xPm/O+u4ngZw6hlQTQNCXHKLczHSwpSPenMGa8EqcdP
DJuoplVgeB/t1INLZTZYoIpoGyfEk1dW+CY5Fv/w1ZDO33lwVMcNi/dz3rnBs6sR
v7k4uJUR4I93EN3Hwhm5jHRnQwih5H9F2yVL+uMBizUqO4RQmjug40nhha/NqIGg
d0y2ir02mE4+GHvv8dVG1CeE/qDKcJRqs1pZWIOlV1Ef2jm51uEZ8Os4gE2EcsCQ
cc80JJpIZ7gJdA2pU6sr1cAQVKyRGAtmc2IjOyGuSjlLRHVmsPOTMuH5CLBb9tuy
0mmdP+ObBe4gOcJ6a3xWnzxegLP/PYbITgDadTrODA5Qurl1kDuon60erms5SUWt
+pqRtenEPCGI21OwhdmTneSA3wpPxUPrIwxuuZydzKZgMI5R8LtsL0726Owfaiwi
ybenNAhqqjBqzl918v8XKPaLDVPgcVD2e6SEUBvZAiNr14gf4aGw+iwmDJnPDI6B
u2gIdSQbiQNr9fmraG3E4DAl90uWD91mMjCgtGHpr247260Xjga7wlfIC9eCFZ15
xRDv+6igNmAw8ue2p4oq5CcfMk91AkkuaUuZ6NlwXNoE0uvetuCi00Xl1aWCTSL2
karJ05Qcr/rE3H/P6jqs/jFepdBpxl2LeDSDGG5l4739lyT0j6s8rcVThmTiqvSZ
crRC+Q7iUirPwiovX31b8UEDDSfOxikjal1oDKrEq7SIwtrQPQGdUAMmZ20W1Sis
lRQfEYaR6MclQjn4Va1DNpnuKT03g4Wjr964/kYH3RSUDgA1Srgl/6StHNTssnqx
uJhBde2KsJ1gYhPHltrzsfE2fP/+/qQ8YOuJG0neeAcaYS9IlfOxmzMC76yWfN0g
FUTK8Oq/P4KzqpqFrF2G9kpBEHl+WiOmctDTEZEpk/JOryEs1J9F8Z2FkSK420gB
1t9m9h2sfAqD2CpDqrkYv4AJVTme/72G8eMcOrWxi9lIb0hKcq9Oz2SyuWSNZKdk
Ye1HatUnB7RWGFR0Ul2mt7A+zYbpFGorf0QZ5RGvFS1xbm+LdndR+FNc619iFynB
Xfv4KCEsq15cUzqQ7GBZ6DFhLLJ53KsmG6mCZ0Ag6FGD38Yc+4+6LcF9nLKfRmrC
NmVwLTaIxltns8mUHe1d66JoZiVXxLU0IajT/g8SsijaMR35RKY42Su1bGm6EEGn
9VHF7zcPqUG7W+xoSHVjEavoppgTUIpIFZ5HVZ7qeElTbRqv8vVbx5jGN3xC7iGz
3yjro12iCtuCOO/r5wRn8/oI+s6So+TjQH7MKA5EuyBxz3RIakOJesw2NmNfjW0V
pSJL8WhBK79FSspaDzWZJV4v0NvmZKTyUlhYa/BbQUMOv090+2i6D8QyyVN1arra
d/srpZh3K61cS96J7DTF9JN8NLuFS6VeNaiQdDZgF9cJX46KdhydLK8/p/yeWFO0
8fm/ABmat1CCpkEx+g/pIHKY+WHIT7GepSl6usCgsFncoANJgyQIJHRtdQtYM77c
Fu/zqjW8oe5rsLn+61ZYHClmKobwz6eQ2G7RnYTbQK8BjRMaQLHZ2bm/ApQcVBMM
mue1HNLVT+vfoFBR4sRMGsqdZ1d8wm88AxUPLRDoGl1bqmmLKv2sHT87k1SnZ6sx
GAseE7wql5wh4L8r/8XBmigEpkTmauB/YNqtaX7qAVg2II8OnsIDr46LbUsy4Cld
MwygFcDFgSdiVHuj4fgO6AHcx4Rmnv+knB+8slJMQj5W2hrWaqOr9bEGwVqmAT2/
K5G/K0F9d+htLeJz6yaWY7GqLPtHTU83254G5S3e/y1IsAkDmmRnwycoqOGryeSG
kwMDhQTfyHYwDRMaLpf8iVDICibuvzOPPLijra0KAhCAykU5lthqFLQRGiJGpG11
hRILHgk8k8yO+M8zpulJxI6IHsoogk/2JEzKWhvKbEMQPj/FDSIj3L68dtle0HbE
GJY88xa8RDocNFzs0tjwUsq3MiESY+RI0clK92j2FYm6nv+SR7b1TLK36labp/v9
6YYoxXnbnHDJ7jt0YU4+QQ5fNTAsv0yg/Vm3a+zvorHao8XdeY/gMW9Z+8IpmyKx
VM/x5vVV+ZqeEBDIi5G/15d3aV/Pm1NaODnz25TarzWJrSq8AgDAh2S1zSmHqKEQ
TsUy9COlgqWN2g5OV4AJoYv2JVCKlUisADh0qCw5HtNyMUeG7UeBz4qPpSvBueUJ
M/iN9GxzVwwIAnzrkrk4tLk1MkhZKV1sKzs+Rq7D64eG9Xh+fmAgsEnn8qVVQ0+N
m87RD+8ptftc1wkY9xkholERJ2umNowoWTKt4k+Gz/m5AikS4u4G/UBkvMP24Ho+
yrOKWRlchAPVzTmlNckbWKB8XdwoMfxjPc1WxZyPTeLseklemhcmunCM88EVTeN5
MJnh5uZbVZ/u66bkW1ECyyyBncCXU3AJ1Q67X4lqiBQ0PC1V9aOKm8KLIsML5tYp
B0V9CW3XTykNYptywOqQebgc+4K2kwMhLRWBFwg7QjH28i/zeiUZYv00tPbVSCR1
kLht6WobAs7lcDDbHvQIWlcydnNFb2guNLY9MbHzWzO7nxVNHfL5givCoQKpQvND
q7IrKU3qav7rmzb3s3dyXESG4aimdLyfurkIU0OPbcHeS1x4nNhkfZKHCUlN7Bfo
xpxjGRlV2D11d4u0AbAmrD9Bc3HYIpRS0Qby+C7TNVRekQokUrMY/VAmFCaK4lvA
UhIxhCvfH5uIpobJK0IbnF04eN/e5MhOy3JxzX0yvmGhlgEfmZ0Z+yEmx2NLcjlg
196vM6y3X/3tI9j4R8UN+ytgUQppRVaVL/7gJMz6SCEXTYigTpJJfU+ohTQ2B960
QeOj4VGLpt/eYjR0QF6tDzBeMzm+YT9Clo7dpHufRVzE4vvnWxuK3klQBdjiABBt
CS+ebJjnz24Jgh2VPQXN1sZJ8+KC5XYHT8syChr7xLF0U3dt+6hyJVws+aA1bBcU
rp2AegXjIkV79+4bSJ17wJ23Bz6X+N2nR/Ueeux9ciSIVYWvDtegYiljgyCD09Zw
b+yqc6B9FJUFJmcVFr/iZwtxbFPtIziTqCWlag6wisN2r2tLRv+gauG916wecJG5
6LHscc8G0EhWuJO3U5RBNTeXWvKVtRN7Q6TsXCKbMe7EpFJmIPrAuLwVeiIbOA4H
XDFp/OhwiNkq8RyadIMVoFYEY30exgyOPp2DqJ7HRjqNpiiur7bjPCj4GAMGR+WI
dhsJIlTlB26c8AVHgAZrL6xBdXY4Ab3er1Vy349VJQUbMmO8G4Zcklki02OwBglL
++U5tnajP0TxwO8xKBfepJylxUIwX5vGVZWOyac+rafrC1xX/uI2iZD0xWFOGLKk
g1/PR5/2Q388JrltSAi4eiJdY/OwD9BWfera8/alyoDRaHLO9WHSZnxUFuj7eCSP
78M1k5WZSKzxcFQUcM3nELD4Q4kOniHlZJTfGLLAsVI+txJl73Mcl/LrHUS1Gtgx
9CVZ41uXV00anfnMmPHQsPjAfO5bTDhtvhPs34oSFRBj3Ja3DhIGa1/tFlBKNTDM
N2KxgAt+u2AiAEiMGFR4xNjZrcPWXFNZa/Ck5leHlBfJTzaQZR9jdv0p7S2W9m8D
EwKqenDABtRua9hbDxiFWZ7edAB3OfTOuGSAvW1UVlDkT12l0zYfWTvYR8N4LSzp
wbPrQeRvsn+oCHQRFUF6h+s6Rq/FUvA0/DC1KDaesw+RI/2j1MSKSPNbIFz7ZPXf
EsH1ZpsK0g+Hyl2MGq0KIyjU5cgX1mT8fmjTQl2vyDyAhbHy63LffQezvkRaDOTs
aHUfxmbaz75PsDBFzPY5EGplDZgWkRysID0RBRQxrplcY3NfGzv9j2YNY/zZS191
VsDXX8YKw1jAUzMLGefBbqCZBfDeqQuFJtEfFHNWxMgIRNfSBEy/lATUPK6FQ8KN
6zqdUGWY0W52rdOVZf6Gisf1rkkyDl2FmcrBAL+Q0wH0GTNSXkH6wb7kJJO3Ei3n
IHwNjaGQfpSpwD39cVdIaj3b1dMw916SNV2mB9Eb2M2etCeeFLOEkbsi/0vMNptt
GTo/bBmxXzL38ti8zUZFF0WbmXVO9B4cK0kw/Mo0IPPLleyrD/8DFu5wV2uUFSND
yssCSUPax3aYbjZt5lrsphlaP2EUmhpNdg+w7VeYN6Sd1ZRFxawWvZ7aJJS8p2jb
mQMRyh8hHyjdouQPhK1H2RsGJv9i3qweCpwQDps41PkC1Ur3c7gd7GTNp1X0IZvI
23qv6jA71WJpX9Oya4uBy0vjUN+WPTIB6O+sRe5sDLnnq0i90n1bHcn9ICh2+ZQI
r9KU9SsKHkmw8+cSA0SB5sF6MYkWUcmPaW4yKXmVBL7sRkxyuQFIUiwE1ST4n7ok
sPqz2Fe/ONO+dccj8CZxDnYHw2et4726kf4Rtfrpq+4odLMCMifJRU6Nlgpp3Jzv
A9IjdZ6WT+biaS9ybZ1GlK3JFQoYUAsvLLyjeABjHhbQ6Iph6jnIUOcPhLz7Y9/U
C9B/w/R6NBKP9TWWjy/q9Hgum0A522Xll32bhyc/VFkVuaz5rCoPAmvpBvhJobQ6
E5mM42EZSPoT7D1TxxP7bDNRRtHBmhEzqUSLxc8pqQCUFln7UxHxx7NPQWbVC0sC
UPQsTWE704zYwx+9H1lWnTK3LFDTYfy1ubpDoef7FimKUVWRStnKR12tuJUKTwC4
UEt3U0WDusGzzrnZHXn6L0SX2edzADmNjcUv0tnOpY5bQZTz3p333QI4jTq3GZ7d
H/amtK2us5P9GwJC3tf2qARSOP2a1xlDcuAyzvCnTWErMb2LwyBQTIx5k4IMkwMl
Vyp9dU4vg1JHkOhL0ZoZ8N4sUPw/aPGmB90Kq/8mEwDSGPHFCX1uhzv0zJIw4wtq
vISII3yfI77dAdkvr+RJP1uvMLKb1zzICLv58tjbiInz8cqS29jdI+qFsYp8wPP5
1VwidZMx4pog/aP9H0ikcbPgHHi6+UNXsps2s54RnXJ+4Gpdi3UaLFlN3RlSjbC2
NNa69cjeX+WRF24Pbu0vHCxVhYEw33EUBPXFE4E2dVnez00RxrG49gKL4UnKrXd7
08h+UjnYGK5tEh9shmeMg8OlqfeWM0kIN6T4Q3MP/cESDTGskZqhcsM1MM+WRBRK
3345yA5w3b+UTlbYV9CR2l2YgaSjb9CcrARaW/8nEXSmer4F0fnQ3C7mnXkW1nqU
lw3U+mGkX4/Jc8LQZqKK3VVW1LSLOxOfyJIS4LeE8cjR2gz7oDbi5hEaY7p6o01K
NcXiizn0IR315LS7+sh5X9Y7dX1woSwHbYq7PCXlr1E9EuMf2iedzaczVE5KAjvR
0oookdy8X1L7u4TC+twwOq4ZiS85HoolXAIvbBQUnxAVUyX5YgFrm3ROpyUor+7m
6uv4BsWZ6isZt7HB/bFr8JSVO5en89vyNduYYbLYF3V6Dq/9e7fjYfUIMijoYkjW
l0DZZmt5E+ux3WRFSnlM1jb00HmctACUGH4Avcy5+ILdLUv+A5rUvoR8apMA+Hde
8Gy/JJvJHNGStFcD151rt089jmTOHbL40QQYJCl9VFuP83ZqbRveGEoBcZYpcqgb
qxtNKF07op2DdhLxtdVDWen8qK9/w2NisiJIvq6YlArO84Dx7k4JB2kDhhJh4AoG
ZyLZpqj+c0HINJeYlXbZmgsxlPNpPwCAbiBTX1DJKPwi4tI1rU7okZQAEOVC5Th4
T0vhXubZ5KYhj975YjDq7GwFlYlLAV43l6bt7yDQ+HRKmcRymlm6qFR68DemMLdT
lbe5pmAmz0XQo4j6U8brmU4NO6YWhZwREDJth1+XiJUGUQ7aOyGDQyMOeCt+vaI4
i3IVFoiM/nZnErFUevN7Qwyw+jPJm85WKUxuoeTpTt5IclHG9ap2eR4aojw0aEaK
eF/CmmYNOgEkLdXXTz7kZt3RotUCy5YyiMn3mFCC10U/PFNUJmfn6VdHTHQ/wQ33
1D1PfDzu+ZiSpuZvNAKBwqFRiZ9OK8rRCZZgAIyfOKPbAtKjAeMLyJi9O2iq/nw5
ml9QLcPnNeq+AX0n9t7nkQt/y/cPZCL+Cmfpt9STaLPwQ3uFvNPa4DFcydSD3L3G
uABjSYkB0l9z3Z7DOVF1fuWHLFWMp7Ph2WIqY5Q7zmy+UGHZHz52prtIH84hXV1k
o+7JVtHPZjczuwOmvpDaDYByKD7bUsiNTcHrdYCT78T9cqZ5wMwzQIIfZ7hcnJdf
xOJe01z/b0289tE+VOGBUeq6x9VsEvat6Ck/TmSFo+CFAqqTgiYdpbOhHQQXeKY5
HQVtCqJ5FP/7orBR9xl+Ke8ktC411IuwZE/RgPCFkrPCcITVvyhNWdMJfZXIH45z
kfia89KOzRxinBBGbcIF3W0txeNgVU2Eks7VpsflHRzHEWq9qZ36LruFpbweQ9LS
zlzwAUW07rdxuYCFrQakvP5Fjob40PnGzEIIMdEBPMzkA+mFvsAZaTGcSKlDdSed
lGf4duaVLjYTMbR0L1mg7+L5wIWkcsBk/IRJlclDoKndIKfhkOIBHp2uerhTYaTl
Slml3sYubko8abyBvcyA0ZWyNyU8SO7gQujfZ5bgHQ9UkTpeKjY3r4yibCgzZS/Q
bqiMZjWJqDRz+mwJPX4YIYckJ9zu1pToFQxk9F6BAST0AhDDlkSl642grlk0FKoZ
oNS/VtKwvKKcZ1VAsBHHIm8pKb1Ru0f9VKOY8y6bRuShplL6NI3ZQpDwDYnwd/Jt
l27Ads28Hu0BfjJKnBLlDKYUxu4rfQEvtAeTHTb6Noac69QIUGbosgQhTX9Y1urf
m9z1fx847zWzQ/3xztH9hO3YZq4bchw+fX7DvaBY6DexbvdnFvrg0zXft6SoIsjZ
jK6jp7SoltgBfzgWJvT4FyP1ZRb7LEuPi4IUweVPxvP9z9oma43sOgaEDT06vHXu
hK88SdBzV2Yz1xGMocW3o3Ro2xb5A4SELyXmv3R08P1vfQ9kT1/lMZ8FHi1uCxYq
BpQVCVmAOJKZxy2Sj5VQjCrWckeNUumvz/MWLvAns93NslSKDHIK3Z6MenGrS1p2
y5gG2fEtUUSEAF/PPYDdn77Y8ynBI4eKgjqWhpOdBeoKdseY3mn9PvKaMbxtvCfC
TA4LI4orOu4AOZM1aGZ11sRDWVy5nC0uhyUpDMRhQQ82/fTfZ9SVv5jxuDt5O6xJ
4LBQMofPQVE8zb7N1+vjmKaKy11Y202l10Vi6iXmpsZCxkTKAHzPso8upPbw6XQ4
ZZ0ZVdoae0OjL6PqP0v79m9JOQ98vRNGIFLp6FLPofxzluTdNMgJ861LMH/zb2AG
ElRmo2lzn9cz0kex5mvRxLMUzCM3ecO8q6c44PxdXdhHO/VSLahMyvSSI+kBwkuo
1E8H3pbCDZOzrhocgHSNeXvOs45Dk5HW6zcRUMrVbyDaI00sGrzD/veVDlD3TmA0
50mJ6UXi/pxsv6MylL6YcLecBbzaYAZC2/8B9s/Qv0UIOJJzCxogOOLmIMhNhUlP
mqefXHurcFZiDR98uu7U2Uv8H7RSRnYv+RrJgtc2kT7CmZkrzYrgxXS72zCEoiFQ
vvScT9E8hnvne12mofAvP+biuWCXVl5QMg8pmfvEReprelJb5BeEhH/A3T8HmOuN
KU/2N2hSy+BHx+sbFGEsUIXq59wWmKrQeV+yDu3Io8W0MYMlshicKBCGdRBBqeX+
m2v0ZqVw1G3K9qZvDBKCyrOtHDbe/pb9flBO5Ph72RrZ7BwpAlkTCqPUCp7grRR3
2/8+83s7/00l4PCLSV8vhYQM7XG6oBTo73HBzp0+aU2gjt/2CAxCUbe7B4rW1WJy
o5Sb3qR4TLUa1fm080NwDEgL3L2PqtOIaPctxFhskOzMUUNiYvLV0CQ74RkponE0
RN4GsvS9ZgegWcyDO7tZEbNGldxvOC/viEReJ66HCp45XxvEYww9DBxHKH2q7Dsa
EexW6zuvHFfhLq1IXL73gxwbnbiBBKSF/T8taFBqbpIQNj4FflNEtiZtvpEy3fnM
NyZ2SS8AjIGFSgHehkRVktqmt7vgPsNUJ48kcktckl1qt9V4WXMQyRx8XN68fFfs
iTbsCDlz0C2nqDIlmtWyLsi5nOqhxN0cAWmJVyLab/RZvrH3HAzkhOMXtDgZ6tcX
0e3wAC7/Y1IFWp3EIiNwXUE53hV9RaucwVtcCq4euwfb8Acdy9fhbavNFuZ5/ZnJ
zvUktTYYTh6R+KjaPb8qilYFBX8yku5Cq0tOYRf0EQ2pw/k/GQFBNNuOXyTss/L6
lk7pYUdU6DXIjkZ2R9CdfbxxMp3nGOwy70uYXgb3nYUr6vdwHoNZAbt2M2oKIzVO
7cxogIVuRH89l+aAoP5vMRFWIvYMRP2thUaeDpYEpPoaZrKD/m6Jj+MLXfqmX5IP
PsJdfZTeKe7ZrNmHAxyzbQSSLVYVMLQ93qTDk8Q2CZKgpUE6Mv9HPXzWFo/y37Vo
ZXuBWPfE/sitnv5qAq9FCcyRSbvWWiNvhUdMJEaau/9W4QxotXpVDzdFKyCKRDPM
yyADtqs4/PBjX/oGYkuWIeemaLrv+s7ghD0BnxZM4jbP8CkvFFXaFH8Ok5JhQGDk
IGODO7shQlcf4dDTSqdr+6tbDUZO40UkvShGjaBw1fCmA9Vte7AGNT+soae9PzPv
CdxLg+oYohnDf6ZMo2fmRhOMa9AV4y8YweAKlJGK9gunJ+zUhVCH+idA5AYQMj/v
W30D9yXYtEHIHPzWYnRQ3R2sK7jkFExJi9phifpv9n3NJqhbYOt3FxRsLStk8AlX
pze5el2xf0pIM+CO/DoxIaX7kG/AVvYFCqYcFquCVhVVBl721cvtNrcniZhXbFNd
h/dUrd0gZtxAZeGZJe3hR6ofDwQToQjbY8r9+TyWBjDkJXeDO/B3/gA/JgnP8/EH
f6nQxIVe+jz11R3750zcIpHPpTMeadmrc9gSHQwPfD7bvyVUn7MmmyuU6Jlf77Zw
CKuqV8BTtp4s04CPovJ1HeDVPHEEMgU5HV6djx7zwYgZv+BdNJSOOkEgVoVL/8u7
1p9y4x21Lt/zSbf8GpejfguP9aA4CW9ib691aRg+ACCTIRyt2U5S2X22VtzTJXOr
OGx7A9AE64hf+FdrNgUbQKY4Wjuy3kJQTum8am+acH3e0w0DsUIVnwK6djotGmui
l+W71F1U1//dZumQS7soNtvp8/L3xcavKDEQR+gQDhfqgMEfb4aFgARJQgcD0xXy
oRkWCOxKLOcbwBegQyYNavRh8weLHX6VTvehBR878dJqpFNwpOuZKWLZcsGkHO6f
dDff7lKSpu9/qeGL3QkYHXQQZrOWrtP6M5UvDjFVCKjh+gtkffCb3id8MPzcXv1E
3jpoO68qLJytjn+2QqTARHavd3Hm9CSijyqlP3N4P69r82kHHVO1Pyn9ySvFQVLH
2xGI+kgvLjzmgyvoFQiVbOFdCcH8pqRcMPAppI2EZsLbQ3AS7BN5qS5ivmBQSGPc
jbGj+rEsbYnlWFATAfiFwiQviZrASHJXnx62ISYY11GdeNZ/8xZ1KQwhdLt1Kpw1
OwyoER/PmgskSQxUW+MI82OZcGBqvsqriAjzAt2oKZ2CPdmSPLgUzAKVOWdnw5hb
Juz/CCzAXXEWLbF0NZlKOG8Epy7PmpM08G+xRZWCCz9JRsX8Gpny771GM4dVOILh
y9AVJWnacHvG2vK0X6IIkq5I47Xcmyvq/WOM2T6ox9bwU2biW4M10UXcB0jZVFXT
JtOxh/o/Luh1lUYC5Ow0hnIitdeRQk67MoHtoTiUJ86Jp7pfewPIAByxxdullThc
+8Wo+fiIA+Iwv8iyze4GCoRrO2Xejumi4ZirRCPmNucysSqPBXZSq5/3og5eKRk7
2hEPgY/Mk4wkylpnfAcuXmS1q0C5pGyx2s37GUpaX9jf1ao5bGovPlbWsavzG5of
qa9MtewbvwQTXLSH/M/SSpCvZIvh58EOzLLFUY6e8OHeQNgpHQh3ydCSoJGJNi9d
aSyeN26ZGnq6XveM7i7O6sgoxZr7I7q47N5gVr9bsMVhJ6Au+VBjEv5OYUATBTBz
Ie9F9BnDdSl7C1WToqcE0KaOw2biEhzTRT8/5yzJ5G+aUfnn2oai4MXOZy5RiNFU
L49UimexgNkZAczmaGRX4oMmhYGTinXZHIcJQkIMZ/WcNwOcP1kLHGitwxOWhlQx
nyVTpQVuiy75isKTfOPo8c+KBhcBXifttT+nWemUIpJgBbg48FZYeyb3B0O6XTrz
V5qd2Flw5loVdHz78EN+KZxSmWaLN1im+Y1kFS8Z4wivS2vwhTEHmknITloJuzIw
8/Xw121yGmejZLptMUJW1E9GaG6J9WZvqSaaHq0aqE9dz7L36KK0RltpMJ9bvapv
Fsh+/Rk1UJY9PyAy8PgTbmGx1IespD1TFkEuQMftFEIFHkgG5el3J8bBxf6G5CP9
n24qdx6mngDuDOax3Snc6SYDatyGKK83KFjTZlFxphDe8g8ZffdZV8VbAQ+snJ9Q
ycxEf7ZHsG805GMWBvEI3n7efRzocTMGMNXqkBtxsGvh6+Y9F4Vx/2ixo/XPtfa9
Y6hIu8ImRAW5biMjeQK2HpgX5wbZDswpVGabe+F7P4dXsUN/4g6cgSjNapCgtNVG
HaGcNWL1djILzW408ivl/eoxTtT4+NdAX72OacNbRvwgD3pdhGQoyyGivBZPtTsN
v9uwGTXkm7olppKsOXJMc5AqCroQl+9XliWqfYWAqDq6feVczWdWHbZsB+SD2SRL
Pyf4Mn/MbIRV+h0FMhaumRfV1n74FB1IfMoLpsr+RAPv0H/Rh4P/cX/OVVcFcSNL
UCktTBcTl16uxLt7C26GCQbspQzs0Yv98WTytWli8IVlveLK2bJos+NoLGD6SLkm
uRYQAHe4TcoapatOLfc6TyK9N2s+FFB0SSEkvkHeAhzNoygdU5bEkYsDEQtip5zx
poWQPbZkB4+TwGC/8mDhLIpesLeDo6yOBlZg4psq04PUU2xzQhSkdaWsguQYUZHe
1SSY/KDSr8EClQ3MuOulQ4tCcjdsI4t5gtQvYAb8+60JLlvtpX5N4K0yUcQH1Vrg
OtuBxyuVFp86UwpxWtqv3hN/JHTZAbV5vYUUdjqDpTICZvsDAiqOo1tD29GK+CEk
4Mh4Kb3qJgwS6uv3TyzSd6zeJW/3uILcgKoI5DdcmYLhv/ZC1BLu/gl4l5Zb8ZJ6
XI5OrtzFykTyUuHX7AEEnRxkyvxhWE1oM4TAzDwVOJoaR2FJTexFNYnHTeOi2RB4
YFWkBd1O8kfdhWIn0S00V5QdfJ0C0/sVHa4qSVtmJfYCpJmeBtjTGAITmu0YPsM8
jBN7pXIG/YB9oGFtAaQHqj3j+lm0F7FSFN0GaY3keHGHW97oyjMFI6cv2BbN5Thd
AL76qE5cZLZcZ+LMOrd5xvkAgoWI9fQjJf1X7UF2Truk8nLYb4r3uNTcmK5gbDqW
OF28Sq1pYxEY9JkTQRhyO1J4WF4yy5NCdbGNHigA0yIjP8hyaUsbRhZh3rDcJdyh
BRKNwC9kcRhV5TBXzo/Ktqf49ftm0Kae0vDBTfoldz79LDv22/Sr0TzvEWBq95xz
8z4HeVBcbvWa4bmob5WSUQY7XftdTMO/z04QTncMOmVqrspTYcD8xyOOM74zAZA8
oCpd/BECErWzGBwr5pEA8PZS3ZcavFqLLmnpqPPaJ9jGmzLf7hoLOaxygXP7Rgps
rgelkY7LsGrh9I7iQ14W8J/GrQr93mLNsVufpMf7B8DKPuSUJl3II2E4p4+g4NmM
S79/UlzUyST1ws+pBXeYCEuymEwrpnFZrBLSOEvQI1Ajmc+T2Foqunqlo14zy6AG
sBv+NJ7rdw/p02kbUgpU4xfiuyZrmZUYJj6Dr02VzvQ+aE/JdYLAQMNGgDQExd/w
kJBHnV6+Oson6Vq7l6qJIShzBUC0a2qMEogZI2iqXhARtTSbZmfcAb64pNfYEwaE
G9yf3SsXd4Thq8xAeNiaLTY/K9w+SL9wRmNf/pZ5qUVNLtTq4wkY8Sg0Ihem/fK6
CuZkDyj6+4EBufUtfZDJt+NrIeSUnW6bf18Olh2YBPzlwdRoGGKUqBjgFsqj/Zj8
QPlXrK4CdWJq+7SDO4z+cQmFhG2cqHCrhcsU0QYHDAc0dCaF/V0tnPt/deEcJRLC
nJxYQon6wUbnnNosGD2Jl7l8hCdCEKl0HuBN7RRHWK2tE2PQv8F/Nt9Ub4ZvCSjj
G0/vKR5TI577iYA8uflLvQyNHCxe1irFKAa0z/DU2yUuWllm9DrVyjNvfA0BRK+2
wunoaB8vGaGYsvMT3OYjlby39jcHR9KHahMQ2GzfKs0mGnfdzEZy5vvMwNJQa9i0
c3fAHJ8Zu2VFeHwoGc8MhZbdcx2JubjdKH8lu8MKh5+jbM+Q3xYoWsma/1XKmPi5
6/xoJfia7V8g7MZtQmNQfE/Q2qlJ0+taTW73JCpM7nkctX9gYYHpF/Vi/Hf8Z+SM
hgm/C8FkIQPqFFh+eOgCA8O1SHQCqv0aJ7JduxujRSCxEZkYhTMmvKccOUbPebkG
u5G6AWUm6UtgUdPteem+eOluvUZHZ7odGKMREBWHiTbw7LGWWSH/EOEqLdhDQwt+
TPgmuiuPVix66Wy8v5uMD7io/ZmACYLF98hs7T17869tYC6ECIAb4SNugR7kmenI
1HpbKWyAia8p4Cu5Woes153FtWYlNftyoxMndgPpbwuU/3+ojDlM+ao7mDVCMRla
bTHc3Vkd75nUFfwLEMmgcqRcva7qccYYvey/Cvk4JCYbIHYPdov3RqWUBcxRYTNG
tswjej3Qw0jHySQwlsCU60LLEMCOy2hSWWoJpEb7s4hitjTEQlJo3CgWzStRh9hm
GrYAREEx++i9MCXLXFl4F4R849OhKZkYYxza6+uajzRLEF1YPANySKemj61WmtBJ
9pz3s4ooovaN/hZ6mMrkye/rXu2MrnuYDbPskv0fgMXwzAX9onElRKHrS3Avzif0
MMUT7jq8oaFQSORyy5l3oHaOQMhbUdOVwvLqr2uEjvy58Nh7whDOBkn0/Iz5Y+vz
KhMTWezNepwotiMVjiucEpi27T13TD7qTK8OsRkj6ySs9yo8AnZZf8X0TPp5bOox
fwhviTkLTLBtLdoOKTUwD51Kyt9Dlr5WHHRnRCudlSvaCMYhsK3nUi2ANm4mpZNx
JUB1l4MP/fpjhdKInnSABxVJbV1U8yKBo95pCpk+6OZtVsaK67O0W8V5DghMBtEV
2HYjVLnuW8T+srfYalA/B/4oanH/Yi74otmAsVgtqnjjJUMMSCm2znpq6ZCYwnq8
swSSbx0zL1Iwm3Ny5Kn9obanTObDymyDppYHvsTVCpoh5ds0bEkGDw84U5g7VJiD
UGz78EwDO7rem7oYoMZ00Re3D0PTWbUVn8DJ+hW3KcQerQkSFTfJdy6NEGGeOTnd
nMtOyri+ev6oz+DIaa1pSyxpfng7kKpO0W0zIfYoJrTnjZYyhUr5V3PAa+nMZb+0
MeskXFwwHMTiA8av4AkmHnzj+wDg75AwPXWep9WxEs0gHIpxvJ/z7EK7Ds0KwCxP
XEBBQN3E+eNdUYGZnlx+D79w1NKU5Pg4+DGqznjKjGE0jsb+dh/7uIAuwgB33e31
mim0Uo6MhQdFG2Q8Ps7i3RmaE7G194ctp6mUymZGryM5pKnYMn9kEs8lihJMhPAy
McvF9IXCmdxVyXV9ooF4q4e7Ehe01eHv0f2e0Oqm6wvGJsiHcqBq3sy2Nss2hwOV
F+e8VPXoF8lkUznsyzTq8Slaj8A1QdmtEnLxltxvTgCO7v06fMJoFpHQIeugi0KV
7VXiFzCfJT2x/dvTQKAzhAppH4vPDy43ELvuyKllN4HU2FpJcvFEmAANSpd7XtZh
frmijxaUshyHHMx9v96st2Xdgd7F4C4mEn/u4ZVUzEHsVlvNv588D0Cz1xfOpDrh
EPgJRBfN28cMDJgrZP30a2W1OmLnJ/Jm3I9qu8mPoR8ohdvLXlMT34/1nI7uBEXc
NP7BhRRCA2rqKG823EEVDFtIIeiNsvN5p2jA354qPi39DD2A5USsbI0s2XNNBj3o
FfVFm/+pfFHwWvttPeKRX7BQJmOsODUsFPbBYml+l1kkeWQfrnJppL3c044VSrbp
chCeKDENcAGQ7qqAwAgY2d5N25GbYS9X3f5RdlsnmATU016MIkv55ldDMOYFELzI
692S7GmxK2ACIYZfs0GdSfcWis8RIGa4+Az41KbXu2FktlN0ozpCyXk+kK7P2Ea6
Hu/mkJnQNzzV9KZgCfPlFl1Y1ESU61qagE8iKBlJcWFj7r79wcLuQZhMvmVLi159
rZ1RpBKdPC4RtKg4aaWT42eiBAOkgrzvUTu3jRx4ysn6iMsm/PTDS0Y9WHubVm7S
KNWNW3WJdpMc2A10YXTT/lCFttigN0qLPnya3GrFbD2TGXy/w07qov1WBWRJlBfa
vXC1rkEFuDGLmCqk/1YVFdS0srl71n0Pa1bIGoSRIpqPKYVq96eK5Gx/uhdWvYdE
GyrReaUO9bIlAOGdquofdQiQshTSLrI9gUKRTBTe+ZkA18rcIxlYb8jOkQPp6F7N
Iy+fxF9NNhlAD4QmO4l9zL3zMzIs4B0XuOar4YKI7vkVY25tsBrHu9serkGqQYKH
ZhzJWkscz/QcIJpojOJ2go5/qPD41vtf+nDAVgxcrxedFmJavERk5nyXT95Hqyln
AZJl2viLisWqrg4cLzi3yLJGqh2mh9d/VkZFToJrnz/RNL69dFH4n4v1a3+McTw8
PzCzm/0KhQ+JsyGvdmF5mD/Le0pMY3dnX3XGJg+dN0AVUDQ4hz33tic07p3l2U2E
434RF2Ih8lVNg6fMv9ixfMNdc5QGMft++ISdSU2GGtukWGtEHGVJlP3Sg6ZqX9Lt
IvEzaJSpZmsBbGRyFMW6cqagNgSLXE+7hbdgDTApOThxFnsJVFO4q01xDmBfiShc
buPGQVFUcpaLBHo7rFXnjTcMxSAk5XQM4mZnzi14YMbH5HUrE5Ol35JDbG/odCEE
6g1hGvrYojAlnozAAH0HFdeptchzZyAl0YKCn+jNhKgjZVHSotxfIm0HA5g0v9uF
`pragma protect end_protected
