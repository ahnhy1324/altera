// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HI9p/EWJOBERy4Cx0cKDxCD5giL5ACU0TEO3VE4ggHPjCDqxpuwfqpyHKzSlngvx
D24KVMy01HkDEN7vr7wVrlWFUTuRGWOD+qE4JdmLW+RMRpK8Q+y5JZM9lXi5045P
S5TcMo/UUHZrMzLgFLF5yLsNs6VEl8tpVZPLcGRPPDY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7200)
hA2SckUUXf4xfY4AHZXGgyFUaK+jYOr1oOZ9bNTLEGxZ6xDuOoHSlFpaAIystj5r
posTX8KNDRdMMAjWEUPPrwqvJikdkvktTKp4nJE9FV3g7DdIiYN4R/lcuV3txYXk
+6962jEmFR2HQE00/emoOWlVKWMYX8UkDg8obLRqchE5Q3ZKGWcWqAk7m7eKCPez
OcyFaJGAVZ+fAAIC9GSyu6lBOeGVCvS6CyaR9KxRXvMYEzGs6EvEhvlaLheQWi0X
8V0vaZ7ISCEWwivUxm74tIpQqhRYRyn2k8GtThtiSDoussBfmjJytwHedp1I7hvV
CORoQSO9tmU0F0hJSIz2/WlfOWxtIujNu0Vu01rKcF5wANEz1OlLUW6d3+PadEnT
oLfkriLEWsAd6caFe+eDlShNJlDu+OU1cJ5/k8xxfp/pbvBxhip5tB6BmzI9l4F9
f0coccWX0TusYYbylDdpmuP2q5J3TeKRdQ6D7OLp09Lo22nKUgCZKrRl+IyThgi6
NcZDOHc0YURlJ7JSjqR3GR9bIlLhm8qYETq/yL2a2RX/sSkQi36Ek952W4tlBsQA
xC2iIcCrKWqdnHzDXHWBPyGWRoHnZW8xTC+hrlpCyTBsTwEX77fdWMXfbVKpjV3+
AjO8EptcPg77eFHGr72j6HJiGni/ECSR//dr1gyESfBJ6wybX382HJyrZdKJJkZf
WKElvKyx0xSi7zpv66dKG2v68CZXWlu2ihKBOGV3myu5IghlkqNTMgU6J3NpCfqW
kQH2DAr2DZnhePtSqWoSxPQn1iELeArOYz1/anl+ftvcCy29pQ1Ar72cYy6hDTC1
qV3nPGnQIi/QAUD+RuyxmpcGHVJtFnKR/oD+kXIXi0Zyhwd4GQR/8UnqRUfOCbZY
+YXuWs56x27uXxS5Ymrbg6gqmJ5+Mh6BfEWzYeLOGdUmDKhkmMglzlbAuTHekj6B
n7KhJdzaaRzeL54X/hmgNPlXsEbEklHlwLAVGJTwLKD041+niChTjLl0BC1AHdTI
DTdcpb00v5p3/l28EAKuMthOSU5wwfVsBG+1EuxhXV1aJlS1ws0MW8cWk0qa3T41
2WwMLkERETXDIzBDusBebGDj5puAQB/6WtIOXXA7psrgB/ObpUDMO6DFQXnIFj9S
/ndwqiqIQY4gvssMA4uGeJXIKOzXjD5+3ocKFtg0ZghqxDJs3JkEitR06jFfJRVl
B+BVw+ND83qU9DEwg/sXFl+W5sWxvq3M+QiWUSJ9+aNSvKcWQQB9sIedt2n+YOYY
X5y0quPtXQVglxVnkBWavjj3WHUjXY0S7nh90sH1zTyzXNZp/f2HbaLdAE4Ho9H0
jjaLmvwEjDjOSJEI3F+cd2uQfVGXh+TYC8DwLcWyNEY/uEhcGPNbOPLlW6yR3nK6
UeUnQ+wIRZgKrUhJUwk6QTvAzN9N0BH4E73HJJouefqmYORrWay4pjYYPB/DuTIS
CH8L54t2dh2DHjAu+c0CJ5440/YXjbBvkyNEe35YjJ6ynb6m8w/STHT2tSCnSXj7
dlbgKKP3QOPjTeYv7puJnkNgMGr30EC+rnRCm7sXkznA9obT/K81AfCUv2BaniGT
jjUSUbDhQE9ENgm1r5xbZld9abJ5SmRHrBCcXglRATcQWla+FjaAc+zyXs4qnFdM
MEAQVx7xCzXi/TaQF0OPpIRa4uQV+Zq8/gLzb+heMPO+rGfwIPsmcvgQhUbypZjZ
gahFYKpsHjheKi6Xc7Csiv4JxNpgdyb63uPVG/s+JDrJ/zGWermMU0wMDX36ymy/
magfX4+1zvbH4RT7Q6ydPCnl+cBBzIuiOVH0qUTplPlhZN5yN64gqw6zLlAO421s
7ozTMIqDcQpwmk5hGxOnaQYV19KgUi4ZUnu5bpyOIFq++WbVpOyVh4FqqUWOMImu
ePGLJL565HiiqqD52uaSAz808jkViEJVl2GMUpEvx5Z8d7jy3B5MjBn6o5jfH+fg
Q4zHtx5DTsn1gzUrgyqsocd+iASGNKa6QznOWFFPT/3PADY60uMW79h9YaJ2uV0q
wzjYc3u7wXOPWB6u9k6zabhd6WfiSpucrAMSdebli+gbFhBJOpSpIUQWJWc7bi/L
CofR4HT7T1UABpc1XaRCiMuCh1F/FKleU9Ba/+7o9wjzy2YK1+1xzaIZly4OcN34
3OtDH8K176znOxLCbzt3ijRSTXXmgNJ+fcgCyZsOPa9fgTmXe8KRkbd3OTuQNvXu
m19Qyb6ZtOZoIW6jL3Jz0XrfdOm57es+0jQaX+HU62GvVirnMpWdRs65wgw3s2rb
Rzlq5eHJH97uhuzkDZz5PyUdKnHK6bcbrROZ6adKsU3QzDj4Hlo0SJLoSsseYcwh
AdDeMJVveSMhsJrX1GOFESfZFo0FiUvRvpeKTyRwmF2uPEsfFIj7FUYf7Av4X0Xw
ER+QvoCk0AR6jH939cWEAh6uf/CIMPV+UcVxotoBXqoNHRn/MV1FBrIAu2H5WXNP
I56pMOT1eokoHiHEbRzHg5pkR+x1vixb8dcRBK3O0JYPbawwQleLDfiz0gWZ8KoY
6QqkRXc1poUZTofIhWl25TGeeJr562C4XC1qfBapJKfjFu6dgq7o8ygkWfEiPdPZ
APDCJ7YME6L1QQ6t2xAwzpwW+iGB8e8gUFII7jyKmMXn4Eq+EvaGarkJApq6RqxT
WwhPwYi1gWkCB5WKSjYY3dWC0DLqxgCCxcQpwVmqmfIgNH+S5PqbqhvY32GKDLtd
HBWJNhW7ejdt9WrtJTngcEis0Hp92YRcZ4q0g3ZKcRZ46WTwIC7d91bM0fibWqP0
wiA/lDj6NGanpQpO8CqkHrzdtg53US3aZTVoL/keu6mTyPpkNIXP3nIapnnMzkQI
vs7zswceIFtXMSR5urcyx52JkyucKcGDR8Aakg1/Rhn7+fucJH+WVfGUcqm082Ho
UqSDhrzzuQ/U+H/xPqHiok3OLm2HCCXSejsyj1OtDgMzp2z8P7XYERowD8v8gDHj
8OLBiM2UlI0Q5Y/NeWXs1x+JUjjuNDuCYBuo8asqdvAPcK9cJN1WUn7ctVPShv38
L9tquyrcpp5i0vbJA5YC7ZJ9/aLcNOUxZOuIncbCLjYCO/4Ryb6Srq3Wfs6XuqE6
2TDtFo7euYcuvop2bERTcODHAL0BjyS17weWcMw5QR3Y8CEZPec8vXnNiXZVTIlF
S1gM71Rgbf+WcWRAKSIK+w5kynYKdnKFLWY4mav68uhw5+pztnO6sB90gfkTQPi9
XJaAA+bJ5ibEzQ3K6XSWOriS293XYqGy61lf4WYZD4XyqJX0uYIDWjfwS/l5c4q9
7jVBrxLRZAaI8i3iOK7LpvtcQXO63Qlv7FyMb/b+Xj6sLHFsKH0FrwQPQsF+4Ham
gQAO1rITBysTGhshMlMH0QfgM45Gc7Z11fr6TcNbsl8Mg/WdBh6ZXxTXzJeWyb3m
hH3J+9YgO11yT6gA0V8clBKpiGCLbk+9zPQH1BeRtRbTdaCZZnH2OkA+p587jwCm
sAtrk7kN1jf25M0iYXl79Wnx73VtuqEgICG83FHiwA8S9eUfdvnOCyWnGkW6+uHz
eoQKiORhhOKjGGXKhmsU5mdkI3zrFbp2fAVT+PfSPgWaX9tt21Af2f3aelcUd+ZW
9bk7lK02z3ssOXISTKbcObtI7Xiatg+HuSshB5WCdR1/kW2dojaKPDegOijj5z/8
Tbgpb48x5x1wAT5VK6MGH4GnuBsbbSMC+mnkU1tkgduSnVPjushKigI/BHD90I4J
F4eShXjuLM9+SrEHQZf2bg+LbvZRhWDRvcwsF6rBImgbGLGOJw/FLDOFzXQgPtns
aYXNl1tf8H7P3z3kZde/AkcHORl1PEk5T6Fuq4wo6sgcO8ZjcGCGrApq26H0e1UW
oVERlIt69a9w1MvuhNmKUb+JhJNyKGffUxp3WUlwsCh/AilrvppwIJmnNtteywCN
us+WOu658+vJjqk0yc7XR0KkVuymGTL/BMYWcDR/VyN//MHz/Pscw0sKmhHzIo2r
LPnXm+dfdWrQsoZ4UnpP5udhuvRncHAg2HHFpyb+hN+0Jf0mNFUDT2/g8bPFMu45
QqgdaQPcNLhmqx1kLOA10H26s0ru9Gwj0qYPKJ0W/E2p7XexuBBK3ZEeYcEW7N/c
D8aq6Q9qJCke3dI4lQQ1ZPWjAR/J5V6RGE6cNJH7FdpNNdkUUy1FNPPDGx5yDg2v
RJnQ+XjI/YOQhlEHO1NaHA2EL55vWPUik9z5+/O/8fM2lr9LxWAQxckzFAdZRCal
GGTyul9GNVquAxZv9cYlirXDtt2EOdw3NmZnqoWoQEuZ8++ROcv42Ml63nwhsD0X
IicpqKujZv50m3vryx5zVEAPa5ZPBD+6RAURtt1VQlVFjJ/6orxkv6A6CZ5LXwgn
f8b7iytqhf6zTBzXKc70v/t+Oi/J8n6mk81Nq5Gg3oIUvQ310uLRR0MmMrunxjta
ZQ5PuacHTovhEb94eRhl7cKaPN8Ydo2+sU+30vyfjGD2YmJzIVmIIQfRav4jYF1R
GWUmWG9flBvKldT2ldfb/wlSxyosAhFynwrxbHvW4eqo//j+x/Ftth0QqVoTt80O
JKPBMA1Pm/rBmfKmotTeNW4Wffng6NSX9F3rF4SgyKPTG0Uf6jp+sIBTDj4shG1r
5Yynk+24PLMcQd0fRfkXV1gjrxmnUStD2o0XIgj+cfGDJ/S5rXTafERItSZR2gVD
PyFo+L3Gz0eqI/y58Z/oAajDRGbZn2uQrQsypUR3PTC1PoLWBw5aP3RVeiAf5IVH
diX899ceMrlUwYYbb+7Z/Gi7kBk2qiP6pojoXzebSo8FxA3YMNzSbbcqlPtCcJxL
kbGISRAryv7ww8MXvg1J/ifaA/sLolmNC7W/e/p97pkSjsYYgTjrnfONC3m7lrBt
cPkZOKawthQa2DCe0Wcxj9oeZuUBGiky6wMmgjhF8PdWDKnGevwVi1ZdF6z5dMwQ
1dLQvkDbBq3w9+5FA93/l0wvrRIsUtds/hzHgtQtyzoYqlWkvlEG4Z8nqREfuZId
KfvSqx7CvqHSnbU6ROyCgTWzQpjLx5cqTLNubxz8Z4hxKZUz7lfAtuEoT+VKY4KR
pOxauC8XH+2hGpgOHCenax5gDovRIeuMv7CiTAVS1qhcr/mQrcZ/esRLG65D1UuW
OEtVTyRq5vJtpqyhEAyyBIfXmZOZCmrcYYqhjblA1Mf6h2cyRDDDzn8dMSgM6Mnk
+S3SFYm9iDNV6mqt956GzhUF/Q8AVBXmo+ddYZnPxk0FdFQtCVcOCdRhRwwca6IH
P2xMoNprsw2kqEpao3lAslnml9dDZeLT+7eMQLI1viklDPOe8bsMq8zy+GtqLeDg
KbM3IyTK5iicX7281KczulhF8654J7RGti6+eIGnlios6NTGn6AOhHO8Gup/sNLP
MHWzK7xNVSkG/x90ryTV0+ZU/eixREmUEl0PhyMii83cYFfPhf/f2T3MLtyCIHBC
qprfSABD8l08Mhczd9wBcF1YlNx2B0EtsrbkYCx+4bRIZI6TE+BZWJ6YGszduir5
kFGTvLPvS4r6prEvWQlpZQ9EB0htfzvepCl51SLjsB024p16Ex5gghd5cfzO8/RG
idAJmWeHXR7KEA07m1JPgZTzFO7krTg6v3jBbXxWacCPclgqEfg83GqtahgG1+Fg
UItFdxck2FPywY7BQWOPCOWQ2PgJufe2GrHtsKE49hGusLS/g+wYMooEr9DFK8oR
+ebg9qCL/wpSay50zAaQGBS1YUWjnyqdWDh8NTmppPc+6wGU+wuMjXB+kv7Z7bB/
wgrSpqMJRU2MYxhJyPjp7gKv/RGa6OoRwzjhrJZswhTbapl3xYIdPv5TxclT1jeQ
L43SmIF9pI8eP8mtMC7c1NToFgONVGSBm/ioHkGs+85FENcCZ3Md6NdmZnACvANN
QhgVs+ycj+IVC1GyCosFtQU8qUJrt8ObaORvJx0ovNY2wd2+6cewos5lNW3K74hZ
QZhCR2b+zTKN9PipIZM+TNh1mBr9oVtPRzRShQZawf0dqJBt3wziYQWvDOGhHksn
LjH2+PrULoruRDJFTHRAc95MiPUPNLodr8jRjb3s1xtFGURSma3f4RQUHmPD87Qk
axbRefZLXL3nrR5rwJ3o8Y/WRxKUunvJWZTozWw4O1+8/UqOqi0f8Gw5W8e+y+iM
yYJ3j7309l/0dHHVf/PGH3nFHpE5x5kHSDzEFi6AWz9UDeOe782xDNk0lD2tErDH
E8FRcgKp9mq3Yj4gZQhRvxwu3ZXIbYkfBZlOfYj5vf7REaZ9MVD2JYvwB3kDEkEG
+J/5uStQTp7dgGPKWCRViJmYyg6dn2Xc+AyzmzvZHFLzDE2rTmSET5bO6Ba7/6vE
RpI44EvA3g37kdKbTEcILT4ducmFoa2NjX3iAUAhkM3AmyNUpRtnygC/nOocO6J8
nAsVi4xdYqnjYJOkXhj4mEgU1+C/2uYGB9bmrw+0lTLmVSQPKHVE4ZiX2HDDwwSA
+VL8jgo63Snbghz1Jg3x6M31Y62HcVpMR7QbjjQxGkGJrHKu5ojs/PmtEfZZiEX8
dEiqgGQZfB6vg2IT+N9uJm9ltH7wCVhVyIN1MtvsBlfJFpNnUUQP5PB7sM4nK5ot
2QewCwJYeQs8vTekq757CHN4BuX9Mvo4PZJ/lRQ7AooQQVW6437lQsOpZIiolRao
1i1sc5ddkFvr2FmiaOsHNJJMaZMgU3pQbYgJJdVzZNwAC4pCIF5osBgpdgAHLwet
so+WDvYpV6wGtnzjInW8px+/g5Z/53SVkk83sbC1qi+dn9GVtk2Gp/HFqsNDfwUr
QRNP4iq0B3P/NI208ZXTloGgEhntS//AJkLRzmSduUQfeNSTtES7gVWSm3ZTHNP2
6tbmgljuQuUHEo6w3e4PKvBCMYuwt6HtIxwejJJYA/9rbaeP24QBBQy57v2yaMip
kaYIgP03+mOh42JICSMjNtrFgVkLIv0BEdV0miu5ibancmCG7mR7NCPfpqsxgsnj
dAb2Ln8y83I/Nvb4rgJ/H24/uzV9cy91fA+c/sv4VtnArCHd/p+sNzpYA/VfV7+X
ZL52U1VR1bhASuhjCC2xuLYfFEVFbPnBqZekCK+ZHIWlL96fs5Vm1OvWBjIIIO1z
rjMvEvB5DSv4UTn2PmPkxsJpGsy4wQ2RmvesFjkt53XJUG2zCpQkEUiWZdZzxxzo
I2nMpT+S62F/uocCvW8b1eWghcrZYvZ95/NNybaDrh/3Wn9qrsBoSflQ8A6LWRvj
+YDCg1EaqQG3/pCt68RlukDTIKNW0NKYOGjBnXO/ZU+JMG8f1APNo8RzPYCWYfj2
1KPBfgOLnwBo4atUNxWK5m0s4jdl0iALVkxco0UcyBFxs5MaaRM3iReJbUEcWr+T
Qg9KHMLIhdywHL79sDGvVPeZyYMG+k3gPx7OWS0UyM0rNKwETr4xZeNkaYYiTU3b
+QUalmb2RBDxC7bK3lepMDlyy29qAhsQ8b1f9FW304mjfBEhXhgEdkkxZhCkgU2r
AKlyJP7dN2J57s3huRC3MN+rvosGOtQzl752Q3OHxyYxR6mhYQ4fUAEa/cR3jdvu
IoJNpHh1/tKhGbGCOPhciTzYOlGskCy+Rh5Eaf+BC+nEpeKERij08PfWGUl7Cu+i
ohHiAMxyDqzbDDEYKhoSAvq5WFpMVIitXhQcgWcSvsRxCysRez+F5pF7fpDm34uo
N/8/nrkieuqcxDd3m738bkcQ64sEY2ABbjnGbzTrHSnBy9yoR/x1vp7lLpAE43Ir
z1TM17TBZ4jpNQa7dBMZzySZSoZW1mr1XYyI3h0uCp6B3/B4kjppnJS1NhjgsEo/
r9qC/4vwL7K3mKq1O4xDKJsqpbHPn+wrdnutxInw1r4icBRVHL6f4E2PUEN+3hI+
zBniZWIj+J8uz3PMPhcmKnusM5tqLesRme5itq85eJUPOefGXDi5gxD7PI27xnUm
oPAwJcXY7Zx2NtDpvHkHNrRHZrsgC9nAT0RBqBwaItKmDZuLhRqtEdyT4P8rX0kA
ywCPQf7XGI7FjxMW6LDO7HjQKA+IhcVXALs2HOeyYxJ38rKeM4QxXp4wTQTx1bFF
hF06LLm6SPpzhyKQ6I6Cm/Xgsff1TYCrZEsVOfFxS9ZlgtS8uJ8VUbzK4rGBMGga
I3+ryro93kUDLeT4up7KqgDA6m8gaJrWt2xrVMAg7hUc8XEgcYjkCmat2dbgDRNu
5a47EIErOC/a943w4BRDSwYkUvRdw3fltnLuIcgRsNmqm7veyAEGbD+xZAsvvJ65
ewrAu2KouzPxnMxw+Ii/MxE3fqyYxj5n1tpAFG04dtMcP68sLA2XrIW95ha+25EP
1tBTFJyb5iUwmjZn7ikvN9FIOiGjezo5l5qfzsqi0ywSaAU9A0Hs42bRPwzT3RNl
CS6Ksy8GWKLDIA+2FTyJLOI4WZtI47+oLZh8OWlPVPnZ25iUR0UlBpGu4jnX3Ow0
uYKtPOZWfoCJj7bsQi2dDba3ZBqiionKHdLP3imLV2H5ZFtr+W0T/1XIqEqUUHua
EeH8rGKyNs//pgVydaf6D7wOjA48upYjOqCgzEaU3tjbyMRua2cgFyCYfR9dAtpi
lxO48bIx9vdrjxUBdjfqghkQ8n4hEGvxQB1Xu9+r+ckB2mk8FRshJ+tJ+LtK1xQQ
uSg6sg9eSuTIOn1IdKqW6BP8pduSakIw7ijDtGAo1H2cXP7uGbHqTIuTQZGYVf3d
eh6mkrthSqSM523t6dVERuOqZViNXn2I5t5lkShE0+sNpqCxFaw42kKY6TLTCqwp
Qq8XjVSlin6Uyjb1IlmVjSti1QxqmhxLN4Y19WxhuMaTdVopTV1G1SaC3VUbw4St
RM3QLpT04ARJWnoCGR6gG2WpSQ56t5BV8QF8HgitHlCvsjbRB2OwgFqYnn2FNGqu
nk0yWvW7nwbg2MZYbDUsx78lI5+ejU1r2RqIGqowxjggtnyyeW4wjKNHcSasdTv5
Ls++X8wSCUxFLkLH456pWfp7tBtwyUAX1bccnwvGoJ/Liy0p/A9uyIkxJtDdwWTQ
N8v2mEb5elCyY1nhjDwRsaA+rOkxg/KTDnj9jQuo5RjgMWoIvsPKn5nepFIW/lTd
bBS+CiLXq+Ac7tARW//+prDpHX2WJFtTXeup+KF+m4EkBhr9y6wbjKatMRc3Y/gj
rzRT+KO6C2fM7tMtfho61dpKMvAuoFF1WoDE6fuRhUUfdaBNkZzjbtjNT8N0dQPf
WJ3k0WqwzrGaT9FuBq7j/Mjdts6A1woz9JTXmPQoAithrBsNyT+ApmVMkhj90x/O
qpR4qb/+bZzNslo3WPsV2y2dXIWlCrQiwgXuMF0I/0XhjCYpF1eSYrmSEF77v26K
cvLFiTWBdYrGC/UbLhbPDp03FCIF8/WbBgfvVa7dWOgomxk/NlojT5mCXA2wqHPg
LPZXNS7qBPvfVZU3zZ0dLkeBbBqYp9cV5IKpd8ALr2mzCh+dcxlEmkyBssbTV6F5
7T5Fo6Pt8GwR2zKyoZme58CjhFOSKjjetYAYBK3viz8ic0Y2f+8rd9WYHz+VUPoS
`pragma protect end_protected
