// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RQRn81DmofkjEi1z+KZ1GDHemO928W4jfPX3S0MBBRPk/eqDSUW9HCU/iVjnz6HG
3ZcSVgWqzNGb1mwkEvtSjWsVTDOjckyx/m9E0OXQ2OxrXWpNwPJe7ENVgXDOrD5y
hq9kahzrl3aZrQO5zZgzfJdxqXPrXq197VDtx0ZDT0w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 62224)
1D/j9n8xGlLTwjpP9D3MasJg8OHXu1MBzgx+l4dm99xvuv0/9REV0nF9kZuK5d2O
+jKUkTVuWF5HF0IZsF48Ypk+4BIUMthlNq4WPHjd/lOoMjN0Xs+yjU1BhjInBjgm
EJsFcYAyqvpUsAYJAxhjtY+TG5sryBzNC5opx2iVTU1oBWopv1wikEwa8GM+oRxU
lVnhNsoqSfTF2HTSmp6ao18mSr9Q7EJNcQi0vmLrvbBJNBqVzJkiI8NtMkHeL2ww
OL+BmZM72GGS87xoCcvecvpPMJTiIuZAJIzItXN5PIS45QtBJ0+S0M0pQC/nnQAT
bG1I6X0BjXNUMNXTes06gT1FnmT1J6gIpzOHBAMj4Cb+5SkRTQfEy8rlWR3koNhw
gW5WC3CPL29ALypmHfb762SkfBn3OZJGiOFhXsmtCPrxkWSDsETVtcEH0Fxkm3oS
Z5jDyQtdJ2RXa9K9YXTrWOA4C9nv2iKq6xfIqRZXMFwFevi2QT0Du2R8U21Mv0sY
4Fgj48JyLVkHnq7gUVHVy4I3xGWERVSU2jCpSpLbMdyMau+WtPWA+daVn9huHZpk
6hSs3th+UywnlWhQuWpycW9LwzxsE7BIzn1pSu87+P2hMnLo5Ux6sI9cTYBRMmBk
NwZAoCx2iuzFiR7XXf6iKjenVVezHX+4i1EsdghMCiQ9A+0Wr+lMXH5c6s9C7KK2
OLSPrHXfHuSWKw1ix3uS6rD44J2C1JrHQ7KIzbWw30+vcC2L4Sp+zmciYpCKoi3/
X9QCK7C7VZQZEK6M7h2tvY8Mx227rpW2m+IxQ+QQNQ9x/rFifxrd9Fo0CZfX+dl7
CLRB4f3j+mr2KwRV1XKa4WQoJvPd/mrUhkpmoWYOAqv/ljYm56DC9LzI6gY+XHYe
EdcWc2KSANjneyvgvLv1CMMiJyGwNex79NAfL6INNWIY3/9fGC/fzplc40W5H1me
ismbmi7wfurWIldYlMmdybVyxBtp7NQBRMXqLoCf8gyT/76h39gY0BlJZbl6/8YL
Q0Iot/RUYbnfvit0jp63HXxbQ5KgICxmfVmMZF5YjMocQbNYfaUGwvhrxPD+Vs13
IIraXR43OzMUNSbzaSJSR5z+UzbBvnsryJh2Qw88krcZIaw9Wipwa1kUL2hCIgeu
FfpZzptSUtv8hpDgTOwMKuDVsJfyIxnp7uaMPLQMssvI+n1NTltwN8Uxi88ySk3Q
QIKzWLZVY+UaD79A9BQXh1/HhwvY3yoy92j45fZFTip95hpWEMjl5fTiZhqKQCR3
g3YmMYZ2p4DXTuhS1nmtYYJG873Gj2r1YW6zxdDWK4A8xUYHCEqgSeclIzXwPTFI
vQiv909hIEd91SIZC0jfknhFdo8R9dMcw1EsAblZB/HyITPvRp/z3cM3z5pV/qce
OZ/qQMcpl6NjqUgc8ZEEi/DMhne74KoVdQIsR0bosNeNGAiKo/kNApj0l6n2bmw/
AkLR6qf46ZVUyUx1BKVc0Q1l47Yhv/XPEtIrhp13PKS2ieUoQ1puOgLNtVI0pJVB
RwJzxlW1j7xx8R3ihsHeTtkgNTMqdO2b9DFXumsA6UwDp87y9d8rNxGFNFq0ivLf
WT1sqAa9VdhIyEc0SoEtxUIel2kYCrdqUghD7eNjP8cA18XuGFYe4fyw05ydd6DP
QjB8rjyeBA9Ikxp0yX01HO7A2lhr+JB/5Ms3w1wr4UIdYmsNWOf920G2oSrNf/jc
4e5neDsaX4057l3SFM7uItNaRTRHMO5I8Douax+7HfOdg+WFjD61pQcELECmQ2t5
WuRyYyKNG8/MRr3lS1J/4pX5B/EUenVLPh09r3blCmm0RICG/m3TC6WOZP1DwcvF
TELh5kL4O2YMiQZxmOV0/C8Q1r0YCKtw+/L+iPDmTyjqiamMyP81hmS/0t4wkn4t
XlkRZwnmC2yDNRLa6INCW6HbpIJhBozoanJXfNZW5Z9wV3BkYxdKX8TxzdJcn6sF
yOGGgy+OuVSzbxnqmB+TFz4Cul0nCpuFFgbKToDmgd0kgegfTzulEReIOuM4Cl/j
9TNriBBfddKPCl3ue4trtY0cva/CvYafTvs6S+ZYwDVooZ0o0m55wSV1tFKCdwul
9G9vRf2/JPQR9Dtc9UPItyIUvdbkpnWEqxL6qx2gx0+uDTtGR5c0NfbPePBn1IWV
tdxQvvItq3vZJFsXwk9P5G3PEolgw/jcTQCt7ffM0S2/Y0HdZKjTdSjpxmxCVDCh
4JWNhRWSZxYYh/XSzL3NKDg5HOrnsIxMtE/jFHOmoQHjTICZnWjN8J4bJxZsMWKk
0I/x4fLAz3YNcXYYLN9bMfOcBkt6ASl2IER8HRoqgTsfvopdFhTNeoZTauJaDAs1
JRBoNx8dKUwr7ZRYZLuXsfpckNmcVcLnIRdQmHCspQM3k+p80riJZOiWjqyesAU7
qdJiuEsNVa3XsdF1n6lYJNTPv419qZeqqB5Rf2ydVm+19bVTsdYl2LPIvreXgku3
W27GUL9v5NjvoAyAbe3cIxM6XK83gmrNTDV+djEr7t3f3DrB8vHDX/SCTbU4fOQg
WdrkhugJzkgQytArEUGFPS2GxG96YeY+QJIZud9iDZf7NqLfzTi5SdraJ5QqBCcx
InWFiPAFhe7rtJCzlGR+1xhlwQwOdahlK1FeZB57J4QbtNIrY/ULVxmm7TBvjXdd
lRw9zdTvU3gisKrAm3rUtHF2oArWi34qFLBVi832sJgv1waDmuGfrc8Qo+FGSt07
PX7UgtDRPL3jiL9uJJFljjFUV3+40f6vKionT3xIQq/7qodewcjCTTk5lTolVfe7
Fp4I/tmFqHFQ9Z2thS3f4k6ZPEIRqjw4zvxOUk/Lfu1TIdkEXOROaKN3EnRupmFM
GrLqIBdRW6Oh+eMPCpCo+lag/xIfL8Jk4RyvxKFAu1OTmR/sXQDir8MyBXlBCpzE
RUl9RWzl4xzN7NW3OBIVnwmzXGysEUoOnCed8mdBsH2gY/3Ao/bpfZw3UCvmovUM
ku8ndiwealwvS0aRMs7VgdxuFzacv4SjO8BkMsi1+PejqcbtE1n482Ca1oTE6mjC
xDE8hMghUj5mBjuHV3qKCNO2KhHE0qhPybFssNQmA/Y3WILwB0WJfvNQ5Z5FFHAj
5fLDtMHqBeLnAWSZk/5kMrFChAzXMqZ99CqTgc0nv9wytLnafn2wh68l4VM9UWwR
7+GKxIn9l0NiMNAWtKHJ0JUL+QGNoXDUBchaLu2R3eEVSAnG8+ZDaTwI2vfbj7EO
6L2hPsV8YPlJ4e2cE0zLvp3HB0aJU00TPJ88vKWnO5ylh4457Fmb8dPlk8pmzR/D
FKAObt+rIeE11OZLe8ruQp4cPnAUF/OaTk+vPFOA7LOEgTRSEiP6EyAhKIPWdDzb
PTP822MhHwmXNbMTAeSGBPeMR7vNIfc9DYpa+FtMT1icPxlcmvXC/BAXYYyQvGml
BFMw+LhAsoYlYjAIWjqjxPH8B06GOhTlaDsrbDVUlLhrDsILuJlTxAY/KODkgKNX
HYtZEuXi4TfDIo5fsR0Ux6SX21nj/C3dDxkkxSVnWSEn6R1m6TSijF8ggOSvg7pd
wppkdSeMf0Pq0Ga67Ayy1b9Mc0vvi0bsWV8DNzz/Eo7QIQkZwsSL6TYV7dTVhknP
FHVsmGyG/EdOPUjhstsrteiq6K15QYvoDNGgBc5pF6Bg36axfJtf2jDgHuMzkfpJ
oz8BJ4b4XWObqglXVDCUPyZ4IEQ2v2RGHa/r1p0rvA0ASdffhzhL6rI2AW8uye1w
gkuAtsBYXisW6OOnumlDAyWde1cIRA8LmNq+7PS/sFtZ3MRQK3JMViXkHXA0oqks
RjfjKyBfaenkGdoJFM0vJJlmHNLwFMFFqH3rbulv4XyCOxoIAg4QyTTq74wG0aNZ
a5JDqHkQSSve1NjdPVtL5dNdCx2lB5UIZbzKxiQvOiEORrm3Va/3O6+iwiseVy2/
WC7JYUohVPhiLLxnEXd7UWHH+YFGLTRuvYAol9QbnmC50KbtfilFhESpEaPHM6Uj
WOrif1ur3I9wmiKoflbNNAF79TDYPrGUId/DBeFeDnFkQMPcJzh40szDBs3Yls7U
gRpgPWXyNsAG3ystKUhqvI1KxClDljXJL1UBycmrl5plLpn88fi+GtED/QMwE6Nv
PSNmjrwKP1kR8XFGbjnxL+3rakeHA69gIWL/bzLGxc6uqyKuttWIy3b0ZYCmI08M
/v1CiBSILiDcXnWm9AHITm9SZfZCG8bfNDtrAKnYIBPK81niW7ZQbwpeimuqz81O
5yGMOhnLXYpVC5fXIaz+090iJAtwevKIjB0G+kAxx49b33p9/9q94TEO2LfPg3Qw
8flk8+fFCWZ+cb9aLrp0lNrqYfsVsd/KCbIVyluMoNPhnIygDsyTpZxEEHs7tU0K
kBcZOkBw9tH9yTCMYsei4debJXkeXk/acfmg0AqekPO4p3f2Z1ul5UEI/erHS+tJ
fK8ek6uCQb8PIEivTLNi3SPwa9KlF5XLmhBd/C9K0vyJth8fXnXC/twrSjqmiR6g
IDPnTh0bIRnFVVisuLDlXuPzJ1w6q7dpMVn5i/dPoQAHuhyhTwQwVomZp7hll5G+
FoQF8zkomoyNIgIsSRUrCqZmjU1R79Yj69VzPDYLnm9gmGbfqPF3tSOrgnU0zQ15
G1mWdMjWsze5ua9WnOSMm/jDYUXbblqgI9p0STiowRzam3J8f9lThpCRl2T9DgeV
dNXyP9e5rw7IZ3GM0oko/JYVX96DXSLLlNLN6FU8IfJ8nD2C2R4rcW1OgBdGMuuU
V+ji6LrXFuwCPtGAm37jGk8l3PfuSGMrPZvFNCKRm4YWpObqqOHMW3hBMhES87m/
BCm0YGJcaWEJHG0hff/izq2Jx9Lg4cRS48T/9TSDTA08mSTtZbl2LvejeoaO2Uvy
FlsvTKAdh9Hn2fOrdVpY2Q81/n8Y9uRR+NmO54USBqPsJZJltUs6c1VZygDQOLzT
jdxzSsOVGTrbPKqL4WRdlbWuG+Ds+zOvyugm+kLD4WKIiw7A+GLlG7SS4ZkNjwS5
muZHYcwxGSYG8LkY3v483Z7Hga9VLpSftAPeih49M99W5MfaueWSNXMIGIn1ZVmT
l5gWSKe95N+N22/noKf8bgpsDZ8G+asmWMrlRqD3M3mP+Q9yHRofILNIuBAgMDrU
z+PWEh3TMF8I2DhBUYOko0RndrrzQqs3kZZVR+Ho1eZX9B26PCuSNpHVJ8PVMZWd
YBYK0WxuAyax5KMbvtMwQcTu8VWTYTU3OZZeVSOiRS6xjLgi2HZH8m6O6PC3coVG
ULNJj4+UG0vjyWshpGmgMmE1eondB0rMfaXc3Th/h+sxw6YSiP/0/49w3yXrV3Fo
Jp1OuRDOXsfO5nK3e94SP3+nPynZVYG3eEwdc2OfCHR/D3gBekMSP24MeMC/6ytp
QM1vNxPve3vChTfqocCS4adoBpP0CklWoQVtgEclzKfvEI5QCG3L8uNcoNgOlnuT
hBRTB0d2FrJMLj11brCIJfWkcsrgNnvnLQplR03IOTL2q7mI5D6KH5aSr55/DBId
Y030zmYqRRolXEsLcXsAEVoyDTwhS5X0Iyo+RcRpoBLEdVM/ytgvnsVvEDbqeKMW
J05CU7wHiAE7QENmmTk1vYd7wGFKlWVXg4Ths2tfZi9AzdWxnlxfnp9Dc9IA68CY
8Lt9r5qjGulcjMkVvqVRcxAr72qfBKiqxKoJ4goyIHq+shqGv6HkbPL9QTEy+r+V
1P86iFHXctBex9xPD4fJTpa/MxjHPPXSArlnQE2EhNq0V37ytBfKEajGyXTEDPj7
c527eSAIpMmjMveQdM0KJcuRwECJbeNwQDSDuBrrh+dBcGCIeinNrAx2Z0SHi5m3
8q6m638eJ9eHlZNocJeLsvpluhDlVJFwzdxBR+9yPJZafq9RXmbERwtW4TXTowIJ
gq07+LIAwENmjK8KIv7xgI5Kc16xt+QCCz3vz0eCHIEyFgcAVpOgji7vTFusv8Wq
I56EOwmsHQrLz6qPmyZkZA/kA16SYr1jYzDyizO30PppJAeSblmHS1AKwmJpkmpp
0EsFemIopqq35KYWGFOggVjHKP+XT3BG68LVWVeeY6K+E/BZLFuAJx9g1BLsjjXY
qqNoYCZ6izI11hlIdoNCLu/NnoySHWOHUIwuq0c5qqSWTpEyHS6dF6ppM+dEnuLe
Gvv/enLS14c9Va+R0iyt4ae3epEADW7EIk6usT4XKLlAlm8IRWUZXjtOFcRfn8rw
24COd3XGAMSNlJxOp6CTL3Z6kRnGAZzTnWzLU3wBFsEPqn2gnvxa4h8wbOTl+P0B
QuifNtsYAIul6q/u3y5/lnivMzjqcskmuRuHlK19n2cZSVM90SM5gwkaK7S2lzmW
JsiuuqVuV8q/9+STCJ8UoLkNCCleAy9HQuV4lNHnPI2iM4uM3S4ZHw1aueq3RFwa
1JZe1qx0Jn+0iyS4GqZSeVTnqkhN+FXCCNhhUb5FtaoU9fJRmnjX5rAJeYuD3utX
apwpfwT+5d1jxyskhoxT4BKT+vfQbUxqS53wKQCRTDmwuhp0GTEioYuII/OSSJsH
LhbcBFaz3JqFZkZNz/r11RTON86djJv5vcdrlJTETqA25XM1fKdgTYXd7Xh18BxN
rnh6Ma5q4Hs1w1EcDR04d3SPIKOYisHwKvuJ3q2kE/A/2rIXp1qXZ6aW1Pqyi9N/
24e2hSPKBXWkLSA9nacCk/XAT0U4yCYoLojRodCqzpJR20QZQjD9Tropn8AFQrI/
FtvYZ0u8zcbxt5GopxFDLE784314wtgnEjs5EhnaxkkZ6cTmULceBNkQBPlFeuww
grwyQ5TL5OH7VR11Auq9OfC1NJg1QO8DmECa3AsFjhqjc3+f/2VI9EgRP8vbOD5t
rSzV+XZUA99zeuW/Yu6NufOPFZjjDeGJxDZzhf0Ft9jn6pPevzgnD7/9s3lv9buf
RYQuKwH4McM/aaNWiQTH8lldOZcRJAbBFrXCngJPQUtJKXLCkeowBLLMv1PkvtjV
xp9R28sdNiRxTS9ahnRe7h9/Li4kxtEhZNyhO2xcaLgbGELsK9CzcqpLitvmql7q
p9sPkih2Y2GITEjvfPF0WERP5f8XQgYktdNFmXet0z0+I45qr4bbsL62C7pE/BaT
xD9lE7N2K+tMax7WdqHgRmscY1cH1siyTBx8dHYCJFykr37wsOoYKPpl4DezRdzO
jBfgr5gIF7BSWOGFzrb8Z3ylBaxfjEA3QFAng4kUQkXuWYd/RpFEhEMyDKHvP4tV
Y66HjiQ/vYtec865pBnjkX1DnMeWzLvBlTB7aIyFQLIiER/xAqP52YLFXylSx31U
hOcMq53LMPgBonBnrzeMNHzt8ASDQQs1k1e36e3DXB8SqVutPS6yh9gPvgwEHE/r
0eQL5yJPhi6LwETWFfuayrpiFTnmCxxpXJMgxCoLq7Cq0pQ0tb4rp6XkDL9oK+hd
kOezCM8uz/EL9b36rXjigGVuyyil64mxkUarU19Xj/qY1LAMZOVZSO1Mrk1WV2a1
/GKaeenJtyCemYymRfvH7/wQWPnGF5OglCNJ4vfrjA5vCi81eEgXJyi5nVvkMP1n
SwALHvq4OvA0ER5zvGfdTgZyEb7PMmCBi1pavNQXOIbbQqLEQ9W2DKRwFyp2alEl
YM0tcDKNkby3FDo8xOPr7pgSMmpaSzwNsk3GnqfODLW7hq2AbJ/qj5z5ap6JrJfN
UcMZwHKE1lTsyt/6GwwZsY+Nz0M0jUfpoel/N11++hyyUxfCkSd3qHLK1f1oEkCn
ylovx/bFAnwFT/XuU/zkYbOw88jM67bENSCmYzGL+9rDgM+BIzDQ8VgJt9g+pLJ/
dtIP8ZwCAqUirlHFsbDy4e3nZ0bY5UIsS58MldcCH7aw3RVSTMZjbfQ9RNAEiHkq
uZNZa7KQgdjy/+jn+a71BB1GpmoQSBt6RBtFAFmQ7D7IkxzvE24eCrvzH/tO/Acj
JtuxI1Z2NaO5vwpA5kYaW0XZcQT1IfWqpWPl8ae7Ck/CHZMAsw7CiHN+wAcjDw6J
lJScB+kkD2F245AplmaIgtr8r6wLAcrEocAYEOeCE4eSjXE/nSJzrRVRnrfgOnwM
mDLIuOyVnhw7HEXkV9TRm1IubLXhPiocsQ29VPmYUZo8pZw2Mq7Y76QkwYLajjfK
P0Zxg6J+ctRlaws4HrkP4P9fKwbZwPFMdISRFHxbYGKBAP40zQYl82eDhzpLBsKv
qSB6w2595zUb44RaTtULdxvuW7yQVuKyfy7kxd5yg/dOISpors2vMZzlQiGdMr/y
naK77lygOOWUufn8RTPuod7iMnyb1BMu66A7qQeVxOwPz4ZhwvzgpV5c9ZbJBpEG
7a0kkWYWW8GxwCUEF6VjZ45KT3o0E1yhcdCYEym35vWr/jserOyOcD1Hrgp5+6y+
P3uMbcPtWQxOcpZYWK1khDxln+BhzF0yyy5xguBo6CjPvm3poQXM8NvPsp/ITj4C
/GLz8CFNUaPh2g4qJfysoJ2UYl9dJkqiIXaxvmZbO4o9H0CZTkuLSqvmEbil0gt9
+sfQ6OtY2hwZtDK39dw4hLbtSpi2RGakzMU85BmxmgTUB2rNOtLfZhVREtTPiKPv
qr9u1oVy7hw0+RCevIaw9jPGtbt6MvBAgsa7/pVlhm9FOT5YJKi8Xuxum23vl+oL
rQ7hk4lYOiWa2c2UExwRDEpB6kBS8JQu+YltXegZKoSTOZI+0ZzVU0OUeYqMdAkc
733UqjO0x5eqJNQfRAT3Bz2FSANJe7TQFWG3FzwxD5A5SAvkKv0qjQMLvQcV9Pu6
ULljUVW3V9Q4ajGClyv5sCJ2hUnP4fChqfUaLXoivYs/dc895dfPdZ/Z0pUncMHi
dcFc/HjUtvGUzNA7nI/kGpC6A/W8zJYi1XSk3arCk7105XVPJ6QX8uD5eF7nAn1a
pivgsw0IqbJqZ5mxnxViWZheb1M0tQfFxKdjaoY+LtvG3uMW5xC0G+7e8dzGgoz7
biqfgCUaDaffuUlT4fclkeo7LjQSV9AYASNLZR6/wdNVGqxKRMPjCqwVlL9ELThZ
FFLsBILTfMYDEdBQxgEJXal6qObdcashqrtHhIy3snhREMwWl2NNTC6/I45eaaak
uB55loC5liVuD+Zs+eaUBiFn5aiwYxnRjTYVJxj5/l6hL9rqh0X1GbykYLnaroby
iM23YGTDgd1zeAwwFW82ELXQELdZcDtOTarD30qEAik422mEcWslw76EksGXo6wA
lFvVSsq4C1rcr0J/GQXs7NI+d5oitCcDmpYw6YBNB146bURkx24Zfjc3p7T9DxlK
NI8vSxi7XsaTS0af74SpZCgMgYavDJQYWv1sWiZTWb3aHn7yf7ELjFOO5Kn1UfwI
5f19LKpwI8QNy6AuRXDViUjRNa9WMCVb9pNpqxVTmXwCLij3Ow6DsPVM/gtW0Xoh
mBNiWDok7SaoctG+kIQeS3O6pgkDlEKbLa+WSMMsOfxCTDt0Eu4yORJWbo/Zmeo2
W+GpPtWI8ceKULaht21M+5Hb0CjpPxxbhE9ZO6a1mQVbO2BK4o66AaGOi4pH6vty
gj6plNKbLoXgU1chqj8kEW8NrE5J6SKN0D86ifB4bi3OyFG7BDxvDiSwF1CeXOP/
Ebje4e0Yc6b7XijZjSrZIcFjqIYlJDXAEZE17IE1VXc3ifq+rwphSBZLpzjZoQuq
/yFMq3j2sBvuDTccm6Odkdv30LxUadECPg7alcu8GqErJo9QY8UTqm8paLBB5IYH
fgk8NqjEI5INy4QGDHaP9t8bjZOAUQmSodjNKlAW4+yMR4SXQ3knv1rHy9id7oXb
AJCElN1FclGMGwKbarxpXzR4tFAM4AaYL9Qc3YH1MtegpEqEBTIwCgsSL6SilKgK
qc+01uQuQEeJZ74plJfeai5dlzdS2fGcsjfT9PDhMtrsQrdfOR2iYCXfiZ/famks
nwN/4fPHgirVtJQPEspahM30Ura03vt964S6aYdla2rjwjZVT6QjSz3Kz/0PVxM6
U56dGeFweEDxvp10jhoOgnlm2laxcFZUs4661Zp++CCno1XECfJt4SLtxbMttZvv
lCaiTAXn2TKf6e39BH+xPutJpwWsU2jqNhAncvjy/w+KZ/ja5hsqxPEDtBkIanRu
fvH0a9i+97+iXI8c/B7elS5ygDqBbPmoRcfCsYs6peUPkXiA7W2pNUtbKVkjG0cg
PJURqqHntpqFWWg4F3TVSXR6vsDq5tMWf6Grjo1AP14VG0JFr28eaMtflCkQ2ovy
jriGzJUT1xkH1vGAu8LrFZEEbtEQh3vVtdJCpIlZh6MMW/eBgusaBvuogCyI/1Mu
QczEN5TT2VCA8ffnygx6YQu7G41BK9iQc+VFid2qIICuu/DOYpnPiRvdArz4f+Q7
5ISZBXFBpeaEi4WtPJ1o2dMKcF7ISBd6WB+9tuRNsJElTrBus3qiK8iOKMvExO9D
PaTWKVkQlqUigYhpzLCCQHT0pJCX5jSfG1ABwbV8tr79xuJ2J3TBtrd+La/uHpsS
9dW3nxa4JxoCIesW9erPz1tb1v5t//tqPhjw0lvK0kH1mR4nQgsqd6FzC/gGxzYI
1aBibXKqsqrMjlTp/mkE67xznQoUj8kZCvbwLQDi6+rTkUBDydVxVOeeKfoGjfJp
gcnr31asE3kZ9mxZTGYMeMPuPYq7Ckvoee01FeJnFxASJP/Me7aIKQV+OVvoNVos
39FhfrBYmKiUaXqVIpWEdE80gCfhepXkbbR5hR6OOIp6/quVjMxbqud8LlbpvnCL
TpdU4bYGFGgBDQ50Ja5Se3rcHyrqMpGQFqdzUvP0znBPTWrwARrYvWzVG97APXz7
i5iXKTBV1Rdnh6ZSXP7BHywb+4tp4kdYmXs6Gj0AOfR9alefFHIG8eTv/BHMhC4X
D37Uudyu0NEy7m0plAGxLXgYALkcVIcvYtuu6YcIRpvv2p/3fN6+s8rABrspYEzv
lToiDGH97tMLkKHARXdDThU+dq8Ejt03gPqLTYkHH2x9EjskkvMyVxu94TVB4Kk6
Gs31dY/olnok5nz1jvvs0CwpD+msrkdkj2kd9w5Z00HvOyTy/BNoQEEpO1hk4Nf0
KMNTeCQT4boQrjrDyyS3rMDgTBqZtW4JPTFe6P9JP3PVX6k/Pw6xbbbcn+mPGKPN
QdiwTmD3ioXN2VtZyLiVT0v8NHQCMTtfD9soB+Jl79WH/D89EWDMKUE6OfynMwAb
XfGdyG1SKTc4szutLaZsOlnB1xyZu3Sc1YSabWuKbBtAVKTj13rthgvlqpTbkR6o
fZpDzYCbTgbsJR5nS/XizSZThp+cAWr4c21NYH8Y1YBsQBxfTpyOfnwXTbYGFhY4
zGwZ8RmNruYC1VL2v7WfUDyx6Ax+DPXyAbUMR7OXVPDQoktc31NcGUMe6aFKNhAq
sNWX8IfH8noEHxke2G3L/U3dqXa1tFczBkHFSqW/7lcQZtEeNf0t+O7Hm6WfVYDL
gIkWk1y6tZhvOFuMQYZ23KZk9AK1uEUT4ghUEKbVqVPPXTE2UHx4xENppPwhVcn9
foznqUrq45MEi9uDacFvOFDaVgJ/L0/YNrgypIeIGSSvBVUB3yeEMCr6xwbmlXqD
LimphSrSbOUA+6i3lXeEYRFUa2qOTZ+YHSys30sO85yCLKCUDH5evGK4eAvAve0N
RwCVKBM2FBw4pMLHKE/lKG8Nx1BOn1yEDIaRYNLbI8XspM0YaznzCY6iz0iUHngL
4pP4WglMONu9+xDqhTd/RvhAHLO2nIOs1I1zibGijIed4BUXKYL4u039XTDzh1AB
A90oRqEIoeHW637jxSzrTof3dr9IsjKat8HX6wVfWm40DpfrwQ4+PMbz5drsuLh4
PEVxf3JTKcWRTxW4lbRAM8HADrK73v212Jrl8txMxbkoTNwTOMcxbm9als2RDmh8
DbS9pnwZDGX3iVVXRk1Qajerh9uYgxgOqhP6wjCuu+/fqTBC36Aiu085Rfb+bqmB
XIQ+JPPJGQ92DpBhGmJ7Bq2ogKtCq8DMHSypW9950N0UWfXNDKZuGjiREy0UkMsg
kzSWrNvyHwj4xaxvk1hsrcM3ewmcZhJRkQ8+Qc5MoQvsvXCQcKK/YKov4TsMzY+e
Fedlxyj28PaN7wM2HJJMNa/d/fHYl6bPJvJU6p7/iQqDmzeqlmlX1ByxqI9fAv7w
NClXFenrtQTF2L9C+FN0ukrJYDB9zcPggSxwXtZPLMgcS1alT/uNumPVxpkFgQ2G
NLr22PHucY76X3dJM1fv5b9IqNXBcV8MuSyYJdoe/TicC0jiATDVTkEWAx/inze0
MHA6Wr2ybDV3qNHMiGu4akVpiW05s/re/7fz/ZFCIotxC6HWDh1cr4gOd2XysyQz
MTDtMzbMxhIoIdmWX3UL8VKBt2w1x+osffw049PPvNINxnsoh1XXmJp8qMejaGss
bB6VqUaIztNsLXDP3z6JnzLMykAmNevh0z91RcFyzj06vd0aoLcGDMAEea/OZC9Z
R0SK6gsz3RyEu4oS80MINc4hl0hJ5G8ozu4xY+kfvpjkgCQNiXRUzAU6hEL8LBvM
B34oOhvqFBs2amKpp9L5S0up6sCq0lyqdcp+cXtAeb0TjeUGS389hbSolbfNO1jm
/1gDiIrNwtxtKkS7Rc+SKnO770i3cHgIVgTjDPVgRRs93JS8j4sJ3Hqilcn3g7G3
q1JpRKCQCKAb7Mvl2yPxAZfNxnzqSIuLkkaUvSKI0FSCvqGLRxIwOWsQcazMLaYk
GMfZH6OGuLWVxg7dlo7ugM+gpD+TxEIpCjvOAmv2czqJWXYnQ/MNvk8FUaqfT0dt
W4AOSNnrXdyvb72yxTQhWNDpWv6sgBGMUbbFN3eSw24hkWx/0ly01vlG6yggPEEE
zjmQs1+A3IG5HRKAAzp8kEyTG1qAmcdF6zPxWk3aMSWtnSF7oYh04OEjzkDCxhCt
xgC+M453+VplmucuOZr/nM9ukoIuzdO3OusO1JYK9DdmM4UfqJv5Xn6yUAf6aW5+
GfKHuavHWHTnF8p/OemEqwR+tyWA0KmzmCe5ydryktjJ3j3vNwmTDpjYxOwyENzZ
atFjl3SP3IH6E/WoFCtdTjlRajum6+WojfUQ8GNlvd5ctJgyMxYyBD6QDZUms8QO
jFsEx04ZEU2GPJjQzNBbzVGJlpCFXLsHSrYqWPIqGFd3opXGRmDIII6C9+sr9boz
fr+2ds8YziS3ayB27TAuYB5WkSyj/8lqdCrM0fj6YmkZdfihynhMZFlmAn14YDoz
oGbjOec7FHdNeSAQxaRYxQ/TZrijLlRsyebl7fKZN3xMbCsYW4yguB7NbnOPOP6T
iErNz7jmOuCmnhQ4vV0XmOTx/8gbHPGMtPq6IAxvTtTrtWsnPHkkblJbtzwHA5OY
90VGmY2zWtE/6HKd0U2yq1pGbdtUmuKd1nmdQGau6n09kxirbXH+3Gp60PvrJQxj
mj8bel86KHiGyzI4BQqbYnEhvd2NO2PTofS5Z/bHuXUasNeEnA9yMcbp5ZkcCs0d
HXCM9W4RTl1eZg+ySB8sUE7qbezk2k//raVfNXdWll/LXx2oAx2FWUNtGpuOfuch
tt6L9ot30G1K7dzvOjI/wvc75WZQq0ngtvdv60lDjkJvxybmDQe2MZ4eX5dTZ+YG
BLU9lOPMFqU2zy1IDpyge4ORx1r0BGcoXd45Sqgsd/2SBTt0C8LkdcsDUo2DA4Ty
JECC3FrepShXazmp3SPNF8vd122cZuwuY0XVL2cpEtkPBw7FPp8MtLnO1FUH6P2W
pfLbpoHqhCxEe/zuqRX0kRKS4vIPB/mg719S0Wf5CvEGhSlyDsBBdLHkKgCwQiJj
qr3Z6CgXm6mNW7cl3MuWWrvtzSHdV5WQHbRX4J7HfaQS8gQe/Ywbog8HTeHNF1r2
kZAfuSGdDQcVb9HUAxtiDztemiRQSxtzqWOZc7K50ATfnDsA/thAHjl3XEBNjDKA
e2c0z9eTKH2l5xRrT/rfOBxn1y6W37HYno656WqyI7Y9DyJDDopZcIT+00FgkOs6
mTI4lIo8GgyJccJqNfkGKOQfTXh2bUmdJCJt1aNW+6ka2srT0urGUryu5xqcD3Qp
X+gGsr9HZzR2YdBGZ+VI4Lf0rqG0sT5J7+sU/G1uabFToV9dxeAdd1jQMZHyAWVO
xiLv++7XnKTKROhSTNnx01Yr19R53o/ZeH5/+m+3CWVX4Y2VVLoYvpYa6xIY55qX
Z3gv9zZz5B9fSWJu+JAuF8wGsTs+1N1+7QvZ4Y1wRPKanAYtEws95WMmY3LCl0qU
t7+Hmja5d8FxatiKLkY/xgNfu4g8+i1UCCpEPY1bS7+m0Ns4OcCOY+2XaCt6VZeB
thzJKinqdXhgjviZp8ISnAmSPoBUZup3zF9ptha3E5y/bPZmCqW9RJzaVyZhwnnG
gzP2PHzgpWakOPQmA9H09AzNLWxUe9Qtr3pXoV5e/j3gFSr6tC6CrP/wjuwR67h+
xBHIU9Q1zTrTETB1yZjxEEJ7BxiglnqMVggjLC6xhwSIrU9KM4i4sBXrsQu/0mVN
5LYGcKR5uEUpODQ+aa+fL/JEhgNsQ4stWN5pNLIr1G0dIosQ76v+ja8NREHmGw3y
vyxpEBdxTaKyn/Es7F3bX6sY2fW5xuV1KQeSEe/HAHJEAK5ETBnz3w29lf/WLF++
B6lSFPF9WJLKsouazLbQ9zfyDyvrmcR5Ji5lqqhV0KoPlklvcnDB8N69/ArYfB09
ZwBgz4opi9ClynbwgrrGyDX8sZMMFOq4iS4dsoU1EKQpp7dWxX20CbotFSrMsBH/
8/PCryOyeTk8nvxBs/0DWAwFgqWKMNwi+1aUnWxUA8hF0+Z9wUbnjgeiwHF10X1K
3O0edXrzbsZnIqHRyCKrKg8mFnu/d5CucVwqq5GWp/PGrXfhkdOtUIaTHesrwYrn
7QeSSvpEeDT+XQkwS8zPMCQAjWPWY1gWqpTWaODNev4zXeTz98eeMG0NhiZv5/TC
XNw7RHx6tReywLRtVWpeGuniNy2TH+Y6skPCJ18JwAWGEpBVfJfTkj0lLjEp1r+V
Y+wIc8dCEjYjozOPUM9eRTHZ1Lhgu0GlRIFwcOqsEp7S9bD/OGquvKBPyceyaQ2n
HFICw0X5il62QaiDTtAQikS3Hq08LG8i60RT41PxgbrIoHWFggjdaWS60GE6cPhZ
sq/+KQouOhvOqk866mopzApFdwku9OjYGbX9EnKdNrdn+Y/eT7z0/ZxwxsnUfqKU
NEyEMVbLI/MWs2wcaSpIamIhMJ0SmLhrkQkq/sdXVFHtVfrdDfMO/lWmD6jiZGZH
AtAzgvyhkBknaWGt9tlX7mZcQUNuQghwbIvSNTLXBvOZPwI1gGlsLpTe9RislCmQ
oQwvllqK7aKCUBqZRRQJJqBVJiGI5J/KO4aEWQd2UOVDrU4aZ3LspK50UfM7Fkae
+iYNHOXXr8U2bDaetsAU9rOlU7P5daZ8zUf07BLV+ptIiR+034FlPD7VjFD26VD+
PQ1O33zAFKmEvVVl5+kRDwmprNQMmLCEfubt3xh/IoE+qTt3GR5axlDB3xn0e2xR
j5whQKzYVRqEXkWPPYOcGHXC/aEsQZGgnv1JrmvOoB/qxA9SlEFisHlURtt9Nn8F
biw74M3AdSiFBHEMD4eqoYnyMEebaNTMgzm94Eyp0/2kZ+SedCXuPACBsOzWuyAH
XcT1gWC4dMxMY+O+duWre5Kf+7By2iAgsnOrBXpqf7ymhNACxl+RMnLTx2rewsxB
Ut96g05A4LsR+moj1wpmtCCCrl20t/rFB6bu2a7d+JDu1wb4rU8u1D6FSTG66XN/
/+kcj5yT7YHKS2BPt0Armc1nb1a2IpaBijHvWyybXOiz6kDaEZgm0Ijp+ByGEP8y
XJ5DB3qqA7DzOLNkNSLTZSdyDChf3PcyhALQUlNcwGiJgZ8IefUlXy1//yg/H8kQ
13x1Aa5c4t9xltf17JJSggwo75Qnah0cPmNcuqflviZlz3F8BUYMC+Mf2uq0pU/k
aTKXrDFIHjwmHT8BvPST5EYa938Tfr9JegxY8oHpCx1Gizuu3ruhL9c8UR2oaQu+
5Pu1p4P9KayIpKDLRcOa3jheqP+qFIt9Zvx7dkr6AvUpYCCtdqVgupbh/1riAhWv
xIWhSvYUW/5sZxycXyEjzPbPt0mJsDS1TyHsdrhM98K8iVwwWduzVU4IOr83eStv
9D6M2TZ9/KrOUd9Gl6Su9v5YqHcQsEEvcPEZvuPPIL1xurLQpqAH9iggjAfEN4eE
QwVMv2D/3tem6bignjalrqy0E4qwAERBZpX9rfeWNpGdmfcGTHV5VrAiTwlgnEQJ
yGelgsZzfXtUqmAlT/D7UYDzzyTVPyjN2dUFhbg9pIQutbyhokfNaL2FFZ2gKhql
PfDEiuCHekEA9IJbnfKvoG8lBJYumTEUdKIM5Dy1moXChRvj/q30Vw3v7Dr6/fVI
adPO2J2WhNCvdUd+wQuD03xPzkjSyVkBRedwKVd+2gac9a/oC5QyCUzgwqsy5rsL
OZ9Xd0vIpXAmaYFzFGTVYC9RDVi22AkaipDzAQIR//iOgs0Au+V1iTYY1j2/zMGI
0bEov2k2Dz8AvBF1hZW39RRD5nZoDUNFLe4+6V0AVNKVDuJROPm1VCszCusK53z/
QlZbqMi+7fm+Ms8CSNiWEgX1mnm0NLt0eC+DyoIDDk9Ducf6XdZ1KU1DHkGZw66j
NTLfSjxHwjhs+9ePrBLGIWsH/BENxNwev+QdzocPjJfarav6npMaRI8zRxA4m41d
0/2ghvuyUzyfLcufZUlbKVYpcvwhozzCwoM0FLXPeOpzZE1NKef6DnAz9D8JsZmv
7iiZycF2CK10Em/X3wTKm2MjibiHy0YTJ5JjQUlvAgkFaSjx98vBLkJIOj2C/P/V
S3ynpVIPz77BzM+GWJkZZOvLC/4ta4n20GUYSZ7SZNMNfZnv0QrOafTYDTgay9OV
RmKGCThUZyCWzBJFb3mWVYrIiwSIzCSiHz5OJstgk+k7xV3uhxv7x7BO0LVMQnqy
XNWNwyQZ6CIXVFEIWI3eFTYtE75qhjgWFli1ZsgFGq8g7WZMt3dtkzo9JizZwiE4
ZmDV5zndayhVz+lVaN4VUup1t1e6EWRZFhHLP3u/93sE6DgpdfPzxZoFfoJh8TqJ
XsRFjAIVy8JP0DIkzd6zzSyxl3u9CMg+KCXfSSysaOiXUyaJp0pAOeUD0rAk/aoY
UC/EJPXX0HVka0HIrzKiIpnOid2WIC+F4gVxz2KywEUmABE5HkVUu8mgoU3QuUDS
VabElu5qb8LXIhno1Gnv9LJM7b8RZ1bEEjyTalcwNDn1FEvNsZsVY7TIMHi2/41Q
jcCLDggN7O19oHPSfHpCfcmHGzj6WZM5cG7xTtgjWJQfOIDYIO5Ak+rJ3fSpMP3q
KFDQquGI88UoGwNZOnjbTP+pwkNbYtQtj9Jeo6UlmOBsblPAAzsNw5Hb/Ae1Boog
Samd3b2yVOIxwj0oZVbnXq0c/G0Vr+sphiAZIFOvT2uHi7uD3o9ewQvbO/Q90gzF
KTsUJWDxlAlkBABs/pb/7xXb+XwHNB7EjO9eJVpujAq/colRHGgqYLRwc+q4Me8e
ko1Zw7jRToJp4qRhkkZ/rZGxTgtL9rpySK5kyZc8wMFLSA94YhRw46OLtKXqdvpd
KM47uZb8Tv8tOS/wJejvOJOgpon2LDlbD5DZM19HZRo+36rQO0lh3hgM4MdQNr4b
u0VMoE6k/MuUFHNh7j6UL/nMKKAlTScy5vAcPu5x4lZA0ji6CDy7eadayQJgR40v
6lgB09irHpnotizzpbm5zlJesOqDx5NXSGV0FzELYR/vIBcKAEpguBExdnXjvmJ5
OTzvYkvvGgKAjizX9AwpODNjTJxs1Nr45CE/GAvcNJhly6qPyY4M7kVDbs8R0IPD
hb4McD/Xyf3e2m9HBP2ifAVIOo3f53MTL49omIhl4mjMFovY2to2QXqSfWBpWIgB
RLBj8P0CXKFLQOnOcr5tKlyr0kr0g0LOvJVWZF8QFbNND1c2/9++0EWHeU9MlBEz
jhiaRR0v3gpYhA/hqRuAQfvEffSZoyn8Vm6QvpU0qW8rhmpXqJ007WtL4VWPLu/i
vO0OHc2OrIWiSVgjQ0VWY5h0SjT1e8jSFNdNfWz3IS5BQjklQoIA24MEDLRD8pco
OxxNHSAO5CDVG4pUrG0WLHgJqi8w0zG6JHO/zIE/aoaI9qJqB2APd6HprMWw2gJ1
wltnjA2FBzJrv30ubWUBwwTyJxKMysSjHpBECTk8ZtLW8/qbiU2xtsVIIElr8wLX
KHyFS7Nj+OIG29isc0R4Q7Nm2Wo4V28DL9rzPsXB0bedT8VcIFm3S2lPeqEK1oAh
tnsYeKZ7/nhAYrMbH6sq8Oj/7yqitjpHKLjrzWkifXwwCb5wpWeB8GXA25eddOC6
4vus10/NXkKksc7qF/nHUvn9N9V6IGq7xPjpxcixNKwOjY8SdfPx5y1diAqzwGAf
S3KAbMrrKZKrYA+VG0GqjM6YFHhLiJXD+E5tVYNRkQUSKkWvg6gJI6DKF/EPf6Zo
iYetQ86YPsqEJcKUoFovq2QaMP/SYk4IaNE4eg4ZCAMuGLFSXtl/0Em+6sMSUYEB
Is/KxCwFKQHsnS9O7DWLIa67rs0tV02K7OU5xoou1jUbVnN07sHCtY5VKtRbXGvD
RfSDddJSZeMHV9d28hpqAGgnVAXU/kpvxsNPav3pyUbpwJKBCBpQO/Z4rEqp27EM
R4SzAWFoisNH48FdzEl4Yb+v9A7gA5w/oENfIiU03aiuHpX74qcZbsD9cWzgimWb
9WT1XUUcfI35romtM7L/aoJpO0vSm3nIF3PIo2tuhh4uWcVtizxMSCGfoP8FAM8y
qCRjSXwECoJR5gWkkLZplCTIAJsYREA8sRaStWWGS2F0W1q00gg8QisLa7JX6qeV
NWsn/Wdk+aXNVAQike6LDFNMkiPnBtD58e/Gt90DA4sT9o7BHIBqATHZLu3FwCAf
r27qJrj9vo3lHcsetLK4RLpyLcds1jb79CTTmivqwy9MiK0MXeiBpL8LOv7Z0+6Q
ZdJEKBz5s6jovcDdYJ8vlMdLuxJjm5L3Uge78Ya/xQ271DlIceN4uYY8oIrInzAB
g1MuCpuIy3qrVATOyzUH8CqNyFd6ltSy47koikJ6oMtAQV5pgBiRTH13UWaDap/e
vG420ixDZi34mICjfFiYOfXFofKnu8SwdtNC1zISldujv4tl2qirpnrLMug67afM
RyQFMu8uJIskwkLXshmMGrve0PBGSZ4aX/5gWiAuL++BNp3eEG2unAzneB2URVvc
bN25viExlOkImzMHcYw3+/jZvZOOxqENx+yIqegHYhXAiiY25x/WasPTMyq0LhuV
Mwh7D25jjcmfxspNNyuk2Cbd8Brtr/QX9LI9D7mif6Wrdz1PA3V37YwsKGe1Un7Q
X9xg+Q/n7PRcLq1zrQiyOBENv5WGK1KpfH54MB6Khw+iMRljfHQQrcgj+zLosVVp
pn4pQbk2AB2Q5QhnY/+XCjCvuRZNVdAeWa1TOQ48ofoQq17FBSbFTZCZHrhj8UqG
4fHOHYBRkDO4U/qoPqzTfA2xVVvYlsF6ba1cbXpBVhueeIB8lXkhjTe/LeqXWlZV
JaRjBjg15qhuR8uAKAS5trNb0W/7gkhIHWbnxztkFwWhVZTltz32vap88njskOr7
wJo6hTQXdHZvi/FPmEUTA8/U6pTw5xDwkoakVajdNZUm41c5RXrqqdUpnatu+ncv
s9uomoOVuXP49NtCNt8MvBFl+srCkIclzltbWFyFRyCiOJSZuf5RKkAJfmf8RzCD
LXxM0YrvYnzWGtuST9XfkONwcjmcbtr7MHkriFRoJWEhu23OjPay8ch35loGpd8P
AbxKti+kelQ7pxkss8CO/KE2U85v79NUoj/8xxottrj5BmNLdv9Qvp5BQIGY6Yhx
s94kNaVkCA7GVoS/oDYAGpvKUpkSUd2NpSEP1spVuNPqJF76Or0+STI9kc0GAvS3
/+QS/AtcNjAgRLObP8CCAkiSJaa8UGHDxjxwPVvG/LMyWOyAFHGXXSmSjpohawin
tw82qVr82FmdrVXs+X5CeKoryi2wVNZ/6ewOXw4NvjI39MLuRk8j4Z77YaVoacNI
eWAx6TVzc1dWqTithuNbn/JOK6gmXit0pZMXZq0m6diFSqmpKTyV2S6Ok/H9TH29
tl1ObaMx2msH9AkPre/5REnXTjPlh33HLR+R7q+fO58AzIwVjyDMXvQobRHxTFt2
O1tQ9DsOcF1V3dlXEwtpO4St+7olOarPXHvmhmbsQRkB0uVgwBhA+2Q1iyBXQItj
17N+JnPxiam2EuOFyGis3lZc3jaSd7ucjeZ2A4IAhjPwXcxmcr6sJajgnTrwsb9u
VCH9oKXz0P9CIC0+fnPS3h+2B5rdsPSo/A1K+9Fv1vKdGmkZSfkTSA0iQoaJlDWm
ZiLUa1R7J2ttuKyoaIkM4eMDLl1fT7JPD7tCAl3oW0mvno3JVMY0tGoTAr4iVQsr
Cs9XmN7NSv95Y57RI4EfZelJcpNpW0EdADZmZCbOPNE0TxZ6QLtE3LuYe8i4OHu1
mPtNSGV98YleFYR53z/pLNyu4r0hSNAJLF7Qcq6xK4vdgkgKGA6z6+etswvRdjGk
oK1JgtsK1Ati1iJGwr16dFzLWutRSRZ1eOmbG+NY75dn0g9UQlE+HZ84VwmPk1vO
COETmAMt9ae3iQwyGqRIDai4nS2d2YR2ASZpddXyfeuMN8OkD1rFEP3wAKcm7aO7
EG6jPPX6L5de0SW4BB45viZVyk8f9kaIXQ80AbXKR+7BUhjXVwNoDXNtiSjBe4nq
Gr02BMKmMr1at04W2b766F8mSreE7ZydUYEoOuSWIHMvZGIJJDGL8ZHFQgyN/aHY
x3ITmH43AhCVXFYCVXtsfwB1PaI5ZjV2zDN5bmulZIF4qx+1Ih5aL77nAK7Ywog+
rBlMBkAMvfkw9bZFpDVIJ24139JDdbgalAdAZuZe1Eu3Zf+N2RXC0CI5P9Z4maut
cz4M+egOCbCOVu04SnvbKXj5cRBR2ZM4d2jzxD2NZDtlQ1f+E0jMXNX3PHZtFSEm
6yThwu2ljb2SsrbOlm19uq5TM47o2E+zc9N9Tm1V/u92YHVNVFPAe6zfFt/iGpsa
QkEA74UYdX4ZpPCU16Rmgoee9WoLwhwliMpGtd1BvpotECEkuf4rDQCM20LoLIww
trOIDnK1c84CPl3m6UkZcAVnEuku7k6/JY2kj5MozppWn8m75d0MJSAO0vtag1wN
/4iKdtOEXrI/8p039NQ4YlPVLjS9jDvkb2cdEDCVxOcQ6aa9ZvDeGE/Vvk3vaEGI
kqWDXs6EDvTD5zTesbCPOOKlLslpmRZAVnkpVzckENiphItEkyVqhuVB+4w/gMaE
+DdecPo3jDZwEru7JgUns68B+P+TmlOxQjDFrZIwVHqP0hEOfsQ8vVSWGrKl04AW
eIO4XQ+YgCXYocTYgEGOu6X891+ap+xXrqHmP3D9gTk2AWuoL46XhTmhMcL6YD92
ikoryQ+0gJUnq5AEZT6QDk1L9onYN0I7PMrAqKDNXi6zwnBLYuUMpojScf2sW5hR
a4DqYdYdWTHK3OBWNG2ZAr7dxC1meOT5xOFRwbQGXfEvVGwuJ5QlYrj78TeYCT7U
efmWfQ+8V//QVhEyJL+KebBrVli49cy65cIOT0qHdtNEghzuI1H2w3+Ln+KrF8Cy
/wn41+k+13iro7TiU6v1Q2W5rK/zkYTarTxMpKZIGyzWtej9rx0My7fqib0pXTw0
qtyHJtGlCbwQJ+uswF9aewn5oXm5R5/BZg6W9H5C83Do2TdZJJBST6JGJ46A0P62
st1Z+I81bhIdFpoHYAIlCz1yR37Slq0VJYDKLzPTO/7zYsp1dN8EmYHxk8XqnHHw
+jVtlCZ0Gs3wRwtH54mBIByoA2j+v9VpC1wSwjdYAD0jGy0pdDGN2Rbw1/fa4+Mj
yyRMSj0SObWDMY3LGr37A02+xwjyOL8lTcpJ+OcjDYiyBrcNNJoAA9kIHNujXAC5
iCpM8aw1nVWcb+hudSXoNYBd8XjIAirlQBw9iZTHtTMhXFmbfaO13czoWZeE/r9u
4bDe6PMsIpIsMsLKUseAe88g2ze/jR9lDOSF4XV5rAlRp67yX6w88fUgJw9t3X7s
5vwy31lPUvGJFMoNlMaSlB0joTV0dDBDcYWqQGr48WtgzjFpEDqlvcPrBxm0PLoq
cjVXjhL+DkIwq1gVm2a6shDSsc7bXmYtczFPRBsphz88KajIv2oegE2W6mGoaPlt
oTo/hyRmH+r0TFGDZI1jcrcwElwOQgGVAIym/mxBqc3Q0W5G4NBLbW+EdJy4B6lK
IihyYOBh5yKyAZnSMr763LbJ7ClNondSEVhMh+Q0/i7m9S3uy65mI6OOLIfL6iw/
R8zqwNtmqsTwpCtDNpaart4bozcDsFRPoyQR7D25qprRhxJfjly8hatFr8C1Wkkn
/UyMqZYpyav335hpEg16rz+nNbZRjceV3xuedJph6BwKge+rLdqAU0VDxsCjU2V+
S3sirSuXpT9BNf7YTOlfRla4tmwimK6ueviZ6I1ssN5Ompxl+UODqWjOl1j2XNL/
Sod6AEWO6n+OLymqjW3T+EuoV0TMofk4kOdjwfvm6zt+AY3RdqgIR1AKj846+ArE
ath7n0haMhj/gOnlY0my4HNecl/eO8CyeydR/8PJrqXzDInkuDg5JqvJQyNgd9fN
c6YutYQPtVP6TEtj0cordK7h/4k2HTHd6+DQgz6skOKH9DX0xdisNjWj7Z/iDypG
w5rRkg0hdDsx5F1sdDdboQBvT9XascdGt3IfiNgH0wwoQnZ+Lf0E8CzY420XDXAD
eHp80SzN4OMbsdWQMfUHj/AfID1fSlKwnqQUFEoJiJKp8uwn5TXH+NbKOai8nrlR
8PLJwUQLpKpTPFCG2kQVl5wXhcwsr2RvR5fKF60z98MBqapch0fFAOfX/584ms5i
Zt9wBkVturFDSIq/Ytw6S15LlZ6/1R5JfTqr8noCKgQRoLQFhfU6D+x7zuRsmx+8
fk9TPsdQBelxCEZFsoR8iq7QZzSaShz/rmihkxv700RA4I5O6mqlk1v+dXQbpiQm
MfkNmaXFwWF++MBD+hkl8+QoFowmWblW6gJRSnaFyGpq2l/PDumYKBlw9bbj1u7b
8UNyb4BzDbhr6K7elco7+gTUiAO1nIs5BFEVg9dNrBtboFWVtEHnOH6zS6C1qBQ+
r3ApmMY2VgfiDwPXzp0NCkeIp/pWulsEnRIGMF1g45Ne0xIv+Z5x59PovmNpIO9p
riW5pC+OBSBcpxPaMvQzCGiVGXf+hRYMwCNYcOSxK56tXN/GCW0CzqbyCy8lfxpt
TzPbj1ac0fKduCNrGtQ8NY82uzunfhpBz715C1tbB0eLABY0Mx772kIYVThOUGJ3
Wam3nCgjE6OybpSZtXkiwMlhepW3Ruqwja1gofH1IorZ9vXH214gyboWilfZb5y0
KlEWWSG9JHY2cH7xIyegElKdE7a099lAcV3WE9GSbO1oX0MwCIig2QfE6tHw4Pk0
Rj27CLnhZnoEnm1e25YnFibkz9wr9kNK9n0FI0w7NBhf/d6yMoMZunhYHNGTJ2q1
ZFRx4xkamNXGq2oHujP8t/cza2T9flOzqICLvaWgpBIWBErIlFx7aC6x1LO0bu12
wdAmzVRkqujui8CQA6oIchhJ55MeZYFhcrFj8flpAmB8EEkLhTO3RsEznJ8Fza9p
AUVLFae6+aIgBem+RXiFToCLJdReghpCGFUJSPpyv1dadv3diX16x17acFdR4xm3
Bxm/gGKsYX+2J1C3g3lL5Wa0WNjGOkJlaoFZQl47Xzqt3spleiEiANMF3alOEupV
0IHBCjTpc1B8XpPUmREL7r2KtPhI+ISRUeI4PaB7r133fAEhTbxI5k6gMXB/8Mbv
GmG5/+gn5s1emfgbl/oVWPHBGAe9X5jWuWTktuFRYEuNqy+xh4n/C8SWGzUtDMTE
LPh2eoNyAghkGiARMPD5wBuaP28WbtH7shp4KYGZaz1bA8eFUsB3nhaDx0wKuntS
80Lvlq82hLMKXdz5mwyfCFGc5Ma7mnVpQCGfuz3AUbaWfgBR9gFPgcvRv+wpgCMr
W9q5UmIinirNJK2synszgUQzIQDhcHA0q4zDPjiP6yauaC7iYOc5oqv5UV+bqRb8
XWE7JQKemYsULjKr0MySzSgpPOGvy70RdnmkOYxItm0TmIjjRZjApWSZtw6cpNTw
z+ZHWlNhZr4TxLkqHfvEDO19OC/LnJHhIOTHFjIeEvAY3bQlIkU5l1OIP9fFdRD/
cmUvdtmQssXczXMnwXf56oGl+Vm88ywpWWEk6zicRNd+yDFnyn/VIfhvyFdl+pOW
Dxn8fq7Ha2SEKJkZ8J7/uXESO4CkB3pe0C2quTAKYBN9B9Uc+QLMfvKGNKMq/nKR
oCvDMVTCZpjcCnfeysJqP+FhlhAl3tYZ0zzzekOA0nDfh+WO7+yOjNx98/G705ek
v9b1hmUY5pIztJjIBWpfzITjtlX+Y8q+wCIkQevMGPtivaNcdqVUW499OScQnMg7
tVcEGQJAf01KlSi28lfFzsgpRHFC55mISUqNHYhs6l38vOIPz7h81U6/7t271E1t
Ilv7bmJvS6inh1YkIHB07DmkaC6yZ7x5nvAUox1BfIh9KOuU7a0aFHTqK7IRd70q
p4SUi1M0bOn4rcdrWh7Jg8siHRKSBsfqfj4W+5sSqgwcFMQuMYr1FXeaD7330Ivb
UsGP4smWN2Mf1dxxH+C7XREjBBZbLfkHmKb6EfX+9MEk30E/RXpNiMQe/a3O/Ms3
aC1FGbcUHMyYLIPgvaIzMMNyTYOwQPTV3lMw+WEsuF0f/PsYJHu4dWicajJzE740
bNWgBu4Oyk6OJu2/F8W4s1HJ8r1CvKlM1/wtbI9sycbqmIQyCqz3IAKyMPA+6tpU
SuxkW6027D3pcbH36Vo+Qi8XgENA0nTOmXqm/biEPEDLHhOtP+AIHyCm0Z7X++3m
Kkw5njc5fDVF+O/Mnel0Wtq8ysUvXZPkITXffuAWQ8ba/dNUNko6bgrHiDaFbe9r
DcVlsqk9LsPzoVh6CgmTJ9fNDTVvHCp30BlazdVj/+CuGdNdT2CSwsbDhXi1Pbba
XoA2EZr2cj5yVI3UA3LiV3J9FeugBhHCJ6N/IMgxp/0ozz8Va67S+cReznm9kDKU
QgrEBrm6immlQu1ZgjYaukoxChMxQz+WPJ+TgKwNKiTZ1WKNFWWc+d6h0Bp6W2V1
TKwQmMLDX0ovxlFgJ5zlIkWR2Qwvb9QAuR7XaXjstqlphiffdiWlHtDXND4AvvaQ
gzGW3vrOm0ID7cn5nsZe6/Quq7IJTKeK44CgO2KBixMHxYg+/bie2La5Yz2Dc5iH
5jGMw9QSEAhdfA4D5fjZXvKbrvgvNOuKBcL37zUV4fuj2IjhRTckCRXhwX0zSW8h
/2Vgj2MCTgYyDBDbYleI7D/aoe7iGHgpDZGC03T6Hy/qHBkwlAc/cGmpMjYBUMGM
6ekNl9+BvKenTUrqP22qO7vrimmtf84uw6txcYW1a1kDgG6IxRtffGwjKh+pM939
0KoaYFiWGCEn2JiJMpvY4LlGVQDRlL1h7nKz0jIe8ThTM7yhldsgLfbDZazimOoS
aznOwbpU+nz8HOKiSn1DsAruBT/b4I0lX/nMzGH93p7dbsjagMLI0BkUFmNnn5y6
Kb3xb/i40cC7LwH03SMlLxLlCYLHnw20PGjSeZHdt8mpWVdhRXTefd4R1sXJrwST
ERcuZm/S0m8zdQ6XCrVseURwwCJUaH6jVkFbYB8rGqJWfq+DmbGtfmEW+up4CU+Z
VC7i/9PkqiT/Jeccoyc4MZoH2ZtLJSObwKDJpvCTf9/pw7aAXgoOQhoDuL/My5nf
323Q7ShqLNNJsWOiLrkRTcVnW3MZHYmIRHUeiCCGCJXz96F8XM8kSWc5ovhVU03+
nGKlOI7cVG6LrQkLg6pLBVQLVjOAuZOsH1LebY80xSQooPjsZXAONJSYwbWLj5F7
tOM3Loa/beMGJcMArPzp1kDGaQi/FM4zvj6w+83mV0YKLO5MVeNG52YiR/ULxEhh
j0JWE9PdE9seBcA2WcViFBU76bd9IA7GdnUslQ+VKbh6DZRtzXjRfRFz4LZ07ZQk
8MBFzoR7U0QPQRhPM0xZgQJ6AIk8gX7CziMFqERj5HImH70RBbuZD9wCv+Aud9H2
RiGx7YvtJX+wATU+l5YLWy0Qhtp8pmSQvXFCvCKuMMPv0BCPP81hmHAZ7esOsvtz
WadY+b+Xe44Wy578gKtOSHRwft+rYobbjw+4X0+cJbpJIE+PvE2VvghYZeMX4zXm
+ySgch7RgF1h7r/Wh47ClPIycCrSKExTdWAkesc89qdi+YcZ4mzmd+2spN0SrlPV
WQ1BtR7PpYrgOF6OjXhSSOAUUutWiVNpQqTyFQje2UySIxNBRNY5JIT7h62kkV1n
dCM55huqBvCxzE0Jgx6UEOHF8WIos++21JpClrvTtx1mvUl4E7R1VYobMxqv2B9W
SUUI6LD/OUMVC6UIzR1vQJPkmlQCJOJt9W2tiPrIGd0s1SbfANuTrhCi9Mw85Oad
NEwEfGhUiXOepdCaLNMzDJvcplKkyQJhj2zyj63rPwsuslQu8HajXH/Z2n4wjeiH
IYVhH5iPDqiTazk4MaAqBajsbhZ+SYwXxEn7882gHg7Z9RA9gi+TIch+WiDdwECb
CyG1N5ugdjVRVL2sCgWZ1Wcdu69Lj20YxUcbg3Odw2ZCbAX+8jw3y7vjDSTWTR9K
FsO/m96wIWmT7Rmt+dMroeTZm8ya0PtCYZYkerYhLV4byez60xOTTPZDkxyUTpqc
yI3pwPDdpYgEjTXnz3pv9UYzl9RbBheUMx15e/UoNKAF/WG9+oImI9SolOK41s5W
n/JSN72kjwShrmG4IBMUJd2sHeSnjRdd+vZ7H1tyVBrVj4gqrHaV4NHmZDleey3c
e0EKsMwwojPYgE3jatIlxPBj2hDz0Hy9mm9P5m3KZEGas2Xlq7Gmopf08trSlfCQ
gO1ZK5XfZDGuFW9PxTTd2/lvKY4x8h+iR5pjp2wN809eHT4Kxszrgedw3+a8VzAV
O80Jim3S/RThukfHkisNZvIs/978ulAVG4vxP2MsXWikoxqKMtu709bwRztEkCOn
VqDr7ZamfviY0lgNmtWNGB+vJ8uwWiJ22REPxgN/qCkHMBZatVpIZW7DrLXnzMCD
WBj2cSJtBnbfd8JJcYA9vb8IOk0BKZNBcobqXeiUmTfUfiUazjSJzN9kyxp0E8s7
xI3t9Y5rtQaPgXDXYskMvOwP/BJWbjRq68gAR2Xf/33VEeOmABKZ822bnBVizuu1
CJMxmkXCFVpSto29y4olWcr+TJrG7j729FP29U5lrUSi56p3eYEYJFpg0lAdAYs4
gXuKhbS12mf9jtl3Q9nkpi+FgRUb+MvnrAl0o4qbfi5HVZlGhx2SCMGVfkV/vDII
I21SQfkE8oTsFZ4FN7RUpeihsMNwFmtnfE6N+tAUTNY6pc6HvgKEfTFoqOr8V3Fg
+k07/vEEfgTGBj9k2NfhAX7S9M5C2uQxcTNlEDUJJvTV8mIDasG7dbYq2SRXkqWk
2j7W586C8/ky4lMla/g5WkNL/X5ox/3e2UNhOKAoo5sIj/Xz0O+60Uv2wRcV9QU7
OZcvqLs26lmA/EWjO8J40w4nLIOutOmhms2Yckb8WKVYJMizVamyr8iRKjSMD3vu
2r7S8ipwPCUio3HPVGvEDgJu6wbF3UjFQ51TcFG8AXOkeP8E9jhYqHDekNnHnNRd
ZhBWElg1RFpv6KflWMjTUoAV4eL25OPGTRG6O7z7V62SRZ1rFbBN3owo8SzDbkvo
LpzPIhHwRWlhDy6ptifwsfifPTdx7tRCk3ItnclOKiHCmdf6mLcfEWvWmLzTBn5S
G1pX6nlYlBCNEX7KVLTLC2X8iomuBLDIivxNrP6e8piLAl8SZU1uCXxshqBTnDoN
ccDWBfjgvKatNPyebGHv8nGuFtyQc0jkQkzh5/p+mLSSjE/Pw0cYpe80miDAiQBz
O2zj7aJOp8qK5CfF8/rIOKgtWjvTqeVTrD7eQdwnSHkyI59ZqffBDrtjcbNEV9JN
OhhWB/LIdOZImu6FOfXCo7ncbAnmlda+k9hKsogJ4m4QU9OwWogo/iJ04EPOYV+9
VA44wiUaIHMg9aKOOYgm/xZJ0GTSwePIwErFz3pXaBXKh0hQJqkSzTvVGWsrNr2i
6WDi4a+nCprWRXkqwJ+NBZ9IhCu7Xz8EYyPB5Eu6rpGWJNGL5AJ6zMIR3+ZbMyzd
HCrs/seRsuPhX++ll1h2paLPQXAnw9eh/nathaeex9aOtKHKNQ5ULITk05yWSn5N
CvlgNY2jcjOGc6dh8aC5ASG0rjSScmlIqNBmSqPMMvx/bN31b/vwCJUwLhF8B7Mr
l6gJjKJBlK9stoCMov3WI4TcaPhc+nfjpe24fZYjVOyRoqrWeQVqfugFAInsr7tc
ylUeEmPC/1M+AQnAN4NL/AszCWJ+Mb1tZ8z90YlBNTOJS5ddiCu+9HG9Fciq7ktX
Wg+yXZqDugDEsJdSBw8FdCkQsiquTgc2q0FWN4qQgzBK+pOEHnQZu/jxwzZDOXUZ
kCWOEjZZ9cQpvxIy2up86yCs3Wm6bX6OxGZGXBKNxOn21u5Is4MC0g5p0OAB9ZwW
90AOI5heZn9spcGDI04OW86U/VmTdRD1wz7PoW6izJFJ2qXqiavh14vk7DxcBzyK
0MC7DLTTr8cPxUmrte2fJHX3DT4ZdGiZa71yd5gL+1+ftuM2nZrO6Fh5CJszuAIN
tLV1DJCNBmoqU0eAzjsL6rCiSsaSabnfBjz4gSTnO+FvjExeh1kMJihVsYvnqBjW
TRBIn6O05qnKpTUeiBVz3S8hO87p9nGb7i555722KuNymOav0Af9a/LWSnhNvT/m
Db2uACYPOqBz9/6vMY6HzVoUbeKVmenyyx3UDqJAKH3wioqaduGmGlaO4/5NACDP
r18FtjZA2TIZyM3uf3MJL9qgRy6sIakd+QclKC7T8u9fUefkxIdtAVxytTfSJ1Hh
u9yT1N5/Yw+M2kiDyvS8LcCIr5qkNKxdO2cl/Ni4b6iVxavtHB27UrnA93xkocZS
VJWXw4zCX6mGuVWhbfv07LGxDgGxfuP4N1ryiMV9pj7KVZSsyFJTwji8EaPugu+D
n49NqsrZcK3U9dzWw/IEpO4jpHgepotb8EO+r0J/GhlvpTOG44Pr97Ajx5mVQtVi
9gjYZrxtCTLyOVP66YQPSAjw7SJhvcqdRq55UAd6tRnSMmfNq/tFB1mZy5Btj8Fd
DboFrN0Sl1EkN/p8isEVqJgWDwz7c/RwLoPwZesv8P7Hrf6XkBsi+cE9PpGHn9MD
j++kxe463grXx3kZ2idX5AdfvMl7OiTFk64e4S3mhRIwq+6RwwpECU3lsw//BJ30
EZq2XtWW8Eu+yQhIoL0BEJ3ThlK33yY2prmWI7Ewv4UiVumKmCB7533FcbBAzQdR
ytrThkSGOgolKLXv6LTh6nzpixm4oHfzhNmN07KJb0lN4BFgbgBh0hd2v8sfpMPx
Wl/vlmCo2sCpHjPeZVfTS6eV8mvX4xozFycEy7UXd4oFfapgk40SCgvDf9scgZFl
k7NOLRHu6RjL2qDvdDkT4R0BX38F8pGndQl/H2J6Ikz744vl7zt7nBZcBpqsw1aQ
RqTaVHs1MuXBx8ONIB3q51Tp5pPhGIX9VOqYDRBxzp4Q6ssObxIUy01kcdWhaz+Z
ShGwAfRP4OM5dEOaXRMzToC7lwDDnnT3pLXtT8q/0wg+NpdMyd0xh8jIrx0Vn+ut
BjdWTuFa4gCHMywW5EfojxmBiZjZSUn8DGWSZZRACk9E0Y2xMFYlpavISlKsIxeN
RwldcLYVTdMzOqFv/gO+X/SXuJrsy3JFGWwnLZYLVDTROwZbhms92VkvW/zO8Gg/
cokj4LBm7UtRtCWUu004QHKvnpn+v9a2wbhHatC9LQBvsAeb6necnJUk1wMHnY4n
GK5Jt/NnJgt52aqukzi8zqYSPzJVhTcCK3rIfJDW32QV3TNg7TKRNd3DwOVHc6Yy
UFG0JPGodv2Oar5oHzyvtpqTCyf/z9hFINa49BWTUJFg2fJNvRuY8CsQi9At3Ewr
Jcn+Htl8szwckCrVHe8UYpvYzHd1i3CDekYrebXHwrOMqRhIf2u8ApGIUTWRqNgY
IHb66WCXT7Jf6q3YrXh0KCbZa0wYfK3+hv61gVh3H+QhqSryIgVgEhug8VnfOWpH
w+daqRdm+5++9EKkVVfwaEvElHKVMFsZKQG6zX9RdqLBhVtGuJNMT8I+fGbixgra
VDAgrSMI3oW/Pzbwmpb4QXvspmnD4P2Ux8XWvbj3FXfoUyD649XHqLcLGl/ZdwlN
flxj6cd2b6hMUCAzBv8FsW6RmyOfQTD5CjYHAXP0G27J3zYdUEIYxtToswoEKI3v
HCEiWiTjKk+V2sklRiCRdp1zD8iRwUiQ8B8D0pDBdbU7iTf5h/9rvAbeW2EeTRh+
g9Z4Kf3DmHE1HQPHC5Jg30m5boe80qgxx533njLJqRSHhSu7yYj54ezyhkKJw8Cx
WSs/H5KwfkkQ22sFE8MpfKzcGqSI2NTvcMU/SBERgHi9lykUNMNU+9uS8+98D9A9
IRIUM3JA14Io55mF9L/AbRvF07oue1RkdibbUTGBT7o5VRrYN5ZABc0X21EdO6Z9
qwEchPRj+3WrK79aU33X+LC1uFsBkfEF96DwJdiccSdc6pmbNDqQzjzMNXTnovuE
Xn6+Ey+Le4hACPUfzp33iaDQSwNBYBjDXi/NtCI0CwZ4oQS3rYl88GCLss/XA26k
iw3RkSi7VF2H7S96i4G47ZZeBDL3Sqdoy6ZCBadaHbgFMyQaaXOmijdxkSW1+d4f
5LpF6Z2Tl8pANs1Ne07d5Vq+036/HFDD1PeFrRMzT9kkPfHrpVzuUHsSwVNVBs2/
6wGza5D6rgRYB2mHM68lM9yxtxvxzRd6sHnqUpJNbIZS+BIsrcXJriBTX8AGiDGm
ntHJItPlMhx3tFKPs2jqyGwNyc+7/6jrO4BPU/vrMEKDeoFqYCs+xRlNp3SjzyT1
OEhxJL47M7vnyxKlYnTGnuR64U17sQ5+4qUWCahO+8jjQA23TUKy1gDxPV7oImc5
ndM1evUULvdDOZB2I69m/f0crra3/nmG+lGQPR9TUasd758M0m4BKC7t8nxYFXhl
XZAMAxuhQUMNfCGP4tFA91Og1pkZjxdnhCwWsPhuksEtpwKF54D0v+E1f0lQPxzK
kH6Si53itF/aX9wv4IDmSNpJejwhavrtZzrmiPzl4Y2IwEzsnHfqwlVNfEJXWGdw
XtuJSuUB7jGfHFtF5ZUzbXn7T3h73+Z8TJoEk9jwqzeSIY0eap92w5JNASE49R9G
Y7yGaS67wj/kPjYuZCgbAtJUVL2v0wBKR1bG0EKI6t0dpCooA6m6BvKVbrF9aXe3
x7llecGAuVZTa+RQEKJWmaX9q21vFD63dDZqHfvg9elL7tXP+q3xb2k/ufQUpZ9A
HtclQZ7p3fLGORX4UEkV/LjovwreKdcXNIICL75Hn/qMmhz9UAl2LeJUpmAoAx1Y
sClRitmAfCpN0/J7QmwDdVK8xB6rJMvK/QA4j/P+3h80TGXgEjdztGdsMmNUY1WS
+cnFhtDiXyi4BtKKmVb6dmyFw+xgUcOJ8eszi/hata2fACJxku2CyWkyBfucSuEW
5eEQL/JFciLgwwMqgsdZttfbntCDL/uL/vlDGyNGgZQln/y9qO/XXdYyq0rmTzZ5
6M5Cbd/DiIArYQQAeiJuC0KGFjcWpsOwfgJ/dcmbVkyOYuPaJbqYZNO6Y1ms+pYR
lvG1r8wzceGmmmf/LHnqODZZayT+p+XwWprabMdQp1tQtDJQWT/qkDpmYBx/D6ii
zSX5fRQEK/cXQgz/2o2LKF0VHb4f8Yq+jdlWQ0WJVvxxWGJp2owE09K+Y1Yd2mtF
DfLe+lq6wUBzcU6/2NZpR2/Jj9xedQrZfqkXf+Zx3orR98URVCISnkDfcD/uHxc/
oo+/GdgqowpzITXLjSzPqqWfqIjqi4FLKpIDI1UYklc1U+ute7T0E+FcBqRHWnLO
CdR1LSkk2a14CJKs+GTdjP85OmAk8dxl2h2hrdYaHbB7dFgMwip9y4gSe/KrPL4L
kg67pL16qdrVQLeReDKM0NExlf9UiFnbh+d6Uf/7X27EH77iYQEtcswzfrqNriU8
TqFx5jyPHKwUSswaZ/aUOjafi3Vb0iC4ObruqVXGhA4MFz9aNfIGbucXp4xKfSNX
W4fD9Wtf2+Pr73CCGjAMxb71Pj30ostS+onnTJzU+bcRnDe/Yw9g73kaEhPAudeP
x4tx68tQMiGwXAhLFj+slyDaBE51c+J76QPD27hhKhHtzlBIX1oiQuK70LicV8rU
phHnmFPMQz/sswgYd23UX1ns6h58ZTqVwooW9JfrJJaXW/8JsUnXJB7k+/UAMUv8
rt8pLZvSC8AtYyJh+XtTOzbDcbL5d2l50zqOfzb2/XoZPz33h1AhY1tpvAH5hL6b
ft/7H9OteCquR4syGNwfMqrpUBQlwe8P3UT16uCk9lHsJ8Yorjk7SK0u5jXOA0St
nrzPUungjPNhF7O3SFjTaqubQLes5FU3cm4A2eYhleCpvO9uQbh44eqjpBC0qb/f
183NxtSF8POS0UocihouSiQNYXJgZtIg9POrY2aD/yqSXGccmCfl7p/2cC+296yf
M12oJysvqc2HM+Kujo4IPCsp26inlSb8vpP/6cRxiEEGWtIyPOJoTLyla3vfaA6y
ce5KRcu1iLkf+/goijNoC9MlmZWgtzeqVY0JsDozoVUkgIjXzMfwgAJOT3mjacOK
7ooXOuf8JBPun8tgkfl5LmIr6CtstVe7PmR1jibeZBhRjNhptBYZQgd1n4Mk0W6G
gcBWWhRKy8y2sZbID/C42776i4jl3/btv9thBuPejn9tQcIqsB8aAYAXAXEbU/Bv
UwK6jdLWEkIR5y/kncmbxGleNs+TQn38SXjRP/LLoiuGtK7qJqM3/DTdzJch8kwO
YKFCW4UCyK0X8W0hsdy6M0pcHkklDvnpm8ZctqGl8fkmX+ZIe7J2Q5YEHU32Ofov
9Mzwry47PMDzpAEX7NkazCsoGTpy9jrlLKNBSZoiT9uVTupoy40SFilhXM5B5the
sc6tqdSeBexrYux8wrAowoVmFSuRbnrBuzGyj/1YzBYWpaFoLVu8JBhwEfMRjeZw
qSTgCiIAC8UyTq4evC7YychKSK0zO1OfM8BLHQDTBjmnFlEpCmgSam93t2M6UOIy
TvBKX2Pd4YwfeznKqK34IeDUPbpKd9TkthFBpFIF6C1ZuV/s/kL6s7DUsSDG1omk
1ZW49uV7mfIEHMzDSP7kE/ZtyMrx05vihWSJtCGFuzoD7kRFTjBJYnLOUJXO1RVU
0yXjYyqPNTK9ktUC0X0QlWto0sOTmdXVU67v+er+EUR2hte9FJEstf9cbvKGqA/9
giAZEC1U+sDOBSCDBoUN/1obfiw2CEe5OhaMOzEN2bO3FZLpFDdWJxJ/PjJ97BF6
Lv8noYK/MmaDicJY8zEUAWot4VlOYB1ZTSAZvd0XaK67oebTnM+hAMOIIJ2i8RQY
OQPxAcY2PJTCMye0AnK7B++6RBiH8WolIh3vmw2C+dZ7takOhUCGyC6I6I3P9c1s
lj0f+jE1etSleM6zLR7KCR+Ai6Bo8lfRowpiWTb2Rt0/lPi0LoJsmS+hFik4h8br
RTBB+q1teKYRHB6lCqkHowdlssMRobEpofx+uw8IzOqj1QZYPR1Dhw/SJELxOcT2
VLpekgBZcETFh4G2a8M+PYnbJn5TI88oF+eWyet487Ri2iAgxMrZJtLtCd3qD7Rr
ymTB0AKdDtSM6PkhFBpp843vlP0sCquWHlZSO6oh5qU6JY/OX/YFOHpwdt44MwIp
z7hhX8t/Vlt6k8KD5RojzY4AIWSeM8JZb8q0Hhof+Allzn9xahRhdv/PTxoagoM+
ciOg/vW3emD1dGJc2K8cimNG3Q40qCM93dTQ9XSsnv4NY0+ELgsiIS8w9cN/yR7e
W6Y7PfvOYoMNCdzlyDEiwZ4htZm8XMtcLO5tszFifZGFsTvQ20KtCYM+0Ssr3FnY
0m1uImNhVQCK19d2kppbav7o7Jhj3cDLsiWYvAHQjU3reDdVSa4Mqlrped0TFRNA
4WUHVEeMU8qtJWwcbWIjXMXTal3pUqBK6J0sb8T8M3DLFMoXskbkYaaV64DYJxN4
9KGQZIfELDKua19JMyxcyuz8cHjbhWRKDvfYRvfA9V+URhzy8gbaGEFTVRCqJaNr
kc0VVAOK/O7v90ezi9k+5+ObZjy2SLdq96T1Xavh95oo7HStaTbM9BPGpCxSfVTw
qFEb+3cjeBUs0HqtNtNZeSQpl8uFuSs6YGjlhn/DWPioKPOlbHIQASeYFf+STGao
FryDvPZ/MkgGIIAJ59YTu1NKFcdAEm9rIUz5eAQn+G27WZ9n30J4UwDkDoKI9r32
zhNQuGRFpkOVNs9eLn3A9IdiN8qK6Mtri9XvvKyNmp9Ud69XZCCYGF+wM64hY+lM
oW7dWHsdeQjuQhqEHzkTEoCt64QlibWn7i2Xts58X4Oa2Pf/M5rCZ6LH4Fh060lv
41on2iZNJEOIwpXWNaTBwgNetsdkMkzKANqcpZJPAOMkDJq9jwZW6W5kbk0lk/VX
w1RK8Bw/zL47RKV+jPT5k9YADns+980EbhXnJjICvHyHfq+LCC0Z/f9X8J/bKRPr
QP8g8E2cHR3griYcJ7nJ/mLFHd6vL66u5NjZ/KBkD2H+3Z9+GVFPHcHy8uKAVmPU
IvEvuLfEvJb3gdJx6uAscohSX9VaXNdTgfCltlDZeARfwvF/4fJAihB/gibPgTw4
atnNuE36Lv0d+8XJtSROUgnni9GN5mzJwXMdVFuTg37aPcCGUK686539OXifJyKE
kbTU+tAccJJ+v4ccDuVhfPA1oSudHatvpeUreze4Y2oPlDtgW9kb67VO8f6hxX8J
Mgf2GCUfrvZsBK6afahLB1Ll9KOPuE6cU3Z7UGy02CPwcdyC8ZwwTTuNtxK570Ws
2+2tjLOV7yPvTF1wbtw+UlHxzeLLKix9Qs4gP8TWo4VIR2Cyx1krTQ+jXPaV9zeS
risj7x42RBB1FpCtxoxXkkzy66gyqD4pZ2Fa10+KN2p1wv9ShTsYAAnu7H98EDpT
1tcCZfzauiSgH5pjwLkBlZt7y9eHLkdzrqSjba45DOjgB36hS4F8lPcIXjr3Aq9P
rtO68Q2GXiojllgSZkyE/aKj6coi/d2xxBV8xQoU3Lmnxj4iXb9Kqx85JlkSIi9O
C1gKXkI/whzx0sbJP6WduBqhOqnfW+hE+OQkrZAXI1OPAxYgKf1VjKVmM9ZDJFqn
d1OGQWdIyvuc79NHBSvaOCo5AQ1anXgBSlkXnS6jwch6rbNznlKSiyaSkzvyggk4
vysy/m8dGSHUBzz5yv5wjv51gOo/BR/3v+UM9G6u80yAiziVEuYLaWypp+6IGE7m
g4J979yStKbwT5dgyvGKUbKXyzz7FHFKCvhntwstyVRqgF6tPN+H2Yx6jIj6ilVm
2/lnXU27h2O5aXgcTO3o8emrQRnt6Jkc+23O1ppZQgG9nCW0kjTfYuW5+B/rGdVD
mV4Z0u6DhySU1KyrZy92LmI57zhekhXka7GfWV8MdMCORGbGZ+3SwlNKbSProXC+
8NoutSSMCwmeSJkrKxIo/la9Oncn/89Yk9VQHd4Ui7RTKozUcIpMB4y69drVct8S
QpXozLB/G7QcYlBNf6K3tmdT0qpDoC7sVho7jNZZ1VAYLpAkui7SJwb9WII+haXz
S+5iMMUGO6kG7LB391LX/0tsATPtmLtLVZg6NOLhGkG5KbIn3hVLYkxVw/ui41eZ
8lWXW6xAZAhXDjCVt7T0qo/RFfPu7R3IcJ7iGelU+eREgoNQcO7TMi3wpNj4ppSM
JDhh6I9/qu244HQcWHePJa1hC7qRI87NVv5hsNX6gKb2Wm01wASb0WV3s6ZAu/QR
63+rD8rf3Bn4x3/qg4MSRGvPuGSZ03NpS9oazSZL59yfS6TQe/jggFumdEfkRZ//
pvwhcYxCt2n2PRgUAkZABSqiXD/DIpw29vpbsbwfNgwhXQKFQouQWpQ9qSmnVCcg
E8/5hTRnAURemYbuEYn/7en23YZSneD+yKVoOnHzGDIOw7ttsg6ymedmSDGCiQXW
3K9RGxircLD7fDq0/M//JU6AzKCZl3aJjvj7CnlCNAj+B2RL9NwcJw/ttQXfvAJH
EgD+67nLg7TqxnSO+K0Qg7gDPoAXvBQyqnFYxKqkjsfGTaRhCq89QS6SBSDYU8u1
YqQUb0YHnCQN+jqFGL1BnLZE+KB8DqA5vvo/OzeMc/JXjlkwwE1XIIZ1RVgArUEN
ZZKgIY46ajSBEHDqsgZ1GIHrLgt3vJHb9prSUrDj6UnGzGvJ21LzryhdY6oKqabm
mHyzB/zxJlZVKoGPHRB+JEPt+4z8xInu8OcmqPPSkWADxAlbTM6pUPEbez6/wltj
q3CaCTL7fvGlCm1lxwqwm49zzf3Vm60/yYqA1B1zUTvarpxGJVh6zBg3aomRjfcn
8qANT3gPMnqBbrXQeluDdY3wI3q/xbUT31l0Dd3I51rDD7ZM3IPIvG9pwbtrEREy
WJNdIoS96zRcnOhoXUi5Okks+mYA55QYAhvKkb1YW6PnScwyCMi1S/9lGQ3bq2uZ
rQq14w9aac39cgHnCYT2y8IkhwOquLEhrBNdb8avvmnlk2uuA3QhegqUc9O4gzka
VxaPz38fDq3aD6jvwrqlzfj3DgRqO7h2PzxhtUyQ7/pg4lsHZjmObGd2VK86d3r3
Zo1nsHDzR+0/Vd7ImUQAoYyOUoYDBai+j6d7nN/olH4NN5dx+ufml9ky1lDdPU58
UcWclC9d1eEncCcD7o/0ZCiDo2DhheX0RvvDW4D1EkBMYYj3lSfZRh065sEp+0GU
UjQggWD/03OhHXAkoVYi2cdsBJLfGnLSLD9Pdy1MCkNbTeJfRVyyYGJMtW6Sy7V3
LUw5oIVr934RB8hBBMO5wNHmbnRTcTCvpKYQ+WXiSeJ/iUu3+PBVjDz073aCas+1
UT9Zd6tXW8eQzEpTsc3/KtM7kjt0XOxXI/ghSA36tZ6sh+N/MPbzDKjkLeDcB6nA
vI82FRhGtj655mvPgUkuw7wy/qp/2sGEmS/UT/ju1uMpDQetq9t8blj5Ayq8aTD7
cXsdlWigIxauNr7zbS/AY8xhG5EVDX8uxpFOZ8DhXMz7Vs2xLmILzzF1iF3Oay2I
ywjUIwvcSz3GAtDnoKBavQdF60pnbdr4kbSz2XnfjH9DaCjoqHRDK2vf4KxP3sns
jdRrZQESABaTvjmxCLKH+1ud91DQb3H7j/ZUz3xpfn+aCC3UltdSXMhHJ6oTZ/yv
UAorp5pla3YmftpA9Z/1b/pev4HOFJtv44NI7yOzt8MdrOBFrBwvlVhji4OyfaJQ
eJgwBBlyThMtFAjNA3G4+EOs7JewHEO8O3fNKgVTs+k0L1qa8IZJwQp4u9JxaLcG
JtMzHmSTraCJdTeBhY8fJMNjMGWBqM4EzbPhfYdu/SSEiWYED2fOSfzSOv+dnL/l
rTzVMrzvo7Ff5qRvY2yDwXE0zf/TDSSMpRn8zFFHJ9whAW5uAh86kJUKaGc0QWmv
7+3puWDwnErNDyUt+qgYhs9rxne/XJQNUVtxyB/60M6c4WZQVRN6+4bZ+RZFlySj
Jn5zOKWPhgUas34N/jAvG+dFXie9FfhLg+zbXyWBGOth2UM0JnQquDc17pUvRVja
BnNcWdd3J7g270MKcTdyOJkzages0il7Q5est4XJDRCAG9ngoeQOn8mT2JmiZct4
O5I95NPAqhMYcUt/RnbHSd9KygSbIyZQF+oyixqAzgmlulYOOe22nuWhF85GbZiX
w9CGRjjTjpj/gCSKzFXgYNCuvm9uFKtb13wnmLldY4MpuIUidwldVuWjZYruJHBe
idRQ7IU2GpnS5ap150Zxs5nlGwyhEpiHjt3P8nKWJ01xnqKM+fscSWfqAy4r1+37
wC+cC46oesx4Go1RUeDdBQyoEwgmtryo8I8sQ7tWmWXn7Xvke0I2apHoI3AMt15G
9k1Ac5po7ElzPDnh5Ut1HOIQ8BhW7FV3tJz8EHKPkIqO+BI5Riy6/PKj1L3waw0g
A4Y3synPMrlwi+e2ciWt2aK+AM6jtr3eU9nYRUkllmwsPbSaUhM/JqSTEjSM8eU0
QszPhQkMA4apPEOs6wsVhrBKAUbHDdJk2dpVPRvSHoH/0sK6hrPJB/hjTK1pVXZw
YN4kMYnxwX5pMv6Nt7EmndiPP+Fopi9I4PEW4jYbGJh/PgPooHrzImA3O7G5sNE1
OO1Pl4WIpNRsY0geNiZ991KfRDL30styriLWXxgAkZa2RaXHd5aT1tnKurxFdfmX
mjRHDawbpFeAnl7DBrkh0RgapO2bZjVu09raL138T4YWteCbAAcusIXCpRmq24mn
SS0aPOxLnz4CZUzrG4488hYrqwGs1vzaFo13cFh4yJEWY0WU5XI0Y04YiTj+uzh1
OZ80ivKhvjmEnvNmmTMVMNmIoLNxgZDVSwliCsmtra4wrRvKtLYOyFv7QMkqJ5ME
5fIpanjxsPeS5tdzxmLxCz5up3pSh3TCLKp2JFZxynvhbk0mHkwCgSidy1IWoX5A
PaqsgyvtydBMPv9oMSd1QcxVgkGYWBqeURbavMeDdUfGkPqVD28INnREzzjXCsjG
5WIBaEEjHpm1NApp9aK7L85N91RuBK2ePcXXp6PB9rOEj/fd0kXfEr3vHMqmBbyH
z4fu+/1/kqw8RwSNwZb0I5dQ4SlL5roNp1Rqjz6thouEB1ByxDe1mV7kxykWbNRX
ON/kGu0KL6x/GXYGC+XutROMnrSvHDb3IaSR2yw+U2vi5Re4Pf/5mK+CBJyKUnGE
vtU/aVlgjLGYZp5gzszRN5Jh4JcV76wCGYY7a6wsSZJHkEd9A6BuuOCg4ExFnBuX
jI+OdAsdHttEsQU7yOAaNPWjtcbqRxjuhiyxzZyOD5l/R/y8bYxc4iOikJchvHsz
MSYjj3Y3+Q/jnMk2Se8mtzvgTjfEcnUraFG1LYqjxk+jk6HaV07acA1OfdDXea5K
hRylHjffo/otmmxXfLRDpyvUgStIfSjA8C6Yp++yRx/rlW9mhrXdKeD7sXziygd1
nP7JGJN2VNZulsn2hQFB2Bnr62xlta+aKevVuktHoSG+2GXZFElXuC9YWcAwE/n1
jpnZqjpxXNzPU8axuyaQ3RmlsWyE1eEyNC0QRoC0f4/fpAUd7lVMwWDrhpG7a+un
BccR8jhRrvt9Jt7xpE+WR11jsncoAUtm8NqfNcZCQIG2+WQ4ofCZO0qfXqqFCEFF
MYLjV7v+sWjBi/eiMtunmTJ7t40nomZ/LS4T98B2dEkgkvy5HHnX/TCsk2XZZMgp
luJO1LHtUg5tmaeygNoW8LYlLObRbDoN7fQKXWMghJGltsYnIso7ZyM5JHsOqgKA
aGOopTEvBnFKk0qyTdzO5/3huNP7F2q5mAcuhIaronMob3TtzzB7MjBFrz9MeMcU
j7QhtRywyGqqEGkulsh7/ZKSTJIWGANVf5oMtkUpqa5ZSXC6vx60vIfwvu2yhc6O
VWAky9HgHPaClTD8BhqHTxQMKkX7TPD22sSRNoKkNa7r1ZiTh2LqcZF8Xj2LH8EH
zsvxZ3d40dLeFDtVwjBYN6avn/2rmCrtgL50WUQmfTAXVQYw7MCvjTsY/5JhR6i7
/0C/3nmcGougjntP2rX4hH7ClSYjGPsvuItrdz3qZjhXETVAPkUbeowjs8A+ADJS
a6ycy72mMln6FLWGRlCX/gCSFuOkjIatsjGZwO85X0U8lXQdx2trxob+ymLN9okd
+LiaxqzzxkZou2MvN/MG9Jwb276HVL+QxPXXyo3DyQ4JrWYtL4Hgvw1szW+kp2r6
fINJXDeH/h5jFbueAZq/0ql0fBNSdWWYtao588oboApoAWaHU8yZust5vVkBZe8S
AGEuT1F2PNZGH4Flt3/iD+N5DvVQrzWtgh7Lbjie5XE8auQBxEEfERjXHwvfuXKN
uMXTZVyLX1ehkT/JpRsLOU98FyQAmLnv5wbH7ZdCQ0HlQ0DHOfS8TUkw/omJz4MZ
OYWiV8MtwBJelyzuAzJ51PEf2wwYbRbxT+r+uqJ4rN/9ttKzC6a83LtyF/vKlUjT
NDVtX6GtBWIF5SK78tf10kuUNspGXfa9sE3YKK6UlL0F5E3gOzPF7kA/jatSMGkE
X5vxBfQ26VjT+JmA9/mat9ULSDQJpqznwRCj0HORXEBqf9l6zXxxWbDVOasOKNy2
FqHMn+cP1lucGpEGQV6cvxn5oyZhmerwtfG79mXoKG+kMupa6zgoYLdhZpcgm+Oj
xYlIy4nItq2WAbTZH+OI6YqDDljvabiloycdMANN/8nNmlcZThSIt/cMqu07zFdt
XS+m9zh8ok/xNw6cBUOggnUI6MwEDFeNAp3K1BoA9d4FSMqkgkgsh1GPz/BFwN6E
yY4oY5roiKxKxN3Uxq+b2aBvs7P+tLKMNb1EStGHTJxjPxmQNIWKatVZ+lJZJJ37
tFD0pDDvbIADdy2rak9PCDJ28b9mEbC8+uyvZuNlrX28F4btdEP3hGI0LzeSE+SM
Yvec5Q54yYj/If4opeEDi5WZAeDgfseoXN/GpCxaa0QgrF0QyvATnnes1rJdcaM8
Pb3zb7YgueZB4/k4CQ+CALqI4IE098v1Gs0nNP9LQzrC/z5lstnGY0eBWTYhgleB
Y9KCmK5+pFS2VXuVZ+9d8Bf2g0CDv5QCuv913Gq5sAN/WOXZ4SC66cMurpkl9JJi
PgK0qiA24d8HppscFGhILzbxc4IufUnHmMm27LNxBWd/KEZxm/tVuUBI/8iCc2Wc
nG1FQao6M5ciad+iiECnmaQB3EXZ8n/aJcqtbLruogjSvSZwRwKRQTOyvg9G2ER2
+I+YPxhA+9KhgBq6ZkWbublAGeEol2kBrRVJBr9gWXbyg5rAxH3SElrPD3nVv/NJ
u/RSnR197ug4Q8CweKo5ZLIASDzibPUCYMGGydCbzS7wA0KtXhINUQ+YnqyGBix1
ngFEOi8wZ4WYvLYMmZfEIo8Xn/dkGHDTI83BXu8LphQS6YDP2bJKYo4J/Ft9yTRg
bXoIXpKAvoGBhjGeM04WdT/qlQQzpO/9MqMofd6QTqQrrlf2Gy6dKIfkvzPhDfmR
zWC/AZG6r9bQMeafXuGYcr9Jfc/KZZ0FGQRyQczQL0VTTEYEwL4mFnmbtRnKEOUm
C/9Q2zdgxQMzimLXez6blOCt9XzgYRW892BmIaTntroPDa8mvAAxrSvtiU0WEcqw
3RCA/sh4vJKu9H8msa27k0ShVBDdjjg6PNgsTPQIzu746g8Hv/CmmVODfObqokbO
KhMA8ZxbpDrjRcbLmJ3tU+/Kj+B+G8DUvg673X+uLPst+6+h74dUNa/p71B6lzWU
kLQ87tI+pIadrw/0wOdUtPa3qFKxPePEL59PgODcLrokzf4rkk6/DtTTF369t6YJ
Cu5FnL/DsrfOeezwxe866AnEAq6FbOdHnFbhz+1RxpNj9LdUaUIxEocqurCLMhWS
+SlSMY9UwQBkW/CoTa76PZNwHui46npbKwsBbZptf1LQV9+eGGaddC/VX9Dbt1Ib
U9exRVgDrUpfnL8A0K3NdQJvPGpJEQFMAuiFregF67n3r6siH390v4RHyXBvBJow
9PvD+2aYXu7Aua+BcARuOTyXuLD1O8/i0VBSqRbIk/VPPASQDrjxLkWVj3DvRPg+
Rkx21FF6YGwc8ICzlC2E2XtOpUOJvwxEQW1lvJkzpRaKaeWVtw8dv0JJkJj7juAI
yYPon44eLfSQIAPyZVILgTjTbwJF5tKV8+fBJArnqSr5khJxzwCrMl8+Uaaz2mH1
mOOOV5SCWk+fZaB0qt3cjWJVRsBZ/XLFzzY9ivG1dY3RiAaCgKmreGeVpg93lufc
pnDZX1Fu0J4QdIUDOwjiePCuw0QqoSAdeJWSIPK/Eu4SbFVdjzL+7St/iRNk32Bh
9mvHbRQak3fM01OO0rZjk9/NfL3AgUyY3y2/XMqjH95nexMxKGYOdvErLvmNm/E9
d2JPpZKfEQ+Kz9LDXpNoDPulYnUWU5z2iMlXFqQyRDdcHiMS9dkTOLu64SXgiQLK
I7pz7acrLJYEYr/x8O8ejDb/edzgJ3walh5Ddz3zNwTKM7Wusl3B4XZSt5oFdyEm
MtvWpbMiPbNygKs/CEUSGB7FBpTwKIRIMeE+VYFSPqWpO9m6FJiTlonlrr4ECzIr
tXpBd+OiaHo82DmlzUITzHTp2kAyKMQOJyIJ/tuzraJ/X9HCpAeVZFQlAOGTlREV
1F4QCIMTbdjqUpTgE0iNBxWrKmfaBL0p7/Ft6hPSgwH2TslWKohlWV10pBt5KEie
gZPuHIxCFSNSldA1AWAbxsL0JdqA2ZCKpaY64WA9oT6Y3jqqaluKg45e+vG7TDQH
m8CjlrJQ/81gUpVw9Zvia4jfai2CF+3z+BFaUyvZb/ImbYNI8DPV68xs1p4QG6we
GZZv3pbEM2V89y8+JUk0Tm7vXeTFNUvRqbOPx5CXnysPd8NlpHhqQ7SPz48m+4sx
4ol8+8qWGv4KAZAEc7p1jZmyLxmD0gsxEKuzQyJzrFvc2/mv8kwqCWdkgtzCjEyv
+2ct9/R5lodHOWpv9AkJ4fhJhheIqZY4VP8AaFZBX5qonnHvem/aTwEcUav8YHVc
KixQSN5rGbPkzUreBei2YlHgUC0gTjhhr6Ysbijbrd4PhG6XUvJTdLdwuwLqMVvQ
e6lTwLChnzAZHRgB9o7k2O9KeN+K9iHWsElmV8K65wLnaE7F6HOrhvCCvDqAbOax
gCcroAdrTnBVD4yCsQp4m2fBAqJYBmMqTiK4LMZJrXf/AYW1/FvIl63aUeM5o/E2
oFTcINePxDEJ9E7ggSM6aEfJiNP1k5JjYpugeCwV5EPM757yBOuw218wr64RCvqD
8kwqU1RLSSlbTFvpxNy5EKmWzagR5FpblsA916prnEboQzitcl3/U9lG9wdw0Pbl
eRPBfjYps14j7p2hB1Y5LDDv2+9GeYTzYHnG2XjrqwASxZ/Tzt+IYtfOzyYhvwAi
HVHRzhHhG/HUR+H+6JEHPbExA+MNm5/aRX5h37HWs0e0mdA/r0SVTFChhlEwXgWh
wQI0RIAVkV40ycnJqiEA4UKDLndieMxS5dAcMZpxjJlzVS0WC/AycuBWKbJgbiz2
9uNz7ah8RSzP8RdVtVxiOZmwwmJDDgcn70roqXj9qJbVKDwpCEgOshKQLxI95u2i
Jb353kqusyphMWNrRHBbtpij6uK7eZOV6kUNVCyTa79sSd3JNDJop438fRn7AW2C
oYpn/RWpxCVPWNj2RliOKd+Im5eCHvQ/QxdTJ4jfD+NLRUDhgpJfw6hpzWReahcx
03waEnXMBZtqLnDxxiQXL2n3Bu5Cx3EnqAKQw4us5sA6dA949Fsy6EV0W2wuSdHC
ZzgYgBpW4q5aVFdp2wTGDNkT8ExDh9MM77tXV5fJa7huM3wPgTCcXhfRm6jUc5Ue
hLIJQVaUPgmfkZDeiocFzbXei47QAEpt04qL5nEqRpUbLX1ugHBPdNfX2Z57kHms
ZB4GHL7wbdgSyIUxyFFb0ETWsWTRslh/bT9HWA9Nh2tOwOTJ9mAw3ONDYomSbixi
z++Gb8tkEnrOoeNPKllU1RnHQKUefGLLIcpxmSzv/3gwjad+hdLQJvWvGMzdcafP
UrrdI2BvweH237CTUQybIXRbClA6k0Y8w08W4/0Tk/SkeW3RrnQ6KJxNzmHo4HkE
umzp2mZvxc8Gh3ci2QhKFqMsImUDAHKISGMJ4PsMxiOyJQ6pV3W58QNKVt1R1IAX
956ua4WSSPX+B7VXL0Aar5UNcsv7uarxJRHIT8h+bioDRMzjPtkYUrCRLFE+ZeJw
3dMF46AtGcVhLNSsdaAAGKqoAasDQnpYViblpbxXN2My7KiFCAcD8zx3Io0ehsss
q/YpkMGjcxYIbj6barxBNCkJhYBsaDFGBZVoSrP9ciikh9fAuH3BtaZK+dLKiLct
noLnrT63PCoQXOW6jzFtvRKp/3E20z/sGBKBREQxC4H2egZjg1k6PYYzQinIdxmQ
NTTmusQ4n4Mv3AHl+OTioRqclUhIIrGxR73Ns+S54tui3Z+GwI97rwUcUodEz4qz
j7Yaauvh1P+0NsAphBzoFpIW4efgltmKMg4v/iHDpVhKZyGLs0tJ9N+zrdFQi5Fr
fxVWmqrqFTx+B3KJjunQH0fkXftjXao8vQLWwGKOGsADbQYByAOtzsL3iyW56Ggz
FOy6PagGlCzM83yfmWBMmgHT2DVNFzBAHKgK3BnwssE4Vlp9noCDAS/gqSxinnvA
Cgswamf2LYXkDPhZCZTaE2UC77jv5iUcT7dxQ/Uo12+yxtF6AZMaiTWZDijoMXNZ
Y/vIAznT88IWHCFxpXcAWXpCP+Y+uv3Fpx8eMLhd3VSzv5EDEgMZ1cCs/Fhebeup
xf60WeBK6Cd1B9lgI2XfIuWt0wz6MM715VFCBm9ktzlH1Nw6FfmRSKYK38Ihmu/9
M+/UZEWjPVvooro0EJJCk8ayM/mx8LH5I26XsQ5EEU8il3Mx/QSCKVbPki4PrHG7
Ui4Q2pQPmRkmiIIuBboEY8oSlD+lbQyNaADprcu0a3OkBjisK2S77KoRUQTkQ4MS
gxxGWRWdxz4U7Zc1bYntUHu20CO7BpmHZfzeNqRGrhfYvQiwDeFJTJSDCcqeyJeg
nyZdTFIx7JBB++E2pUMOeI8Qrk/vSgr9g+6VPRNeHp9vN14MSRnZvvKhtxFCTz8O
VC0rAu3+7f6M3+c9bIrHvO6dmJ1CtGnZ2/kXGXNvU/qxO74wF5qpmOJc+Ta4OPib
DQwLgJl+c1WMlQXL8q8ycI50+N0EVqxWyqFHQmvtP09JHMb/QCpvXy7iMJk5I/Sd
wRdDalWqztPuXC+ARr9ulAGIYE78AQ50omKEFD2wpUAVbXwLeB7nVglmAL6IRnzq
X1FazKU7hOh8IkjOj/uVHv8TXlTbVyZRDlxRC9wbsDhX+yrwf9O/tVBAx+7yfQRG
3TLlxNMd2ayreoDgY3k68ylFoClS72YO/OpQVpnmT1dfT76wJa9NPHNM/fh0vC1Z
lXzxJAnab0eA6KON77iOj/odl9reqFyymKFFCLF8xD5nXqkD6kYNlv4tJzC6/+aA
aVECOX27fdtOY4yzPvdpapoMD0/M2U308ZGXdeljBFuHbC8v66k0VKMDMR376Cg9
aKwkcvddwzhPQSyGF6/qcM5fWvciPOFGuw6rJULh19jkH9xG0dCstXBE5qI4MZZ/
ohjJNdgQ4zLNnKH3ah/WevzOHBAOvOcT0Mx5awDZNH5AQMMSjBo106m/SS7xBlHq
6nE4ZoxqZpkM8XME8F75pUcWKIONayZ9BkIW1dqHXkoMaYHZBM0OhWSbZjTuObe2
Hkv3FCjzfD1n+9rcmUYt9mNpRQug8TXtMfdK+qLLUD9pus9UZrqNAs4I8VQE7OT4
WopOAFwayUaL8rnvXdF+VWmbVorqeXEoDGmuT9rXRT+tvYrMKApRL7zo57L8Wg2P
K4a5argNTDO2l6+lKfm+gaRpCws3ntCfeRuk9HDrwuBZ+mmzz4YTkaiwKs0lCs2F
ovbRX+rxvq3uFXw3u1g7SmnAzAmK1IwWsp1HIol0IK7txZBK7fHqiIbk/hzzeyym
kCCbOj+8JnVfDA2Ho0VYvktnyt6VukT1gEswzJv5lQRIESUu43JLvcaM/bWa/CKf
Xh0yAriu0Ke4LYyfSn0hM0YdodeC23hLVHFlEtXTZ+GM0d7kOd8a4nE2aMvRjeeP
gauoCR/7FKYVJb81EfoYys9b2CRPAWQuAngN7+rOj9bCCydVoGrz+J36MGPqfc0h
R3vjomBHgGnfpPntaLjfMdKIrPiQDZOvqZJQWu3Ti3NAecNpqAkm04raqwN7zVmO
bfQTne5/RdW/3Tz4EbIdMdMJokx+G9WzCeUUYYSZSyRB/ZvwcBWGduPBuSNlVEbo
u9EovO6hlg+TreA8bnqQa2/bpc/syI2WPwXQENRdx1vXdUvkBonsrpoHoEvrgTqB
Ee9rlvZPdi6PPu1o+MPpJsJvtf6AoH39QPMaLbD85xYUdShvXnNcz690ErPVRowX
h8Fyu8KOY48ULWqBto+JF2GpcskNJ0uB4q/loCYceQ78RT6nGPm/Uf+5wrgMOfkj
LtwmyxnsSMSEPCc3zfurAJPnPQvtLf24AlgC327HHhlAHKso+gLbAlYM+Pr4kbaK
SWEr5HL5ZnuFNL74QAz9dnjyCfASbQzOclTC3PF4rH5JJTiw4xCoHNf9bp4YHBC9
UKRVLHJMhdSRlGHJsfjmJf0HaWaqyBFOKaExCprwwEFqOdPI6YTdMgGh59rMRkDt
oBPreFvg7UOh8YwROqXXKmB4+aXBXM6Ji+Ag1GS3vNLorFglA5avIM7Liczp+O+4
YaddIfY2JaLMTGhncUEZuYuFyHtqk/eaSwwN9XqBmQ6REnMz/htV/kn6XSbSCK5J
ZmFMAKXwrsts5uOutM4yyOqXHVzRFJYOEyy7pxCL6q6velDi9P2vl7M+1zXZV5iV
/22MgInYTXRAk6sSvO+IpZ7B2ZDvq9vvCWHQWH7uiLKIdN4KA8zZU7DQF5zCag0x
7uX6EPwMrMTIP6L+M9bw+zTaGrHBMP+BpsOlJGllXputjHvwCsf6ihtpQtoutwAP
WmC9KjZOXohRK4k6SV5DJhwbGfFL0FFpfiPc8sIvH6owK34/78l12xp9wjFYDfLM
WEnQ9+kJw50LhPEtSNDnYUp6nJqZwa0fY8Xh/NmJEvY4+IALqNj1sp5MhQFUynhH
uIWgCbJx8W/WIryAmkja0ityIMHKDygGexpk0+7nz0Lrb9SPkE7Pjm+BotJ3EmTB
tyetNIf1xdP0unghiDkdvZH3qNnAzF6UVR73mkWd1fsgdm92sbKl6n599/9I0tGY
oVAy6m+qoL2iZ1U3ShB5XvSz6sIXItLHoDzXG52bnsNho8ml40VRRZZtdLNz171p
ddkWK98BJ6PZ5YAX1gcthYDqef/CiZIXRLLY5Vkwldkl3kOW8blbxEYoDOEX2hCc
UMArlUzyoVZrPlL36H1wbmdP0VCyez8TmlqffOhD1MED0/k11Ik8h1jeYW5l+nk1
2Nb7o56cgex4JqboOFzGxJXyIW7LIpTqwDBe5glVo0Ng7dP3eO9OCMyRslJQ+91r
2HCB9qYaDxNKr2zDWpC4kjPDTk7uSImqLOmNCCgDQRPMptXLlQ0q/2cb/2ecWQhe
NeVisozhIUc6Aq7w6ndGWfaXBxScuK29oHm//4uWnmHGFBQBZzU8cmtgKFnf0FmA
/Y+5edmdgrueYGHRRI5aE9UC8XB2K8uaLKdwW3JoozYv5qM3l6wlPQok6lfWW9ql
tFNyIv6QiFYFbvPyA+kVryPzCYybHpuTaYB8DtAOy2PrcORVLe2Ej3P71n9XRTKm
QJSFmXm0eHD3zEhzO80kjs17aB4OhwR7ES6zedxXapGRnWDQVL5/frPQ7B7K11EM
nH21MXmeJooquC3oYHqD010LC4Te/uevhf62/2M9BVeWk8WRnv6R/UOuM4PbDmiq
FFzA8KPS0tpF1OVdgpUG1hcqo+sKszMR9+JBhAlO9qsaCvslewS1n0XiaTHNLbBa
Tz5M7gMyxBCpif77L3xc8r4ioi4+5I1m/s6F+1IQJ7NqgtMCviitKCeEC9KaAGV/
DYrX+6YxbnLTaYpq18oLnj8fjs1t4ZoLupHqAJq/wvgug7NSZ/Dt4/niPjg5g5g4
u/8uu1+acGkj2iwBnFJJCSsMKWvnHpysbzwFTJreXgb19yijEMtv7jSuMDSg+UeB
ngBDIhU+S3otm3hTxgFo02FE8kHfU5YhCY6/A/53TKIyonMDpjEov8qJ6r9LEcGG
8vzAffLhRar9n2HgHgMiNE4LDW1WphJFQT4R79J6hHOfgwuJ67JR6CxxA3BVdT/A
c4ieJNxvbBsba5ha01q/L0ccNpFqaVMXrD5nr7P0fN0iy9DT7hA/WmyZBiUjyLW9
YtAcLHVUnOTWEBXDU1THaPNpGaS87TaP3eHksyV4KHm5vm6vLe20QCzKq4RX0HEF
om6jTeAvF4oAikygNSGFp8zAlefvmAusWVBmxV1pWNAC0w0To72AmqqXeM9Q0dvc
vuIbR51+6Ah3Q/7p3Y3p0oTB2A03eyu8cPkekwa6K/3/SjoZuRwMVB7/8HR6p/Sz
1RxXKUgPVnTrzP3Co3wPsllYtVoLgEp31rVMg8OBzLQdV6r4yhouy7svxpJmNW4V
qbwdR1W6D25jLrUHfhJ+pWFvj1KfA0pGlHgojPdyaqrAuqPzYQBNxlurNs5ht8At
j9A+LojkaTFnMdVM7UCtnvug260y4gg+mh4nVV6Mt1KSNToJUfv46bFskdsjvwDI
gyhBcKgrUzknpELH7S//mkuiYqJBvL68IdcIoxuHO9ZwJBpc+K0vSZQm0mh1Egyn
FQ1avu+7/KW7DhEMLw5Ccp8cIiSlgnsLXBvqp2C2Bc8Euzp+zQhCGrwZT15Uoo0K
YZ0fWaaMXUERDIyA38d88bFmcz9Qa7+h8g8VX8z1HMuKksIO5zCUqgffdvacaEus
EFGcCIShsaOB+E30PXMPRmSSyw9HUlObCU6byQnQDLechFoZAf5xFMVKyUjWddy+
C1RdiG1+BBJ5kLp7EceE02ku1DA8+hw31cUlX10bbTmNTXeor/nNwRAtZ20DoOkw
DeNZCzBOVZnLPPMoO2IbeEeQALDZTIR+/85aWQHlU2uexPh/JiARnRQXl4BU5FLi
kqjUaWCNORP7nUiAEHlNhK8R12EHywxRFJXj0sT3shWi0LUluMav8G+6DhiLkX1A
x4iBM5FsRLJfQGfOUhjQsp4uUJLoJTMzSkLi5Yldpsh4Kh5YXkVIQ3Y91xlKv3l5
bUPqC0gamqLGfV59XFESl/mJPBEOsZZpFEq0QUVDHqbf6vrAw9gdt63NtfuY4Gto
xo4pRd1/SoZhWL+00if5gyAXBnw4n5N90oZQf7kEfOP7eewHOYzfMuJf33VqOLz5
U4f1cLSxRHNlKQwl4L2azPxEvr/ZTNuoa84aZYUJr4ma2A+OCHTIznOOVP9eY+22
VbvH2TFErbAL8jnEEBRYuLDaNgvzhRYPDoGlpVCSA+An5ypL28PrA1UZdnIUVNSF
0TGBu/drJddKCcz/HQVeeC/W3o8v0zoyBkmn4paL86Vstf6mDWBb+L2B9Z0GvsfN
1skCbd5StHUoikPB8p545iJxKtbnvog5xzjVKhsTua390XorPA71+DuzO3H5eRrK
wSDZKmbU6EtzNQ4cR+avcr3jUn1XsN+wp52c5A7DFbfa1G8wIEpwL9X3PVBhb8ox
WAnvhuKTO69yV8V+z5mH4rCrybExQgLE+FgKOyKmEmTMPgRfG/+V5Wfj872AEJ0V
PqdJZ+A5z/Iuw5iriA7iWoaLsyutZvvZsp9Dv/HCjE0iC7uOV8p1M6mMQc/kxv1g
VaG2bheZ5W00DgHlp1B8VM+SAhk4uhKcVxCHeFl8LCShm0AqQ3vZJmbcxGFZ4ibS
nm0ZiZ+I5YPV7KUf9Zi40LprorQQ+yxUa82e+nJv0Sv8og3HQFfWi6lxOf7mERIk
ZrJKe9d1Wsq/DkQUPkOAPcMcq3nXkSezw0OjzjIfnNVqWINw52XxUwwEGoB3w2kj
hisaaPA0TQykoydAVyKhbVe2jDyE6BryTWGPD+sx8w+DSqvD++kCWSOymmaZMPCO
OT3en55l/pgN0UkGrf244MrO9weSmfhLAhiWhTonc/a3psD5twrH8EalbjNo7QFB
9dvLO5jpxwM8WIhL2IViVZF66VnvTk7cN3sWN9c9/H750xCCcLf9D4enoysxc5CI
GZi1bmPxrhUHajAKUgPVyr1yGESdl9VerFeBTHsJog15z3QosL/XIkXjRtfPGwir
jxr5aEF79W1XHzLzvBy19lz08t4awvCsCuob36JfpnkEsqFPyVP+WJlyJjvwmIst
xlkJt11ovt/giKTI4kD6z2HdBtUJxTEYVxF43V1760sGwnUr62okocypxlrNQWqv
rU2GME+RbKc9RXrnucPJKD7ZuEO0li335EDmhtaHiwjP048UElvCP5mccW+6Go/4
RrG11lAbYx6pPg+CE+nfg0WDvQO3VcYZoXxxI/02zt8Xce+pYV2nHJ+M7Zouj+Rt
sD9Ybg7R8Hmuu/EgiaR8L0qe9yxTWb7DEiwnIkd063PVMzlWfvN8uwjcfG6xV85J
f6Vq+RQ14iGajJyJj+ZR6obHdIHdkpSg9TrIN0MiNX1cBVBVQjWWgmR3Vo4hfnXI
lF3GVyKdGEA0kDhgLDW36EOJ7HNbgwfzgRwQULZslMDZBeqyklP6rHLH+beWihQc
caklk89l13nmGZHXraPsA0GsCyOGPCxeOKODBUOD0/iR2LrGozoWX4ZyO/PKOB95
urxXt/6ik5UvdDFLLi4hJQ8OeWqAPmH66HRUbt1W+/2yTTVu8SPmU+gse4FWpNQf
VdoCllcLAvdm6kMgMw3UmcyXrV3Io344qxMGhDT5qENTUNAS9b29mhxuCcViwLHv
pkyTOPsn/BQe94pHLOtEBvr+tu4UCd9cVSnXCSo+++Gz+/8KNIqAKnStXgA7zqFr
SsjfWEghJeNFLunX9AjaB+TZuoQ8YafusC7Ry3l6L0Zew+XmBgKP14vSUbnDCD3U
MSdHKLlK+zJMcsALflaxlbP8+lzGoeg2s/r8Vv1405R+q3wovFJM6bR0vtUtUynB
RYYJrTLrvz8SWmiUG/2J5bUd97ZOOmOyotK15OtSzkqaGLV+Li9cEGmOgSqcqu9P
Uk8JWV/3rUgdiP6IdMzxX1OiCRH7teXsTiIOahYBbPxadr7zPPw0wGL25Wne5gRo
/mL6JBBfkNFzRgLRQSybg6iveBLjSyBcU3CnseAk4e7vhqXKPDfSbDOaDr1yNxri
FPV6I0j+vFtXnQoGevf9U5r3Yrmkz6JmmhbpBQ9V8qYnpvpINI3umyrvYF2wGQb/
cyXs4d8tegpMPxH0ybjdCjTcSGBzTsES2Rtg/3Wa4STeYar+RHz8OmFrBFTP1s8t
Nly2oB4YHnoj4wQOhKrq+Xf1mFq9EtancCM50IblAbXu7tEBCB1vj4ObWhhyly3s
89Gm/VQSlh3od9NTWkTzrsoZAY60MH5PRo+HMuiDza60Hfnsva7cOrWTFwkM1cWc
aY7p4zB1Mriy8yE4lm/2Uvd0VGuCIkV0xgCTqURD4ikVBAn5FreVfSI/eUJp8+T5
EcpjDNAX5banv9wy8HfEOkP5LIpAaYEZYi+JWiNTA5OdkSttgNiIpEr3SDtFNuMw
8yV2kVTqu4ydJN5JvegdTqesQA3kq/JL3onXgZzwVC8UBhwPsezrtEIi2IKsWj41
hWDNc1Dde6ofvdF2j7VQn6NZL3S/SM3M158MnoEssqz4xSbMkATfz5OxwKg/bLbD
AvZwc3EDpWtgxcN6FKFLBcJtQxN2DUmdWhZQ6xV7mlwZMXdMIrbCSsjzU5wm+aw8
BoeNL7TAXI6Jfalp6Xz2vRc/L7nvLukWchRTrXKj8pHJ4ZJ5HDIX4uGepfPmgwyW
sbLWDuqo/kT3GcX1xui8CCdWlSu+WWaTgyisSi6j9HmQecZ+wqhbwHJeL6USrYEA
Rm3dJF7TtUzcMCSYawLR6fQddlnJG2N9p4ex9Zz7Ofd9YlR0SXEIW+eNsUeQRffx
ZK7q5YLY7g4fWP85/MsTvs8yLAzucRaHElJtt7ZY2BksFTbv3UY8iTjDUW/MN3pG
/Sh31ua/UeC5p8Yn3Qlt6ZPW+qF2osHdo1RIXtvy9L1EJQimxlVHcYcWoe6dkV0N
Z6jj/kktIeI8LhK6sNhz9PDH3q++eqZhJ1wmgdxFpFHWdkEyFg14CCwapMh2DLud
ONrMrrCieM07oKJRiG9tJP6210RDs/P7VRsFgM/Vegoak7MhMeyqnLtp1oVRFy4W
j8VUrQbGRO8JEgTCt9Ob0JUg8ZsqLJwyOlO8Yy2dTqTwAYt/p/hN0A85HftAi1Na
2HsxZviTAy4gPbFzLwQiqm/8zI5wZxvxw4cvJmPB/AjQsS+Cbu5U1uN4kOglxZqh
e/XW3XLZa5Ker0l/KBjoaeVRQMGDVRBUNEoCLiz/0hyrIw7mcMMspcAgjrkQu/EU
KzcLiVK1vFn+sv5gIMeOifFGA+SpK9E9jLSbV9uYPECxArJKsLEhCOGuddmRwNM+
70AzTnEs3T1eMKSthSs48otlhDwwHoqCpA2LUY9Tki9yp0zitUCQryptOoVrGp8w
FqKGDE2Pr2ZqdDtP4KsFxKr3FeKqLqo3tt7dAHxjB9qFMj+kDTZPQxy8mfKznZx8
lq8oTbPlIfHAbKQvKpwSrTC6+WvAJ5tsrtupbEoCxO6C1Wvv8zhJWTaGB3N/Njq8
w0NK8WVqCsOVRroypQPN90wE8sGaNW9VRJtRI728SRWPZp9geTVkBXEyZlYSMqRr
S36/N3OFkMZiQB80M041GIzkP6OOljiOiv+BhObYF5+cTlxO6cbWl43wTbkBwQCt
d/9eI555jx0sKylmChRmBbAQvs8XKfVqOQPgukJwEIU8wZV1BOD2rhRvOq5A17Iw
SlugQQfGRY7KBEa27/YVxwrufVBHHWIG6C29QudwtQF3PzhKlUBa1qVHFQS+q1NS
Rz+jHfvHhFXfJnEtTaPmyeNHXq3Ux4EBzuMzqMCo0vDgJ7VGkb+2mCGOXTO6YClC
7QUUxfHQ0fzqPRwJMNqjyI36P4/CtmtmynMv9ecSDmxAsurgaYMT0Le9XFonyZRP
nPX5AmS2JKzjjnnw/FAFUZv3CFX9OVc7Lg+5kX2HTcbO19gvEw3vOYnUTOpflxZy
YLvKEm4f6WkvRlqHQ2IzCZhUTgM993wYnClgOnBOFqu+PSJLKGhVF8A66TjTTGOX
/Oqx7aW9TmFaJ8pMx9j/RAGDWYWBDJnG5TOIPNayb0YqJl4Z6Mgg+ws9vKZEHkzL
sxsY5ViQOim5VEdOAsUdne2RFSC3BYhFpLwd4Xzsnbr+ZDMZz4N4km2fI8x7A+TD
gHXf/rb1X8L0+wAOyS6d2tfgVnSKSJPXZ3qu3kV5B6fcYa6ypdNZVg4UYZHHruJA
fWR2NfUXvMRDov5bhuGVHKtAonE4+IWbPe75nR/+xv2iaNBE8loqZiTOaiF815Pa
Cfsq6qWYg/YeahmSlsBQ+7TamCLpRSizuqC6fwHGl+F4P9Ofa8o5+zWcetbUjs9e
KMoJkqqU1v0yBdhtA7qheaf2Hoi+pj25MOmFZApkWv4WxVO/fekIdv+mA+u+5sX3
K3mAJBrpaOClxEtPcicAA+IoN61RBqRbkFWtnELbUIHl2sgpaVbve6IpypEDS/gJ
4wu82VkrWxX522o1ff9i4BpidE753rRBU3qwh/4mYnq5Tx0/S7VpgEErgYzlV2k4
RrdjQRNvMGUCVdeg8wDcegtCr35v6I6yuJIharPPLU/C93hMIjVb9HkJa/IwEWG8
38Rv0rewJXvr9nFUlv23XxHsd+MfWJPQz6MREov23wH5GaAZzxC/hpaAUWq3WV3H
OspkH28w3pEj9djKogftjrBrL6kb/6WncvLZjEJrb/zkmfGCeuIrcLtE5If4bnCR
kZ+Zl9BAJbRz+JKDxOzfUr0FfJSH70QjDWeG6lX0QdsgqNvOghJAasPbIbSwpIoN
fhZJl2r/4tLx4xK4v+y+AmKhV8v1CVIe+1s6A42XZXf8WccD6dClMoKCdVH+HVA+
8eMU82gVkaM466I9CoxKsmKkhbJUSWNlQYrJLmnBS5wVPX2uiUlOPzX+cJlJO3QJ
NDmswuCitYl0Z7wSBidE/6P2pt4gxLuDY7qgiW1Ex2GzBgOHaeQ9y86w9sc3uBjL
gmyJkf18nsQh7oDCFNbs8WiCZzgc3zln7Ah5S+O4fEKDA52vKTWjiAyq3bwFcdQ5
IlrEcMBTG/ndseLnAdrVOHLEfWBIacN/BHjhT7t9lkkh4Ltw2AbsguvUHpcG/nYQ
6Zv5Y/2C67OFBuBXZegq7p48seicS8B0xFsBDEpD5jMGhFNQ4FvkY7PKhYZ9ABbj
DsFqRTR7uWwbXYJ88pJBO5r7+98cxskYVW4JLfM9vOdL5kvuagBNCU5uXAmQE113
GKNEh0rs+r/+VjdYRUGa0XdNyXK3RD7qEbRnmD8fxZpOQlGUzbr4srjBmvn0Se4B
GSyrXIBJYrMZRozJK7YNb7g1ranLGPUaYUlT+9DK0VjRbWPeWWbDLyye85whRPIU
SJXJT47cJLBM1/XU7MBh+/6/IZjm5N3RMaVBB+RrKrjwanLidl42oiWhKUczoB1+
+pDiuZJVKLJNLRfkMoWKd8qcKej1ZV1laPPwef87dfVYJTkSUlk9AW/a6M3euI0q
7XnucYvxu17xM1KqdVVHZfHIG2KA4UXWFrfty9g+QP6Axr8iDETWsGdFhqppf6Ag
odxkShy4ICMKTmis9YLXiI1iypXMxwocapKLeecP4GUcjEkg6y1EuzmVUJ43Tq4z
uOb3v8T38l7vcskp7lm+ZAPXJndLLtTrVlO3eI3Ke/Hamnu69CavJWdwfy5wdeaw
r0L9ibJQ0zcII12xO/p8n0gGHEqTGH+m10gz30/oOBd3TL5fdwwtQws/HbrtGSL9
nxYLWlpf4hrfhqKo2M97NddXq7v2J/IqfjLQR54sD/+dAVt9Ju5TxVSlkZIYSFWk
IfoviDRf5wKPbfThgebGhSc6lQv2dh/vYRx3i6TgpZItsBd16Agts8TGozGtHurT
4c4WeU9z1h5e0FJXLa16eVp6rjGyYsxR5W57pfqD6QDwMcqafWZrsm9xhbELtEQX
PKpYxFVXJ51eATO8P97VcGyPkmugrS+kNarqGhy3Q/LFcdjjlDQC5gbuWc6lGZqx
8J6wScAzCtVVofuFO1boXMCZyKKHuf8Dh8jgn6DNh8ScjeAwKDCwy7oelFV5DFXd
DqLmjvKipN0XPnhOnb02zRFR3tFjy6AzWDtADDKL/0YMh2nLWT/PPP5ibjFw/eY1
c78rHVop0t753jTwERWDC5C/hDYsSzGmJSspQJTTZXxv6rZuBtTqVy8Lr8FfVzf8
GmBX/Xm97nP93XvQdkh+c3epkaEw8SZrfDs1k9sAZbPYEzaBnBZAgnT9/9W+11tK
VDju+QnXyOL5hzUmmwanGxLsLSuFb3rzI3CwnkQ2EC4VidBkgi4FztQK9e61ITGA
nB29AKTQFTThb7oSBwJaoQpSPhbjOCoQXEw7C/QptRFsQzC58zbqvYTX0J+T8lal
rFiPz+loFmHntDEQdF0R1I4QseJwjLuYG3A5CswASh4V9Gvh+bS2TtuS8pSxhK3L
ZGJ3sTzSKqvZDHh0XTApO2yMA29dTrsFcen6IVJztvHaN4pfbDGF0cPz/KHsBrZb
HTTP4hITqxmFoHnDtPrOQBmRUAmFNsz9KvQE49OnC/FA6bbkfwfEQmQTQiQI1y3r
090K2s9zUM252X4vcziRCLSX3up8B1vHfhR7GHBxJLZWH5WQBguIY6nbJcGcXzIc
WuZst8gLBfAaItGEyGk69R69z+YaiMYPCXkd2p6uDgH5+NRXLDrZKV4ZtU74bIdx
V2I9RQ8WPoSsC9mgbDlst3EF9VEs5xeochviY17K1udA5QdNOw1Aq4W3ylFjvqbY
Jp30xf63YB7essQ52zyWhWyoV3djfUFckt2l2Lc4m/7ljN/hK0eTaMjt017Fk9bP
jHKIWOcc0uo7Ox8XMlwqrUyajcefZOy5Q4y/3FSgHT44f6nH52hJV3qTZBlM6Re3
h1ra09VIuG1A9gYg/cLB2vyqT1HpsOGpWGImQQ70JOWvQCvls6VeHkVqvECz2UX/
r56GJAD35Mc4fonSHIaupTJpF4nDrSgO+VMpGMxBGfkup9i1sZ16YRO1xQlYGoUo
wufuBjjGRujGJgA1I9z/BHxMmZe83f7I7pWv+/KsTARnuXdtwXm/2u6wgQ05qltu
PMHHUNEw+xWeL72xVQiPgPSJhjJyApBzD6oeBIqu/49g9rizSob//N1S9/rOULZb
9MPoBNitHxPMUscdb6vMPOL7bXAEyzVrmIJU56Qe6iiEHaJqTdwPvDySHdhVGham
rZCJ+NFyGHDKKoVUwFzpYA4RZUKtjIq93qW0PA7dSP+YY2PQZfeVuiE3VCD8xOm7
EbdBSqilJVu9oQoopsM9NvgJK88C4ktFLTLbPuSNO7tAv+sGlQDmsDzZTYXbKmey
P6gmyjTcKVC5YtoYThFeZf45Rji2gNu5pyF/vgjL3xuYZ/zSV1cSpL/5bLGhcema
ycZRcUuraFUfv8d4Ve5Y160a7bGiyj4H5JzOrwYxl/XfxvP1kux6aEatIigs0HrW
LQeFts85IVKR2OXeKVfKihao6WAIy8TdW1JMDrUH6yjE2Jta3A46FTdCpG7NEXDp
8FsMlADhyy3LYQcb3BXPBGE4GlIVmaQwr8Jdtsb7IjRYjvgzTsHoizaB2wYLOkiC
Kitrz1fZ3PGE7F1G7DfgT58Pjeb7IaQOhde4RZ1Zh8N3SDaTz9PerrOnAuz7Bqpi
FH7YHc3gFAaD5nNZs7a6ja2nkG7jfBRk6ckoiVjmB77hv5miyJB34RvxddfLCx3Y
ynwc6hM3RDHz823wiKyOJ21Z86MGuvZ3JzROCmFa9ts43us3OycUtygshrDk2faQ
ZomxV4Age93vHhYsK8z7fkiFI4fl4pXglzEJeKL9FUif15779Hj2syTt2FQ2yYzh
aCObzwctiiR6EFUfw1QYsVvJnKIpC/k2Voyn3yFYO5a92MKf45Z70Z01+APD8g16
F+HjqiHErkjyHaKXI8lGZcjVFA3w7pLSQ7ZSQVPcBmcwLQTVp9yrvwljPAWNw5Gc
K3zoFBb6Cg0Nwdfs+gG/qVEVrEcBSpt8Tb6AB5bUUHHE/N31Bu6n34Z+WF/lTzaX
uAjPs9PpTlzPUTUz09cAMHi53jEo0qOfELDLxoMOF51YtOzBDrHmMrwnIKJTLqRS
m1FzoUAeVDpN2HJ8YqzaFvgXUe4zieS52o8HfxOTU4eiBQ7DLitCsYSS/95o9UiT
JJ9APRw8RT8c5eQ1z0tbwP0qXXXS+68WQTa05za+YchUVt0Nh069AAN3nc47iZjH
3vobvItsozOV9TXdeGNYgN6sSuit+0nLFZiH0vw3R+LpB8nZQoOgZNhV3s9iMWqV
JWX1cRsxG1BEX2TgMYrDbiF8/59hVa7f27CVxA2xL1lPl/eK5JJIsWaA8tM/bypJ
PO9Z7OcwGFIg65numElWgjzS+Gqe9y51diULzXOp1cfNBUMYsS1mSCw4WSKUJkyA
fW3mLOFrSWglw31LQB2fWpc5GMdLm7KjhEiEhoV9TcHxSsZdRlPyncCrQJFSK2fK
nwAGASF6my9nUofR+BfvxdmqvqvrTCiSp6R3OA4V6IA3sw8iW6wsICg8h5pGspay
u+maEf4DFUUkuA1iDTfVcF8iR31C0+UWNHSg+230xKTRj3bKzpFAn727EIne9y6l
Iz6BLmM75Gv+5zqZ41we/vU5ivNlm86i+KuILfrJWMIFMAROlyzvE1/mfTYXP14A
rLFe/l3FP9zNyL6EouT07LwxID3SnNg1VG4Wm7Nz2+VJQUscTfx2ouWy+nRtoqNx
5M6tsqiptF9ZvcTNKJbCKhWqsq3R1pUl7b6tSOXxLCPgBgGaG2ZLMAIZ9enFANz0
k7ICM3tQ4Y01I2Z3wK+u1yxbPJ4DMNgw4+DBEgYhEEyvb/ojkx4wdipa+fKsimIn
+k/CgwNUqChDFAs9/RWHfwzVwnD1sViaALI61E3JJFPLXw63hGXTbgSx8y/DVEnw
6QxahOcaSvmS+BfwBvX3IVnI5yvMwg53gItazlYT481nPXEruWB3PKzNhJSnWvGw
4W6mUstNXhJV8OMwIkwvnNvMMAbgq8Pku+Jkowyh7niFiG4t4l+U3VyPHSo9W9Z8
481CNfDOv4YSee1E38sva5w8mFL0GzBMiXXYlZmfAsQUxjVftFhrlBuM7JoQZWYe
s9mdeRxGrLtwVANkaZcnuoKQNHVMsLagG9HGwO9lMCZCVHQ9gzaglXrwumbPjP4f
OQ5OZspGFg0PqrRT4xx1LSbnh3FYBPWNqcrrRK+SP35XF8xdFtAz00EpKGVkAZtr
PSpCgCTyoqWS+GWsbgegmuodfcc/Kszg0frrp07en7AQH5HnxcR8k9CYlrK9TcKO
T3uEWnzyR5+DgJCX+CHqbl7ZeiFW8Opm/RYHEWhL3V+YMk4a6gATFP+7xFlGc+gl
qys0u8z75gQelIEhxN2/t4w+rUh4gUc/KK21Gyu0YRQmMPhA1fhtR49/u13agGnI
ZT/qDQk0K8gYUDoXY+GPCDDbWLuBTLAItZAKiqAyG9r9h0j46jaf5DpNAIDv8Wqp
NPD3M0sazdzG3EhCtCMEtNknMg9Vgpbypeijtu/ni10gvBtX1Kj5RwkdhEMPRix2
EaEHt8BHz9spkzGLoYNyh5ODEZnw2QYHT0JxtvN6A2JstHxnfApXYTB4yJFweoJx
s07WHiiw1BX4IAnTGcitbh8PFAX7tgSs4yO7zTEE02Nh3tFBCuvVkFJKGMC5i1JL
NFprL9fdvsnK6llYKuXcmJDqBt1CO7L59TK5n7rUomtIjMl7YuCTXoym5sGu4uBG
I7zPQPkOqnCTRf/n0PB0/UlKQlsZC5zafs9Flce1RlTjIpquGH9glfrLlMbdH/JM
JFG+0t66Jhgf/Ir4Nxrdx7aL7q28XA0J/Hy4qNss/SFAC+LnoAmg9WSIpJkznUP7
rL9Vpzui6tlGBD+xsmJJ4Nrlg5NBSqd5p8fPuoUD55HV6IHxhJz6c4cReCdSkgtT
V5g25QKGTbapj7N3C+3Xdu6+jlBgZ9Hp1CBV1skeHtuTnD8go8Hof0sjIVSsXvy6
Rd4K2zD0XMaqDQqppcIXWcGT0tLJCrHw1yFIamMoUTJ83kr2v1IGTvvv45w1IwVx
Iv1h6bwQKSv+Cm/CloGKxzB0aQcSMxc0woOdnuD5W4OMnAEqVX1is2S1G3uAv01C
iemJ12m5uIMgkd7PrqLHQ1d3BUmXpg2ktyg5eRnOLtjl37crrpcvKvEqPYMgi1NI
P8bQNLZSAbe6ECPdk091Sz+Ix6mVNaOKjI1U4r9S4josfncW5mn/MsFkDTVEXQzg
OowSrSjUxknLTFhBgAy+HPRIIlkRS3kmqXDL3Ht/Wfa6E/yGeOObcIIMNmIvxd+D
R2w/mUFbt+gdN8i2wxfFR7v0kERmKyPHWILrV2EX9JcAjp+t3yb08ZwiC7TFQIza
MpM6JpHR7WIHDwFYuD0LUSnHJ53BMg76QLsqFFj61tmpJ+2QrrQRAOfaqWYoXg1H
iIUaPUpLaF5T3n+n8fGU0a6W/SrYcfC5DUGlj5WFfGE2A8pHmG7/OJTuXSzWIxoB
Z8nenT1o4EffZSEyV+a5D2yWhEtQPOq7kzkWrqylmsWxvfTxpk+vdVWOUq6qqKQe
cXNmh6HhirLypPJHTWL/NWsi2fTvdYT9jsy5GRJl74th83MMIQztsyTknwNrCMNo
uRAncmnhuS7at2bXygCSb/5i8NicH0I+83crPPP2N14UEVqUtF/Y/V+UV2TcHV1A
XcyXOkTSvAcPa2kT7AxB0XI6oDKm1b90nh9bMdxSS+65R9LXxL3qv0kpS1HTx791
q0h0JPN2t7NOmQHx6CYw2Fdw9oksv2zHMSP1uIrnbLaXOjN6fk4SJcDtUmU9d/l7
lfGr4v/DZVz8h/VgProBW13JyQmOZ9SX7tpbh8vK8auBKPO1eQEM45UZR0ae83fo
iNRkRy+LEA5F/L9+yU1tx2oA2KJDPw9Ku/3WN4waIBmOqXeYJftHkV6A+giP8xeO
GO+Y29Gb2jIp2Cr0vBYBQ80BZgsWmVQlR4SQQTAmDYUVL8DPIp0kBn7CblqSauRK
Tj79aMC41SgrVyRyHhdt2YUU4LHn0dSx0+qeUC1FZ2cfIfF7pZKrsdiHjjOKw2yo
csgXg2gatrD53xWlYneD+pgAzGbK0VdN0E0k/AmF1Q65pKbw5n/DKP1Mh+M37ako
VkBCIu8MieS3PiCXjrUgwEQ5T+VBbeVv2m602DjoZYOEyJcrBF1FCKN27ZD3w8G9
ZKssxom04XgVXaK5PkyJXIu6ACQiVu+cTT8p5PEJIBSrL9zz5tGX3sYMoOMlvzIB
dE5U6YbfCoPjy1DJyj8Mla/TLOgXgtfYO8SZ1cZzK6+crkl2dJ5XvvHkAcKrb483
Hhf3Sy5eD81iFoN7jHsTpriv1RiA/PjDCH2dA3g8hZ//tzuXucqxXB8Zrr7qKaFO
GKjVlJpqllRnSuEsPtrIAUx4+CgtfFrVZPAxuP5gA3dFkXm6naWeSxwD2igsCq3x
cAftHQSp9X6AiwYLCMayksFyb+NoIQwhY3cb/I44ovK0QtJ1xKsyOmLku0U0NdTq
8vEDctuJkcFSdEkq7mbJABvTYqlPa5KZQksnk2s132/gZDT4a9XO19UKzmN5YxQm
iVK0AAjfcG4nTq71Ta5iYFP4RzXdUSBrBMJPm0tI1YKLWWMN1AUDJfWeeo6L5sNu
V/rvkF+luyzRv2SMsdNNpjpmn8cBJ73o3/K+3uF6QiP4IMPJ5U9leVrIPNYv3fj4
5X+cvv99EhSFbMJX/cmyVAFtKBA0KfrWKQAcf5aebTXbMv9a6z8DLBp69V8pfjF3
6e2+QFwfJfAxfzAg27Q6BxPy1OHWPLwqSu2fTg4kbi1rcJ5hA0tOfvTJsg2OOmY7
r09TOv9Hqu+MH0Y7tFsFc8LsJPOeYTXa05nIQiSR2ioyCcLu24/frfY5IPLtrwk8
IB1H2KHSY/Vx4M6qalP5aNL/PFxNc8UvmjPh039r27041v5CyX6vrsAkDICzbW1t
a+aDVi/ImLglJRMDBuKuTeMLpQZICbE+m53Dsq1U117Krq26VWmoA2j4Y7rZdLWk
64KAJ/fYOGsBf3yPpt2AY06mOukJWxbC7TbIw4oC6eRfi25xUgWpRnuH/nq9gdoR
B1G2tNVC/C/ObO98nMbpUfNWBh5PL54hAu8rKmv+NNZac5nTNBK2pYQ39PMuFkFw
KipSjyqnsQ5qP3LzqunQ13oTYeaSe/A+2ybP6l8aLbaTRcSJ7nePhpmw1tSy6fZH
Cf1Lipm8nDZkV4V4EBz0WR2ac2R3tkSbtAVBqJ/dEsHV8baELCA6b5K/SNINz4sM
2elDN4Qd6sT9v1UleU78FPu/5rc2ehi4fxDZTj/dSJTbQnQDDaRazcd2kMa8pYwJ
ynhylafZGRigSkIKJwWoV69gsiUTFoec1W7IcU3e6Vl8sW4aSmuRQM5u1SeZkFH6
y8qY3DFrKJqSIdJNKkY6njRZW2o/ycHpJ/76gqrL07jkEZD22SCfAb4c5hwQ9s8D
2eogAFfwF0R0JqBHqIPr8bfsAAaNaURbJqOH8WsEWAzwBuITaWV505HThHOZgGGn
CY7CpZLhsjaEIh8ooM8GLmf1UkuxZ8Nv9zZ64sgcaBcJB5UUATeHCte6MwZGIG0x
Lvz3bvheLiqREYgJ+Sm729YSnHh9zfmhhUQyYIMZctEPcSXx0C/trNCffhrhe0Ig
NLdDUqPfXfpxL7uIKU90uRx1zofrXIYUvdQxhSLLB2l5r68hfCZ/Wdvs9eFhQT1o
YyvlvlUUHYL3f+S+cgo1itotcGLsp+BmxPHkHp0+33oHnMLdjgk7B34eP/7cqlFy
fMlymbBmLoaYGxuUxzQ5pcc3lMWsgQ9cIuIFUBk+32OKen+u4Nucps+b/B+IeUpE
GNkcWUiaoDzVTwxJyB3fjreql0+DsevfCcrRgJ5kDTsnpaYFFeN6QtPJw0DAEv+S
350wWc+aUZBQuGmtxS/2ZMS7A4SXTp+0EKcF9mhC2/bw4lmvbVrOaaHlfSvgiCaS
C1vonDN+vBzmeYz7ffrlsysFkZp5XMheEiHzfKNpLF+NsriC+s9Beiw2pYzqWNoR
Xy0h3KdN73JjqB9iDqame4IcmJ98NRGyZ+zadJCT/8tY0uIqcIPeuL+xOtHvNzCZ
LS2knkm8NcwuiHpKs3CK5nq+UFx0sZ+QHtYeLJuP1U/f/9B092cyDJOSSL0yEYY0
6MjB/+QFbv1lOPpOYnP3/CVSmp/8UxtGyTwp0eS27quqZz8WCJ7TSishIeYq5vuZ
Oe67AMS6S1ZBfzJub2/YVQreAVxksGH3xUrhXqUpZ1ETgxAPTnuBwkx5I0VpWFYs
kU8P3kTuJ4IMBlRKoB16cLTHLJ0TRIkfoTTIPRJS5HZY4e9q4FHY3JgkkV8rp/B4
o5Z0zO+V6PfKFYfHHfwLSNjGIQr6rmCUGHsfX3fQ15T8tv9uxwMSbDO8DN3IZIu7
X35Ow6XrpAdwZy0Ex6mMdWceNVmFoFPL9x2RDLRN//v3DuNVGDc3kMzCX6h69Asa
PqjE1erTpMumUwziG79/2ZDKnG+OiQq2/N/u9RUNbnFCz/L7/wJNSBl3MBFxy5BL
CGrt8eblVPEoxUGjHfNg7YoHjMZy9uNCg57SSebUwc0KbKeVSfvhHzvovKEIR2vH
GoKr8Z2/YzzACEf/nY/wuTr2hI6DcuQYL0gBveDOKFMLOjfFowsKECmQmLAtN9C8
SVUOMU3x2GeSXvpnHoVJi9aRTWFd/gPB3TS+0TTS06aesLDHk7zyuOvQZl8eDik6
M9onVNhCuzSjcHOSTJQeUSwLB2HwMa+TY7an+7pRcucRU/3297fUnrktU7PuF+a8
0FEuTyCpEfPYIG3+rb2B6Vh7ws62A56Lr1+Img4B4SQhppDcq9MtH9hHm/V3QtzH
l0BpDoudL+ZJtWLFWKXYpZUKaUOr29L9jdBfmFCQPOSgNDhm7B2SHFTWfarSS9F4
EHzLFEaZefdLcjqkMa4aZ720tBXUuwJoV/eUlUoHEQnYSf18CCHnQxw67B5O11fV
ayjPn0hqgoUpktlwaGQ16+QmbqMmIDL0CfEb3MbQbBeyy0icQC41YPibTbhapcy3
tbQjqnGVMYSIMgeMY0zbABYd8acHgvGSdIJ1PSLXNn2GceLh2apnXmRJ615G48tp
NU3ajCjeoS97UblbyXCj9Tawy1UgD2dfpJmlTwP6sihNo+zJr4K0WwK8u6sjgbLI
kam/ShCPuySSdZ2HKv/Gs0pYyeOIQ7yI7oYf0k1wrCuI99Y8EjDnRwQlKxgpi9hb
tnC4716rkax8F9XgiQNKHOgulgBLfuj3mRbHjkSh+yx/iuUSPT0sCkXI28nRzJzu
uIcHyt22ZoZPRyKkA6bsJpg/d2Yhz73N4+HjfcVpJkxoWvikK9xkHh7NIU7XL4ve
k2LzcruC7N4vWkomM5/E7NEo3ZiQFhtoez4dSEbLMsByJNG9N4QvneTOxx0WIBL6
5z747vl0xuM36YtZhKFlK9gkZIy3XBSPLOLdQi0lCleBUb2d7ohgARBMnZwVC4Uh
aLAdMxdmiKluPbfr2t1VukTuRCD1cKeGjtknVw3CtdGrozBdDkMrb8pUtpDUvZM7
o+kPE8kHsj+XoMEMr0tehGtQXIw+lwQepbyAmMe3EaJRt1ExO+Qn9OEOUYF1JvTm
HuUDAN4gNKLPVGEqNQe6b/F1QJFt440xD1Dr24FLXGTc9ogjE08qMeAYt/qHArS9
lA/atlf92LxsVq3Erz1KYKBRbKIJz3qgZn+GUU0GYure73DxEBV1Chp+tk7HuCIB
DYo45lQxd1jUnA67GU9q21VvrWTT2evfAmdZr2lPFx6EgtoFAD+5VHCm9JIrW3/H
lbw0E9XxyFazPiOUTITV6DRWOs3/VfnPxS7erX8MlKtVk1qsF7TZw60UDz++R8z9
6aOSbtUAXEcYWCr2RiNUpQwxyeCRAc1mIO37SvyvInIqIfWjPTJidi//VZm933fP
lkrFk4BmJprh0dQYGPYX1Ari86KBryadxlNq/3x1RC6nAH2N30yZwYXTKqwNM1Na
JQRDg6Qu+eX+80nZQQWuUIBPzW+R9/wsUrELtqZVcMKbf2NZQ0jegBJBISG3dAtm
fsYfo19VqMP9CQ3/6hSyBlKogJffsaeOQLimv79FllwcF/PZpaBMZgRZswXqQdRy
0i1bn9S1hFr2NvEQZREwgBRy4J7dwYtl9YCDUQT/NPFfRG/RUIGjtsiEsJ6iAWQq
WydGnCI89qN6Mn5lf+kghx01Zk20Q+efjF9O4bKI9BazYdqZK9kKthFiRIB7WRZx
+tnn1Zi/zcDj/3Q/+/weP/UV15N/owtbT5G/XwMZuVMfCntO4vSd8Q4bwGQWtvGu
pPhTi3GTN0/pyy7pQZGABC9p1yf4ua2vSe0DiNpwhJacLZX0hKb+GqU5aK6+UYKp
rXA5x1uYVme9tD0ylxzM66s5BduhyYF6ad1SHy2rjttwZqAYueXnzy0s4dUyMBdB
lvrD8uiF0SlaMkZgrVRk0oTT3RsOTdjwMKfsk4xJb4xWE2uaEWq5AaDrc9efzmQX
kyYuZS3WjWSNxw97Ux/osdhff0hYKK/94uyO9FmOtfp0/Q/9C3HetsJFSV5AtlGp
wbFUiJ9dXsVcPx0ROFeMoLMw5T3T4WimeyLF42jtfrC8Egn2LFrTORiSrzUQsYSs
pXAUbDsRDJwPueY4GA2l7ledVQMhZXSaKykWPfQpDMc5lolG/0riF4O/+mSgCz55
4+hjonQ2QE+GvxR2E412ko66Z/fQsxyUjRKAz2kdpVpPKfFNLGsGgRdS/EOPpFrC
EWl8K5+4CnyCVWEBOKA/kAftUljsO+IcCpRUPWcPgTXj9P+h5HwWJ1QLBThGqpMy
0fjA+/NAzctVJO8JKUXmDwjOqFWyHfokoa1twWDXzR+Si1u8g6Pt4HChEyP+3693
Nu9XGidYHQsA7YOh0OSYVlN/+N//scpBCBvveit18LAwdDxQRBs/l3AJLfFbPaZW
gJKqUbxN0x+WsGx8Bd/OGN1OR21QWkNmxgNGi4FykuTcrl0p3Oa6an0pjbuYzUfU
R1ylRmKz5efTiOesOvIz/H8aKPu2QlGDbb7OE/Ga4zNWOD4OBraAW4A7HKWq9VMh
vOcChsYH0FIBHvTI/1ZHiO9kdEEaTyCD1y8m5gUnQBAKhzgwjULEOeONiVmMqsNL
txzkUF3ekxmz8yhuWedYmijttYihzIpNe5qaVpRjJ9qprUEECJPxiJQnf8wZKX0C
8UNVQwJSSmxxWDeyxSos8rUK6Jt1epaUQbXRzmCsP8z+gUiFUPnkhcA0zPL8Bwhk
i51oaGc0yawpLinV7QYQW3HxkJby0FuCh7Vy4zU3E2vNcRm3+1AADCYiiwKHYdyP
VYTMLkgkPGu89g1mJGJUeSNYBx37Gc2LuZFGi+Dgwny6+lYJx+YZNQzy+lPBo1DM
M8HFbpLEe+ItbfuJaCbfLTZcJrSVppxTY2g5NvjveIcivcpvOyoLhm/JYa25rjCD
6vfWbk1NYb85hEnXGzKYMNWf8ay5hdken/OGYPdyY19SRaF2OIkuOLFuo6WJFTip
ZZWY2n6LyRGeK9V8nIQ+w8JWrTdy8IlK4AdpDUVeZajxR5lDh7EHR5wql/liSqzy
/PejhZM7z0qAuF0bFctIyDq/f2R6wHLtP7Cwt+Enbng37Hsg7Rsd2c3laGDFXYhL
W8VgD1U06xWd0Vk5sHMA3q4zCOOVBQDDiLqtmp0Dj5Xn4u5mfP5Y+gM4x42LQ6j/
PGymT8OQhxygE58t70CiGhvcOTqHDdsoltD9L+ZNRfkwS7LZ2PNRNqWtPZV29vki
PQ/uEiqCTqakjJUbI3Hkiu8Pm7EYk6j9S3ObI4dSTb2BpLMMrSDn0H8TemfLIDqK
q7Wvg2Po2p0oDnV8mQg9U9bUpmjvxX+0H2S6DjZ4WAU/ldPOIm+o0+kE//hP4TJT
5VAsPEYbdfeTU2vuSh1r1VP2eluSFUIbWlwzufLo5XOA6T/TTJIHsVqVkWg60Cim
tyis5rf9GEVmVSTzZNcbhkOF0MPFCcYxsRtHbTIIIJlp7hNH6OVfzpw2fElDnIC/
v6taUOjD3Bswh6SjnMIuuL1z2dWx3HryMELzNCZhdUEx+QyJPljjfk8ym8oPtEBU
RBnL0ZJzEURFhFQsra5m9L9wQe/ztLnULbkPRerWL4QoysJuphLAioPTFFv+LTGs
DqdecINbY28Q1PZt1WYESbLVask/g487F5Gybbvkfsl0J3N06gyI0jIXCw8NdstJ
DabtI4i+imUgCOf6CTcvF39sYwWXG1VGe31xMMpfk6AsC+wxB/g/MnAhw1VZmzJP
62sn00woXuA72txJgkD+iAVoG1w8Oui89Htevo+LqH2qheojC6dmcS/CzwLA/XGZ
KR3hk5owsqZJq0I1tHUHZBAF6NBbgIioSnBa6zUdtNtZ6VD4IKZTeH9DYttW/XUS
F9yqS2cHCCOmQwRZ7VcGHDsr0I/h06hIgIr11TNPZkvVnksv4NscErGjN+/qur0Y
DrGvapp2BfOb+QMNiOFKxeihO4+GNTI4SmhWoT4+JDv2yEyKzwwhAtlx91YT6tSU
wyVUS8gYPb9z1z8giVuBXQocnRpACRUWIBHKJJHudjIFtHyySCVlVhfWTZMkCufb
2VdWIkJqtWTDF2pvcYLUIVqRziUH8I+qiOvo7OtjzhJYOn7CiFfHFEoN2AGe8xEG
/sGeLoT4xqGE4/TOW44MAQKRzPM47N3tnez/QlY7P4n8IH2/9Etct5UDa7kbkTXJ
OMsb/cExYUeVbfNK62DAIgubAVAMK9Y0wb7N7xATFeNE7+F6/n//B+7OCSV3CjaG
6T6O2GdQQNrDgopLkuBgzP+p3goWVKUjEAxBs9xozb0kSXj5ldFSt0huWc8ALyjj
FG6oRw+2VUKTz3Q4kAqtmFtuerjQcgzHM0nUJmypQLyYwsBbZApLY6z3ybhsnlaC
YtmU8vwX5HT+JuIOTn5zEhZUsJpVGP36MSxlud1NvLVgj0fan673IjEhjha8IJPh
wCjH3ZLFVetPMfdVbKb++/3hoYhZOoLMtRjwrAwvrSHl46AQHUaMj0xi2xBZTmK/
J/UFiBKgEGZgmyxjo/PU7TtGATZSyUzdmMRfb6L4iRWqcS2TF5R1+iNOwSfi+jjz
O7dso4DQBc4kmnAvK7x8FvkCTqqrdqWqOh5mK9kdV2f+fNV8cKHEA2hSeCRLcWQv
QJ9ZlvayhZXko8aDASp+G4ZgkrgNCLafjTIsj7iagxSEV2ZtPqbOA9Gzl4OLUUF7
wQuK74oCwArRokoXHLoFFoBGx5fECwAWAUI98H78LO+eWINMGbqmxEuEWQRXKYqK
XOxX/iCtVDlsHIeZpqRkbhWwAh6va9udVOvoGrgL4TNIiBxpjPcIN/BjNjLNJTCP
cPTl4QknI6biVOsCc4CZIwluCyraWpqlskXB0Lrq3EQ5F6OChl7yh88niOvOldd/
euW+lHke4h6WZkkCsHEs6BuOx6Uz2wpgoby4yzwvI8hcr8xi0x7gBMfh5aBgs7/+
jzmUC6jZ61xk9naktQ4PILbWoZRJbMHDeuG4sL9cDAyyJoshQVczpy0Lk6Ph6u0T
rQT6Xn0/q89t07b6530T6vlL7i1bDbl6amO2TIjqMPdswKNo+dC0FLvuhJmSFTFT
DO6M3+624M7V1CRO9HWrw5FeTaD11keBTeww9JZUrLlRygp87KV6Ugu5wJ93CG5Z
MZvMQEGzX8ghyUt3rGM+z/LRDDEw+i/XG9Zc8jrcSt68XlK186UMGWawb3j3l3Ph
lFBIQEGX/r8FGDLrqA5879yhc+LctW2PHK1BfIhi70TLp0v77tsxO9C1RnequfND
el1bJX/Z5+nLr7BQIc55geLgfI4OuagxsqyXxqZyBpfYZxxMAExH46LTHp0TjYyz
dTdSwTmcJNueHnnnjbGyCETlUoX2p3SFX/PgvcWxHQKM9/KO5/dheRPQxnIXKeLw
RsktLznm1sYBl4w4t/Yvg1QRY4JkF64xnNNqHufFncfzY6MX+8slPDIC9bHbKz7g
vzbntJ3F3PRE04Ule8ILsMraE/UKWeuwI+DIaYOUbMPaVBjqiF5Dsz8b8oAbpXUE
0AvgXdOQQXmuXcBmy7Zbwzm1KNFJAG3PYovcO0f9o6nfF6DjTv7lVcdCAyiVCG3P
ahLwdSd6NPtmk/6/2cIJi6jr4BZzZ0vj+nZwi29T0uYAEh0PkMjO5LY0kpAS2LJl
jVjPCNZl9NkqX/P2d5lQI4jy5qVBJkfR+wKWQEXjmljZzEYxfYOiHURy/vyLpeWH
+tLNy8ccDXThExTXIbTf0twBf8oA8eQfKGT/6DADMG1gAJ71xPAmg37GI6H8x9A8
ZOpTH6XkOtu/s87wnDMiLET/drczjbFV/LlxSMDrfOXe4C3UHjIwSmFD8h2lBW92
US2MNGwxQCe93lSNZNNfMmBETvQff/M9i8Jp4cjNXQJE/y8dc4SiaKd0YbjuphgF
FkCIsQmPrWAJm3V/jmH/PBwuEqvJFNEFv2ap2q/RU3dUUkASGBc/8EmHmff08QnL
dKzMHsP/xWTqJXLWN/VpYwAEDJbHYk5MVC2qWYZ+uiyPJZ4W6O+cXJXNG5bYhxup
IcDuCCS6/DXB7ShyC4Bv0QrscpE3YJm5rVdz2iDJMRmmiaK1lZQWp8PzcKp/IWaL
3XO4avikAW/nZIZoSVsDJFzie+B6mEPzixf17rVgG/CmLs8bs1CPpwHbQvj9Geht
fFJ48l95c0UDNP6m3UuiZiOn3eGlb+62vZEv6abgykhXQciTfWE7Emur3gRJFWN9
XgO2TpgyNhLSNhIGzQC7yDGmiY+G945nYW3xOjkrscJuy1/gTzYM9e8qDzQ5I41Q
3b/g4W96Qr+XZ/9G0cK/9ZNTxItwwjzTuTzkNwHIrbH179fbnDURswoiWiIJxn5J
5kuadL82lWvGHOBcrsiX0aCdt/larfUsCx/MqQTHpJRGwLIFiIPHknvSMGF1waCD
AVNhvi38O0tDNCRMWRIK/iJxlO4W77t6SvxT3ZYZVFizwADTu/0ARZWZs2vzYec4
Bjsc+GRKFHlBPdjMZtYPapMxKsLa1wnrVOXq781ME2Z94UQ7bmIBDe4glt7L7ZUm
bQVbdabDVYY0QuThV364cfjmx4Q2Ad51RqwRKozAIx30KjRNhXyuBS4ZFr85S9L8
LSErjgKAAmqGWDHvikeH1GHQY4U2J3IQr8tN79PjQVQw9fNCgAg+Rp/y33Pfpx12
CqKEZkXoOoebzoleY0a7qwqPINg9H6XMoBP6hTK1ptbp2NNFEP8fpaTc2NiwJeXz
673P5Y/Vc3WheB2kWyr/KBf3ZTPUC7yik2upairqe5SvKrNA7UgdZhZsiUPG2ZGt
vG6mIz/5TQ9aa/0L6WBx3vUXIPV1DpJLCLSAuL9ZbxxgJ7vsbvDV+W9zo3whthqM
TmM/XftfJ++U+K49ytMYYjw/53LrCpqGeOeteekV1BLv9pjZahFZZNKrjPdDVRnP
5RBANk2hHAE+RP+BEiN/N7IIiO53q5vyY0S5vlQLLRJWtZeKhV4ETya0lNPrhDLi
JhtTjfOotVdlVh1MI8Qxsw3JT3VwoSkhPrlP9fZtk8ykcPkXDqelQ3mxWk6xVUaD
u8WNnDVWwtri0wxxQtDXDJBo+kMHjzfVW2AAH4uz+kpOu02d2EMG/cu2x0Uyeoor
dnWpGPUYM4G4TSvEyNnJ6BHgzE7/UH9Q2CMMl7bhQik+M3FCp5/L9uC7wrnq2gzp
2Rhn9aJEw4unNoE9W7KFUjxsvhwKSfsZZ5k9sDcfS8p0YLEneDlW3Wh6/+OjgHM7
uNfdoLYBDCWX+JIDBR2o4iipiZnL3f230LGWDVCdLcrCyXtB+We7/7PZts6Q6f3w
kQI4o2E6C40hO0Y/EUxdsWIh6vK99PYntsBc7QmBpA9vX15Wt6iNWLPw26/WAh3V
HMXw9HzSoRxr8S5mQJ3X+3DDdnA/Rtve01ae7YVzrB7PXs+iG/6qD6qCmg+UG1tZ
XqNl/djEM6kJub2PhKQspnLMFOlniFKRPIlFg3ZH3nl/NvjgOOwpXB2PAGacQ8kl
x66/U9v/a08MHXBXMQQV5adVtLE/nKTBWLH4TKzGp7sndFq9qn5LVPwzVy/6MX1u
Fpt0NVmv/l7EZq9TQb4+EV/8RRWpCq/cxL2/IwmdLVTVl4yISZBL/zDYI/xwG/km
LCdGJmWZUVqUIFH1/Eo1SRI0riJCWrmDdX7hd61+5km5EnbHvDJpNc/UEAYnF395
chDflZXaWN5hwXJWYKjSAnDiy0moybi0H/4n6YSLu2lBYyULlxwWcsxYt30ruc64
Y+rIGJhfxfMB55wm/uewMRtb49mz0TdYTqvA99UCQKS/jvL0dCWEdzrCXgVxBX2X
+POlpcFxo4dLhLC0WYUQfqcxJQDyOV1oPiRq7RNDiNbNdPNRaPO89LmLumjlu0oQ
ApoPo5WrNnkuFcylPaOc0FuPROqe+KGtrrEAI1BtTQZoxGHf1UYntXaNaVpWza5f
peDmOrDTgx7APGKSylDrikIXT7oKytGyrt3mhsBNX/mwKwJ3ncQgi8PdnkMhoURl
PxcLGeRb1zomoUeNdQEKXHO3uNWbSjbnGL8qgqIBAPHxCHPetfXLNSq8t6CoduOb
t8khsL2r47/F+kQkTY6T1cg/6SOPsxA9PpphVXWtUv5ehpiuFiSu28FpwMOqfTqf
J7TqilxxPW9zk2wjHjkR6VisgdiQ2EDtdZxzLcEbi1O2Qt30LrvCjrMMvoBNAfQK
+MZAN4Q8oI4s0xKntM2Acu46kR+k7i0Kw/it5MPE4v+t2NTZFx4Xhs4UKP4/yS0+
4lmHyBIUEVHsXiEt+PQssaTsYxwYx4CB6QNZ95bpcPL/ZztZkYritsptWgE+s7v2
hRohkcM4HcPXglhYU4EI5mUIacYkuQvPH5nDE+FUK2Bvf1IZp2RQK4X8mTjPiZRw
0sUE7IDloRpDmT1Wrv8m9scXDtPGuKbpzlDSAjg0AUC0EVZSTdwwEWj5laaYX5Uf
Flz4uySk7gm2pQtCAdSlKuESpAj32C5iKyP+EpEBgpsP4n+ROivoVyZALTI8rSTV
5wSuhkuMQkXtPNPoqOsDW79EbtwA96hAXAiAn0R7KWaKgvOOUEYbNikAJKoRSDut
Rdcv4u7Q26T+qidLqj1N5W4IBr8tYDx6PUloqWsvor16+kqzhnU2H3mBVNIzfqkX
CYOPxYxDlSgkBbsUP3jPXrx1yEyBQWui/fCTcgqruHFf1VB++QYZvgpficESWKs4
cKZc9Ncmb+aeSjROkt6XR1imY0k2UgcgC/4MVzqsYhki4tcAd0uFGkc2qvoAhSGM
4zkHrShLVCLlLojZ4p6yaVVpSndBSNmo6niWklJy5KcZh267Dhhu2Cv+jwBzzh4W
M4EL8fUW1euZoqDTKMU17xwh36nHz9/gt0N4TEb3qQLsOyCnr/0debemyiqXIaUx
M+6d0MJOF5UynYuXWNukMH2iQZSPMP2kbCYdZ2yM5b3nDW7u63Xl3Rand0kOgNx2
zxtnQ/kQxo1WoPrt+kdbZ/7kyzsR2ewXavSDV++6yvcPpugnbqreyY97vIQQs2W1
OM6VW3pSeCq3o43n50Xpjvmas6lQpEVZFD1gvPjnUN+CTwRUTs59T8VmY0Oeu3od
4Kzg7VQK9OFq2aIxxN6cFYIZj8F0C9uh/TaRmGaIBUb+tRbbyzh501DRUter1fxU
Vjx533YDSpSm963jo8FKUsEfgTjvVomC8DVW6retPpabfqDo9OtWpMQTJsi14lFi
+uh2xpEktm+qemNSj09TDpXJro6coLkRd1svcnBpjEJE0BdXv7dnhXfFB3iv41iw
wlU2NHLYwPZgfr9MtW/MOROjmiur/qKSCsEc+kY/PfUQ084UkkH8kVjwLTjP+8KA
kOhoMWRxyUPu3jN20O7BDjvO1n4zhJAwrMKl+ZaPFE0z/VHCN5NvKEN8RoIpnvka
jInpx0BfATDO5BJoNtjuSmv7LvRmwrylxXEege/rJCAnx0JopHOzTVNjRv8jWNUh
MPn9baTgmgxjS0hYiHi6KteB3uyM1lJFRPyyw6bTJQrecETGRLbKoTEjaVsUTT05
6MBLUFcGtHOXyoddp6Xtq8d7m178m8ZlQmg2PRPLynLmmRkUaij+LhxSUE/f7rv6
h4k3ljMdRWGgRoLgn7RzMecQNXN1kh3vbHSKaj3XOOygDjfA8kOzG6VNTdPTDdCd
Et6Mj/Ma8cj+7c5URRnLWJaHvMeHFWUqyy/0ofQLjjWcL2fblSnv41Opf2ZiMObv
1ksBOCkcitiejF8fNxx7iS840C0ajSX5CiZRak+3+qVOHqXf2PzSFnnrYLW1nDd5
dS9YAf0NWDsumU8ua1OUuQzPq+lEndO9rEIQZzN1r4ryYWuK3ebB4pr34Xj+wKWe
LasaPC96uyTOg1fykvwYd3WMb5iPDHa+5fG7yXostID53xPJ4lFj20kU0bGXBCEh
OdCVYxolJm0rmVPhBg1uwed2cGxK11SqhGtTHogi82+lOwXGoj8obg7DIWLMnPKI
Iu6XnnoYPy7D+jls/f06DQnG4zX5SxmMsHbtMECKRlplMwl5p9KDBdaYOpvbu70T
F+4h9JZo7AvJae9zs1jxu8q6GrmXH6cQgcVRa4ynZ7VqsjkV4gkxoVo4TODA21H6
uw9cvDpqmFbr6+27noWoeY8SDTNu4CEeQx69KDLHQIXEVn2HEOzRSVCIbSXUmvfH
kQ15tZARSW2kQpK8tLLT8jZsySZnmWy0HG51e2cVCdqwpVfzfe1EMb0zVnSg1q31
Djd1qZYlb2Cn9ThAXOUvNGVzzjPlamOW2Zfv1Bpq6s+e62fnupemtgmfJLKk10g0
pd4ZLKiEak2+g7rxQ/A8Q02wO7RMsN+eZRhGDHbP+gf6ihz0PPvXpXsY4GgMBzHK
hC0Xr3hZC7DZ6TH1HVaV47PvWNOhNZ0z8dr6yy1F5Iq3dicw8MOmxse5E1cEGCom
OejHZtiwFuaHMmlM04pWL+FNzFHFyq37M4WcsfSW2Nbd7WfYcpD+uhlZuqFRVFX2
ohip1GaQap9z9XduoPXbjEWPPDyNEBxW7eGQkc/e2plHiNCgyTmV3nFjDyUinbn7
X0yoBd2lBUSVQPX0opYk4pGQ55VrPJgrK7+SJrvREL6ZU7s1mdxAoHnYWdOi19jr
MAzSp/q9vzGDAsXtuqubA1RIM9EDgpWd0BEBSGgNGuTzufjmgL1qBdqa15JNdgK0
VzljbxtX2bIkO0Np/r65n2v8EhbOK6YbdGS2J8iJGKXw23NO9eijfLdXEyHEd+fP
xpwpI89z45/3bp6Y7y02ymMTCCBpJxn6P5ramQSxsVlRrk2Gts0uF9zzzIzaSeSJ
xevsS5h757sU1im5eer1cp4mMvJJSlkezBTLiIrEfv5a74hzjShmVb/7K2MdYeQ+
QVmS3K9Efoo6g/z3CPXRmr+dROCq8HLvoqfUc8Nq2b4+rNehhdAtlMY4wi6K3tgR
4Z24pUcwBIAZAsYZZkxZoHUig+iGNmQRp+jmwiatRhf7ozg+GPLWeeonEBEJTc0x
H5jhBQeKmpsbAVGA0/bfX1+BaG4oiT7HkYc0Gx32tQPoMYOrGQLaT0WRGMsgxQOG
m2EljbsIxCum39Jb4iIZAhdDdUv5gtGrcfaRKNb3uvj2wM3C3E7Pt9N5esVfRgrB
kjlcPu0qy1Mu2q3ENtKz/s4Dt/cn0zvoEZNqxR+ZZGkgsph/yYd0IZCDVIGy/5n8
m7v5WN7hwrsCqCJ/uWSQ+trCwxyc9/0ko1NLO/s0qmPd6Lx+fgj5xKjcLjl7hgQk
GbpgLzawpM0GK7OEwgdFGO6ikR8RPEzy9RypkpRlx3y/L6OvlUUgnBssxMTKbY9X
kKV9oy3+R8fFp0xUypiUsCHjFg5+iD/QUQnFBbGkUKdyXWWmisgseEvFmWRPLkFK
CdBa+sCt6vkBxmoJ+fb+OoFfos+zWVN2ev0GkCABc5PFG+nAHbXBMh/TcFLSVO/r
Jz1LiaOxJaeSM14+Kt51sE17PNUfiP+lBcq3iFuyzY128GMb54NkLVw5Jah/l3Kj
lIllnSIoJTYdCbaCo+Iq9wLkqAKL3R2o532GFnoFzLHAxwDchw9Goj2USyaLQEB2
h1tlqChV74CTGByYfGBeyLr6LHeENlGYop7iQpliLv0n/4PGl/9btEuCNzFZhjAq
Nxg5sZ5lw2LNhH1PUHuW+2kSbjX4+Cl/z/boAUB0AjPALVaeRYyXlhu0vGSVA89n
cpH+t0kwjAz3SUioS2NP9FYc+Cp/4eIyQ07danARFWUgW3ZL9jwoLoVuORBp/Bpk
OhbNqSJj0XW+6UGeKFb+H/N+17iUR1HRzjcPO416qGijP9EiA3a44yCtDDMj77n7
zI/VtnlsTlta5jj0MtCR+Mwx7XOvcFcQlFxA/BOWlwH0pkNKUg41V4Rv2YO08ik2
LJaTT+vChoOWNxcjYUiRS7botoqIF+jnhZE4DpImjRme/mk/Uxc2ntEi7ZRqldh+
fzln6Qr7XlXPtKI4Km/EmUvDrFqY6YW4iAafLJ0uVH9U/99mzLOrM4kHXD8f0n+i
TXMKt3HGbaeeSOwAn3uEFN/Lrd8yroYSXSWFyBUTxk8lDrhXVg8BOQgwuQ2vKyRl
vW5HDm3m/c/7M4HvhKUlWgm7Dt1F7QggzFHL+9xBVhApOTMUMzjE783CtAH/D6aG
Dfx1ByrBObAykk0MLteiWHVDM5FvWOomBkabRSHshPL7FVbkrVwd5UJvsJiTdDKC
5JIJ1SvLDdW1bJDQBVuOipGNVeoiBu0KrvhPBF7qIVt+p+uXiM/rfzsazdly275d
cgjBrHUxYKfyWIe3o/v8sjcKmkv6/3ngW91dTU+uKexnrtknKd5xAa1GWOWUt4qL
sRCJRda5ofSrjEBN3CZen1D5bJBlYXhG307pyIV+Zy6NBh15qwIe1rrYRLaA4TKG
2Yr9tctcBzvirlwRZLUNYx74ZYf9NJFQb7cKY0s568pWPhlMVwvNuXzH1XC22rQw
PvH5DdyXXzYaqJxbmi2rdX7bCqMhBmUqfEBkeR+wWuBO//T4/NDZcYDE4276x13u
SIw5C4HmCos6tNoCdVHqqB9StlFc07T8OPMmVASWn0aJYe5MBnwWneGdjDAUq4BE
XNlQgkPeQyUWxuMues3iJVV2uzHs6CJbbYgPMuj0Sh1RgS/Oe9lEB94QSnQtxxBB
3GcYTZ4vt10jEmY3hWCfRFic0JbBsKVMXQehsqqdyDDJ7jV+IoMnOfGquwxVK4rR
2SXhJT3QJPA2CtBmWfqJmzcKLomIiMqxLgyAq63mDeZL6tGDcBLavCSya7A+1kma
Hsz1MgwNbnundTaPyyxDYWzb9aUAJhVXWH0rYZUh0i4N1sRTjPlbhrVpyqwLa6uH
ESY/2w7pdEhn+GJzj7Jn/70xYcgqSWBzCJ3fYbsmBZw25CSVs3wBBMCii7Qvd1Bz
NBEWrAQ8NnZdDwDSk09Ady4kfyokpHelBjqYx6/jaaa27nJ4fzXh343oVAZHNd2X
OdL3IefOSRLNddyq7lTdD+BBHCJvtmaEIqaNtD174Kcz8c9q+pKhnDc00dTGdDhE
8wWnTwPuK+3eUdECy/ubpv6KUqXZj0R/SN1NMFbZ5v5RqG28xvVqrJUhB92UQ7zJ
mtfO23UFZsmrfApc2VpCk3t8jOK5rG9dxzOq58fRbFzd8EuPUgGKaNlKy5B5DS4p
/tKtofTW1l4vturCtXy5qTS+K0zGsCrKO2UYCpiC+ykPSAPJSASNqawZb4MJO+o2
pd9EkjWL+yYZebccLpAurHxCGJizpQ7ZoCSN0kOWA5Xj3S6L8rmQnYVCJnmeUeSy
T4VT/nfVTnd4xXLTjbojLCkZUS30Pjycsajns1NsHEv61Nup4udFmJMB9lITNcqC
qz7lMYX2grpK2aaPHhdPtfhCGQIs1cReNBetIG6Ep49Wt8A3OeNT8ZwZGmDDLAKt
kNoLEp6G4v91m4qQw7+1ubcpxdYuNJuOROevjcZnVvs2S7fBSoWVGUA5S+tBZxcQ
iNgVqiXM8kvGLvAKyBRzfM2A2cSeGkbpzr7MwLHUQAkOku1bjeBJVQqPt7+tVfmw
f9+/BGKxzONEnJb/+9n0V3dlIN09ed+gZNPzlGVavSE4QQhsrHMqJ3Uz0NYPF6nC
k1l8+fhkJIXpfCBGqO8OOc6nji6o/r2hPmfQVDjMwqW3FqYql6kwQTVAWyHb3PhT
rE8BWaeQdDqKFIJ0lhpvQyRJCuGddNdBUsvls9AfhuPQ1qhoVuQBe1gC/hsZSVsi
7hHaW8aaOrL/mMqzjMrTVuWblFoyimGAizats00CiCD+I+Mjq3hw9UI7NT+2rMqU
tyvrCnJ0XrzPdiRyiovOdcRowJL0LMWti0YI01npf3KPhnB/Z2LPTiKS97VXilLK
m5DZpw/2pUGy2mKlPHfJO+tqr11vw16O15iVCK7rbw7cxlj3Eu0aoS9yjvLsVGG3
00CepHdnUaA17oQsuXgsIrCBAiTNkukJC8YfCcxD8e5iStQWj5mj4oEl3nESzw0b
wVBEGsHwLyd34mIdmJ6BYXM494oIBDNMsbXzeaCS7K2kjTIeSjFvezBrrUtLfevC
5VHK1P1+F7+XaL4dF1AtkTPAgLgPA7MAngCTjH8CR6TZXyMZx0TPKme8MMiZ71mD
+zPbTXW0rltn9jnOG6/vWf3TjUKZxZ+SfAL0Yu3npQkP8k1NbmQE8HfyLBo3Qs2v
vlAof/YfOEP2QuQNUet6IvrcFvFLDDr7Ljum8+iex7sBPAKDm7hZ+eH5rcj/0RE0
AJy0JTuhzMhB45Vju662K94wmsGGTSjEx3rRVByqQLBCZuMjcQpetB1at6PWRmWz
HjOhWl9o192J4QlCkdEg5YHEXNROY4oCBYEfxWr8zALzQu0vrzo8OhFdCubDdbMj
u7EZmoyO6gaurzD3CIs0ygbdJkGh+rSAcCWFHSl6SBgE93Cqyvy36kGnyPFBXFKf
+ksHR42r7F+l/QdLPHvm0uEv747OliG657UXuJ6fxyqQzYbzlKoCHS236sHeKwsu
imbZqy10lA9cZgu/+wRhlPTvz+J/VS5h7VAWkl6hTsaH4PSIiVkOFAr6gS4ObbUA
QJ1ps+Cvycgl7oALEphD0J5/IKlzjqZLs+X4fnSX6u1PGWiIwZ9B8Jkkx+3Gg902
eEnLaqfCh/CyJUZRZgydk2ueEla3bJlCKAO5ObRD3xcGw7WqMdKH+PlbC18Sv+/W
aZDk0Zotdi01cr3DnSmC2puWj0uKuH+KjThrgtftW7zImRyy0En3jvvHnaYPJibz
4FN8+uY7Yncoa7mhev+AseCO1W8r8Uswki4qeEEhNGOD6n1Zba7123ENbe2XD6Qu
5iHmVYB+2mB4rVNFCYbMsNW1WdbKGsK9BCw4e61i8E3EkUV0cp/tClYRu4oIer/J
iGoRFjZm0Sla6fqf0enPg3N+/8pulP5e7fH8rMWSCgfsGmW6q8KIKPCWr3HdqsfX
Q9x+8DGl/w5mCIFjEpWchwQH3Zzuco0SUu+roWD78m8ubAhA5MhbU4k4aHX62Hsk
OcH/SOglEUF0O9VTKRFRowPwJuEROpM6zW+6dbE+FKrNqhWZVazOTMiQOeo+n5bn
TPiMB4nK3HdFKgkT2FNNbL0U7+R8uiSJk5WdWusAZWzS/yFjWhLPyTb0K1TL5yO4
29hviUYJghA0aMn5OApCOOoy9egIEoi8SZFgxRHe6HAI3VJE615nk5HWZhOF93vp
D1p3lFLIIFsQEdRihA6Al3D4E7tWuDkZKGR/VACQOEwiQ0Rn5Q4foMk2X8fwvajI
VA/XSD22Tk8EJXz7pxgLW2Cfo0S4G4RMYXepT4CW8NF+Un3VDXV093hNj9C4bKvi
nwf0Kb7CO8IKT+bvHxpE3YrMBqQUKgGTktIWR99UjcQmwt/bzUsuMO8kO7HmAoQt
G+ibk+zAxCojl5JgTWFTHz4NKiZ0Lt5SFHH7rJKZFwCkvJvmgVuf90eEfDbMb9ZH
pwExzDRysfnnrkKozD6PUHWaCFzAKb4fbYo/GqvaEJ8OMUHmU+j4lh+qoZsh2uWx
i0tOLbG3RJ2ntjG5vUWm6cW+7hzPdQf+Pm0cqhaGk8eJaKAhEtZLxlOeEMU5sULl
o/4tmeym+yz//Pv8QHt4sBqXyi0Pslt1MJsG+0nLoVZvUG9OMpsmEfaRiUXSeK8D
fI8KthjTJCcJF275QiWz8/X55ixtiZhtRRzNul7+GNOgS44PUEaZwLla3zr0XUNy
0gAjzq+/EQb0ksZBb9j4yhGii5W+rIAOaX9/zKhVn32bbLW/ubjqPQ4e/CKBhZYn
J4NIqjGdmg60NgZF/8vO9gTC0m2zKveajT4dNKXw5Hp+MOsCc9ahUYWHigiQOUy9
nBJas2sbCFAYwIGEhKZ4M7gIaGDfUTDnD9if1cqGsQt1OWDeMSHLND+Qvl+gExZS
DHxV4MH+cpcNB2vvDL2lrz3N3bYwmeWYcv79lE59hzUWz4pl2Ej2tBC2TC8XI6TD
yb+y58tyRDrbaJLMy9EvhNO96oNNCYzjDg4sIXbs9+ro/3Hb4yBUI7JuKf1Y/slj
L3Vymw+uUbM9pZ8VmVAL9YpjdHJtFdMe/tw3vR+YVZWdQ155CgXjIR19GgUWEVTM
1OcrAZNC/Xvd3nbo9X2xkC3oIZtNJr/0FWbR7j7CFsKzw6baNmaxlU3w4mDNPL8n
qKLJ15BhkNpIhb6wNcHm2dPfQMj3k15Hgr4Anszgg7BrI/1PTpyrwxiFEYhWR9YX
vF10b87XaSpqgQxb6X+fv9m94kTM2ooL5aBgv+/oOEMtEsQQgXfQ2cyrUBoXQdNO
cLngBpScCaDmYzfUWeck2oWNRaAk/VnZvU5Db6TykIOSwEXn93zhy6e8c8tUmwMT
Z0oV1FvKq5ae4evmRgfHbPPy5aVoRcGpWEl4qYJOcbzxn+qwuAnX0SJpQlNpQbr4
GzlvbcMlGYFHDUZDJULfbyyu6Z3eP45Ibf+G+OOnYiXJ3e5ERAErbPQr1IdLfMZn
mnXcwf102yQ7xb7m5excfi4P93wsD28AOCVzGh3NUD+izWcJU/Xx0wePMfNkNfht
rStqAp+TMdujsDBArHBI+fjsq1k5GAaDLtPcY2Vc/gE3LNPYaKpUdoQoiWO+5CrU
9mR3FglJhwBDPqGJRyXqgjUi8qfrbSYlyFOmug60pk+SrefF/+yzow1104dC4CSl
74CrH8mlf/EB8jt5/XCKzl7Qe7Urfz9C8sa6b/Zz2CKQxGZ066ADO3BcY+JgEiij
D5FVVZB2IwUx8pcZnXjBTyoVeFrKEroa5FdBDiokUO9GJeAgLbt34I3v6PFLQuN+
8DtMMbm7/t2SG+ApEddFhkql89xLE7Y5BfnKO+v9hq+yEbVh9bPU6w0V3mCwmExm
Py5xP/klRxtec25yjetBB+rvRBqoBmGv2PF0HSTA3GVepTkhgI5UMAtuBTkSBTdV
iIPeVoFQsA30hxsdORcotjbcVgxPmtBy7uJ8Lt2V0WHmbbLF5B2WsVvntJj9dCaU
evqJlPZkadLoLYPki3zzR/w3HGGC05hGApKEUOEXfGF8ibbii1EQQ28dLafOqgsF
9v2oy6IKHKsugVGPz8hFybGMSGUh14GC9lMQOxbYK+KC2v+33mNbOVgQA8/QLXR1
oVUV39BppVSpEfLtyINvfHWphrPvqF+hrp8RtcYUl7cGJUo6w9Y82lFpm6Yjb8VJ
0Awf1pTm0oUB5e8FmzZbYx15nsIroG6earrJ/o9hmg9uCfKBreKQ0NX+3UqXaXmt
Vnpwdw8AzVQfa+K5oglLvgufQEmF8ToOjYBoFTnQEzOxNIvRCbVLvonTpxhBSKS9
vEz/ft4jM/QUN0znsk3rhARECShANuYSYmL1mFT06ZzQ/ZI6qeyjB5TYO+/vOQVP
rNe62w7b2YXR/zXU9E6BI48wclSjnEoaU7lcum9ZUnsMgIbleptsZ4+UzSBS0WRI
izT6Jj8ZXf8KGTyT4WoU7Zq24GPhwOSuXu9q8u0FLIK1HpKEJtf4FKXByS8G6IgY
3dVzSNBKXZhsCGFsX9RB/oaX6xdk/K1IIjzS9hC3/uFi6YJGhvzv+He2lkkUT3+i
ILi72HrEc1wtJPJStONvoA80RUCfh6GaAXBzvn8E/1RKoAo+M4qCY6HDfLyxluyj
kaS5AiUz37lXEhy+Zf8Rkcf0/JHnFgRUx74dHctqJw8s0mrDC41Qscq+AYXx6wnL
yJlG3fXDZEIiB1sdQ3FBmNE2823Y4hYSJ+E/ljp14hRFkTBp0tZQXU9bVzSrPbze
XEbmpEU/zQTXAJ1//igacOOaMhD64lLn5THydeQ6EUNO/lfdILu4LRJYQRMRSSMa
iYIiNrwvA+0UVx2alO1yC/rIg0mB5GDCMN4lam5wdUAuvxYL8ro7749OKlLxduM6
nhf1SSMcaVxItZaXqj2S0EphNw6USs85JZZA/aL/AL+E0upO8xyag7NTp0HkoAGx
Bve3K8ZTIk3Biij7nXr3IFH5x0bB+Sv4rZdMOrsyOVM+bi0/Og8XvOVLnXyIYeBg
nzcv1NjbdxCizfvzlekiJncTCaYyeMRfq9FJBAVP/9912pLjRdManeOVxvq72DcJ
/sOq1++jx6K1ddg5ISilEpPGzzNhQeNpdfDjDEjJieSOnlT7FxhzBnkFzk44JhMO
1pVODDqSE//QQIk4GuMSE7rtDbs5mrLJKen2vnnZXLFKwOXWz6kUffC/Xs2LI9I8
sUAnsEOkX6WSGi55aoFBbRj+/aN9+UGeMD4utVw2XpD7NwC/cH8eOE38b8OHuoSD
c2A9k2aXmA6jDQaEZYs3Zamungj0rFUMtwbpkc/rWR/CRyXIovjT6E4+Y1rmDB+7
Eb+isAJcCQ+ThPQkFBLgcA7R5lPzqFROwekXyuqB5+Vmj0UEo9+naY/5vHEfnCQe
sMzMMqyIqx/L8hVDJITGLhUxwollNpMlnz6f/PhOD+/fYuTtqy3dgBAJUzkyYq8Q
hNPTMRlkpEa6WSgX75U8VyV3QGn4cbYPihU203WNQc5g+ob87BOqWhgmgi6s5Ukv
n9ZjJP3OJk/KFqxu3SKynHey9JX3pE5M8WBikxfghm0LZ9q0bQMDtfonbVIg77GF
0bqclqWhmv9QwI/B1g/zuBTkjhW1tyXaTe2SLfcap6UeWhI1Odw3MGwRZ5tbTGpZ
x9suXJ8PsuaNieUcaCn4T/DpCCV3K6QC31A+g1guAqW9CM7eiFWZc00pmdrj15gQ
4gQdJiXlhrbMWNsSGTfVw+j2rXTL5+ucCl6f6ORpNMkAblNN7TwGeQV2uvP3e6l6
wRPRdMz+SRu0kl2fFrs9Ut0h9nPD1pykOA7yFeaGjN26Na3lo0WD1/54P2ioVeA5
QzU8z+eFpkz/YagSHsaBT+wvrMG4oDouKzd86/plk9JLso0B+Nm1v/mItjqEfLoP
YfcwoeF5/Zl+xQ6l5aeu9VOjnWkgECLjpJvOmiykmp3Jxy5DsBOsDGlGwuUBJB7t
yPgoas56wvzMDLgJ3QTvREZcUxe4iYvVZf4NFf4oi/ZcnaewQj28uixcN3ACZ/wZ
IMgr4Sh2k4JFlmvJpzd7Fg0Rv5RHyM5QRBJ9Y+wmVxc/QY5NDADnprMZVxdYUyvq
947rDXovsQqK1Ac1qt35zqNs/tu7dtF4lUXIxszKQMvV2aYlSMu9ljiYrawTzv8/
BEG8qFAWDTzuiJr76sPtQGsDIX2mNNQfvwGqM+64f3MEcJJBnAGzXQbwRKJ8aO5W
ZJArJiaTQRI4ISuThy/62PUMPpXr/RBMvdv1ddVpce552LA28XyuD0c9Vg67W7Ry
Ld9xMkP5GXBlRPcfcrhCuguaImj+QHZpRzU4KBnpNq153jGQ71sDYlmNXqQrD3qS
UVWTofmi2WLm//UUE+3YknNLcLJqoxACqR4GktQR9WdUtKKEuhr1Os6n8eBt/jm9
lj67Ko0QzzeQo9KxcBAkZveP+1auG0NX7qVovLB6VQOkayPJyaMZLuqr2yRmKybB
Pln5yKuVOu3+l9DAVvhGaQqeCnjzrf9vGvDB99N7xnKob6bgj15MeisKs1tpqXTC
CAdo9rQOYvzMijDAevMomi3doomDsB9duI50THb+YB7sNh0Z4k07ZYNeGMmwEEtg
DXwhYdZiv0Ct825/7qWKf1mvwNAC+uq3iHooN0+X/3Ipa+ySv0juo9vjxgSV3dKl
AFSsZcv5uY+LJFLlJnaV4LqZc3E/3tqflGhpKntM6RLnoQalr1RUmSRc2um88tf1
lTbIeoZDhM7tsuVp+CsOYXEBe1epV9uuaTpx5Bs8YhuB/w0k3uF6DPW8zDTN9Cwq
GzwBAA+XgnlCht4Wclft4HDhpHBQeYRYXOqWb0GZ3AvUNdNwkrnwkF2ZBa2gCtMF
PFlkhDSrZTq87dImQtvZUA==
`pragma protect end_protected
