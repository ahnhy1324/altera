// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
XEyRqPr59xETBsbsnQbrATBIoGAeAUUZjixyFTE4sqs2pQ8eeIvVZIGt0MZsUNr5aLs52kI/b3Y0
wt9fd2OaOy6qof+lkEeibJgNkEnfwghp7etJCILp+oyE2Izz7AeankWq5iHXd1W2zK+pq3h2iKxh
gtfToe2lPc/vpaQ66V/vcs6gIDRBcS0oOROv2Lk3cbohby5pj43csWmulq5iEA4yGprS4EckJ7Bm
+5KEHDI9z1YpEj4PJkce5IzdbsunawLJZhqbTcYkStTK2o05z+BBaZRWJ8pygAfogR5/Yta9RpdZ
hVqistABGW+Pk5Am2T9ZBY8ytD1nVt9H7DnBrg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
r/pqez53/4HAEdLxHv4ERYjwulCqx7avC+uDn6QHNIlNVsKofjRdfHS8rpHCEHmBa2RCLXX3COCZ
J2VYXEC/kpHILO8nl2qmPEFZpfA45Tdv0Q9BjGUVA29yHZ7J9Ull3BmMVb8C7HvwJqBXdmfmSb6F
OLb0c3hB/Fe5kw+jjwot88bvzRkwpHGoSgwfHUtCfzQNLgWEJhgzJPk0O2xMw+ZFYS7dkrewSI7+
Ed48K6+ecOzPyBm3C/oDUcndn6zyNV/jeSAXTb1aILnGB34Xer2NeICJFJG7mpE53s+/GNoIQxtl
MLt0sZ3kdMcQ807ULTaolKxf7JjoNIkq0uBzFOq+Vgev+zGUGI9C9cUcATYHJB9YSpVXhO9GRaj6
2Ozo7eHb56KrlCi416irg2TtDgaHvaFyGDUB4nAX9HnVYFATZHceM+CoMiv6o3ED0uq3YXsMo6cq
yQESFDxBzR9vLC89UFV6XfaLmjbR/ekw5IO+wfXQO3kf8TC9TvZiQFlQJyR3aqPaGyT5co0kkWMt
B/pz3B+3y9fTKOotzwPCC7DGN7Ug4aYj6WkcbTSrIqyy/1PJml/ENagVrkmeBEOAFxgZ2VByIixF
JYsLwmwNV50JgcUJw/xguVTh3bEo9pyv6k+ZrPdO2PNI63U7pJdrCkFDBo3KpXrBYCJFNPydguID
+jqoLWWX15Q6b+TUQrOojNgMjbAsPojYbcXv7IG8EAMvg4DzYq7Vb1vWEGDnzkrcP+kXvjp56PjQ
qY4WbmIGyL4N2ckBP/wHNEZtnbgHslV/ImECuumZlFbhFhB4/MZqN91H/R4N9ltXa7nFf0KTA/qV
3mYQor77k6lLglHmt6fixKRzjaGM/NSIGoNjetrZBdkI4ks48b3qvfuH8qjw1tu+2XDrypufme7+
nR479fzHW6chpH6IY1tk4N8wi9bU8oYAa9n5UZfts9bwhoy7ynowyKet8sG/+BBr3A0XFCY33N7Y
qKElzOzjHy+/OwZkQ/HHeFfvXY9CuTEjFngMyjGZWwVEEX7H/ZSTTL07otL4eBdM0y/bQ/YsRRHe
jSx4owRo2veKMBmw+HsgmZXAlrl6KDFK7xMkewhylZA4B5FP6Uogpq1rEaq9AZ84hKMbgbG0rem7
KBDwK/y16K3dT5jfOXgE31SmQJWxKoa0DaQqordYh8mhLLLzWk85LEiIVfidgOFEh6m43h4tIaIM
3V1oYUSsyY+SsZrPLCMkG3F3+DAbCcOpti7KTe1H02XQYila4OeCRZHWLhNMtQg2+cTEqx/qH6tP
ReT2RYXs+mj9IXevCM9JTdK8TjK9P1CXqCOlho+aICA9n931GHbMoil/lU86i30h8srZB3JGlnmZ
9nRFvpU8DsKH2TLmH6D+fPhhPS+MHejPI9WaxsW9Q+hIssFzSWHkVfQBS9SdZgGKTM5sm3TPk6mD
r7FqNVgYf/cnCreS2yQGXXLFFSs65AMiTNLLGIp47j9SXQm/1L8R5cm03bDvTRJ6uboInsuXoMiy
l08/7cGSdcK9IZCGoQ58D2h/PHrMblAfVWVysVRTB61z+IN+qBtYBCHKFDKjwaHOpvmhhk8UKmrh
7Es1H57cujV4LKT4wELGbfFBz4InUgxd5EmqeCUlc5juPkSd/XKXbDO9GkUiRHY1YxT2+mVpZ3Jg
dFUWpfiKjjeLYblcAzOV1Wmk2CuUV+2Y3fR50jr0RqbUIYmQrVPNFylFSmjK4SIKZrTjtdQphNgh
acpn18PQIbjH2EBa+n5RnCR0SbyveDNjH3oNfc2/X8iyxLZN+apKxbipxOWDNZb09Sh4N485O2Zu
fuSG4LDN3m8uoF1VO/3SuPcwQs11/rtqwGrrj2hB+OAJ7it/O8WBqfahAt9sZmgvpEhFyV+qxqOM
ZWhh02RKmz61J3BEZ5fl2pbF8u46FASFeJgjnt1k5Dniw1Sv29g7RtFYMQUdAhOzB+Zjw81CANDE
FIIs7evlPgmcJA2c39u9W0YlFK7t8lZLrcPzv2KvwGuNoVZ1G1/hs9ByBVG0EhxZ6o3J8GMoPVCv
nRwJdEiX5BvwF7sxQykv3H/UA4zABqYerPu/Kq+CErx+X8j+RZAMYi1pLYRovxPOjVxqzyGLStbA
KZWQ/FsM/Ue/WUaMlAK33D8QHj+DfBa0oEeQqbWy70yB73n0Yw1j4Zq/v7cAbOo5jJWgrLvTPcmC
wlhbfuV/SZhodh9tFQu8wwnGz24HrSy6hKjQmEQ6z/3kMndJ0R+O0ais+IzTBIB9sc2gFdbmzoI9
lpVIODCwZjO5pg5bgULpTZFf0VNmkdwLephhGEDjV7ToeCVFTNXQyfnAFH+KsbQDpI1gz8kJOlM+
guRMhCU+wZ+eXtno5iKXkLk6JxBv+0b8VTOYscAcvAHYtcWsPuY49TOssi7DZLZ5CtmqZpcDrheB
zWoraEzvQvCszzrxwezyOikJkjLuBVLeqkVf5/evG4sMGSEclHnzAG3qgaw93BKu9cltMpf0oFLl
5SqkKcRjNi5sIrTZ2+8DCBib50hTHy/ipIGrm/rxZbhd+lmlPNLJKdRWn0o0nuIkx9jYP/Oy6PYn
xMUqPpEtKFQJQBmSJwl+UkO4lvelyR2pbnV6yTwqcIZEMKlepVEYONljzqIRGYZRlyC7BrNVW2f+
Lv9LUhHWppAKd9QOseJgsQol8vueZqwifEnZld3kke+rPL9ivnjB3+BYyVl9+1x8FkZku/fAsvDg
ap3it9BNgvdItFcAP+3YvcSfSD7lPvX5i5lpbiEvVbgK7us55oNrOWCUR7STxudTz1aDkBvaYBXA
DZq+EaXqYEx8cDVSfrrp1nh/qU1oY4RaN9yawV8FM+ktgC41QSm6LoYVPJeas0KWKMTnis94ATjc
HPyb033se2L4hGfiPBkJJkN7noKhCGECwnfbgN9osu1WZDbxiwlWcj/RKW1Duver1vuhwvKDyR+B
7+iJMO9ql+Gs31JIcD5kuP+ASY8czw8lYCHdazKvAMh1ECHkx7Sgy7k7//Fz5tK46ypUhAB7OrCU
xTci4/Own/8DWKEx/MoABc8IVIzN3UXKOLrg/1vPWCA5CWp6xWAD7BadDTmC3zqxl0c9/VYruI1t
yDgHkIEQYr5ns54fRJEeP55bcw3R0t/qLhd9WQazIGqnRlIHmC+XoHx6qR5q92Z8HlZxaWeGgCed
tnTF5Goly5YRxX3QX7DpYSj8xTZdlLXRPQl957hKsll+iq6iWKclR1zfseEQ4ypPqZmjDzL4iACv
ObJ4Dul400JhzZlu1SMrvQ1sZOedSFODcAlAtll/yycVh1i8UW1ju6co6uRzNEcldSFiE1Ps66Wu
hdIpyX9DPPPUWD55cSLvVW/puEsvJsxGCi6aCODM5yxX2fVvPj4vWW+icgogL9IhieNmnMmRmDGt
y6ZmECV5TKOHJlIOTlPwmDpQx+uTR0eIZx8t4qsjAbpFCO7b1bEyd8yEihaZlp3MpFSsB/MQ1WBV
qfuj/hjAVdYCEn4WcE37AxyGPr8pHKOGL46Lf/4rCjicWLRIVhRf2vD7qdqLciP9ngUg0fHo1YIO
vwIg+vR4UgSMXg6DYVARFHYU4WkQIOmlSa+5tATtPPuerawjsoBl5CiG0ybmtF35GYlBE0xUGrJn
M8WAxzh7tHwb5pEN5Z66J4y/JaBq6yg3QSS7tWvVYvCuILN2c8171QMVdgF9KwO7fYVJRwTs4lU5
s9O6EIfJdpij3J90TIR0PkxecXnkOF8D+Fr2JpHzlFiTSqcWVssiLK1E/WZFvMVKiAOnBCa/+b9A
PPKgl+TSs7Oz2D8dklj49OHSA+DDv4eEZZvBDnu2k6xr0yLjATrIwd6GzrZs/8cqyXAlx4cwNpE8
2sfNtvqT+JputPo9Sh3skWJVIqiVU4QgfSfaFMfxI3DeRbMFkIfnuk9+kt88rslElHjcq7dsm4nm
5bsQvNRa1Mc29YWZv4Qv5Ql3SQb6kRX6aZJHpmsnbf1FMsWkMhLHqg3vuSHAI+th5oYVZMh4m/Wj
17AUpGKL9lZiuEYkFlL4WhRUGK72431IWvt/sR3Rs9q4kqxJDE1PJaxIOOcfA52VzflV49SldzQG
vpD4M4iizDxnOPXE8+V/r5onSA04kUMMlsUW//snfZwAuzPlbCcfF7O1GKh/8xjkb7rNBlDMTU4U
OegBAcPBWnYBXQv7PFs2gueOQ4vrGRlezvfG4f2r0OhKeyTyXB3iHo2ytSKcIiIDxlnfNSPIZnuI
6QIIH1qjYjfqX49EjTFsUzrXkTdptGJif/O66KI+zOlHMZldqrhghbQXuRcpzdsRfz3k0owe21NA
EoPsip+dSph8mw3w5Jio548pLf8FnaFPFCbvOvba+43ENg1tGA7yRb5mfCXIvjwXkxTkzGv4Ostr
DG7Ljh99ICQFbA+tXMMgzRHPdfcz0tE13k/TNDPuHH6VNZSvkdVobu2kMDxIPasNRQ3GOhNK2+gH
+RS8TBDH7A3Xt3iCUdq8d4g6fimW1m48nTK/JniGuw3/UwS2wBK13Wiw/oQBJvK2U8XKd2r8LXSa
VCtPcERZy++QNlqrUxwvyEQxZSaj4u80Q+YiV35o8ZpBeEQNCMVEP4dqHEpeZEn0WcTqH2g6y2ut
BeopT0G1kR60o3rFUhon0i6IeUreH1L3gg07mIyW9/KABMMUmDzzaN+OKquTjsN8yC8jMC69gBxe
FuNrn1DoocfhmKVHyOZrx+NzxXw4mqErJ6PIT3Me6pUo7fV279Oj5gShw/SqITSB7xBDuhVUyILl
k7xkpoNythD+XiHhDjQFhME9UL271RRFLxW2wPgUN1KkjWl5NHGuw1lzIKoIMD2ll987Mgg7FH+H
IcwCmQ47JVPurqNf4+OABH9mIQ/NoxEEU5pqFKl/YXzJt9MCqkqfvPGRb1mMU2xwJadnuVqQ3Ey/
D3Nv0YVuLqzA8a3VzMUc4wb72mH45jG4qPPB4IYm8m1xonR1lxIb38jcTfurQH9zgBLnqjVI/ia/
1+iIcGWBps1jhboXTSrZmezsVNhO90WXH2qojNWMl0impi5Qqals3wswiZ2XkhproLszt1USe4qT
2T6nbu8RnGHpC/P7gPhH4S6Aw4rU97sfGWOqMNBOVKgVraqC9xGHb6ifEsVOd7lhqAfLoh83yaxZ
0yEuF5mKKvS0YDYt3mauX/9IyxaXehbvTzmRDfyhCCErq/TvvyGFmVcvKMZZWq2/hH+1cGntnb7B
sXKUDqTEG2ujHxtol0LNzR+/xn5mOCbDGDHnfLVMNfgei3Tdp7M+9cQtEbFYIQIPO7uavDbc5vWL
XGlNCrpjbky8h+HHMUyUMIpFEO88b2egqZHvuIEFJV9Z6cDSHbRUZbVG1hsXsgAJfgD1V46Xd0g9
7nouViS1y7sYEdf8S1W2FpuUuJhmnj1TDVawf6sCmh12uT6m/JOT+JeaXVbro/ROIcmaqYulQzYB
loy3EfPvQBIHhOkQHAIl2PGCsTb77eXe5McVDzUtJheOQv2S+AZIVz4AMkO/2twf6DBCjSwuc+uD
SYEXoTdiP3JlkvycoDY/lTL2P2VRJSFLLQj9hAGzh4NP3HBZ91woDaESURZNhhAtGferzzwJKcGZ
m+n5VkFVK/qJ9//FWb+zPwFb+FVYBOVf1iSqywvm+ugC3H9dIWmc3xjEtyeK50egVrb7IzYzOpUg
zqFpFWf3ryY95SVJeujyeecZgLffUiflSTWGXM4i3YPDo+qKdnrpDNAL3/Sn7LxGjeYQWyy1aBy8
/CRnIWzJDsoviRS9HZo4GK1iJzU15leVobL4i4u2HvWOrtFgVTpDc+oIIFciy8i29bAmUH8z6cyj
BPIBS0+6i4DVbAjvJ+eY9mA/8SZ2VTFBTKjv2/osTRo5EgeJEe4U3qZoOMt9kSMtJk6me5X1hdbI
pnFw9hYZIEmtjWNsgUA5V9XYo2wiLkFhtlPvBy1kn/Xd0QASiQ9YnD3+DGDe4SylmkNljfK/VoN+
w//FEzt6RxwlnzHAxWRUQpLZRKmuvjAMwMVA83CJbqust218gxUDXkgTqbLN+yKtqq/U/I2jrDRY
3N8qqumEUZQk2BRqllcqhBUU+XyARB7ZqOnPFJwwUHQCFw3yB+xIysFmAf4kCkkhh1S1MMg291QA
rJdJVs9N7qZk7sTuH6PraxpoaPL+RxKtUHvk13HOWkgLt5R06xIIaFZy43gpjozNUOcWd0tTFRIw
14N+bWJ1HW1k+F9GCFgViB+9nQYS0ygcMECCLfjVeRUa6UPCliO4/wTRT7mVm95xYUNTcU2GG7MF
QnoJYqit9lrhcqzLrgrJBn3c2HL9noeZlAnNjqZZ6S3u5M/7PDKQMXs/jl1vPA0ImIU9Hiwj3v2g
xfUWbytzU6Gw3UauMw4Tkv8A7Lh1vLcRCTolsJ1lJCvKEIXx9kD4zBK9xEjIRYewr4uV9rW2gYFw
QJGdd4r8kaG9J9dNOarViGy/gQ3LAtK125Vb+c/mdafzQw3clfbSmPdPgfIgdHLGQMQ65ekejaQe
skENwZ7i4z3GLiQG4dlGcj1fa75+xB2jfBeyYXwFuyB3zFeR2XEzy7yqHuKe3W6XuHO7qIAP2uyx
2VwDEtNdLMZ1hP8VeggtE0QFqI/9AFYTnf/EaJ3c9Z5XiXDl6vbBDAdhyCzdWsHxkmRH4JLpcN7g
Ua00e/PtnTDUrQ8Z1b7U0ELQMh19pWu+6ku3ivfuk3FXD9LC77qUTya4cK714gTmEC9OBm9+0VNF
wO4ygV6xzZEBO0cj2GZ3XShFK1hvkitZuHEJwLPmSHWU2LTZG8rBO2uRpWuO8umRvmh+zm/Lt62f
NlU9xFA0BhhZbk7oH6bnZuSIEBJTmDjkBKwdBaaVWNNg6X1TbACjEy0D97fP+n4gQOLPzYZNR3q/
jGZJwNzB+HOyY1D633yh887vUov0TcIkxNqeUhzAUt5Wy6fdRxqgt9CLn/SLR/yvsETAMWnob3ye
P+Z/NT7u4PDVw/TouM/QfS6WGBChUD3AD5mU5ZTJUU9Qf4yqCDTVY1Rn3G8K5SjmdxBulvFw89sm
YYQQ82rDc/AxtSWQvTuZlmIAF0QrJYhizDl8kivrQV3N455Hi6t8nXrwn1BjiXaPve8fP49fK9gm
2aWInaLBLxWhKis5290gvA8HMCNLp/7tXshKQyE1rko3fXN4oYClYGvs75wK7/sjgcTQx3rzX+yB
u8CJntizjUQwTk7gasxZKBQHyI5bZMjgkzzgHLqlJax/vJTxYzxgt4B6Nf1iloNGlpqFDcA3E+La
PIzZREQuUpsHRAsFTk9JiuDSkix284oazxXf32lFJUwCqHFBjz1x1mgGnWkukzqOWpnZk6/5e9dn
/JfH80CKlIM5B/vCVxdGfXMjcDFvCTLfxflC2MM9Otv3QVIOuKhN1B3cqERDprMwCLmQB5BFs42c
C1ON3xTjP3P71/fH1p26dzs8YUzhT32xP5CrhNKAzH2yIJ/OkfzTYLOKkJash0bR8SaCVQzUOV+i
XntJWsjekFwmfwO7FwjXjRkT+2KRvGNtJQJDEtodlpAN5Zv+nyGGqfhOYCv6yJlCZ0xp+06vdqPe
gZMYJ0PdiphKL9yrhAmwNfChIpNXwh9oM3nA18i2z2ZkJcq0iOXL4eErYJEyCBJ3yOyh2BM56mzI
PP67pnRFQbPqL+YjIpWva5+5yWwK++kxwaw0ZZFa4lV8kJuMnk1RwFeyFpGJzniCKTTMXkgNc8HU
6D/rBDTekn3PqMga7ZKzAXqINAYlpESHGO4ED5Zqf391IuYXUl6TWUBzKIQns6YT2pGvYKpWroZn
VTws6sij4TiM/3Af/CESeJndyWFFwP0v0MPGF4mKFiR7VTrlwkZedTvZ93HctQO4R6KQb05rTCVS
/rz9o7xHaeXVMEgMj6OXrvsRehNKm99t+geBxENEPb9Ke4sZOQixhUo93ZxbOayGPb7xI885xWBb
220L6IvnZlr2Q8mNha6Q9EYB+0tsU7gUziW1LWkUyb/IAyuyZrItSsG7GXWdHto/drcxcroNQTea
/lduGgrFIlvLhFc833b1ZhdKmRO4mlpi+xF9kF9MnDi2he0HCWnfjxC4DB7QLLq+7OfMoH+UO8zj
M5CXD4BocywDzSxAoBHoyl3rUO6svoipzJFIdO9Z0yCZouYL3S6icoH1F0C27Ri8vvZmEaEOMG6j
JLv6KstQCOjm8+Er8Kmr8qFjvueyTBmNhd5H8lBFfY/v5F4NXyOyKMxcaQmH2noYYnPZKytj4Nm3
/AFSNDHUCNGrcOkl/7GnPp8kO/Y3uqwcwlN5Sy3/J6FGpS2b6D5EA1khdUl0KFdoI3Hdrg6gRD73
aZFC9CAGt8RAQNPyHuGOxlawL6WJTFGBVYU2LK86jCxVRPMlUc8Gzp6NFwtPPgu0ILzuO+W2Gbul
8vu/7YOo9Gr9MmUflfWcrKAT200eaEv+Qs7nuk/mhuqn1s6brTOAjGV9aC5LqZOjTkuSIxm0PlAx
FX5lA8FtJ4mu0+Z8iZYYiWcnSiD1wWipxjpeaRS7L8GXwMYZWMehpwgTG0qDFxFwRpEZVtjyEgrR
GV4kZiaUmbC9mVrWKREKuJtZMTX6iVtU3sKrPABfysGPGDy5tQ33+U2SIACC7BtYqQdB172lH8SA
JaL5fggmIzcUbRkPdN7y3D88AqJT7r9vPL2wscwLQs6++rch+azAcMbh0+hDzCXCtV/Wq6UJVwj5
VECy3s3F3jlVnWwTwC2QgKPPRBaRHZ4yjk62OlT3rK14jKJHmZZJ4VfzHS5nPQEzKEB8gBEZRTP8
oMLLYGTvZqcVKoKHzt2jaKcGWkenLx9nPePjxAkNWWCO266xx/bBhNaFscHjbrHcbzXXXro/qsZn
TzOyKjI45oe00fDcLnKOPRPq6vgn6ppWXFq1DaufQiAVfYy0gKQLKLOHXMn+ZKxGPhQQ8fKUi2Mb
ay9dbQqCTWVdTnShHI+8x+j6KNpY2gcVbrSLeFDTLmKtEl43vnCVDHwaufQ6Q7q8bBbEePabB8uf
KKO0J92XYQYi0bPRGOIrYe/5TaXCXW6MbxnG863Sy5MZwvVwNqXaLuFLiw8FvcoEuIeSYeYSZlya
y+MBxPbX5t1Agk6z00GgbHjG82ZEjMYFBjhhxXKtxyHKZWYiJJB8ml/Ih/nd3oqqMUopgaZdXTFp
Fph7YJKT8ti2or+qAB3csAemdYlElf8d5RtlqgcOHhyyOdXWtmqJUfFjPlSl23GW5FDqYS4JLOUK
q42i5vUFeNnPEihd+ntWiSxnIjrVgXWrf55+U47mI6H9EKpHYZ9Re46EkIhVUF8u2Pgrv+YB3XLc
Ua2/+QbzCs+NSBx4ZYBunTdm5U3vNzYYggl0se6K5rsZuDFdtEgoPqLCmcZ9Y6Oeaug8u4nO9cgp
jJNo8AHHkCDrF3Be7frvGoI6Zg9UDhEl8MbJdCstXn8PW00TR11OkfGnqz545h3C91mOjhI0loVa
Zrvd5e9fwVD4yRrfAR1kT5wPzvadd32rJgdM6/rsUVeiNDqoa5QaGW1OvrMNsuyDNta+wj4nN/GT
459xa/t9+6HIzJ3fxh17wL7kwKfzvJAND3RSHRQqmdvt89vtZl8wmp3lBDQAsT3l1inEnPCUhrTR
dJAPhU10NcKKjy7sCGK/WLkAuET9o/S+8y4TRdHLLLfkNgJiOXk5Ui6GdwYbRgJFKRvb97LjTECu
5cwSLKDShTB/oA+2vYIrhw3mKe4AGTdy9aCv+K5cKXwaQighWFQgjHcmfGqMMuVjgFULny7jLSoE
VpZeqOVD8BH6+u8SLoC/X8dWlmWc+gHnFsSHw1esTBTxmric9mftHk23K297tUfQ60GR8nduiLDf
btzAS737flrfM5I1UFJHPiyOFpumGobySJ0z3tVz+O6JNg37hS4N72CeRcFh4w0vjX/ij8KBdPMq
wUeUCBlj83sE8EGol4q/C+FsBqWkXgGvQ26nn0Pup1iy/1ZEntTb6gzoAIJEQ0tvRWOpOqCOeTU1
v4nAvcXi5MytFEpq2xDLYktWk4c5je0OMPotW1pQDr9k5GbhApbY5YxvPCT7R0E8ynNhkOj8JSaX
zlgQfvYpol6+B+vwg9Qw0yewlMdGnXmrX/nHndAH+9M9mREgMnxCumdKPo9anLPrKWkCmYyA/XjC
S3U6KSomdPLmF8ChmddCePkFIEAgSLDBKwaIiRI+UErYUj6NOwTbxGetTPPwlDS8xK9xyi/8+JSZ
iKdp9iN98cvb91TuD9+6BoSglypG/P7ejmpM4ayvR5VPdBu8XXFa1O5LW4dlrW+e1kydLBPeWdhC
PUOY/nY0UDfamTje1Rl7nGLOtpFdWvuQ0XZxR1UwdpgWUtpyM10EkrvZevqhaUmMTtQiQ/QJz0hM
jC9gJmOhYT8Y9DmvNHXpP68CLc8rCxz1RsOVmfi0R0G4MRefs0D1VVaYGnBRmtzmn3HwZCAWldvH
8Kd2dCbx4Rp/mxyEXaJIkXDv5XLTOMYLp8raoYXmVuNpSROvuLcA2dseafjqsIVIcPPBCaHY+itn
GBCznrEeM79si/lf94ohvZZKBrPiLb9A58KjBTWDeZ03b6OGjN+7W9w63YGo0Nex0oqDrlrfa81+
8e+hULEy2nFtdi9jd4N7YefMlx6obt0Bu++RB172gK8ZUuloPji8BT0k/vcPaJsRt3KmhnrQaFpp
GsMSYJnGo97Rl2x7YRaRnwyyb/RHq+ta4Ryl080komgPUrNqjSGsChvXMI8q1L/sKd3XXUTr+NAg
zeBXhXZpCkLY+C2d//jZ6wJDUzb8a3W24jsDTiJMfqgikrF2DvlBSldh/6j3Ax9t4taUgYfXqBGE
zOqFzqgYyMDQKET7qvtBsbAQdJnGH6SgbjZLpZBrKi8Pprwx3MBd948hbIZvpLOAeWG8PM/80Hk0
XRrLRDnxNh7Y9jbjE/4PMIwETA+Ft/HrhyDIi2AiAoajcl5rzj/JRl45COcsNfrcdt/Brl996MtK
YFJJuxdcz245wTKvk4iefF206YHXfT+S2LKDtEYuekA6wc6m9YYW7FoHyc2zadM6mVw+4Q5cx1Hb
u3JBpaYMJWVVKe5rbXWZItYeDgY4eOxOr5YKYjqRTQeYzygqsn6y7ENEt9Sd7tuaLS8aDiKx/2X+
0ycRb7lFW8aNShA2LWBghKfpkFNEpq5Ak/7VkgX/zz52bbZ7z+vyLpXSgGYLA/zAQvxgccNStpkE
/vtTd7gN0DFyAv2cClwVEOIELC8WCfibpFZTQ73G08VPwFxCeAKLo9KKH7ALsfXuXDjwiibEtvK7
hr502jRInCwUc+AraQwNbT8Akoo0Skpe7xLiQ+4SrIcKqraq7cUfztOBBKqRehYFt2BNoWox7Nlz
qB/WsI20dczQkW7BIby82oezWZJineJnQBjxA1Yx7P5nXTNvXw1+UwU+nHH0GTTQX5zXwxpTyH6E
xzhaLjOLgm9vbgNFt4L8geAuNVqEHH8DGXQ9HkeswlOzquiMjOL/emGrdFnjU+Hqy0SNZK+WWov0
kkeIpzya0hn3ORJQCIPDeaJ1k07tOD+Ovzi+Fh3n3fq1p03gJE9vvrcDpWtJOMkMt3IfzWOWuEu6
MxYrMNJzlI8h6WTwXl//KmLi1c5FAODE/pJpZEPX9fwfNt3/CgOOyYI29pdpODc0B4UEUeDKt/O8
JB1F3rx8kPLX19bCz1/OgPey+fM8WbJ0QCw3xPypRpV1eVn1EokzYNd4MhBq0ndyhiSwIhEK4Okb
5mmo4uywtF5hHhxXr2QeLNPMq0csmeSC0vVNqqysqj/tO94ZlXsjgE/A+l+oWSxjSBeq6NAA96q+
y+/6x0bYRb3QN7NU2fcILSfqXFLNo2Rdh2CHrugmuaW2jgPbKU4A3p/u5oA+X+0Jh8WGl00XS2d2
vc2VSGdVYTHtfZSua3i8U9utnRVYBYxFjq5Dgm1QIwGj3ZCU9MjzM5+J0aVhRh9tc4uaGFSIlTd9
k8C2kWxPB+3Exl3pHiGb0oIZA8Q3ZZLWrgTePKlsUmN/q/TLbbXkAPjyMVqnLDeDc8j4nlP4UfTs
onDAtV8jB0FoLHcMLrA9wdSuS0rJ8bBbqRfWWgPNbCyqEjpwgEzE6gEuYZ1js0d4U+4xtntubr8p
22BE5IFLFAY2f3CWUBxCBQsQK2FIzftXpUFRBMNCn1jH/ZQHAKrI+ROC1nLqn8O1am1Ai6kvQPU5
EGHxn8jcxXtcFNJYtt81tCwZ8wPn+d4x5/IV/q9xiI7GkNwbNtiRIdOnhKtmpm4jGOsY9OkA3i04
289rooZXCH/hmVAX8H7PSuCfMboMr4DQckYHXnk8Cdm3oa8hO9EaM07eshY6wU8NiY0jJIglrxhb
UWoxk5+YgATHp3BgMClQXI7SNa+r6VefJO94vdMucjuUfRQwOWUgny3RFSgq12hPVyKjncdForkv
MGY3tlj05o1KtpIf5Xjt52LTt9xp+NZUKkurx50Rz1kPzjtcSUTY5qZKgQjtnPuvDxXy2ix06TPm
KOcpRBABpll5FYYmWIk1GeNh+1av1jtL+UM2gtoV8QjXU001jCKYEm1qyDnlvH0eqNr6+arldbrc
MTLVtKG3flwSdLe4VRcIQNbzF4IUyxpbQA04kGRVexFJ81bGhUBZk2m+RwU3/25bhBBGSm08uYDo
Nsa0xbB6CbD/dB90ixfTBIvgiOkLKUSRQ2SHr0ydIgEG0VosFOufPTVhixj+XXVmjflvfdfOU5Sm
pPuAjQNr8lM=
`pragma protect end_protected
