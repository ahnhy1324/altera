// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
o9azebE5N61zuNtcc5WpVUYntpQK8BR8TsV+hg19kqqLv8cvdkA8pnzlHwTVr27P
hil7ioAeItFTpTC0yqJJm4Sp4djN7BWZDnBqz7EtdpCPmck1MKs+Qq+1hG6m/yti
ZRUcRgDB59Vg2x/x00acQmlDnLUt6WRcEhbipkhS5/g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9008)
ZZiPC571gZfIZ5l9VH2I913ZW9c0H3FZZvrUDROBd0RNvkZTLesYrtkk9YO7/Tdf
OeVMg1B03OTcFPK7bdk2mIqxoOmGMoVtHiPSQ2T37YMHPas2To0t0bdH37AnSmyh
tNz8YsZ/l4LbbodreYfaor7cAK+sC6t4S/o6KZ/iGUd/7ZjMZSWE8juen5dqU930
VDJ/bGpvfIa4m9K+VreTEDBTjeCdfJaiakDihOf2n18RNnXlgTDh96o1oKgU/80R
TUVlgxx+UrS87k70jCCG9ECa+uZUh/bLVei4Qgi88KPVSsti0BxlOCHk5ZjFBmSw
5RWaRLzZbVj4VYljsvNPKmnDXzmJ08IP21RHeUKOUj9+gy5X+x/aos6llSgksbbB
bA0W30/84PPfg4gD5PuthHQYXmTZfPgXZ3JyKjIVc4eJMzhlLpP7bjCnbv2EogsI
LcRn8p8mOgbC8w2RXnj/rqsDiC+e0rtA/pdAd4lETUmW4ocAtTk+/c6DCmxG+3Vr
mD3nTlNZO/e3wTvbpuYlt+PPO3W52/7du1kDs4vshjrm51eqidQ2pVMmz3VzXFcf
//pN8/i8Z+bFJoXOnKP7ETrs3avccOGI+Hhjp8/9Zibj0u1fvxsJXKYZXu0CPa6y
npgJhFJHlWQ4ta3Vb0SAgHV5bjg1TkNOunLF8ZDbSW4sfnvFWyN5Y9cjvxQqohjf
31157D9lu4zLNG+05/xb51tCNHRFIv4hMsbCSMOtYx8FC7/zsmja3AXlhHY8nFAq
bbbyXsSU9hQOnYGSk1CsjHMyHyErBDJWM078N2sEaWOqFCjv3hROneo8vVafU5OM
3f5/CQKy7Em51yjwRuVI+amC80VE6jvco1BwpufFJlYVO4TvdRK3YZuXmRE6kHcT
tDs5mvRMZEscrSmh1oBKY+YmSPyEIRaHjGDAtUWKwp2xG6UxBD2yijWPNfPb2f9e
xgeR/KJb9f7Os1FtZPg8eNNuhQ7SFMHhWZu6cTHkKhcpByRhr5oWgb5eBN1of7Xc
ryDi5N/kHdEcpw7FFEVI3KEmxGyQbhZtxwOjDSCs5dT7AC2S2QABDsDyOtCiH69o
038Cv5ZArAYBN7tUhm+/Gxi80MuL1A/Ha+1VLfbENPY5eD1KRXtWdG+OpQquTZyq
4hhVEiOM+ksrbayW0U4Srw2igxlkaUe6fkgLIoCykcjGwWXnyR2XTySEcFLAsM7+
dNUt5VAY2wYMM5/lqBwsNtDhX+wmNJO9j0SnN/GLXcN6H7SdQAYk9V3ypz3CiTGX
/O5BZGTClj+hGNraT/HQYGSX/XGDE7pVDws59QmKJDMtO8jbeK/p4Sw8CrHvnh01
ec9Cjwz6RqL9kwnp8V7ZC0+G3t5DyV+Cw2O3ptAOTE6+SI+Tn4LG9KHttp58Jwkl
qG7Pv68bVXVm+NajswEkr9x8Hr0HPdAmA+w0q3sE98XOiCX8LtFGJ3DVuVuSNSQH
Y0fgdZ9p/+1ZyQClPn3iAYQeYWNDBUJ/FYaXjOxzYGIxR7UnrldaBqiUwQIAK4Jp
SmULFgiptnc+tWR8iYvTvdTffYIe9/n3dE0S4/wrVVbNPHsbm1TwZ/rxQVArdUqn
eFTBlxtRLWyB/vK6F6xUxtTrWWAtesZN7xvyl4K21AL3Blrb9j2T5oiHWTd763aI
zE+W1PzCCtaO/2k1S6EgJLV7h3mTkrZoBGxN/ub4oudVaXDvBxOeLrPtbCiw4THw
i9M6lF7ftWLZ+wG2G3wWLhgNCNpKwQzBpUA6I7vgId4WJ4QmsdtjaGq0YlXfseB/
4ERzayIIrxWPqx8Hhi3MspWYdFz2umWifKxllelanuVjjJQeV852mVvgig9avczJ
Ud/csl7DPRy0rhln20SoznYXJk623pecUMxtEQWXIC8gvKOWXvq0f+8TCvslk25B
DNTO/t0S+KWm1jkuJMDnjWpa/dKBuHNXNg8e9bKDIWCRjsdA5OphzSMLSFYgI6tZ
danKUlB2r645comwEFYx2GOZyHM4EMLXHpX4sEPM6Ey7pVIzaIeFl4MQ4bKP271T
SKSw+O568gbVBYw3mNupLcNt8xa3WuyUvbDkPC3H3jUCnNtDRBHSVfQO0DCq1xoq
7g8jhWLJmnVYHGPf9gkJUxN/e8Oi9cGzZpbwzHmjONzXZCGKLztNhEveVXQUtevl
F18Oiuvn9jxuHAeJRlKcP8F9QNk7vkB6zxCzyVvkK3P11dyRfKCy8YAWIkBrBs36
Ixgc48d2DtoHGiLHwBovg87CBcrvmdcgibmDFU5ty2Y2iZcfFyQVzdXcPG++Wl0b
EA7n5b0sl5TCmyCJko2l/oCaSR8Cs6J7H6YXhvm/iiK1sdJ3Y9IrrIHU/wVJUUQP
q7UPbSHjeV/y1ctU7KVfzoe45+MXCodzxVSWbIAx42maMXOFv8eSp7/6/tWOGbQY
Phuwi3il6UybI5ihioSzasaM+YRqXpPsfunvAtvKudbiKnLTUQDTSujj/fZ32UKv
Cm0ip/X6ytxi+S1QcrULFaFnAnDR4bCl+KEMwpHhKARGUCDt5o2vMvmte+rf1/dX
I4oyCphJISd7CTUqCBHa4CGz/kTcYh5dirEK+KR2VpjE00p27pKeTf/s2osHPj+H
/WBiCZSVt66EgGhobMxw3QRGfI420BKhJd2j2F8SgkQTte0o/nbd8WPdyAY0wkxH
pZDGfPVzZwCrsIeFV0ZqTSmMI33F7j5uVGBIoDm8g3nal/SPnx2b1baCQTuKfMIt
ZEPy+uPbWpovywghvwxNLWvw7hO0/F7T4AKUrLVl4PM8EaksBzOcXsUysg+uW6uc
DoafIdvztccE0m78ja5XI1HjUkSMD8JV/LEyLLALHTUanaGLPlalXRHDWiKuPhQv
ogVFpJT41N9xWDNcBgT8NyujHrISYuFlx0kjPwjGJxbEG/PMUAUsPXQCSORcWwvL
Rr8oE7fJV1WXzmhXslySQW9TqD+50UaWpVOH4t7J/gR+573MLD/Jt3ohRjSLBqOQ
yFe3knvQQadONhF5Vpxog33/8KzBzTwLMbm5wWwqs9zJBvNBVrjcvYQicpMd8b6T
CJ4KY+KZBJPnPdj/N6UBD3NGWX9rNENH7gmQRd0mMPgrPUdCHqJnVtQTVIuAKAXO
kW43P3fpSfx55y+0EP+HzZvbBsKcAmq+78kIhCed2mZzuj9muGLGTfMEgx3+QvNe
KVnkVrYQUh1bnNGNyr2BdtMOeM70Y9VZ5Gma/56hUra7qqwKKJj63pJvDfReYW0c
078brEVJetNGqmuegYzIJwGUs4rOcoLoArOHzfR7EJn4jhN4joHXaR+WAm4VWuA5
FPDrSc8y7+vsXVv7TjpGjey7Ecem5YK8KWadJC3Y0K8Z3jlVGv5pk3RfCvNLSTZI
tRBG9LKpa4s81y1uast9fn6vfu0vJQWwizxAtk2DHqIrmXmGu5BUMAA743nMPp7/
nSW8U9YITCIPRKMFQr/T7SnH7LjtNDva6jNwJ6hM8Gzq8YU8D9RlQ6Y/gjkqHQvt
ijcTnWQhtkyZTeRP5tgf+5dHbuE+iLslvv9i8UiDc1xCL+/a4sW5pxR43cIj2Ihw
qunx8UoCI+acC8AQdPSCtNl0nam82C6KAODZEHc/Cx3pMdfT1zywPcLNWhgYHukk
sUm4anzF97JseZMmnQPEUIcVxiNzA1iEAzNvabZPumc/3UseYLje7JeJGjT+twLX
AUohFTwJMVP/syKX8wRZq6ynRcuXqRM0w+LX9z1YaUIUrI8LoKEmMZETfIv8VRRW
PEVUbk28bFgWR93jSIkbVB9Ir3vaWIyOG2CFTo8pkVHoIxlRL80Uj96eN4b6LVF1
7oDWfPbf8zGRlkV68lN3tkoXsMLvqrgLeAtDwpPTRbeoP4jovhpFGR+RV1M5MxQw
PiluJqQY1WwO6uhtQ8JJ90ONUsQjdmuQ39Lpo0LYqVmfIZnTgHOvfcuuIBl4/fzp
//E+o5cTO7hwwmGdi4qpY9nFsZsB7NGuuoYGiYk8EGZ9Bpo+tNoVW9qlcFI4D4g1
y84OzhhAUydrjbwUmt5No3uE4yz11Yf7dwJJ6Jqk8CuX8F+BSeCFA2OC4dK4RmY6
PVFsrhjOrfhWCIb03RtOeTTuw1jGt91gj/+QxEQWEHmu//BIYJbhcsU8WGfUqpT3
NseLQAd94urDz94y3VUvAhBiQMKee47np/up1V0DvLTEnBYdSqrWF0BXu4paINdX
HL+rW30slLvb416TYxwHbUneCMszceVd7M+s7tkiydhMcmZOpQzUjiOL7n8BJEsK
lNdPSH+8qOVtfyncqUbmXr6ONQb3fQUCDH4fZrq432zHQ5kcdh3eYEePTTmFDRMa
18sFJrOW3qY+e+qpS71PPYdJ4GjZNkJYCVBjjsaZA9pFLSzIjAWILLDe0NqYe460
ZnFu2vVwSNq2kEddCh100v6t559GkteXpl872wG/wSsh10L6blnCvKhcfRPUTKbp
dHpkHi2oJBjw8LfXb7Tgr9Zt9dfhwUzArL+ETQwJRL+ry8ZWhGQuhGtyPuMnCiUz
qN1m2kFOqTqu2DUynWVdUfLAI/jE7fjUQ3fojHrB4BARQkksgsZAjIaBN2p9LgVY
/Bt23kf0eWCesLnNjs9NPQHx8OCyVQ07Xqx0v6InmSpYkwdKTHymrKwdX+n433Im
0J5EKpUvNIt5RZ6H+XNUDMQtVxPbex+pPNUqbsRsEAXpWHRjaj/zl59E8tiZUpR0
OTiDfOjk8UkvWS1FRcjE5b2Zl/eH0YSf0C4zhk+VfPFkZY2LTRVnyH7+Tp/KjRFC
hkJM4/D54NMO3V/PgjDYHtuTOB281mMXpUt1f6prhZlcsPjRzUg4xNRvVCpyNhMV
hITqX4fUJ96iL/zGzLmbVpYN9vSuK+HhNBnmWVOT2KGTWNB5fFp1Gq7Hp+Wi0yEE
/DWHWCWboCDoG9I9gdXCAcJvqAOFpZM4uECSqiL8GIPmRkYwNl8Ad3wYSgxg6/NV
EXdnP1IFc7xwRpdcerirPIUuQDGhaUemzkdX/KFkS1YC5kKILm8TMA/fPrJfzZfG
+ePW9FHVdKi5QGLpS3zdR0ZUUUnl8V9fk7yF0SvIFEsF/yLidAGpYpjlOhex64uo
Jqr8geDxSKidtT+VnM9Os1QMEpBGLFBUcoAtXx2/p4Zax/Kg6NVOD+4tRa37ecra
acDci7zm1dpOKd6wtebUambWFJVJLByfi5Wu0GA6goaSl2kiP3ARG5VYNUuRSlLG
1kdLz0n14q2ZG6OPoILsPvh9wUthi+v7pFchTT6D2G3gO2w2uBvxW4I7MzOBBaSo
LrIDOfmmsjggEbTUsmYCUcNMFnaq/JayHeJ7M18OddWZXDVVpn4MrC2L6kQMmvVi
aLr1Le/ZTouCav00xQl94Jf4W+sWgMokXBaJ2rTfrC1R9bfKh2QndGF0m9xOTWD4
GFPVoWmrn1PegKLd/W00IVYvXc43vLoaK7AcRkPlHn1Ei3Qu8bslAW2fH5DcN0kW
Q6yXubwE1BgPXu/TKFhEQa3L3nyI6AF7oLJkX1ouTf+EWFTU4acc5v1BYbZHYPxw
bSNkOlbe2dDYFGMM8mxUWxUt+TiThVYN5tXLZFVIufDaMyowSsw8Q0HPzoRMXk8j
YcCzTa1dJ1bB1+6bSqXaOG8KUrpSXlbP4tnUjJcQdWDlIV8RBrow9iqqcCP1ezdQ
9fwyHRgaUxqjI52Oaga/yLD9VokZf0mV3oiW8onyNqB/4GJL77xDzlAqcTZ4AroJ
9f+lNbEKbtUNoIq8vBr3FqaZI4qZocFzkKcZYZhdzhs7jswTx7AnYWj9qquAPlRl
eT38BUvQD5wHkxcxIGrXkHExxwHt8+eCf1lJqozREJiMbD6EY3pGy/OpiSF/V9Y5
88d+woupuEQX33loJk8fcg7Yv6QjRWeh9dEeSJmqVbu1NSTAeajIdJBlhVqlUjaM
gBUxBQkwEJ8khd8ca6EqKUi2BGlGNZsVYpfjnSd0GXj6sRG8Ff/lB2gHHGoIsrjH
fGINS76YXc+hFl1Wr2APVoM+OZc84bkvDy8JQu8+kiw0ubA0SuPT08ZywEq0Hce4
Hjw3H2hidEnmjQ3QhnMCU+d8yScm0aWJsg0iqQow95DKK6sPcuG5WhWiSRn3ek9U
8Vzbmn4vZjEK0z3rDUGv9eSf9mjCHN6GkN27Pz2CZnLCVX1L+FpZT+2tvcTT/0iO
Z4C9GY2aV0OL6VofU5EYvr90hJP1zbl9rVME1ixhaE/pWUoBriCvyhL5eJkugFlt
s44j1zYE8ZgutsjdbsNATbDNBuLB81i6ThN89hPKZjqk8oxKxPnriK20WI267OXJ
T//4fah6Yx9T84+XqlS35AlIRnDLI6KZ9s4AuU4la1jc2DhFfdsbq46JVbBGIwi4
qCia1G7tZLLjqqh2zgKcEuM1oOk3Hk3mm2omuGUB0iPGu+rLwed+ppCtZxa2SV2n
fOTzGEiuN2GKYDtC9hkEolWUaehLvNbAA+OGle7CNbZ08p0+6L4A9fK9kPlpj/tx
f7KxzXhbLIQm+gQFLRkXKvxxMTylIrJGmkdzeZKaUr1vhbBNDIA4Q2hs8ujEvstV
PdYw7Un/R75fb5scBGqdZEXl5uSuHj38iIZhdQMOK1Z9n32+/nm88p5zAPWGCHui
fvp1udv8Pyq0SFrxx+bZg9Ezx4c0N5urnGD8uAp3mrKNKHQHkae8kKFYl8re1sF6
9d3VITxZILM+tgPzO7ngB6YkZgt77yFVV3L6MydIR/cmjv9JjGy9jZwH+c2gGuou
nZa3QvSrCfofwcIT9SWMoLh2ck2eq3N1KRABPM2F2drIxELyHj5omgpNjrMsPYIj
sUFhLedjIdCo7uIqsMAze3J7ihGltOY0/N6RQoST0P84q5hX0aZu3n/30L+Sbt3i
UeNcm83yB0jC7gKd6qVIxjQgd3vtXavrWKASA1A7fDeuzixDpGOVs6ja/MWFrgFD
eS93OgDDPVetWn3Z/dYRiUIh7zZ2n3D+k7SCm4fHY2eAu/+VwV+fHJV7YGcJVPaN
MqEo9A5MXegXO7SfLa+JcW+zWgH4a4e3BVFfg5U4iVL/RPVCwuXaFeIDcgM0Akks
OwDVe0cIRy7y+sYLmLC9meN2hZarNtUbSQK3Me3JJc6j+Nfzaxaz8o4LKAFzHpN1
H6IKjGHFXcfCjBM8sYrTDArLMGzB6mVRvE/xOvReNHhyXyaLcoosLGLVoeBYpcVs
e1eLVMW0UeJ410eo73uMzf14lVZLGHXm6XCBO1agb/tAd79aDiFDN8MwFCyC30kK
kudYWUZT8vyLsuyxyzSfZ46IxGxf5Q4RTlgCd4ROheenRMEa5kei4+DRUN6wr7gM
f3ExZFTkOY0vE6QS50wBHXaahS6y4KsR3RPJLkpzPOEtnXma/qjk0pWK1CibvPCf
jAJ8ck8Dw+9eYbVD+jD3dYHgXSUTOXOJuAttPtr4gqII2219/Ho7H+xHCMW8+3jv
hs7Q6HxDpAkPXS8ndEJHZiPZ71Bec9B4754Iy+DJXwvmZ1ZH12nq0CB+06P+VJIt
oi2VSyirDCrGTZzxKzc7GkruXRT1eri5YpT45IrolCnFvjb/0/VMoNayeHUniGc6
K5s7ra5Joa62RoBsrwv6DN+FrLqZOg3FzglSbtItfsRwBfOrgDz8zp+f31kAV1q+
yoJClEin6hD3pxbBLL3UurtXn1iJ4WRqIfxjEyVwRRWLtQAUs5UubS2K5/cZ22l7
AF2y+RtwODIum4tsMwMaS5Q73o1NOw79hZEN6lpBSPzthPCPocAdEDKuvm+9Sq0/
mmXAQD8zrMSBynR37IBYb040ajIz67FtYztMx4EB3Ks0q23tkWlu5DKlS9n9k6R7
YJpGD4R2aJNm2kbCQP4IJaB8Ehy3mvyJWneTtG13rrocAw2b1RzRa11kNP0tYiTO
3V7WBwhIEOB3CSLpFw7wh7YEnV+EXefdTquT/ywPZ0isJmGsS6XwrpUajsnMNK8s
kG7SJcNRLSa3PZKP50cWIxETG4sq73IhwucRxATWEwVFkM83Ks3LzNK7JqFNHz4x
ROOsdPDkWVbIfSTLVQIeAGT5Z1lg9ED/A/3xqj+iPvo1Nuh8Z9aT03ufnM4ToBPV
lJYI3s12ochZCn5oyPZRAiBuHZXOJ2sEQyDbLXWQZSO47Q88waynTci1yoUcKkP4
azt3t+bftAviYw6A9gEAjdsUENWDpPK0tOQ8PSrhaAegIUo6JCNAiOiwEgXHbOgO
kA6aIDoezV1zXfxuA+noQAxBxwT7ooE3Mkiab35pQMVplkMuBC+4YydJxR0Nr2Ve
okXU4FSjtCfDynnYYkRJUbmtcJ+iGl/sTqlVv3fgGh+jmYl4qdYes/HAiMcCO/rk
ltV+BGcjDEicxOnwKBXpH77eZSuGhBTs78+gIJiPh6mcb/PPMeS9ecSuKkg2mgKn
A/7D5QL1rBxvvlPy7KQU4jQB0k6l0dsp3WnNUJqj3ngmjHeRyM8zZTJYb6PW2bnW
dUsX+u6hPWcejhTBQ4fRXKQcwWTFgx0SDKi3499HAxYZkxBjJKvOThzVuKZPgIs7
vanX5eLkeOxmUE9GwkKwkEEDKO3WhB5odoCFIDJf4detmlF0Vx68QSizrtCcmhX6
V00Im+bB+gVibMJE5z2UM94JUbDZBShXF43gFBM0Rs8D51KFz/vkJqN0b5Qi9cI+
YgZK602rywQruBWv45iqTTUJ8HKcafftHp/N96KuSD3Vsht4O1KYa6e5miM32gby
KXVKsvz+XH5LubcbiWuSBQ+cE03UFgRViWKrZ4nlfq7JSINQQCSaDNrJMEt18VOm
P7MLeH8M/NtKLIVYQfMoWj4f4Igb7ohBVApaSY6eJ0ydhkKIsK2o1f/0fjoKngOF
297TS2sA1gLog02Dtu/WkO2yfTcyT0TMKOyoDNuvbwKAa+kz+0pLxEBDkL8qvSHj
lwOrGrm9YbkIUJGd/VnmyaMCwO3Li4g9VV5u+GyId7pX1OUKJkzdHtcJoNIsChjb
ODx6u/8Tjme+ecqBQNbSS96wHwCP0fL2VUYOLCODGVOfOgjChC1DO+lcr9DsySmg
H21AXDDGkuRZ7ttz5+wxqwD5eBzAKse33tAoinHJCfwOGS3N6BfmfjUlhmkLlYsx
sxnYCl8K4A+vgmia3C0UkS/pCm9a/Rk1DtmsaBA69cxxoPQSLqLkWqg8qkx2tqE0
L78YOhaN4YePX1j794jzpcxH6FMF1xF7GTaAIl0HxGPJyFgIVl+qHaSOxaZTb7oG
ozd3F2pDS2BhaA4tGo87pnlIuHi5Tw+tO1g29jsk75P9kZ1J/yUzFsHX30Wh4iAw
Q31oP94xUmz3l5G0I0Znapf8xnoSWPitRjqaxuNP26oWI+bgaaws4hyFYwasvR0B
stNj1dCGyVEyQj6Png7z9a3wtiR67vdbVNgPqn190VyjpwbKUT0JwKUhOjFUptCs
SLfcaLTmbMHv0qiAfRmXUN95SGrwPlGRGiL/U0bqe93YcN1JzdvuwPMn7o0GA+Re
fLZGf9Qnoq7VihUemQ7ohQ/Z/qhjkyFFfATaOlNSfX/hGH0m5IqyUOY5ilWNqY7b
0+0hJJ2Erlw7MeKeo03U9p1UA/EWzz5KoayRH5s2BrPNcCreXELQipWYEjmJTQSg
yaQudTX5L+a7tkVM/UXujA5aq1BZDylkNDWjF+w0P5Lx8wwRZss57NZsZIzI2cma
vjDtnr+kWW9dOc9R/q9cIAZB9kRR3T7ADX+IID4qHDAC/5oMJLzTsqbS273u3lbo
gyehmlOaqZQlgufCKk4jKc1DgOP0zgYp74qLKtTIdCwTHDNhA0OiL9Q0Rd8l0wfZ
TzYEdPXwkqyI5TvABiZKF1EQIwYXgQs/pJIwE1/H8Xzr84sFRsmy++DAP9xoeVyK
S3929JmQjDMhQUj6yRI0fdy/DQ+av27PFVhzek4OQFVpE1yp1nHdrDSCEpfNnmam
NvBoiSz4Yl2b4MGGQvM8YOQeRqGFZ3MgXVoFn7jjGunJrAL0ijGvn1Or1+WjjKTh
duZGLMZOWlDmN0GGvjlR1+hrkqPm2aoTAQ5Svv9aODj7O4kPTxhrQG0KqilGBZMB
MeEtkXx9PlPJbtJLv5LdXZM+jcEw5j+AdSvWh0mieY2ovknDrsxddB6Emzdg5qaw
PAA8lmlWd2GC2frbRKgjS2E5s6EvonG3vQwcvqym6iK1BUd+5u8XBxgLuU9FvPNT
Xy7xJ1PN70k4cKlmUds4iVi2nO/HW2Vn8uRRMcURL4Phj6YI+QQGLDgBTDEbTXfG
EJFP+nqYinl7fZGik3G7d3lNixDb5yGRAtW4c7koUk6bB46+HW18K0EliIQOiNv7
XAMRJKZc2BIq0OTCVEYZtAoNZdPAqAs99QPjWZNXPUgXakDDFh3CaYVh93F4DFBr
hXP42COdAVZvUhlNJzp5B7RPwWaQlWIOrcS43EtZtMOCOt61EWY8Z6A2QSyhBj7A
uAKC+BaWybkpbM3RoHVDFAT/5mI6p1SKZOjwcDvt4isjTyh/+tu8+DqP69G2G8Yt
DJAyB+pw14+8qm1GhP6eoyFLW6hKsWTGpNrkw1iQY9TJ0nh+E4vb4Iaw6osnJDS3
9KKKEahPD79qHKXctBkgxYcpN3SKoLjXuMus8eEFzeSLvjpUafQRZ+FgVTtP4u0a
fOSNf32r59yx6WmkLm/4MMN9OejkNNpQUkyZO5IDf6lKE0v/0ovBeddDjn0BNhLT
ovhHmLYKyVwOqXHbXdHqowqOllV4sAbPR8Yb8px+X5hvSmhhLh+apS6T/d7/AzMQ
CfvtlP/EyrGBFxTlQDM/ugYiHJ70V9GThTelgqHTK08BVdM6pwtXeU8InQDXfdJp
KFaMacwxjUHU+a9bw2+BXPowed+98aJ5ZHd+PVToEcZQCUvBRX6DU2M7E6W9EQ46
ZmQS2RMBRTgWAh/CM3PTra4S+X5qhi+oWWZjjRBnzC1m0KAhr4ZFtIaWL5M+o4Ty
NfF7WMI9iEDYtcCXT1KXRTJxnJuLWMfreNq/Asw0nwyHn0FWaOuWEdnhNd7DkO7p
WQlctne5gqjlpgnbdfHkmjvcQZ/RaQmUcYPVZMCQ+3NnwaTq5HmSiISgXHGsIOXY
hyKQejQJltKNDH+iAnW1P8o4t4dfIjBoswhix/ekpeRFmxhxTNS0jCs9des2QJRQ
i1Fd/yqPBRztVClGS9zTc99QZfX/6/cg1/iPtuolFssLP9YUmuVY2ooedBbR9JJr
VkBwLUu+hK7pLYlKJ0Jr6YON7iUtiWlXN3d4x+pTo8IQBR1Wm1m7pwqt2KZmlzRQ
QcHxClhb9b7xSVtqSqWRhk+lhV6p4m3DIO7f91052v20m9Dz9QgkCplpTAh8yi3k
aNeG+Ga7eAxF/luHqb0lsiNwE+F+Qm/qVtrdFKusMwzXJgJFrxfOXThBIesDfin7
6oUrPaBeg7BdXuYWBhAD3UA17okbgFgl5cO78q3MFdMk4DpEpt83UEa3NqFx58Tp
VZF1yshGy84Cqg00Y1aw1IxSajemrto+PzVLjaC726lWcKjrPEEFJw89rdXrBNvf
Bzd3tCyCo+vnp+tcRJdAQMQST3HtNFlQwe8Ted6RxAp0n5EPT+RkyCSzjVlkquYH
97kZCsrORP2fsDtjaTtInQdLkpWkd4pnpydf+IDvpMi/yDc1kz5TAdoxeRLFrNtU
phLT8qzbgaD5DkydUhRSm87n0fvn5HVUSM/1W/PI5hF9HF8g9Pq/tXrY6Xycqo6m
WJJ1LgOlLB6xboTkk/+Q7E8zfcIgf1QkV7jUphCVZeiG9PWv5n3Vmdo3qF8Y0SWb
Qx1YwATdDLDC8EnEfcECTm1iDmbzxbRpYA303Nq773AS0PrL95+bR9NxHyzpdWAl
Kr85kZ7U13Mog/PrBCaAVyfPsC72RLrEyG2SkuymiIKrrPAToNkQNVFWtG97Ph7+
dnkVrfxUbFbGYCdQDwEpHsu4gu/wM5ZrP1HZRM7zI74=
`pragma protect end_protected
