// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
fK5POmnffScG1TO7hFVDgicyVcXgaNXxoS8N6kl48LJvn7BKpm8IyyZipbu0pg048PhN7soj9KTg
TeMx1TQxCpDqq/OdE/vL3TFW5hlS5nL4c1Bo8Ewr96fBa+Q0kNScNOBRUe49Y4340v95Ks6ariMT
yeoRqEBWF86KKkroxBWDbkRyAPj6FKucjfF6SrLhgqbd6sYyYIW7DbsOvrzBJBoA+UjDdz6P0yIC
Gk3OAfevq4LHdcLbeDtlPlE+FTgVxXYdnUKwMFxu66hwaF4R6LPjmMMvG4c5UcBEe3I7H8zHVIdI
wIbBvliP/gvnGELwegyLXp9gCMiMEIlZstWctA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
2yK7DEmWx3Lak31c3pZEyZpI88qNgZS0G6CkNBJ0SQjxrK7cK7CGMk3p/kipm3D//TkTTbkcqeMO
AQDQ6b7khJia9uXFLmwwzThJNXx+B+xaKYaRvHfYk5ij+rhDhPnLNsIyFkkw/bPkMJRL6BjuA+4V
LW1RJrGu3rxXknZAHyjjOBj/CCuyIKoKVsUJap+YoAY4o9PV1Q2h1TREhzCqQCSW0Yefx1eUkcYS
LDCQ3FkzdWygEeo+4CXzEvd486wroaqWZSN4gX9OaEtEBOUbYYdwAlywy5H6SMYeCpfHhhvwmCrM
U8eh7wFC0CuFW2kx287G3rq2pyPq9TqVnfJ9QHzH9nLDJdjxNt6G4DmsuCxdKsAGDX0iASl6MYvO
q+u8uBDGAYL3roEOZsbruT0DXZ/+dtHJU/ma3kWt3Q+2cFDP90SRCtVVb0TpxVFT/OiFF9xg623J
vMWZzPO3gqCP1izRRpw5XaiAg139IbfhzkqNOT8RdF3jngykZanksZYHwirLc0SLsmzxMiGvSLty
v9nB2NidlTP7Hkk9xnNb3HUzn4+cuH7oku38F2ah3vht+Q6jnjLwJiGSuLhUYJkjZwwMZG9w8/Y7
fRIKkqZQK4mv53UcciKEqjarA6vniyoD+3Lmi+v2ARuvsTJN2QxGWB0RFxhhuC8WsgPH5+iFNCLT
1itiTn4ONyW5cXIT7i0IzuuwD7pem2GHTRDXE+MSUCnKBT/TZtl+b3HYSEkTvRfpI/fx67li6llL
B5h7i9wzHVTwMhGyzAO7hIJc0tmcAqueR5x3C7+N4g5EP2whARGm5S2lH0rZ1Oo6fQRXwAlRJWkQ
66cDPAV+gz0NFfuPe2qC4VzJT0SMcASvBZa82Suq70CAlSXbjPCgoELGRDUv/oPNaqUlJ/SEhwoC
IkKM4ZPqGyqpNy3p9/G7+wQfR/FFC3NS79zKXWM4YUntYOQ7EIXwyvD2AaBcPwiOcOE6kGcOUlzv
+6i/VpQ5/lWQxed8aKaIMs4Bz7UdNAQKx62E6oh/MWkmDAfy/GvnNp/XCkeYGgADMpZpUSwqTDjb
hi7uR8DTThGEbie+flDRSS5ZLvawYMwvF7SVpYCpqWBAybJOVatPfD6cF0ynsrhu0XpCMSZqc9lM
DowTGJ3kSFGSyy+Qbj2AfM2Q/zswwperytXrf7tf83z4h/hl9XBLO6ouQnckB4smh3nATiydtup/
pZOsTPrlPhDeQmAHsz4Vk08ud2WdrqF+mFHu8BrLhNbhLDLbTbfrRnMB2G1K8ycOM8A7sx0z5NF4
yjToeQDsjp+DjAynL/NKiVbpGTdBzN74ZX16ekZxjaLFq4N17a+1+DBn/v0rY6hPBMNL7ok5kEIE
2NwcVMRNd21xQ/LzVTmDTEvSDuB2UAzONN85wR7RJq/uZsVhD1StYpYkWp47LuolxvbPW/lTdm12
zLhOYnMKJlSPpuog64twM4tYeWsWmOZ1tprup8fcmc+MORAPekGLSXynVEejdO/+3kmsXBEUmY9/
OrPZWtyGfYXeEzoN7w6Xh82uFNuTedInjAjyEQ/D2VXQGruYctU7ChcMAYvY4qhUVvWVaoQMrr8n
Y7Z9HEau7LxSRDKhY4cRM1d4SS649EI2UZEBUcbYAoAGOkutWJ7gzFA5CuePvqBRKr8Dc5KJn45o
NdaBiECVJN2IEo/N8Eh8PvQXrLDllV6h+L4R/IqKNHZfVN6Qmzc86ZFVsEIiUqfJIr92oYVWOG9m
iA12fZkxZKor7RqqLDl4pqc2obv/pCtmaVT9jWywwOfyuDsENWBgvm9A+I7XEn/fwmsOzU7i23Fq
QBqfz8H3Ng4+YKOw+cQ9/s5mULHC4/uUgqL6UKr2hpcYgSELLaec4ciwgK03RBWwMd53Tkllq7r3
FXBb29KoBnbo+C2iI76SxAdQslNL3FnYuQC/F94Y0oTBzpw9mzIwCkuxgHDiMs/7LTxWwT1WELyg
NbMhK8QY1dFqF2y5aZDbhrUi25uAhLId8AP1ggkR2Pg+sC8twUR4Z1vyXKkWXSMyuPEAGryjuvWQ
YIkNL26IPq8cdoi8/ChyZGlej6tOh3AMXQe92/f80+GJ1ddw1sK3NGtcXODBEs3P8g2o5FzDU2vi
ehMYDEN/tXXOr9Pn07DPjR/E1sk6n4cbnLhTD5NRO7LaLZ5kfoxAa9X69/O5O/9acR3bhH3mPrAM
LQr1i8RSkUSAHQEsoV3ztBVIkyuZf4r5xOz0T+Op7yKagry32h3tFudqRhQPxRKbj+Fg42AZhKA5
cU6jfTnuv45OUQxWPGZxdxzV3U/oumHlzhb3L/hKMCSmcM9t0VhPBSZUvNilzJWIcnPGr4bnkZFq
xnI+j0cEFsDpzJ0wvL8QHtelwu6DFvvQrOQgOtzKex8vPCTMOVZbhkkf+ooUi8LLENdzSzZnxbEP
w+YnMg1X6+BMUqx650LDaK2k0sjjXVkPQRaQb9RPh+aiDSnlaEESu5jW3o31RRYlaO4jG4EKMwVq
pMPlM2I1n0g+8wUwr/4/4WhWDXFn/xm7hFKdsYGjBfwIQAE1cdGVglDi3Sn+4vq8D0y2Ayxys85R
2AHv/IbsZkjs1fZS3YleBrfxv6Lr662hyxJ2tuDHdjm1qy4g6S0zMINAMN6CKcE7td5CjwVFthuS
onUDyr9sl9kD+Hf7JaOXrPScwgzMT0GxzvS96WepyzatT9VhavdYi54TjuAIggtYUMsY7S9n7he3
ePaAJ5iHOcyx3oC1gysiJ3ToFjIPEJtS1Cujio4v+R7izwap0KtVBb0X46SrpVIt9RbU9SwlJBRS
sCYq7vSnbjjdYNFxSXPi9VpHYB5Fj+RciKEbXE8fgXob0DdU/6DPJ3VOU7B6DU3OriQMLYWvYRK6
qGR79C/+joocmQ+N+hjBD0/DXcmrYHrerauBNflP7AnvIMBIxqtFxws+qroHAxowhv4AGD6+4B0K
AbecCei2gfOKOnCprnd51DkYkQnN3SojPGKwFwgaY2GnmN7MHslkkrX6G31/IRCcGIHI2X7Stltv
MxDuID9tR6zNx5HOB40K58M28Hqcnh9yH3qz7uqINIaJGUvoU6CdAP+ggT80d/oZHE0xpCXJT+zI
+E5/zBtJp7QTS4SCaP69cvlWGX8nF6LEXJqATPAdLerD//jN5Z/TB09obsrzEcvq6TYOguOwgY8+
w61NUFpoIgF359tWtTwE8nqaa80klxIOSH0WqoHlCwOmS9gyA8B4UsxJn+sb8A9nMiCVJoZ/+dRX
2NXlztoRdQ2WmDPl8x6pAl3Cj+NYN3VERRGUPFaSlOSrFNO4IGM6wR+NCvLizJOUD9MqlUrj7pb4
q9AYWUYiSBSv7K2IihjZMeQe+DfJp+un1tuIUxgXIIupdXKDgERDSDuIz2e3KpXYk/e27L/+ukcZ
qE8IhWxGdaNvjbjXc0WBBycv5yf8Nw7fBvisQL+ur+HC5LR5LbAZozkUW2omBb9rhwdekBeVZYoY
fJ11t/LYGFvcIEtpgRWObih0bQdcJLyU+nTVmyWo4hrHKZ9prrh962WxRvYMvWw1XJFqvj4NHuWS
0VjyvqfdheALnZ3RrLLM8oKEVGaCnkPq3KKqOfVP25M6FU8gzCHCprhoxKfC/5RI9VXsCwrOeyjb
MYwJweCuXczqqOKYz8IiE7BrenUIazc6AeABDzB5S+qys8yWLxn9Z0EbcTDGS4nMLJatZTrmMAzp
h5t1RVNt8sDEfhZfITs1dlO8eSWMadAT62AIWZvrreO03dmaAUS7TEjsZg8FJk5dB8krIr1st5En
e7xre20AG7NFNlW8K+2b9f7jVInpdVMCCbl8GOJOw9pYzpqCpvOAhKdR630Una7oPABuSck6tXNT
duJm2w1iHHv6uA/9eQ9K9kEFneFM/nhnAKMTNmXqhBoZ0jeHwT7flHnUXIHiuZaoWiiRxUXSLvtW
NNDUqcO7cvYaPhekycEBNJrG4kgpKFVzpaorEDye0Ekv+y9NjcoKLj6+/FnyFSlYBVraHr4yKt9G
7eyvj2ck0xjDXPrZeKVvfad+/LmiAouYWqw4jPdHFzgGFiNl2C/0RWNxDvxqOmfwf8Rb9RuCZObz
kLF3wkefPMgkPdB2Gnk1THBIy6MMCU9i5dbaaDvewmFoFzXmCN8A4nrkw5CDtT40lWEaN0QbYTDN
v/50j3Oagi0ZtMLdhcRKSws0OOyNaJw6223eRTb9zszbmBstBB9k7GNlFQWhWrqTJokT+Nsqu/Ng
y9Vp5l3Xa2KTkYcsSNFDD2ESSqPm6gAHXaHKFIQHOrpkDSIv4b0tdXudyR71Ssw3XbQKkWfBqLUR
hwjKP/E3rNBtsb0x6rPZ0ODHqZiJB4at0IZdEQHfcLMUMEP54VcTo+YiufRSRcMSU4KtRedkR4pE
P0bdZGgft4PlYRQRslbcI8Q5qoXPfVwEPgdrYLeeg11p/rhrMif2v1N+Tq1NAiasInhGGeHxg+Im
4QkxyLNybQMCphbLO41xi2nkvFbfAUcDlFvFyGmRA9EwMNjPauatwKF0nmzuY2ywdIfaPsEWc58m
FY4ViUjHLXlNFGbgMdrLYYMifSAkMrxWZr/vRy9PuHXNOXuVmZYakzIe/OEKYtggEXAKBy7aWJ/K
9sJBamffMTf9vmf44ydK0nVJIMH6g8WjrvZvaF0sIU6flY8X2RyV0hXE6fz3bxwz8af303tAd4lo
9xXWgVbtQXhb2ZUDvxdLqUcUYyPxjWDAXCSIkxfn0mgeIWNOy6TaZjqaMCQGuhZL5Cqr1T0uk/da
xJqlT4cIDsCJIKxMDFzNavONm5SyrqV5GHVX1AZIPL+JKVsPDxH19YP168Sm17UTuFgacG9/47h8
VNsL0A++UAFrDLY08shJJVzdhpt4poOEUWQHQhuMs5ZxjonlA1aHj9ULThzxKzm4OWj+dkPuGy8N
ngDbYgOjBn1FQ+4anAqQGhrJesI6IZIKIK2oMO4GnZR41/3S8NJS5Fbzk+ScHQjgFkkEOJ2d6Tsz
dNFetnH10UygoZd0Ehzs22pTfEqMcE5CecS4JphFvpdp5RbuSYJL8upgcwboR2lXheYIK2BjEpej
r2isw3IlSRZbtAtedpk0MR9vgukyU2pp/Qe5v2lm71CL7n6zsXXLV47GJXgbPMH26qKkuliiIA8/
9LDhrL533kxaVmwUceCEf+0qgQq+kPm5AbaePH1qJzOXSkjBSmqV1UPJa5K/9327heeE7w3h+sVi
1W8IKNksAUBeDjmHez8VjeFcKLAnPRU8akJoh933Ht7r1z+iJQolDqzxxY9w2c8I39ZGM50tvavE
jIJHqDwHpHzrAJiaBHGMc0HobOzYD0DPEvI5Q+larHjORLlbZru+5sZoYdCKWDuAkAI/cDcPKOeR
c9QO8oUkEMaaNgwt7ZDyFM3vb5vXKs/gSSM9+ANb0cOwW12QUwSpQNtW7tNqTfj3GARnLt2hIoPO
SjaW54B2e/8ZCLwUjTdL74VQzz8st3/j9xvG3cAIr6R2wsvYxygYBN56fnz54d7j4VRJoFWYRLjy
pZzakc70UmJUK+joJuJH70/D0s0EXdNo+lmwN+pwFDqiMdEiukgUxxHnq6pLvDeQDkg3b3OeQ71c
Q+rtfzVWCETgwnmfoHqhmJqAKE7ZWjU7Vdaj6ZVs4/vm6pKyyabmfBZvrk3sVWIq9pqlBgauNkTB
Ya3+3Yl9APDug/CKE42YV+nTZaYWKxall48BKiCUuXIX2/M51ZyivIqCg1jgw/PBvvpRBWg9zHqY
vIOmPU/gnTdbg5ETL5SFrwjqAZBek4Y/Iky65noThKyDOGo6yheuUjx8/oNLJP8VgSgUgHweOXYm
wxCObb94qXp89w6kxOCT2bCTI6tQjKvwuKegdqY512RtelwGupG8kAHn7TAa8pbGfxiQQdXnkq/H
dgVeXfWWuKxHSvxgngei1SQkkaSuXI3LHiQgmUppb1YnC/6OZtINqaIbGcMKWAOGpicMVcQuFg7e
vS8RZ1CIKyGz1pB7ikb/Md64cP3VOmnNSr5a23wWlyPzV5cZW1LX0+a4kMSI5arl6eccW2/VriR1
QLVJjyvi7EVhLhQw7IePhZrMg/835XSYhBCnldDiait2L6f210zNoEOuivODC2hE1IbqLEV34DTQ
NIN8jC/N5fTpzkGd2q3er3gv9vvxnCCTM9pAgmS9kg3QVyqiCQwH/FDBlvZHqLStwhakXYaHLWEy
sGkVoX/gp6cHdbtvyUT3A/FMDZHP2BrEbNwvdmpDvADmgdIsX0dgDATwJ62lwlnxCFiTYjyI4Rmv
bJXEBzo1UVFQ7juvoVZJQWEKBq29u2vX33mUhhi3qVRPNxGmsAdMMBISi3fzzCgc2HcPntPGgbWi
DcR2cCy3WQHfX/tKrUEw+XNsVqjd5mnA2bN4Sy08rQvYScZouCxZ/P2H91V5Zmy04C2b9slTVdPb
MpSiYOc56ercsK1Zv3gsZb+2d2stnEmZYBpuqSBiSS58a6aWsecbdlS/UjP9zTLrP1JHjx+HXA2N
Giv97CIpvVe8Qgjmj7rx5Wdx1Tsdsn5l1yLJa6B81FEWtLn3x4AlSrn0VuK5we3AbBGqTRJY7jjk
Il0WWc11vRNAS/fS8bQSR6huWCDwV4qzz2dZVlAxilFW8BOqaraeQpp0chQDjy5U6FiH4jw5iuWd
rC16e+jkJfOsB24zS2H3oyY+JHqc8dcLQuXaq4m0kvkmzNEiKFEqYLBjaCO7IegdO/VC3YiEoekX
/SfYd5c7EXkfrVHqmKgix0LjabS+nDyCHwqtuQU6jBFuuf++SNGFW1Cn45wCcJnj8VxFYHv17RgU
7F2MC88++G/ZV00WjHMyBGSBKAVviVTWBFLLxsTP3IwPCUEMsNbF4dibyVKX9xfqPiQobghSpjsr
32fxakMVvurYGoXA51vlc4TaOjCF2dhMdFCw1TQ7aIzN6bo/+5xuAuj/r2paCVtt3KJdoJu9jI35
IP+IJgfQj3hkd8JIVbmCIYuo1mtKv9KQvKPjNO3KhMZhWqzVhnqf6SWqhGytU04bxHavyDKCmv3b
EYTaTPRSwcqfEpeZJLgj/R/iRgqvzqES14e+VPq1AzpIveEvZmlBsi2BxE+uxv4tR7Lc8Vhlx3c2
GXcqa8VCSyEWl1Z+Qy7ZBUZ8TTMpWjgfikUIK9zjyC3am8i1eSdvD2TKDXkLl8TDGH8WHXxTXQh0
mjwiPHyVenHwGzPKwbXqN5vwdFM9EQioVHKQy4u4iW6GzzAd0aVuP0C/WTr+6pFYxggeAaO10ZZX
NTGVKpZaHJMl9JZL+O3e8OLd/9w2hh5EqbxPGREoLgmEm/RYMV6ROHn7nkqTBQRZIDScZ2JGzGgC
Wzudj5YAYs9nKd7/uR235hwxql57yWsDVQU4Kr45Wa6bRVWLbdQME/Ui4bFlvvH0YtmXhZZip/qi
XBpcqYxIgmZWwlbDRTWFQHcsLlRGv6rHtuHQwUVH/42KETOvy9Nwz6EOW5F3crq6BB7r8CZZxYCI
z7US9DKz7NeJOJkD3dlFisStJcSS8u/9RXO1M60Jy9TYcAma8Rvi8G/Xk1qhJLeWyNDbZDaInr/x
06x7KPkEpAZZVNDi/en30qvap6nL/DsoqvIZbNEkY/SjGiduTrypbGTri2oggCZl42anmZhKR6oB
dfqikqtUoqAsOG8Kcm2azNfuvcVOVxzG4C6bdxFEgwxLRUoWxchNo7tQoETQ0O6VJK/nA6vlFdSf
I13uiHOTNlRH7SECpzEi4kE8AaM1XDOLDvj+wmLmx5X4V2BsFL6Z+NF91PZG2KhY9kbQN9pBlRiZ
9Nj8HWhKHGns39I9Q3lbEcwfK/rWYMyanBH52jUFIHIFsFCWNN/DusK1k9cLyd1/pe6XMLAmQu+9
rubygy8ynwO6Tkk74XPjSNPtcklBR8VGY236xCoIvPKHd2iyGyRkZi655fVbXGXPY2dSjtI53L5I
CH/uZ/J3fzUKzwvmGRZEQxEwJ2z/IU0MVqslk8DeizXBg7S+MK3EIWPUuiyrWzSebkZc7+XPoRlP
kVI5c8sUSCtf+td1z2AyzYRLHWhFLU5ZSPDi3x2IeRBWOUGjQg8ku9JBUOqcznc07yFpiraSjsXE
g8Yj1fgFD/LfgsRVLgC9z3T4zmRTY2Mw+I7rFDlKKIzjb0bL+qTFcjSxU5vLCxLO6IEQlMtuxG1N
+jLA6maMH7J/K5pH4su2DInsDwLkUhbG+INDoxCvj7y3tYYWZXOm3lBrH9GfYGSsUUR661gyA7qx
o3EYaOCk8g5lAVLhpFBqgW1eXZVt0NKjiLBPRU3gMJA1dXd7Gf4LhrnFguUUBSxgcFI1NL6cffPt
IYMKpdVEFiBrD8zVCNakHP0j+k1tlqTeu4dP2q5bRZGbjlLhct2tlaZJ92RnkQJ/ZQ7T/lbRWaGG
I1xUgU/Ibuxl+lFU4kbCynZ5YXIbwv8Oc1L835m6bIJXE9A4mIJijmjG2aT0+2Q/v7nhxnvlcdZC
Rzg9qj6KRcu6Cmsrwogc2+4ln/rhXnSCVpHAXhrTCQnJByYXuZlC8w9OPVOhAwtifKz/i1rGD1LR
GqUy1w8oU1OALzfaiDYNso3e/f6eHuIy0fFBilK3GJ0SIhhOeAvutIz8jwu80ysQrGlXNxomMbFV
U9GfF14u5jQztMfh0qdhI0hI0ZPk3OJZohlsN0qh+m0isRxo5D2n+rYtClVyfbNwMZUMLjks/Vih
e/OuY8VH3bxZLMZ8WZgNbeEqFRQQrVRPRIoZnuWhviWlJn8KVd75RuDVO983dS3Ip6mtzwBAV2JS
+9lLY+ABZblmx6NI3RSRqXgm/98tJR0B4E097BNkJQtAGpV+XzUfqfTPHmoy9f+I8swhlHp6DzrN
DCrjrPh0nx+gGhEy0QIMZ23b+Xu1c9guYDop2I/J/o2yjvs2HGYtVIAmKM6YZECVFX2bEb4WUn6B
G823Hj30SyaeTKiVlzZtAsFLnlxJYCLdfrJ3pnlXf2K0SYGkFLTda4HCkYQKHYUxdR9CT6Yb+Xj6
dBKzoFis/JgDdRHRyzMSi2k=
`pragma protect end_protected
