// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
I4JvDh42uJBjD5LzneKCmIy9fNwS4mMM0MvbQjkAYjFDLc9otpf/0EkrkEp+b5T3b5MyVVicZRFQ
A0QUtip2YxuHZgEgznguo239dTcKJvpclyp7C6xam5pNp0awAXtMJ2lrQ4TULvi25CAIKLhq/bzq
Bs8Kbjpz89tk4yfE4ExWbbB2h60XRjBa4SwfFndJsnom1gu+3XFDKjbdWGPg3FHaQJ64IPxWpXbU
hhc8L7nwjjLYvKL9nd3KWWy8dbhyV00vFQff5mvwX/5Ti8mx2uFLdSOEtyNwLiZknQv8HRqnSEt3
U+xxme/Ct82nno14PiYg+j4RdCX2xdKbu4LiSg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
OYHLSBjRRvPccYOsOsGc9yAa6w8ZV2w/suZnmGRzI2GNL2t99QgbTJPUsFIZgWngBOyJLr6J2kfi
DJ8BIthglo9VVa/+gAK8JIjrN6SDkKhqk4n75qS5F3Rwzb5S8wvJ5NqpGD6uYJERLFWf6/59aCZB
eRb0Tzb2g5sIF73CL1nqKGve6bPbr5/BjJjM/2SWtUuh2hF0dsWk5ysKwbESOOZTydFLyS3lXmjv
3wsrIdRIo+lHDRQ2us1McNnajlTua7PCK4ag56S+3GA7D9YDFobKKFrlqvN/RuBq9BsQDohKutFy
LZXYw1rZZ92avCsm9SgR93of4n9vGYS+HDYpn1fVvwBPmszH1zjKLerluWADvIR843Uq5+lIHh0u
HpwliHuG6j1tUoWPFJtzHAuzdUkmTSs7y1Hly0B8Slgv7Q9cw8P8c0hs0q9ePeW+JXVa6P8KH6v9
MLpYBa7ZtmMEsbWMB8CDTyiOMBG84fQCPsQc9jSYFkGSy7W7lfHrcDTAHQ2id7Rl5rnAttn8M/4+
ltJVLHEAdMPd3V7MZH9EmQhAlnbOHW66A5ClBsMGfYsDc8uqrEkRpgsNbeo21cPyx/3ZD5fzIvSo
kanMfiLkkvZfCfGM/DNUQAsrM36oZq6QfTLf2mdwkdu3HxkS5fhVTPe5WvRjYz5rGDentgQ2+Ef+
CpIk4tnX5iJLFU1Oqql5YeXgDkQ3ZKTQnDXnXF+WTd2Igr+iBfOuYP79ozOt8n9sYZjhCmgHIALJ
OuGHUau+Wh249Aimfjv6fJTqLQGUDsO1F2YThIPjWY6vfbHDX6EwTqfLJ7O6rC08nZ5ApI4Fesx2
vbULsg2IPQH2UDCCssHM8Y0AQz83ogg+TF28ht3HooQmet3f16xZIJy1J3M623jPPRWQn96eFqZI
xeIpPvYBHPp1t3zSWlGNxivnbZZcIldxfqxxJg/Kc4aP0du/4WPbIexikR9HvOmKYupC6NVkUQVl
rKSxOp/h2p7YGKgerfFrFNDr1qhMIC9treQ4BQJH86n9YedslEptVP3+qUTf1X8gOIi/EHZllS+a
xN2kglFvyLJZCTVsan7vvrX5yYg2J4h55j2pe2lsYaE23BSabnOaHKvFoh3TJX2Vj+IVA7J0bvK0
le6fArJWlJnqPurrFgfmH9jO6UMGjtEmQKCWTxG/GDcKk6KNE0H1dS4cy0BC51MKthakfEqvi/6O
BdOKaxOLQ1IsRn2xpvaGAZgzra2+eaL1Mw0kT0gC2HjcEMiBmccgSSBnujXgww00TXwFs58M80Ef
AGekv7GVfkeTeMrMYZn8uAaK2WC9rWAgmJgPQCjplaYL3SuqZSOyD55X4wZq9g38jr+tRukp8uJf
T0f8BYLQnqGrJz9K6Jtz110Iz29ayxlNu9JiuuiiJonxu63Kc8HS+jSGRd/vRIjVL0s2Uspwremc
zvFLBBk8Pvtz7FYJ6MYnjr41fLhu1sxSfIGU8sTeHA7u97qnMnAUnb/xxAJjdhVevUZk3l2AhUti
4STRyOAA+TymvFKcOVHlgIifcvaBbCruSGup8NnuGy93R9XOUd/Chji9j4cxdRZesN0yxvUX8382
teD/pH6xNVR5ATg6ESf0OW/AT70gOiO1Eq91sD2F2ClXwhqFUCnM2jdCObEYB+xT24YrsuoBHSKx
YVGszqBwrD+Yv/NkswQUI1hBpzPQiviyt4suP2KAt2XGAS8pNa+LU8XFpxgUHdjb/IWEEuUKOPj0
9s/WJwFVFfEhwXBtH8KKh3uU2nNwDxCB2tNIFHbpJ45MvPRbOVEaSHah3AMwjbLR2j7x4YoNpBBD
sCPJUHzRSA1W2oUhpkL93xkaR3sK6v+W05tSUBBbegVWHTDgCXTmNpwxquqCSXn6AfQDu9cZaCaD
YWjI4Ng6f8p6La6uEFraB9icsvIu/n9atDFbUck5QSe8PuTtVnzCG+LU3MadCyRl0YU5Q6TQTM/q
Rh/t+b81t5cdniugTx8MwIA0mxl5DeZPpY+tGGvVzXS0HD3qiU9CjhUmyRrs3ttQXCmtyK4mWRG/
HX/erW0XW0feEjMOC0P9cOFNxepuHSL3ZXO0N1ZC+EnrUODCX7og1o1XTLBYpzVJoKLKcOdpSWkL
hD7a1DwWklJ4BOVKWWbvoBZYy6LUJS+mi0uimKNiPol1D7bG189nC5ZD0Ag2ZJXLu5G2IWbRx0fi
B43mp7Ypk7s7SyR1S6arIcrY5FTzlOTfM8wbvHRZI9NcB0FQnbBVjUKzM6/ziZXPDubOauNjdSxT
Y4GZ60hssKwJ6gnYBiDsi0iYgsaWzrX0K24zz42UKMHH4IZW0w2b8uz1M3CUSYT5ebaZwnFBRCe8
cyAgPrzF1EUAlX8jvfcsdOIhbL7kUqBkNwAUgwDrCRYmOb0B5VQFL3hr6CF407jhzqxGqt+m+Etc
YGyDy2MikfGCE1z+/dlkwBnBCabxsDM3LI8Y3XpEI13l5R9hqd7sntuIxnmcSYhXjlWNXXuZWL2j
gPEGUeYiMs50QoiZ3Z+1EIaQxaf5lek82rIMqTC8DHHUhhk2VgC26ad399bqnalq9Ix2nNUeP50E
YA4Yyd21oHNVwtvelNjTJ5vpJy0ZJWBHsteYVT10KRX/2zwGQ+Em+GmmLEDg0zRHPw6GQWXaOe3w
lDq36OZN+ia2hA8t4wTYZTfJSl1lPYsPRkkEm71iN0a8kPAhDhE6xaAHbkS0CToaGwAIW0PoBUq5
Yo2G3ISwNQeUYBzts+17XZn4nf9/T1qh5aKHWMXqLBNl37/tCi+Z+pMDUVCAbLQ9RfFym1n9XHAQ
vGN0LofOqst0+PI8JW+hZvbvCv6YYQuz48ZWpoDSgMHw2AXQjhPB1+Loq7ToKyCnKlf9gHBKHEM1
B8542sVf8SKCgY1ey8ltUnU7g7FD9QTh23lLwxQjA2EwiVmUW/oDyXASZ2FfY5eDCBYwYRjQ3v03
Z0Au2oJXwJqQxnm8hOcx6CyR4Y++WsHmpVAg53dJKNiwEuznBmrmoKEKKzRg+Lg9wM7jHWi1b4eg
elYbI2mJPe4FF+qD+8mzV9SRWgZNdUccRkxl7AMj7ZLEWnJH2dd2Tamijt44kaqpj0z0W+saK3uk
1x8do29+eQI6PixRSKY3IaN0089nL/cRhBOiCRBn6DvL+GFiRc4I81xmUHXfpvhXbwy2Anged2yN
xrj1GrNqjJEJ32euLKIqVyDaqqmD8O9W9iuq0k5FWSNOANabiDu8j/djbif2LqQOhVbrLRS45IoN
YaUEBZG+5q7fyJnyseeJvDRe28HyN8smulefpRW6dGzvSH1HyPHqjp8bUfHZGJ9ItNOVe2URUOe8
Z3fk8vEQWnOMRW+WRcfrlBg37R9q49AN0tE40/1YK8q344lKndI8odgWSDNwxjDKJptvItfLScMl
/+iA/ldcKNUJiQ3/oPwEaXLMPZyMG74+5d4f2sPT6ceUPCm7keMkuvasBWTQlPDWxrb2mDQy1nEv
zULx45zGyIWk/4k5eMn34p4IEejLhjtWEy7uEJztjT9dD7o5q7jkMxUIhpx2QijL7+UtiPJY/y77
0cgHSYgh6pkk81lzXsW3qlRmKRGnE17C9opbeb9ai9DPl6VH+WF/SWmb6u36D9l1et+uXVnGiCAc
Jrci1R+aL5YeBAscKwx70G4U9fSsM5reB+38MMzjQ8dNTh5mbHmgAlpWFDcWQxO8e0ewUGemKYzb
YcaGkUmS7D0tycvshHRjG+rllJf3bwqXqWQ7AEv/5vt9619R7Zyxye9c9bOnjof18U77WwlP+eB1
Upfyr+7DoyP7cRc1tcevfuoQZrM2lLFMto1CJWrDv2G8W6Jcp+up1hkpPpGlsy5I8nlYthcq9Ef9
NMOT5qaN92zaOz6UZgERNevoY89+5GAQqc8Y6gIhGrUizJ6witVvtVwcljupyNgp2blyqlUK0oIG
am0Zw3KB3Ojoc3TCGZFzikJrJEZQ1RmgmBPP2drqJd+z8Egl/o1NuEHUkGl+L/DfEv8Rc6eMcR4l
8bEwMytDCyGqdHOK/wwsR4awvjUoRQFlADF+1b7J6u0QUrRIfl449G5FCY1ZMj7zoKJCpwsaBeEf
DSZBR6M7RArbMaHa4pUhTCSTMNXmqGj1is30IGu31sWbWVDsTY533+4MncG7B2QknsZcMXyjQsoA
1D/ztAYXnzA1mwCL45JL2PMSBQcg5C/4KjEP/ddPsU682pgUtnS6ifcX/grKgrGLolCxOb39aWar
p+C61iCtRmn1qoo2XE61cy0ncSKaOdOigHOc61hQBXb40P5q061QO0u4zaP+D74d1PUWVMSnFMnz
jFd1Z+pv7EnZ5S6vusDwBZ21b99ghyhJw7vbI3tnnvFvGwTdd5tKtPLyyXpSuvMD6XBOTBO/luDi
LgsPFvPwBftBHABEDfmDXnzRpWloqG1Z3l1fLVpHD0eW0XoEWWVj5XOYs+m0YidXxoNq2uOfLbKt
WqCrc6UCy47npsRvlPX41ehOJ9AJ7Q9ty6vfoPqQ5s1g/U9+RUH0fD6aam/zTy+30J/DktM7wYyS
j+4/hcNTsUIb/7la86PDALomW1m7khBKeozqIrQIGbQh7xn5vF8RV94pFI57yAjBzKOVIP3lNREH
5dydrRT19U6r7Cjm1r0b3NIE+pmqEa7BypaGoRrr9zHDIaq02F/xtgnDrUdRMI3HKKNnhCOfAKmq
dtVt+IEdBi1ysZJaWvgfrH3oyRBoqN2sx1aLMo9NggIJFCE7dgUFMrj7oU3QoUma78qgVLe1YmiQ
tPgWZJt/V2528fsfG0EknjhTy0HxVe0m6vt3vrMeHb2z03zJLK+mJ6zSf+uHRyQTI1c2d4klF4Ye
iIYfvNYdw2RIB4LU+b4bxtT7FzVSZd53f53elb/oszn9/MHyUZJFDLNSh1MewubczQb8Q/ARtgpn
IsF4nzo2iMDaaFAKXAYvJCzEPuxrL6/DdHNThiz1XtK5Vb5p8mZSNbGrwOBgd2Y1/JdWxxDOY/ki
xSvua8MZ8fF3b9P7z9zhrFnxRkNzKxEn4Lv76nyc/eWrSgaMmvikeInJ0VY60zgEXy/9hg+Xh+lW
4FeGWnHIPc4YyLQzMiBk1PLUxNGbk8qsxID6GXE+FRXLEpM2EIqmCIkrnkvHas8UX7PS4vlmhBMs
VwoNIi+ONf7YNbgmT1m3xf6sfBZc65JIvs5ffVzFPXmtjrsQw28kunPKiqtN4AYrDKK9QEEJnk49
ehGfJnz5cyZEqPZ1pduRt5pNXrckZbBXJotGlRIy2JYAZ3Gkkd+SV77aPqkTGr46nFJP8b2V6psk
dN1dTfpUBTzrfQsXttrr+iccrTohKtbmryXB1D8pJuJMc/VnoZxnRT1BNInK1w0O1libVCebrCzf
o8hqBR9ar2KRk70sAQVbp+4Tkdl3KkMvSIiHHgYi0owBUw0tPAbhm9Yzn5YX3iOk4M1XShxn2jSM
NWnaaBme/g+5ltQwo5GZCbQoFOT2ejHkkTd2KkuOsr101GXwNuLKqPEDAXLGwihpeWX3SdZiQZND
xnTYOvbzLM7zhCgFx6umnKisdJKPpWleP4uUEbSJOK1XilymfWxtYc4VTBUgI5xculYG7PCCDvDe
323BIV9aIB4i2nEDeVbnZIir6hM7TQzZBCJ7+zYsPb/Kr/iUobtl7eiJEfi+wUDOfxJbZIKWs7Vp
36RcT0x4yuIQMPA0qLXzBoC+oISj57YQu4eW1lFEJvZRbvLwcZnMBQz34J7ebouhwJkBE5hy8NBT
SidH7Q06RyiK9Koh1nOgElp0LmlcNi4fmWATbusiotgVHiwGB0xNfms9iOgULNqARrlZz4er6w6U
bNQ8kLqpHU6QtjSFazI092pR5X30uI2cnNyVBdBVfS4aXP3qqCo47ohPgLKMeWwCtq08r7rMgLgg
GtxGoecpms2vnHMwrSxwAlaIWLSiFqkvb6grLH5VI+p9y/u0DY8rmA7pUoFm/d781ptLGHbbssRa
LwaJ3zc/QS0fsRT7Vfa7eU6o1q8PK+m4JHExRGVR9/Mj5OBgwT/tCN8OhQsG4if1eimpjtaJdH65
VKVDc9E+oXrryro93kEU0zQQh87356dlctigxBVGhF0tEdAq267rKIsHQ5JwOxIRSbxuosWndiWI
kDleBj3ZZAmmjRifACyEWBqAjqy5N3baYXuTooswZVzGdETBR/RXXxeoNfaL2fpvJDAw8aIZxVQg
bHHIH/JTgu+ZRn1ReEbeSfvzCIFbjxgGC4iV5EzlaWUyk0V3rH+2lqIbFbNMeCNxDU8ph53W6/tQ
+UEXobn5M4y833P3Lt31VzMQR/iVN9C51eyR1CLa90DEYji9xv/KUmgJuGrt0HyattQhHtFN0e/r
tT6FHVul5Xi/VJf4t+5uyCNXsFRDGUXZ05Tta3zunm3k1eKh+e34w0SF5NfBRaVXVXXj6YJoQ7eL
s2bDGTXHGQxD1XNC2J/vHZxa77A8ga9AWLQYPnGdUMow2ylCdQ1O7f6vIZqrwEWFcSymbZ9vMs3r
yCz2Ra/miKp+zw1dXQBlL4EM9Ov1MBkxbX2gGkoy/u6M27KRFgUaPDvr++N+5/Jy6/mSIO/x4gx9
62FlNawvF46GEuTBeHAV1hd4U2mBDw2pJfCmr/Ooh9Josc2rnZAshN3kQRcURAjtPTM4UNdr7JS5
c9r4aQA9RoYEUA29OeyPzmbiMSdVWIaGlOoNST7x64HL3QbKD94JjbjEj6A5Z/H5QlrQBK0gy6wp
E6fXnfb0elzeqX9aY1pREm3VsrujobpJc8OBqHTTqgsSltz6cFttjYsAWM56d75X9c7L9hzIrWFQ
0MIt0/W0wpKl8b2V6c2ZkPkIjBudQk/TnyL45/eCG+QPLlY3ElznIZx+8GMML7+XoQtfSjr4ZuGh
ItrkwTEMwxVr843ZxpNN1NxKItfTtFy8N3PAZM8wM72zGPcdBxnEnvl5gx4iEoxTRPWAGQSY+O3/
OhtrJsK78r6t3bpXaAbtex84KCn1fVJPJ56utiyyt+Tn1LK8tuefZcxFxH3P6gjJVnyoH0b6ytD+
4X+DFKN+GAtqn34KUBLI/qPnPaInzWrHCnNn1s8CoDCEVW+spFWHWKUcvkRGSMToEavoI7rcaBST
haW9E7xdL4RLvR+irwWSIhhbEAWPf9YjkhtyfBRK/Rfgqxyv34MaGZ48vHUjtS69DdrzIyHe1OPy
U67C2Tux8tW+BblDLC3HUWz2WqmFDuzN7CeIXqb2oQ1qPtI6iBBIg4W6OKCjbT3awZYmxQCAeIP5
fLxc9KEelkooFz1X83qiRITpzpu6ojlCRlac3Wpt0IMNbCtVXRXv04/A7rb/paKGOiQlnrIKji3s
WoVjrNaYy+rNI7lcX/f/0w4f7mfInCEgTegtT9zlkevk/2LmUOnulqYfcantH3soGcEX6WUItbzD
3oQaMhHRzpswq6tn78I/2NMXto0eWG3ZLr8ak6ambDIrsfJEpOXFIIjro/iN3uHLDTeRKW2pNIA6
1Wy8S9h+LWBAHoHPY0j1plWrU94Hfg2MEJAvkAVO9jX1xrOMU6LPwS+Mo1KuH/5D16syEho8kxx0
oghxgx3aWvdFkb2/W4oUappEezEhKd/VzA1pDlOT8f84tmHt4WQgotUiNGuAHuQ60NXaKwiMoXaF
clZgNCQonQ22TOaiMuwt1s+VaQlfj+OkcEg20a3WZwC7lY940CH8mX+QxYqsPZbQrJUd+SzZ9GW4
hWhi+kXouNt/8mC1WITyIfavzQluVA+YX7vNI9/5SjLhmA8mQ4xVXz3QqquiOHXuvY/1mgd4gqIi
v8nt9Hyd0FU6905huOUTZimIkYF/GRSFc1elcfFzvooD5gH1Ip6gVkFoYXZ3GcZkDC1OrRczs9hT
+aZmmIPWoM9A3NTBp3eCup/Z7kWx/WycBCjzdMcs5rjmnslL31zJqR9DOSfw8xv0wvd9XX5QD5bo
CypaW4/jBiNrtwno8S9EQRRRhxKKFNvFzWWy+EAcvXmg2nsvb/t3NLbFz02c5sI6dcrAaktFm1Sj
2F+z7k5YOIpsDyQL2gq7YM6zROoT+XhYBUsi6vX07SzGJc1tFeVVu5mxZgpfysMNHCu0FCubRmgP
nviN8XICbnTHCRvkUxSqZEa2n+MOr7X0xD5Ovt5Jdh0rWAhH55x2U2u04C2YjNcWSd6QN43iGm/R
EDmwdrPz3vJH/LouV6YDgHF0KQXwGt9JvZ2vNRPSqJrllAdHwdIT7eOFK35d2jjuOH2wSnCwbrxI
GVbu2995P/4IdmmwoBXPdZeujtCbjTysRaFAyiTCLGC+GQ/udntmvQE+kUACsBXVwG2l7hvD3Swf
GUzYXPgBJ2PWr/BcwQy2YRjO9WISjHmQmlBi7tiYz5UWP6ENIMgVtsoYAt+rJQuywCz5PwXfTtLM
Ipq4YwNTgcBgkxePZCJ8HsqXJeoiqcUy1c3BI4RTM1+YyBCELWaDu0TPA7WZTD9zGG5OHDpmXtVd
eHZiHwWEKr6JKhDH/NVTs5lvP1OX1ymbDDE63TFQ6Al1H2a8g0NG7+ibpp7uE0hMLWbjrN4ckR6D
w0ucy/hffoYkgZC1kRITECv5pqKpAAw6n2pZfy07Dxfq2xdkDf9zQJSurMQrO41re/GmXe3jLeJf
iAj3GE/5c3Zzkbloar1EsNVxziB8A6hE6ipbbySr8iRWq96sM75HjOsk5auhW2GH8qSRtIxU0eeu
dBvdYsqbf/ea0WmYnoYm5xmshbjnn/nDa14tmT8XT0SQGHEw+8cK5naqlahbxvQISUQk/T76ELJF
KTMop/+qTkMbxfCfF1hq/5KcBjquubL40WHzgy1pu0sumU7VWNVOELn03GcNWdvjnM6EjJkMvFvb
VXzHDO15JGW0O9lb8V/5+WQ8R34MzTgX8OWWCrLcqht0Dh06Fbu3yy77xhbcl1tKi5+S3NI+2+3W
XNQd88Wi3lqkz8ruPGDnDbm3slmRR1TDslZ8NURfRYCKHLXApYL1yUZmabmIezcp87dwrDP3iFjr
/72RbpCeWPrco7cNeXENxtT+tP+IdHwehtNh6oiZIDjxqBPDIxgCVUPmwJKCPMnc+J7YWLUPINZ7
tZcMIXHzTq4I0NHfgQ+Lbqd/x4lgttRs2mTgwJVPmreHkFS6qEyCoqoA9PGICkzLM6aS2LGHSq8C
T/gJsRKnFBXdkKL5NQ3QQJ5PbCdFnIVEZQq2A4JHHEPKJfxXqwnaaMTIs/LEAwq9qCwEVUakW6Ag
q74uJrnsXTWs70SUz5GJFTi+OHebsIfc9DeTJGyk430GIbljV2WgN1+JwiUfDJNf8tRu7tD/rXLM
Z698nHXPw/molUI4KBgKlxMl0+zrbwYkExhdg6H3YWpJvchSPUoQ4VA0WctfUF198+g4pBMHLJ13
ohB+0ue2ZYIp2mPSYfXbfuLBqOth6RQy2/vnv/pQxTNQaZ1j8ELnecs9p/y+us+W0GsowHkEjxsy
ChLeQ/HX+vWXG4a3gxVzcpEBJpKO86+C0TJsfjobg7bTGNTgTumTYMXk5CH4PUkQaQp8mIIEdnEQ
Jo6yooXK5ID6KpShq4g+JiW96zfXCntcYKwQ2cBpjFcXX0ORImyQspcFUCZa4LrBtfp8YFxXyj4F
Np4KbTuTkP+wkodxf1gX88swx7L2WV+gnFuuEWdYqqS2SYmkkyCDOInbQSHNwth2vFtyeuGPqKKa
xvYeOnPfTvjVVaRuikUa3gQ8CR4nr6U4khRJkU75+xKhVCosBgTWYk4q6F/E34TuKoA7FoVuuUnT
uxdP6ws0SjH6rQG2GFrKgSEjfEqLX48RZ8SPeWX5nRHWD9wW2aEZvmqy4cA/8Wr4amub+gGrEUob
4l9Yc9WzKqif9xiCP3nbL43uNCCmSLzIXEdMfXMWvO1s0ZquNj9YRh6TzFDb/7G4qnr/gd1UgHjE
BX12VYx9NdRZxY5vej4DA/lr55XunxuhnNb00KdubwfYj1J8Z0DWZdqG0KwOqKh4ZooaTNTNylX0
SMowczeP/xCyjSRqk40IMM1p8A+dbNKay4mqkdA8c6fItd9wouWpqCgg4BgLKjbZ112vevoX+zhf
965NVD1rPJ7it0ADa+jBrvXSZatPpyIgvlWeex6L+pcZ5QgxmLhZI3ABYn6BOV7UmsW80OhCWSKy
kkqCDGzd1b7CusTLDg1fOJ3g0hjgrUVsugbYMDox0yYtB2J8LYlUwEOc7Iv0Uh1PrqMcfePGkppa
3otLN3WTA3bOPVNbSo60T8MM0nrZguiMxaxgtO77jLC1LNxMVTT8b+llUDQQ2mH2UHwpsIROY0J+
1FNmFVjNnqePepMloA6OOfXXaLTGCeWAHx9BOl9f/p9f6PH91elS/JdxYLCPUjQ0vMRyt8N+K5TJ
FWIVwgXV3Hs9DQyeqBHKlmIquhzLYS7z8Za8H7vrkRCpZfj1QFFv5P2jUJUsGMEArhYWW06J5E3y
vU4SHnpRNOD/U7d2UZbKkF2YysPlwd+zfQmPWH6vwyGaLMKp57MlhmekDr6PThefd03kz2l2GN82
eCHiX5ah1iBelWA2IpTW7oYvPOhhRe05OMW5cPwUxh+x0cZIOT7SDA6mYERfnK4eG1j6cRDFSQvE
Qf835b5ShRLyVH27BXE7f7spvnHRuFNe2Oe72ewXzMgm16ErbB1TEdqBHCU0UO1yg7SaYEYgVZwa
wqP6UOE8VgcJb5vqklXyEzFa34JWla2l3VnlMiOLWu3vcEqN67/OdFCvhflrUelRZ6WF7jdL6fQa
q03DfIMVF1uLG7qT/IIYUb8QqmOqnPFLjzxCfSLnjh2IYp8OemRrVoOSgY7sJQitqpw0LG7O29jk
PaW0K+/YzcuUTbDp+dLjC25ug79I918vXTmQfjNJ8vKQ/9bBEuBHaCwz7yFlKA3Hb8ip3SzksJ9m
VltxCPoLIB7+wn/dgwhs7Nyq2aqukNTngO3Lze7C4i4rVAHqg/B3dqx+sQZ0xulQ51gpa2g/o0bv
+2Sosf/ZnJy4p+ohrwMNNTz24LE32nJoBbgV5uxpMMIM2IF9NMuKrKPQZKimWuwdaaFS0/xzd9cq
R0AXSf6za/xreAqbOkz1P6GExTxkBHH8mNiBUxkTK10GVafHPxW47ydYO/tVi0RvEjOBG5uzj8kK
YPt96CRYD2zTOJHURqc8FAlydtHS6eQ/jxUvdh3HDJUB0R0l+s97/vdQcrp5owOT3FA0Rvbu6xOx
q8Qtn7x4pFKmBd6l5UAFkA1yX/GRJ65u9Y3LR1GACG3S6XimGMTKOmjcM4wGOo7ffepadGei5VIY
346o5pZi+bM4lRV1qC6lzrn2Q7KTH1Y8pz5HJPTbcPP5crJ/G8K0rTQbHS3raymupWeYleI/2KJk
ET9phR8939K9iaPpsgdh5P7VgZggPIlrPh/UYSW6l9Hy+rv48HPsxFqgSUWfY+X+ykhFIOjbZTlA
4khUpkCc59uQSW39ZBDijAICLwRHr0otKk77aCnyHHoB72fW3vPvfKK2CFTqNpaIBE9WA4mYu2Xk
8pGUHF5R8k9H78oYaliOfWo/uOAq8oawC6vScARBR6vzdnWbqGgeFD9A1+8yrbgmL5P7ThWD0pQ8
jNnTZwOfzQXMR/Wk+MrV9OKchd/7yLsIEcPSbRHECWcrr+VoI/kc2AuiTiroCw8+FPsM3XVZQBMy
R89lt7uANp2YQf6h9RL3zENOgO/RLKQPVuniUjWf+PuHjMgYNCWBigtd/VVzoGG0RWHYIPq5iYqt
wPiHOoK5+j2y+NPJr1AVgDsemMy2YE9PX95yKm4/BcDDZTI+Y81r8rUsAr/opp7Jhyw9F/ApQwYF
+fLorYjsBnDxBjL2HEuo5SB5xR3Lx/w7dPsSI0OJ+ZpwulvWlM7S6b0PfHCRTUmZpoUdthWMvV8G
qfasxmHyUxYF89DE/ylURGswirOA3v0osa6WssH2Jvr/2n8aBjqo5RJTPiLYTIwSg0MRWnRlEXzY
xH411vFKoSMgIcw/TRn+bpiZRupK/wF9dSh+04QF2Uuz+7kU+tcGu9t3P/z2QN+jEclzqQWDqagN
T1ICbWXvT87eR5JcFFhqRR9BdpI4wwbOfSNQDMzCzPjzqWinUckNLLD1sffAgZcRh3z+vfvFYkjn
UOD9aVhskUdK+u9HPh9X61Zby7S234vSRRF8EM4cf2a0WwwNWNkUENL1N7FVt+xgJydX7PZJft3c
MfFaHUPqJ+yJxwWjAAZGvgqbGUIwOkNg/oRD7ndygI7vMo75CyGwRkiYIGSkP+vdLe+4BJhsXSmm
pzrPZ5F2FCG3Z6M0lPFaKpgq4vzyMijhIC+s+RuyJM3/K6y6uww+yunM3uppkqo5Jri91wxbZYmv
nRO6aWUIfmwAhPmEG/X3XFAZzd6ntc1UI4b2kVo1MQaJJpQ6SIOnAACaVAQWt9S9ij2W9lFmgAU6
SQXxi3IfXVicmvQBGBYu3Cutz6UY6DnJl1OrmIlJAg+o7t0mbVP0eHBhanEiKufBEd0dA+sMm3b4
S7Hl21rYV3IhFrnIabS9DRdia6Pgw2hCJqB+qaida3W2WvW7EV7GQSCh/usyHLlvuEiT1geQLjde
hY/+B7jpHhKcp4oEGa7Z+d7RxDdLgPEo/0y25jPfk1LBfIXtIymhQOF/OIxxPeLSOpxe6aLLmHeR
o2o4dyIpo58WHT6HVMesRyKSmZ97ORDaOvMHXfBPzQLYD7pg8nRdDuDy17xEftLf+WgPahjTBq0Z
CzV9jLe4oq3wEHCfui6KCbk3uv2ESqfpC2HCsxbgg319Q9wCVodBz9rzscnEcX8WQpB2UYomMUSc
ahyafZqiG9tR+KWtkgwJNZQrOpvunZlCDY3qdBQ8AHjES+BtdRnLJiDelEO3SdrVaeqanIm5gGE+
OJNKmbkvvyQVPMKDoHDiCEhYMd98eRh5qgVFsFvYWCV1Ek8GsOSFBWg37uW7FbVvF5zguV6RxBvq
0nha0H+bJpz0nY7KVaza7ZqPm0xmp1T9y0rE3F7Hw0yhchMr/H4EX6GWk/+OUu89d8PzUdjGShHU
5pAmZL6SAuF5tLYIR8hEJGZlbB0RDcAcY01dmb5/UOWvkryaH38Naih1p4cFNdXBqP5Xkr6ctxTP
ooWXM5A3rf65MKOlPj3W0d956jo3MMh2vxCPDkGsz0ahyhPLOJ9sB/4JG3z+ojP+YM/ZksxqhZ5a
035G0BULJSXyHH/L07pod1KDr1/uvtO4HDKpeFZDj+toh0MPQoFzVwubxB4JZNE/jJWXSqfOaacM
JLn1YaM1ipaRi/7cJRAXwj2wp/f7msZYNNWcm8io4un1DKZhNE78vyzIqnf84zQg/3SSQ8YSa3yy
hLbjywuKegQ0twaZcij1fOtpnNBj7NyUgij0kXLIjoVScJssF06jZLZUzour2sKtnTbiFI9MGO6w
qLbTNk7LrN0ODuBTWkeUsR0BNjscxb/MtohT8JhBlefS9qzNCteja1MucqOsb592gH0Ru0Ju2sFG
gtJK6InDPghwU8pIJEegOI7j0sgmYQJ+vOeytQPXuNuvde6I37dAxdtbfro4quTNeHeNSa+a3aYQ
+RfWkey3nzf1luif98RD/6rsGec1MVKgFl5iiyYW0bcASz1EFeSJtXDIKtjAOAAymIzQG/lOeM4q
U8ruXtwo9wPXA3bEvuH6VWLErr1D2cBaZF7/EDK2+rSC5rmENBiAQ2hpWZIEl7QdRUKoZvo/8L6j
ujmgiJfIPQScggj5CzrFHel1x9R8eT8VBDeN70VJIZGBHgkb8Sp2eM3VOJ/y1j01l4dVLlhZliPG
U1CPgb3FtxM5MxAOQfePGTeEmL2K242q6/jKJgQx9PbrleoicT62emVhW8S5ExIAnsEOdAlHe12y
3FkxjJm3iIOq63XUciB8M5kjIv2dJHlYZ/dNglGzDBz0odNQxDmYA8K28HFbcHW0p932lYlDVLls
xbbMFIi9crmWdaDopLYyfc2WTO0Yz79nKpMiPZUHHtLYPhKx7ocQi83TuwP7YLGShftWMaf2duOf
axGLDOVZ8bPXcGOvj5mh6l5N84JezZlYSY/5v+bX23N6uDItfruckP3JpdPfdFWLc5bI/VNswrLT
sAmWTgjkxJj5Axqzlu5b8FGgdq8Li/ZVYypfU6zIkKUiFFMmW2uD3CfHHWXt/67CjlHlpxSr87yT
/7+Sw0C+xkBmyO7ibAaR9rWVSYgNohUcUktUXi6SEawJl6q/ev1ptILOWJF3vmUT/fnAaWbKnewt
t19uGjN1pq3DtdJAYV+5zVs0jpS1WLx8nxHzb45yKciIUZQAsDfficmmZb6gY5UC02HzksDFR/ks
98ENC4ti+zjLELBMay3AKHwKnvPbjkTSMy2wkT+aWrVofcbFOrcILq4OF78Q8XFz+MoxTcXWADHT
Jf4DNZTAkYInlJh1owmnp/Kk4Zc5sbAudzQzgBgKQfx4nQr5M1Xmks4O2zgOQh+08t3zMzMyVttH
auk8ijel4RZNTgu6tiLV1pzWNdCo0pDCF8EyphffGzGOH4xShX/vlDEaVU8Bfq5saooCkGrLbj6s
/nwj0bU8jaJRE7WMBt9K/QmIXg3RspkdI57EeQzFejyeh//JhaqYdfqMPKJ0Jm35OARuEOtRm7R3
bh3nvhCxooN5QoUXD5Bx6NxnfHE3UyKIZPK5a9jiQVtDsDNRuroEpXE/EkBW5XEwvPoXrTxI4XwL
fly4BseXxAFZwhc7DEOxit1s3EQqtqlhvc2z41farTBKatoD+ZmYS6sUEQWwdSzAKzaE53S/qqvv
Hz7ODFL5CvtTuOlJ03R5Fl+DxA7YS5ZTbLOO8PJO50BxuJPS/LLk1gal3b6Mxn2A/+rP9Vt1CrIk
be0l9WYsEI+EzulxwLDbx7fDSx1dRK/KH2Wq1RY21wUpv6LSvRm4boJAG2LRSMDDYuTG5VCuyuk6
SwtSLqm3F2vF5G/2A1oX+w0/a8RI7sSfS14Uuc9tyoBpQJm3YkRe3xOUHrTVxyYjAY5umva6lRZH
cqjhKrLBGnJg85MaDwtjLGbPV7uc64FUGB35t+31oIrwX6oWeFunOXTKXJCcuG0hcPhDibooixnD
bHsxxIGpXmnp4m78O9KKkV8toDGloIbT/YqceTpXSUbqOH/6uJf8bkouZ/RqrjbgVg2fEcO+adfR
xvblv2gHGQzlz3vu7AcVifBLXOhFb4MZjzhW5XVi8Oa2CXHoMju8Qnilpcp5KeS+sxZBvdqP65Ax
uGHSp1rZrN7o9uqaznPrzyTI7n2SFJVGKYICLv4Fpp+6Hx1wFD2rIA0WLcA7wJd7znmbWkjPLV37
oIktLFZFJZvBKBBc/BeZng6PB134j7GNQyDhuz+Fay7MbPQzWLUyBWeweKqTd80t+wUhEpH3jXXT
IBxpo2S4SjPGTbpNAmxR1f09GMgNhu8XFEikXMtJ+B2xXIWUOCfTqlf5SrIoTQUBTb9qeNyAENJf
feHAg9UDZCQUF5P6+VoxV5epabe2FGyAaVDcbeK5OEUehzBNjBeXEN0J3JMuNbSzhIL+H9nAa76u
jg0UpzQ5J31aMXP92Ue9dvhNiDqvEETJS1KB8BMoT6FyaDWOyiaRO2KJJzMiNEtbVHM3i8CzpK7Z
tncGqP/y139jG0J3PNuFKtyb2bAz4l/HwKb3Ez5elEzJXDsK+uah2YsQJudVgmO8tdTN/lBJpEDf
erB6errFVJNgscH4CPoMJAQuqIdmzp870wV2Ymt3yAB8OCbwU39Aax9JXp1wbtkzGEBebgGnWl9g
v8tHW3xr4U3PNllwF19M4uTnNmzfoGVlWKDmwxLgSZ4xmMut+wLHSZxZAwFTUepev5iXsoQbopik
GYzJsD/1eBSArsHu4NmjijB+yCDVg+Z3DgxRXcMD+B/teDzjx+PrsuxUvz+5HEFmi/BM5VeoUM3M
EpJG2InBUVqcwxS5/1UcoQjuEG9URStHqiI2YUcKvshNjAIt6cNryFL84IeXdt4i0OQY9xNyE2kG
G6McspsAOvU8HT7mgZYgpvw6GfXTGVqCwDTCqpBH9udeR9V4ubeeqtmwxaJ7BTHZ6xux2ghSw2at
7KxptqdMwM/nYFf40Nqdhv2IQU6Yv0gUwu6/QPcz06VKf3IdaQ+plZSSZ4DPd+CQpg2EjzzXC17V
4hYKQX5j7f9so06r37hLqy2YjTd6vHpgbFPoG8/qfCNShVPsxPtpBwsYqNQiJDvsmssSlj6mioJ3
py4TZLDR2L7sFf0u7Rn02zlVx8bfPqrxEZzYWq9ICaiiiRbkXYOUeYOW+T7fo2ecfGdCUj+JJdVQ
Xc6XsLubAbFdx+17wQmMXOj1Q+q43pJixmFtbgP0f7Ve1NorEF1sVYdznt3ZXXMZsxgX3JBDG5y2
fTJCUWWeQzJ3wvUARAvbDpPWtthSQ3vAsvEwNPmH/eqWjHBsVH30RMYapyELtopUwUaztm+Kf1yM
VncaLAvQH0/DqcsqsbDhGOq8xEoxyh+vhqkAyp1SmoJt3I2DsKpyJCu/MhVt1CJe8xy8Zm+rHd9O
EVsebU1Du3OcjVqbUx17KXLns9lKgFDHixJ54POfu0TRpZkWFZmZsBNri2x5xKZg4Jlzg7OXORZP
XfrAL0of6VKa8rrC6mOpBd9LxrUNQ+KUWooTPc7lcJQBYF8fgLJ3thy0WyHH5X5YVWX5Kvckyu4Z
JzE1m+9nfBcUj/JWJioh5J24jDc1ocr9V6OQF6PxIxqAk7pUdv+kx7PDz0CkeZi27BdwasBIg7ji
3ZqWEX/ggwytxVqq6IQ66zrmQHCy2TuNPs/aDd2Me5lTXxusjiQLeb9hDtfUYunMxHbsl23UVes6
SsdVlLBOUZCF/SxVSfm1ApE7e/jdWLGOyPznOgoqwxwOvPiNly2N/2G4E83SFRtAkTysegeR8JLF
oHnkyb4GpcQ1z/iNP1/RHL9ilfGzIYi4Uw6u+KZfUfvbxWXlmjo45bBai3jWoBIzPMdP4CJ5jVwi
6KKZXH7ukXV/YrJWx/cfpMcXqJk6EKEfkAKH+fP57ulu0mj8IuozHMq79xuHdFKCQFzDD0N6RGx5
TsSAV22n6jls9hIGteWnBwQHaN2+Scb5vPzHxWE7yRkcSiZ1yG0uenGPZ8sZeL8NDr48n5qDJdpG
U4HK83FEKAg6wDiSLP37GXp68CZHsfdUNHOMEi+bs078IrnRDKK2a8VlHuES153yYyzC6/ZHp3Dt
04K0p7NFgMfSNTmKJwvSq6FEIRNMsluuiJ63bpvp6PZzMkQB3YQc34+oOECp7527BZwLS5iYxE2p
ytP9ZHZg7woJOVKkSuar4zzp8xsyyBEtq2/eWkNWmlqJQ8d6W6NY7LduQcfBPHio8DD1MyQtBbnc
sgYz5knVR4fa+QDFTgIDOMwoSvDyL+eWt+FV2gF+gDmm2A9tKKtNBHf+Di8UwkfntjJ8l1+qBpRU
wOZLjiPqvjUCTNj03BCMmU2CUZSSe6T5pgWmZ6QHXZrRCzoYSByJp9UbgDZZF6etQYFkamOWQNM1
sUJ4vaQSeKDbZZvI2EvlpQwsx3hGz2KmD7tC9joIQeEEYO7FZkLPLzY7925+IhrrdTrh+hOt8OOs
hgXW9ZeWeGZsOExUUrbwGGsord2A5ZrbXkd8AYEWRlC71FWj3i2GAQLK2+K0gE9T5mdPoQkCQW4m
qLS1yOu6ODaD3mydf8MN/2coI28A6p0FT2pH7d4e8VePWsJGSOHnoAdKHJExTiK/s3seWN8w10DJ
k3ZNYAyca/7SNK4J8ancQHu6X9cG6pxSahijqOEFNED0Rbjunbz1CUqWllhIhmkA1y17lamT0Tyz
OaZ+NJrgHxYLR1dGEEnI3pSe7gSqyeMYwU0RvC7UEslXaLtcIffOGuaI8gQAW+4QoAPm0OkyevkR
6lr6WV2zPyLKahF05t3G2O+OEAbSwbfox/pXlUSW+0Rh9aSbG4PmCXINNgdc1PwHOKmR0W9di9/f
h3+MUid4wo3g2TEdNZ78qe43qAfHmh2nbTAx8+qOWdFpig4UROIj+7D5nT8zj6pxCiKKdZxZtkXG
3IkVkK7cEGhS3gLoBT14jnq0eROx5I51wXckvk6RxQLncnk9aCjdJ9LTfmVodsQmLhsbLxIaL2Sj
LaLCAiMffRxmeGkfs4SLUIRYNl704vi0QyGBiVTQw+FC67SsJ862h2BC+5BcybsuRqcDEd4Yf+zL
nyp1HpEKrCKX8GxHQrEjV0xSW4aLgedUETQSlXd6W3hdU9+xbyHQi4qKOv5HzyhoXU+ftVfH/UFE
0CLlaTKungHj3WNCiSaQoMxvUQ+IFwZDble9Q1SVYxY1bV8MvLEsHDqA2R1gyc2tcupanEdNemYs
Hhbf5xP82NOOchH3kx6BpxLtYbvOYXz0Y19ZU1CHUsGDGxH7F7f2hQCUjZg/OnWTFvdZhPs9dS5a
ALnOfE4xm6gvKHkzmCPFej5Qd8xc/18GAh+BPjAtzU2/9upgDjb1wCoabHKtNpwrQFaDDytYQLxR
krBFx8wUU7XlFpwZLDSxj5awU83XuP2Z1odL32gvOfI+BXi2BKALMfzHTZA4cs6XgcKhfX0crAFz
2YQjaRHpDis5rKoon5bLLxDcmGs4j3wvvpv536TDlRB/pDnljgXiMBoiv4mwsTVrEGlXlZdwP5l0
7sONPaTaZK5pe5AWwMNGbmFRpWAH0IWiZYFqB95N6WJyWjWDAuwvlYdvY/oZCFI6XttzoEviqzYv
0iAnAanZ5Aa+Jtfd6ZdZUFyI1s3N26wgZIooLl97ho0Nmcc4CXaCu1H6gPcjTZK53sMJRDG0PAFW
I5Gul5a1RELSFBf/egdDMlei3b46mp2L6HUp4JLLjHLJDMETUn2JlwoZykAmsJ+ka16QcQTYYnrz
peFeSPdNJy6GRbA8B/jKxWMlgXEhCm6WZabRT/wyuanIfZVnzMS0/gu+H/VkYoCDSmxIYUkXrlSS
JhtOZcFDNprAV/PhMXQLfpVldG/Zg0t02W1nwWemQIOHVuCK95+jjcxZ+nAXJ+EKLFBj1aw1t2UK
GUKL4ebr+rkX914futLj/wdjbgwf8Dz6TvY5dp+f6i7eZF+82CAWD5c6Ce1gXh3QOrfoiX1SheUO
8SCiTmjQj6FTrylTxn2FxSUiqa1k4bEr7XsdKOy2VZk6wO3d8UGJv4ay+hUUkQsluoJ8t2l23SRV
EelevVwY9c2Z8yRaDp4Tk2Be91RFc/aGuy2kmmbYGGkxP+kUO2z5+TEEJS6Nh2p6/La8M0OtA5U0
oBS7ylpHtfyD7mUVD3uXs2efNaA8s9Kpc9VVGJyz7iiTpax3ZFveYl98BFUw6EhRdpBUcpU8Xt4D
iRPIDzoyHPqaBrz8VN3QlBSrcV8RnX76khuS9gMjrlVKp41CAqSXhWwr48YpyX6sNg9y3feX0+Qo
WzFKzaON3do2hcX1xB1fodkqprsKgu1VR4xH5xRIImdXpaL/lKI07ioE5PwS8APj3/qUs+CANofI
AcvS6ATDPoyz13tSJk2s74bwcczf06LDwcfT9021Ro5IPLIUAVwvpsQ5a79o+G52xD/7TlOmja3r
fmG4cdIScPLkdpq/z4cZQTklovenXv9sXD3AuicFEKiCT0sVA7oPRA+3fL1LgdbOb9hDYLIVubYA
qVIIc6FG7ILzfSbi61SHPaHgtvZwzz+Dtb+AZoYYLzLQ5SsG8trNzh9X4iyhtOu0X2ob/c4yiv8/
q9e30evt4ICj5BgZVKVaOiD8dJdKS7mY28lAV/f2x8QJBZy7eIXHMfg4csWE2qDemYnKPTqEEd3t
twcmiX7XkijP9aMLUgKOJ0igj5TYeeFrhGUFIxOjIhdObORi9/wV1L/5+ZMauKNx5QhNS4uaXl3a
qFN1kFtKZKJ8WLIBSmlV2HgVSUGvBHlDmQKsZb9pPwMufA/19wkEFyC38qLRc6q7wpsl345h2+3j
LHnBy+WgKQxVugu5pkpeK0c2biHvVjLQM2TNzG2AhbcdcnhSmPZi8HO+8ZEkxYRIMMgJezVZTsD8
W4TlJvAGPj+A5e7QkyODyvsWHJTfTc2lXQo7q9iPJjnkovroFU7JhYmOmTEXqTXPaCplOEl1qDzB
ugp8yYybo2sqbccNKV8ZnpQZyW3Leks0rFpPgkFl66a+nzmHyB/wc3nSb6t8+gg9b9sle/zOBvLT
3Ih9zZvW6tmOBlfJnHOBU9+tQ1kwoL7xZCsR+QwBft0gVONbJ1h9VTc2aF4QlBHoX9sG0aZiQ8ZC
0doRBiCo1r/jzaJ7ToKbKfrSr8237Hck5VaWNpknv+Nk8GDVUAMkHdr8MQslD2pO0IVXWEXT7IKt
l5hSGmeNrrAzniWLRv053kQa/kTT7ksgBApVdvSFFbJS//ueiRt3xyx7c/bVOqB91F0AtsnguheS
jaWJ5zIU2TMTkVU2MkHAJlcfJ9AdieO0vVNg6VJqRd0p4Fo1la/QKYV8bkVAXRepdTZkhHDqGEDe
hBXXq+9L4Qr5dhvfzLyZ50rozLXR7uoT8pt54mHMCmhkFK3/FNsDIGJ4aGGarTmjgpurAWp1Xjdt
+kBdK7I/iiHLos7gSXKqgTHgbhI3oVZ4GlvkhQO2Cto+vmyLJ20d/MkXOmbTNknpVWoDXNvuHOKM
X+z+le8fEYTwfEjZqx0dSFei9SFXMSzWF/ny5cVZgUj4nKtIx84VTdj9YemG3A5zPqHleT4hBap4
pgKNnHnSBQJv5BerQpf8WLZk3mjWD0KhC5kWdgDfuxSx8n5O/aYKZ7wDuh3APpw4GIeiguGc0Pxn
rcmyYxUibDp3V/vmD1esWP0v6K0uQjL58vYnAs1gScabe7QjPJDuVD913BPIoXNGKhrSAh1bJkZ3
z/RiU3DtovjxfBo+82BQPKFKwdviU7uQg2j3PPmG6NFDsmD3a5QumMf4LTtnpGvxJbMEFUpT6Ev5
cjfu72l6bT6/YHrqrjUfxtEhtih56Jm6+jiIdjFtzVnFaAbgrBEN/LfdBRLZtksAOFhEr8VPyV3g
LMh61m5EVuMvzOKGHid83n93ngqlE3p5+BIERYjoaPT9aJfrmcpB3mpEs3POwv8yr/KfEg2eMKi3
5bLcaQ3n1VQi3tg8qHYCTeBtkXQMZkDcFBUQsW6GdDHWalAKI93tYlK+/T2ejtHjLTHG45I3Z0KB
0mGNTwXlSNiEZjUCye1whDdoAtEs2OPvvbtCjae21F5vMjFCX49G3BToEdGDok8WomDpCoX1BFhP
1mfipqD/q5LOu0Ftl9otEqlmQ0G+SXiQT1HEobJe0rqCO0vIbM6nhv9JxkzBjwCUPh42UE0ZkHBY
mNnusTKTk3VqC0U8Bvdxq/CQuuhJPfSgx+N7TzydP2VkVvdWPZB2MX3+AvO8hBvrAh2UkDAF8y0q
CnWwOq+jAkkDkY/DwFZZIgqF6I0HG4vK7tdvLCDRtgKVvYKe1E3GLoNbHGWfPbYwE6pC0YoA1P7h
uo3/HWc25KPALLzu40gBQjzhHCPYqDlViUmbrwnw+eXjt2Q85HljGJoJ13Lx4AHJmo0Usmfk4IoR
oyufHRUfRPEXUt1de324qEyGbrYY7dG4JkCmZpZMKu3Sc3MtjoJMr75BthvBhV0TdA1ZPa+Bb+CT
6zJ/LLOnoXjD/ScNrDBCnbZdtTIRmstEAPs2MifCQtTbQYmNfQPwUkBaGG5k/peKdS6wt63uBHwP
EA05ByrTS07bRyPU01OkESd20sZph77I9tZLDrCc4Gh21To+oiOUpIxeuBsQTZabrLBpVBR3awov
4MWZ3RS1BC9ZxKh2tF5UqXpMjPbsA1uVpyMz/vjUVab1rPdFBfgsScemlp8T1lVHY/gO9pCRIk7h
5cwMUixXg5z3/f8FjKNXnWVhMOcz4CgHki4ALBb28FlZWAWdEpJT0ckX8xtaGiXwaCRaBtoDA/bI
zmeeGrkEZxGUrdGhBJ5ZcYui4cgEagNgN73emvULINTmSMbJUMHjTbIzRjhryaNHTEFf5eKhSyd4
UBlXR7t+SF/N8V3WA0W26uWogaxnHEFyFAIWct3/ArxC5nDr9B/0YzhGxB4EEl/MBv95ICxH3hp8
VAgeGOaOaDUJqqtn3kA42HiwRMTw9mkKcQt5+AvqLDEfwjZ2Q/kAhvtVn1mpuNaDGN6u/E9LGj1H
X+5xm13BmymUjyWCG5DI9pdZz4YKE8RvzqhdHBK+ghx0F/+PxXs5yBocHeGOAl97z3mJOcCc4Qzf
ap6yFUTkcvUaDAc7TER45X/fwsgVboGeAONZTsfUvxCzMql/Yt4SIhqUV3bmNRnBVsJ9tSd9YqrQ
cr7XCZVy/HpMgKE68EQR4/IxWoRPWiJa6Zm9Yg3uWNeQX/ZtCUY/ZryizLFiSfWhK/GzZC46HA9Y
5FVq21shpxgFuUrHbfm+6BFITFBs6rdyq0M5vKv7hACr6SuwuOsRuCNXXlRdL8KKE6OX2gBJYjLH
a4TJpGBgx4v8wpEZOi9bPZ6zyQGA8UVeIWk8Nagg4VT5slwZS+yWKglSJnb//2FLfHP+higJxSuU
ZR0TkpZ6X3SxwbA7neaV2Q3Ha+MQqBS5bZBD/rLj5r/bkFQ1MJ/t2yWe2GIvjGUvPEKrFeVr1jY2
JC+uT9zpx4zo8N8kBqURwGpBhAOT8aBp8lKIkPrDNn4xkKO97zoWYs5Kb1nPjSMi++UimYN8RdbJ
JothTy707JXsHA237i3kse7eUNbi4X3rUiSqxaWvglbV/m8RzCelAOKMyXBWpBq0bR1CpFxuhxGQ
x4AXX09g8iQ8CRMHwKdotwg6eqjv6eZR5+35xes1k58a3+CX2mpIjMty2I5cFZ3JYn01Q9zS+wYC
BjSuD9r1T3EIK5iIYsStx9dKCVx6L16uPXO7OCpZVG+/mtWRffl2zCot82hdHzU/2roaKM3a0pfN
2FXcnQx9H+cLvz7Bwozq09huBoQD/vVL3ZwILRD18geaAa+rZmeofvPlQ2WqMXKUkcrUGyc/XlxJ
PjDMBEicEm2OADUk6o9PzfMAm7dHUpK6yPauPHbCpJKDrj0MCLfwF9y/++88bnKnDKtUc1h+2eWA
2vAQmRMs7I702i3HA47flO7rLKOUz6ccfosrHeJyuRNUxUKlnzHWGzeJsgYt2WDNkvPsyezb/FtG
FEVmwMlNLj1WSX72OsxiHJW5gQGOO6G1eCIN+C5cS82rdj31JEzvNVuwOQeJkDkO51dUl7c7yjBa
uz8xMoQriBIE7ub7cqB1s/sJSPNux/xeUtXdfXFtxX5XhQqV5Q0qAbwrmh8W5jtigI0mFF2eBn3j
8RLChXoJ3JwMU/9AJOsUCUS67J8LxWjD6ViBowYroXfuhzE0GeMAiVRG06p5TuJ+jDOWj/yVX53q
JMZGe+UJuoBof64I5ekjuGPsxiuhsKSQ1o2rVcYDdAVXPRRzdHSE3M4fdPtV5Kdp/q+2iJZtTccn
D46Mkc+5KdwSCw0K3JErwiO3CsLAisBFyTRT/5wVwJcZNhBlXpqcbpVPzrxPULSDlbx0d0f3lkxS
ibPwtKnJx7dRi39HxOvj85I4BOKU/4Ah9gBYYMMWdMR7YDq66xy1TYQihHRpAz1urGisFnVNiIak
SL3mWjv4Sabn0n4gHrTBgJQjBFUdqSonCAnkfpTgRsp6Nh+r9LMDNMfP5Buth2j6tn3sbQdgszU+
XVVh74ItOtApWpskInfooXRWXtg+UKRrv0UaQT6F88lBXO6+GCYtfLfT6fWcvwAdR/pcc2IeF7FC
+2j7DwuQ0brPXm41fFePwo2iHYvszVRP1XtRmat0btHV14OQNbMkm4HcNFtsr1peiTPhKsx2USG5
HF6Yrbllz7ABkYojzvWjAbroY6hkgDkskc6zmUufIwy2JTNn6QgDQGoi/QKZqv9XlhX2r8s82U62
czmIA8XkqmnhaTG/wDVznxnLsPVNLiCdAjZ/2QrBLt3yDgivpIru1jF6Ao/Jw69eGqbjjj2mq0nc
E1MZWobctvx5cX6j+/2Wpb/M4mqDy5lX5zJ6Vm5GfVVi1KuDdG/Mw30sF6SNPxbdp5TOMdd62ktV
x4PxSU9UrnGI6MZQIA+KljhLqoC3WDQAwObVQhRvTaMXGApsKeZy3A8MiAhi651v6P9Ho/hzlr2s
uR/Y0lfraPaCBujWqld9WMktfob1iwa/oylMAVTUaSv3kZKcmoNwfWQ5DvhBqNHQ671P/jz73bij
/AezBG5Ei3BTaqqS5o6A3BdTQJDYlrGqgdTy0r8e4xBY0UtcrodNxfEdNA4j9caQkV42TJhm7xX7
Umz5EUjSRfQ4YgTNNWAnXgikj1V8lESgkq1TPL6OQ4JmBPAiGxm4X+ZIExQOrz3sc8u2mzyH5gHZ
bhv7vGyaFDe4H9JP06sf1olfhbUoAdQmoUTvhrcrgVSn4noUCa+E6Qjii/nQcamgDDaKuBUgjXPQ
xdBzcUZ6WTs08BBBpAYUhBofrXVfQ4mAUmYG2hLXreGH4DAcvvf4R7lAL0zJC2+FNf9gXAhNZ5Qg
JboiHkHNJ5hqRHm+Wp+FvuFdgDmhp11WdwQrXg+3i16/ydjWCp6wtDzgQb+JlGz6qTJsYtlyWQVJ
113/yoN7zIPxjqQlJwJuajRA0ULl+EEHbYTRiqBjWZzXZ8+H2nxINPMfLXdz14eos5UPCFpM4wDB
e6JMc4pzGBhb4SCCKCynsUn3WvbOlL+bFqG0Lm3EXB+h5N1/o/8xwhJiTYT3MSMj3ho7zSEQbtGl
UHRhBMM/ZqNBaou2mN7+O1mOJwBrCq9+7A/T8ocM/y3k55sovIMqUKJOtJHbUxDD6McNvSOR8Ke7
UOElQyB8hzgzILwPDz/oFB13AxD0GBcVeDtq2V6D/BVyPwHpfwG/AxPwnwOMRN1T+7ck3CTZ47DW
Svu1dGsngMDEN3KT3ZUEMcw9yM9JES0oiLDXneFyDq3IUKQY8dpuP/kmfqAcVKKHKf2k4WzSVEBE
TROe6DsFL3cJMxYDzM+gBAXjSteVlnlWyag0G6aySSHKq6Vzzj2r0cN6IHWnT1JJXBNUteb1d/eZ
94UnjHrzxuUnzQ//LQyzCVLc+j3dVY748ncHamTmnv86tjGyZK2AZG6w6ga4vfmy9HxEbdDJtDfN
ZcUmduOjefnAaFUn9+sjhX2zI49fLhBIsEGKIc7tC9v6erhsjp5CegmCtFwYm2Iz+Dn7OREeu3ig
RPFdfMK1+hgBxXl63L/3L9rB9LeCZNmr14JDXcLZbAJwyMnFx/q4S136PLQ0DSysNX8MyQh3nfnP
iVXY3cAj8ieOT0xfYb+kf4Fl+KXu4zDuHeXwhUsTXX22EKGXiSGe8N8+akaka67lk5qDgnh2Faf+
uK+RDjn09qtFrkON6ARjmL6KMwpvaZUFCoOuu0yb+XSi5SMDAaV1IB2w06AivZl/2wjTaa9dIGmk
Fr7rDqRe2yWtyXBTdgl90LpFXhSUIWxeW3uRJs6LuM5upuYer84TY59xsknDP8++OY6IFQsXJAdK
brrVsauXM/fxf3e+hJNYeC+/BDL7Ct/WnnqeNBfgbArv+EgpJTh5FilxJ128V0ATnGOw0NjFB91X
rFQSC6k0i/4GVutPL1WGQLVhteim0h2PfA9xCJYn4F7meAth93GoRiRKir2cskZaOyBJIxbR+cWf
/JPKudZob/WZkAKQsiRleP/jXlihvZXl8DzApoQW2Z522LJQJkemLS5rmLzj9hI+yjiEK+7V+CWv
YqxSZt9IP6RkXhFDgmo4xRxOGu/MzuVCflsWLZWZeNpO0Yys0QMv1pFf4wAIbmmsNP6N6/sUt2lS
MV9tkm/meuhXw5W5OBDFqY67W0t4JZxMcNLNvPQ+WeWzZG4+O3U4FH0rU75Qb3hYSk7xXASpWJvJ
bfq8yDmVHXZ+GRxrOKuxFFI7i+Vq9tTdQFsjMAr05BAy5BaNu4T7FqmIQAV4XeeadX1qewHj+tjf
AQQV9udV06MEZZ3I2ZqV7hxYZ2OY8wfx2r/8s7drS0N7Iyuak1mwo1yGhQNuppg1KGggFkJm0TgP
pzZTWh1CG5k8BV4FmMVWvIRiX4ZWiAc2I9cT1uf5CW97tVnyaxLCdvnv/OhjgDgbgv/QcJkEeVKA
JpnxzzA8Mg+SdUMcXJWqhj4LM3Fpdg2bKwdhS4mdqTLg0y61vaZJwxXN4pi0KuwQ51LQZJPeMbfH
x+d0kT9PuPvgciqaut6/N0jt7TjqB1LgZ/Yqh6LZw09hUQcRBQWi01e7Gp1CKA8gBbyUYKK7fORf
5psEVjYAfOm1/I6aXQu46/hFPsIuD1BbvEPzMBF6mMU2Ie8nkjV/ALPtu7WeoE2ImDgrK4jV7J2/
G98NFA/1tCh85qqUH3zmAQUr8I+Ioudx9BXnC6ALPUU1+wX4+xr+Jwclue2DxJhncGlmIsRRIQrx
Ms7MDVGnq57HOYe+924jOGzrG4vJP/aLet7pwDlmMqJ9amObk+Ezcy/6ozCaoGyC8weYqyPy/Fc1
S+aH6lHGdr6NRaQSA35rx2uJl2J6Y4om4AS54eaUOs8nyojj1Bw919Uyy+UsnbLFJSx6AOPuDIls
HtXKBARdkz8fSbj/VeLg8blwg93Km623HtVPFmKFivuN1BPal/uDy6iyX4Rx1nP9QlxApuxdezws
n25rdz1y52tEOEodqLXd7pDWbAL/apaG0r1WYMZONfbCegr8EMgeOr7YsLlr5u7n/Jp1dpFlv+nB
LrIO1+JRNkBT+JTVqA3mUuM6++8R454Ak3JR4J6y+D25UA8YJMgYYhtohOJu/uWVDeJU0UP0sqy9
SryTBAQvQipxcE3g+XwIk9D5Qdp20wWCVu87+E97zECnONvAD1MdNlRrnK8EWepub6BtzMPTSMbK
C6YlyJvfCrWEAX81+ayLB/aiBxnTBiBkf+9/0MGDw5YZZp2+S1Q0y7tPM4GVyJbUKNDURJmZiJsd
Tmt2M9bXniIqjX2njeeij6vYOylanewgtSYMMPswdFuImfkPfzgKUhhjIaCoj61DRCKSSqXKwSAt
VJmsla/nK2fPMvr/Jn+GPnMJxtDQapZQOMKwLHiQTn+Y85HmMflkjbIs+4M5IRD2/L+1xKbuNOU7
1LNyThrWLU4aDu1h+HSQE7pTcBX5WcZsi0vt2w/H8bVBAFvRlTadeBDUpSoCiX+naMIPkArEbvBZ
3S+YdyQXsa108MLAb+OSyBs6fMJSQKcdT988OCDvHerzyZIbeoy3Y0tENjpTuBe2e4JHw+pAWktn
k0tbYFTwfhSp3FcjOuvsksaxPElysVS2RWn7vXb8gKXgkUa1g7C2X1k2zkVD5g2Jo3JDsAXCGlt7
dStb+SO1zgnpnEe5pdblHVBBdVdBxHuC2jltVJkWM5v2wgpksfhqyKX7RtutwIHP/ZgLhDKb/rbk
EuowASCkKpY3r1aUbWYjbMSxkk4s0EQzE3SHdVNYWWkqo9Pb2pE/KCJvLrHv7SPlhfqj3fNX+wB5
LFdReGN2dCkDtid4HvGHMCBulwxUFbY+kezN20Qfc05OF7OjpK9vTmkxeacPjPDpqQ9y2LepmjXV
0RmPjSzEK7/M2rHr/vxtYj37hxhyzHE1v4kah/0sCrTWwyzVJ/a3QJApiDWCWNXmcYIou60xoDtt
53uyaUeg/n2Mn1vZyvzTe+2ad5EsE+58aU+mlNRxqJJhzlNAOY0TAsTss/h831dY2Qvd4rZqJpkq
oSaOkEsHpNqosryYvN4WV2KiRmlUzUelRjqMTXETZR4S0pnKd5+3VPXFIghQnAFxS1TXEg2bZt3A
oRxN/is3K2PJl/lD6Gk+xuYFcVcyqC4GTYYDzCTe/ayhk43kI2k0c2xe97F4wiNIbos6NNHLgBmf
8eWO1v2X58/03fT6Cd+g3FTys5is9TbS4kk0vlqjSiFeOlUaednRP7na1ck1dxlHHPPGNDjKv/rr
dOcUEv1Jp3P6Xz8ocjJMfAFJg50Kh5QwRyosC/VI1csQ+5b6FOQb6QaLDJApLODiKFD1gwjrPBXb
+fYnNNHT0f475HeqsfgtZuaX3AGWankcrM5a0R1sn09PdE47px6isYkIpFA+Da5lg4akPMq9BcnC
6QkJpPr37KGdVSXbN1vBs944pmUB5v+gSSg3Akhg2QIdKIhfTff2QgDoFlhVhVzVHkVmG5XmJXmP
ae4vkkkIVqf1ItFnC11sszwQbugvd04PL+u+K+XHxypXOVxR6H6Gi5vTkt+qoUtFMOi7/6dPMOZS
9hGmfbX3nYIao0Fu03A82LPjG8w14NG4qyhYa2DTVunF7nTFW4g+Mo0UhOg5E1dwjTcm8dGAPHl1
dube3Kj/bipoQf2f8tu1+C+tMTFKegTyW1o3Upap20Y6Gi7mZtPJ7MXT1dPF6Y7yZhUi4FgcBil1
AllUahl9RP8eZSukvz0+xB0xaQMLwzSEtZvbH4JCXKwVgFJzImdtH2EJMqPPBbTu8vXvtAIqMEav
c74vsnB25nPhAmr+7TDbaWOZQAbmfScJpWhwtzdRLEdjrdV1tDqEmGSlCU+f08G35RsSn8n0SLZ6
O/r6LlYa6/veBdnhr7aK8G3Qy2jaFWz9bxqt9x8QeMDC6E6OCou0rVmPAb/8jdCiQc3X3O1pJ84f
aD8WbMr2jYlNNQF3elkGrQ7/Y/MHdFPKUuUHz12GQQn64OTLfjkpP3SwkgCgNo3GgT9FkhjzIUc4
B6DCTByMn2U8PcuYrqurvj8f9TX7Y5AMunTTy7jSyPkzQWLb18j2ny6scgSfpUNvdeGUykH09Di0
WkoWA6MA1gunFxUfz/z6qRe9pWNF3mfVCPiUfiTTTQZGnSdfX3oax7qmbo2hGNZl/Vh9w4Gf9/Au
4JBevBNMpIuBUhYLoGPQBVXln2jfm6lOLKEcSNAKq08yQtBRveXxcrEES4Tc/rSV8AGSrFImKfaq
sIy5UNiH24ux352sDWRERaLUxyIpvJQwvXQ8zLDMFRSgeXtdMVDFzmuBAkgcMWzn2SxFGlCBVLSr
YirmS0JNzpET9csCQe13IiXK38Ld/hI6/6I79F4frR6VLlNOk0tISF2Yrl23A/oI6SERcF28qMA0
orisa5ppERaW0oPkUcPDpqEeDlO/NRfWap+xoPWiCU+kqqgZinYvaLSUMe/w8P7zCcWnnONMmE7X
XTp8UdC2dIZ9cKwzfQPcI9/9BgOi6q/HWCIMQfCOiMfpaMjq8oYpNXXlPvgWonUoj81VcjAeo0g4
6Mu/gcHjv3g8F2Yn4qsfZY+r7Ba4WaSchKFOgM7G/eGBWhMkeJJB59lmFZam7g4esW8Eam/q4dzD
KA9Do0Mf0eymkscwdV+Y7GV9Xprmrt9Twpfl71BVJ1RPlWXWNpxWy1t2pEzxh5V4IOA5pXy56nIu
/dvOmDkpsqpnMjLXsn/vsMyVXZ6n9iL+Ivu9qI3YEsPvfRzo0cvuXfCWuyFqlwKz5+BjOUKBvWBi
0rJ/CnClxVtCaBdleEAGvLINsjHcx6uRpJK3BtZt3eh6U/ZiLSRNoVKtNEmKd/CjxKsiixLgRi3r
FzquDElcqCa2r/WOMpd7hwXxwTt34Gk4hp45tHI07o1EvPge6jAjvuzbiibgpUe7OIGxgcJUVJ0w
Tc0MafdKQJPHmKn4aYORyx4RfQnymn46hhBH9Svyvov7NaEXVrVs2mBJNNJYTAI8jy6mvrs7cr/z
xe2u1YiLp9zg1Qy1QFB5IMLVPsVoMsOehjzbS5G1S/tDUJ8JEq0EcQi1TMs+jVsc1FvyxndT/nc6
qFpwtTwQBq4n4vPxhYo2PttTAgnY3YX5HuuEfXv9wxP2LixCAtZtId6icr4E/h0JI98U3bPr2nHc
zDnEOSl48wc/egvIUTpzuFX5WXIty461yfyHmyhre/BwiPmi3adYuzGwiMW8FZekOCK5GlfhzeuE
tPoqYXispv7hYlChM4BCWiGLJ1k005pK1TSp4fJknRgsNNX2FxgpA7uUDtIQaFaa83/l5NZNrEd1
HHrRPfNRkmEPik7mRrHTjZK2cmvLOPwG/KFoYXP0q3MRSryQE8tlGkLTlxYoK9uE3eysSdh9zafA
wZFSxAnwO3QAGoxmknOw0HvWMa8V1fum6y7qc0SsxgwOXoKE6utPKKkXqAHZhXLliY1IMicAyH+5
o74SJVVtwEtXRvr+T2JyZI/FU6UUuOd+F+9hyDotiXyJN75JWRM3mCD6iXK6g/AOnn6f8mjc9uw/
dki4xf1EgbAeA3zVO2lDtgWVzSr93Y8+2/3y+VwjELfCVNCeUzMljOxqNR/ppEF7qIkWk1BhCiR0
E+IGFP3D5cHBCTtaZZ2l6daPN2u6F575rBW4upbttSfS7XRYD7n33WrfItWWHf+ldDwWsQAA+YLA
7/dMuy6cd3NLQcKKk1B37go2BT538EmDDwsVB5q0Nuy6W8pcZ09K8orpxBHP7gI5/l6ujr6lpss3
duCtC4U2oAZgs7aQNdx2fJ1ApQuzi0/eLCsO32DXprltP+a/M7aH9frzHmPdrYdRnQwvSOkIkz/D
bJ0gjawdzDV4U9wwdYHqSrctmlTRZDxWJOrat+Sm5qwA0yfZTSayljQCYD7q3PYvWthY+8ccqLme
ONurgjJKVcZ7Dq8vOOo4Ezu9DDqwJ4blpAhVIhf4aFWl8efPqOUKbr7jPheZD8U4BB1tmQ9IEhGQ
qDH4SGm6m7teVgfY8HnEDjto4NAyDn5I0KuKhIbh3QKWT0raG9DbvUyOCHP+Sz8TWT70KmxTkdCx
gLSF3Vb1OldDXgeTNIw+/pRUs8pBtf7duPS/D8kPFHaGSjJ4BHo4hQPE2bKE0nsQOAHss6r1gg8K
naGbD10pn4ULon48lLo9pgCQ3KiHPCaUGbcuKooYdob7NhzD+VJ/065HedZ56OQymg2hEA9Ax/Sk
ukhOPmWYe9iRdKuMK9C0TdWiAMjc+hd4CcyJknnFOolmSxnZfxxa4ce52EAWNVuOdsCC0bfYG8f8
v0GyTUC9lo4sitaeSICVZ7XPsMJwJS7QB3w2UBZHY2tks7a/dNkZp0dpxoWMpr0fqUjLB+qg7Y2y
3PV0RDuXO6FmmZ7REQDxvALfYbVZGcIpc5ZLEfQzXaBxfchFNW1l8+iAQNy/x6WkKz/ahN5K72hj
iDcGsh5YYTkg7K15H4Q2Xxa5LgMNvyJEQe/Y84MDO702oeDYXPxx9v9GCBVVMKvwU4u/lsN69Vd5
bKmJaDlRYZwvJZXM9BveakCap1NFh2ak225lEaSk0f0r5ZrDnphkIfte9PrpPsiBcgEv/wpfAilc
ppe88xjjLeDBPezxQskU402cM/+TG+xqJhOPCl1rr6ajtsWeE9eqHFLT3ET4hru8dItCI7DG9wFy
DxHwiNtr0DSSNURJagp7SBIxB2aRXiwDGzH/0jpdOmxPO29YbG4Gu4TLXFE5lnQ2qpAR6duH36Dz
Z/zMu59sTKT1/V6KxRgiqeM6UnjPvJ1LJhxeful3bvoVz3hrLwWgNehWNhmirj/bMzsr/5ZjIGj1
VkdQBpU7wg2hbNh1sDALKSKiNB78blpkDgzn31aAMn8YBNHtLuR2Ibfg7QTE+abDi5nIZ0wA3wko
I2wCPgEhHgUCx10fQ85BY0xz1QpcAE0CGlo2MJt6n/kwef3ceuRnZyRJrg/tWDV5ztMiTv4J/PZX
dKaTSwlTRUQpuGqVasJFP2n28i6D+Fyj4R7GKLJTruOsU7Ry+uQD6fHhjSa4As8EobvWfzSbx/co
k0pf1i/jiEBQPaOgF6c3TsJl9SXUmuCh1c5nA+v2hGD0mZjKjqfSu3JSWVEYHC2qnOhr0Reudqe+
rQ+L7vZWcnus7mttkQFTU4vHyPu+J3uuvRv76gLQ1bq8XB97OqvyyfOuyr3PckWd6k7vRjXfrDpS
uLO+j/2rYCM/cTGYIPIlHVFeknMHA/FrywHtGmVrvftG3DGCIAR1yHQ1WLwXrADqhmPr8IBKs4+f
uHYllOt/rfGfQCRaVRGAFvCedieY9p6D+3EkVyESWt12y3lFYvoqcr+IpIG+lwbGdwuUiGlSMcCL
aTg1iBTxgs8DmS2QVSI2wXKm8o0nQmcZ63+6L1/oUNSWao2Oo9goMmBLQIhzZgt09Gh0K73rzFWP
xKNJhgm+vlmJGxeLcg+uKqRd/VaQg5OWOCDgXoc3cZ29y56Fw2HV/sxAaqE2IwWUc3dczEvtxCSs
ANExKk0bJiqa+GJHivLyjtHUYWaFest/AJGD7m6XWH3awKeOl43OA6DgmcVDl2BHhBhVcoAEJY8=
`pragma protect end_protected
