// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NZ1NnWcXcDE4Jsvf4M62NTRN+wEJpfdFh/2iOm86w2FBV9pY8GzcNGYmioF+C7Rx
CbYUbdf5qCqVJYGrtmCSRMGG6KluMnHJufcY/qn4kWopLBZHPnh1PC1zDByiKKFL
eI7x/+yW+UUDCHSdCSVMstFTcHerSeEFwEBFv0Xlk30=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 62064)
ME3TurL8w/yfSvMEQfjNZY4B9cu81BcLKI9IJkbNOyhuoN9DZSBMdfzvolGVc+cO
Das/Gfonw8P5GiAi5w+PWAw9cg+pCwlgRJ9uUsGYmIcdgLfl+DSvWWUXhfWV89PE
n6Rlb1dffzIs9uDO6PIFxnE9jSYx49BQhtXCIMugns9mhnQa6wrh+2bd8hBYkVQP
s2A3L6ezXxU/CrKbxdP2b3tJSdzJRt1Of9IjW7HZzNePWPCv0l95OYLsZp3EU10P
M1LKW6Jn7l0oFCpHekDvD4GokKADmMOLaL7h5Yl8FPLOJ0kwzmoNLE19vUO0YYiM
fADwgyQmLg93Nm890SK09Tq/lsO+J8C5YJaQyS11laxKydYC3Iaf2pVV82jhGlHr
ZiLSxk04mZBhMmobebMWoFf4+y9cVLlyWDcpKCuPtf0Y0x/msL6/BLccwZNO0bhj
hva9eWv0c9sz3g0KkvpPOGKEJac2nHcewNzx1ZAYSSxBxMWU88pfyFXt/u1Iux8p
X0+Z4mg7flTFngv1++uKc0j+P0mwqjTKzF+Ao/f+oPwetW1mb14jAJ40o5HXY20/
QD47ElumT9/lZ220QNGjo0un5XelRXEPkTYjqVaqYbJ1rJ+/9n+YXja7KTgMIIMy
DwtpZXxeDdS4aUeS/89TREKecVNeEiXoxZB0YTrrdmUcemhR365iYbAvhl0QwkR2
LtmwStn4t3DfqYxNXASxWeUjn1nhWIeced47kf6G1b8Q3NTwB4hEYLOt4TwRAH2U
oKaW6JC2xwQ8hE+Q2sLua5is0hy1iYfnnud3bjK/XA0kU5ZQ9aZlsh5Nd5zE0OCp
URPwvFH+oame+GtYjk/CGKdPF5Hw8ycv6LxeS7k3ATnOq3KaRbmAiAHaR0xuQ8IE
ne5ab6D2cXhb7imM5c1POpnOsoQxhfyo2ewUDnDi4+TdJTnpJdiO3wO6urCdW9gu
YX6JKDWfjnjkm3T8MzhMqmewgE2P/WfRCbqtdpvmV03TTZCTMMm2KIjFW3S7TV/G
K/k/FjCMpF4v7KxSGTJ4t6zjtZeoujtMOEYpQr3wZgQKNDwczCD3k8D6VtWEgIHZ
1LYZ1gaVm03TPCqIGksACxWT234RAYMaaVs/ZbZPvBrfcRtdLODl1tJ5HbDEhEm4
V9t9zWSI8zzyvs2BW+vE1f8+t9IvyqMFFXCUYxcLDE22UE88o3eMON3HcWuR35nR
KHMDYIqct3L6xJyjXwyvAZUNMhvYj0nSa5foq1+LUKVgj6v1VC9se3qX2g5jrMP0
a0/i1wZ+oYoyatWyV6cnn+ZHrPe4cVdw+NmDKzin35ZGW53FgMpAwQ+7R3Z0wfOo
L0/OZI7IU55qmIK8Er7OD7xuhSZKAItpveYLHWkpZ66zHWwD2ZjKydTUri65fv34
3E2o25WDS3s0K5Md45PW2nnszHtcpzUK05pplthiFHLM9nThStJeRLRVRVIladhV
+FysuBcycHktbF9nu+0N3yZRX5mqWyZxwW63hnhrUDLtOg7qpV/nshl6yyqA3KxS
REqPIk3uPZjB9MsKxgEKjX0oGOqIBPbIhAeTOt+sy/grbDhZMc3T0dgT6KgzjJYe
0PwHOez5wkjK8jdCPJroex8DQCmItBA6E+54D/nEEL/4NpIn0HrASu1X5yZ7Xun+
4YqqQVCptLdjcJQIj3tLPvTfvb4Qowl2h85xgSw4kOCVp6xvoa/vX4gEqhueaBK0
rj8RUXT01fJwoZ+0Xo2BiRULlNwNBdYlk3acpyOtOmMv3DmE6DXcPbShWs+DvRTw
bMJbERKKXD1k/DQ6UOYok55u+6jueG2jETqY/T2NlDG1TB35/e9c3PzUk1NIQ56g
X7buR7742fiJRvMripKetwaD6oNMqIgDZu9lgO+KiIxSg5tOzPbxkSRP4D6/yLNG
Z8k+qlJhYEQHXos883NLAGTWfrNU4PdYk1rL1WSj5HHjPQ6iX8MDY+Jy3OFppuD+
2ZgF3CLmLqvOyWuBP8jbK9VdGpT3CjHb6TOx9CmBwgawsOr3FbFOY3ttn+1YNW/N
vRVXOWhcn1zgkVJF3IDLUtOXIuIBcqcHmTwDb9xFSNCb7rbKsRHxT+d+QjBkdi/q
5NHrTzxLM8pS+ZazYdfJ9NOb0R8T+t2NiyNMR0bRsmxR9XRdvGpwI9TFaN1iVpaH
BLuIW5XAiKqBxx/ZStsHDKByUY6s8A2czQIeVgdTTKQtzLgRxYqxnhzvxT+nlksz
cyVjIuQa2/zRN9guDYeM36+hSXn+mKEvNvW3I5jhJIvrIVAnvNyo0HIhV6Mn8k77
etPUqnA+22zPxPb9Pp2OOi3+iL1QIdlgFdgDtC+o2vWd/lZ6Twrdkk/WKhMrf2YZ
JRx/qgBtrY0Yt17jvrmgnDB1sjZtxeT0O88nNaodI8o/wT9CsSAh8F9HUI+WLYlw
SJ8JfdBW5Y/dSXRHee33f58Lmm/48YqWR7m5vcTwBioyE+fIHiEjvhhmcW6NI9na
s7eu2G/DAvyGIN/v37vFRNfWO2Nfws0hjn/SpD1Y4EB7FhsvJTgtZwkLxpWqSW/X
FN7hfiexpx/LXDLigB9y+rIpvPVq+je8vWYWLkpz0pmWgGVyxxy3sM8gSH2oONia
Ke7zXBBJe09b5ToHyVDWJEoXvenun5/No4fJaPOMqSXM9h4HRYtwDBzU9+3Db0mF
LVL3OQV+fEeYtUR3G9KGxmHNU9hWnTFCW6EpzCggjAjVs+fmvx9GPdmkmBRPjORd
l8MLhi/L2p3taNgSrOI22mj4uI44C8zBI3/yoIe42t0BJbusw+90RtH8cbuZiljG
YG9HnfusJ+qDuXngBHVXZe8qNchfoWbmSzpCnDaYjKTKMQpLHHC9r4beV7G1b3wk
u/magxRZliW09wheE0TBlb4OTpdcZUIopr8r3tRASs3Yr4cg+oPT4bbvKY/73Htf
CUSUPuj476KDMlAKCtSyeDJXe3ip0hHRjQ57LS9LjUmCrcjhvRdWv0l/ZkpS+aeT
xeI7tb8L6dqriH1kAdPDlOCCjolx3GCvj86ZVvV7Gy1136iCRURnDk9ZlP878sGD
Kkm2SJ78c1BaPuOfEqtHaG0PFDZMXnnsFq4cwYpZvvAa0tnGZwF4mqjUFq70mpfX
2dsY8IL/rds2fMUUVM+k8YrWM++TBsRN13Uy7Gz2p9vXHqGBIIS6mBWbJc3JUmqa
b3D2edIrkZG+MbOrHjLMj6hqEMx7YxmbIubbohJT7pYFBTQVa+Pap4jIKgVF/8x4
YnCFTVAvcrJfCrj0ZI8GBmlM/66ESLCJBC86tDIH2T8OEkI+nEk65VMc0/9cTe2h
tIvNo1cenJLPWeK3wqbiCF5dUE51rmAXn1ZQJ/k1YkUwZF5l4b/JM1h4P+eC2+9h
0hlX8hKbr6rmhFyhhgvpAz+whq6LUo+NnFl1EuXqkE3547gK7DMt3ONbFixcTV05
GQCIFjJINs/Wz6vUpL7xBvzrhpSK3nQvHMOkdiRIeP2J2H8e1ZUEYZ7xdXdC/M0y
aaHCG6Fh6JAMTx4akkHNuRHLL0kjJUC/yLIAbJFG0sH9npEpxrQ+RTE5M/8RZ9DV
8CbsCzbkozR1YJI4UBRIMc3tEDYb4krp41jHgKdZrQ2Y0C7bZLJcjlarYXGfTd1X
vqZsfC2kU83YC0+/RloTrcT/JAIoCeYZUnr7bNJ/YOXMQztgbwbckQu3zpEk6/nv
ZIR2Ukyx7LvLXBME2gXkJPwQxQsi6VKVgoR++wkUa7HeuYhkCeBiPrjNAl6uRIYM
/g8eo1RzRvHtonsZ+bh2DSEUd5P69+SRjQl4SkK1qPYxlSqePpP+JFfI+ryzHYiF
UogqyQoGLx9Jho3iERLUWl3Lfq4qSUQq4sUuYqhp50gKuDGC8CQnouE1xZCcyK8S
Ztedjk45DW2Ft9CVTQFIZvUg3/Zi+C7XJDn7muKBrF90Z7xH0mHvy6xFPrggZ7aC
cW7BLf3HkFxfmcWe4h6eEcAvAd6QOJsOlO6scGyZV367ubFinkh2j+tLppHg4ThH
xHwOjJs3ZGi4Zga+0HsEK7Kgzsg5+WKRflfYitVFLxmbcohzkWwVdu047NLLvLW0
O3319g0ZdOvMmMZE2yItWB6wp94RAkyU6bRmfkIAdnuGam5bzKKgAO/ADg3GkGXJ
YCDq12Q7idbFuv2iU7+ok+BVeYjoeDc9uDSINnzauj2gL6jS0I6aA8I0sjIUf0Zc
sFiYWhyytbDpSLAcUlgeJzp5CRiWCI3dXjcsrbVsmejcTAoRVXjxweXdzlzXnJlP
GC+ZLXQPKdMOqjlFamz6uY9/abpcpYnB62AgPk5upKFOB13szigYgqnAKbpiGjQE
cPgMqqDbRGn1m341GW1GHYam5jLDCByL587mwjx1mc2D6I8I9htOlu81XDvFBRK5
DEvIADsFuzDp/M7AC5xiUppKOP6+bFAxZ9P9TXgHK8mFOc3oaVYUmloq2NZXMSfC
g6uV185jPmXJ9cbbn7u7mkBSNouhKGdQLCrDZ0lF+hJ/A5J7QVrEEVvH47jEMEAc
7GW0ReE3mEVoD5CTpUeIaT43LhMSPKU7qETy/C75IzufsOLNgTxnihjGhlI9dHCs
5rkKcfyn8uAcR9xsB+c+ZHN3Q/AC/HPHgqWgYFQZq1YCaKbZ4CrOij3lGboCfnrY
toVGA/vsa0/3t7ZluzN1e1VOTAsvlFXqOYlbSvXeXLL2vBu6Idvqy69CXK2Wx+SM
bjnSCfRUNVYfPGVemKsYo0MOXx+nP3K+oLc6dF7b9BNcD06WR7erq/expvOX5239
Q/oXkmdhX86hs81ChdfnSotn8rjBMwFsHR8Y/ucn8HaAFQspvbfbgCgM04sl02nR
2aJ3VicvwZRpWgd6exrpEVOTXj+C7rmA3vyeWO0g4ZkZsXJmnAz+VICL+Cxfct16
/J2YzASKZ+epGjX6fTDf/Z9i1z37JsSpdep5Nuj4t60vrXorKrVa6ZDlgBUlwOS2
LvOUbu0c59lweAtWZJdfbNeB9lhV6BE8xilaechTS2So8SsBnmNW16k1jA5R+fuC
jsd3qFy/RbovEuDwNsIlDY1gt4wbQ6f5eoriS7/nzzqZhOmErMuBD/hNSETIm7dO
qnCIkZ1BclPyrzgtY0Qq3NHDPscGIWQ8HbzrfNDAU94PmWT31t+OzY8lUwdkOkK8
t/Hb5Oz1FTuQrTvYZ6ZfJxHAOKSDWzoyaR/wYk3jSyHAW2XEnNRsU6su34lXcm4g
nu6rMvJcdSq1AE856JK3B3SnbNgTo3gANhq6gXP7ZIYqq34F/MUhgJ4VS3GrRpR0
3YA/Oot92+Yk0HrVdp+m3pHAF2mErQp2R7SJUFtyIM4kN/IPTGqKeNVLifTOEwug
NfCWqoyxwK1sE4XJ6Tj0HvcpaRQiKm1oxZw+t207Ht25iiZiIIAWXhstSQ+C5Yq/
/91Cyv2PdWIZAaUks+fq5XF3e9FCDKLYutdzCychEIBdNYqlAZCzK0QxxLUA2u1p
OUvgsOKuNeqv/Uw99adDrRpInfnjf1I2pNREIzlZ6NYCEki2nESatWK9KZz7HhzB
1Edlo9tKnsJzmIZXVuY8j3McQIY4H1KtULuZwpZMzlUf5V1ly/NvQyg12cy2bJ1/
4D066KKqiwWu9aU+XkDLWSSFHGNZvQZczg9i6MiJXTXPFpM+amqoOIb5z7ahEPrY
u/Ptm//AU1vyHIV8w27Je48/1i9vNpY1b99HwnnNXme2JdMlWkoszZYetWciJb29
8wxloJS5VrkCSLeMWyh47gqMC7bbCTOvu3zhdyREDJc5aOFCh7UfV77aTElAcP83
6lyIpnXE4lhMvvDXdVNkC50uCCwOtFXXlKQus9xt2jRIsC46nGkV7WZ5hereFoTT
NAXCN4qtgNBN4VG4vkCIFNsGkufycbpOGTFmlcXvlB3D3vddfKoNjPbf39dYiIEy
/j/l+2QuWFw1hnhuvT1MAGukjpP7wyVrT+SGS3P7X+VdRnftKItuKCVG5GfcUOl8
Y+vc6dqCVn3Ms5iWnk0i6Zk/jCw1rr5kJ/0k4uzxUSjhNbGWp6rZXgLmAq3ynAcp
WQEXn1hcN6m4zhxyfTnOVdZ3SrlJ1xM6qX+efmdZQaa6Yuq4SjJ3ni9cdUJ8Fs3X
KAbbNOvyu2NEk4DRviqUBj9gtccZnEMSPCIUKWDpj9JfNLhmXHYkzeuJjig1hsua
1BWPCbz9SZZSsbXwOjjiUezYQzd2Lq5Thvn3VaiTG4vRnTyKOzImE4vjsoRy/Bep
7MkWA96jXwyK8AwnBUIvfd30Hea7Lpb2S1+JNrzUZ2p+1bazBebnbEWScuNjPEoP
zHb8AB2u5TIH+2jvh8u/O0TlJUzuoyVgrjAITImtyZ4WXH4e9zfHnBRiRZ66zCTr
YOlkRPIdq4BS5g2PZmE8Vl8rs3O7isWsId8kTYHboMdL24k16FQZvTD46j4mYDmZ
6FEYhmTmPzHqpkFpesSbC4cLO5kBHMRRAPiFJ2C5yt5xOoEZhL8Kdcqku6itktdi
mlHzjyU0pJ27nDCfWl0GXUE8MvBtnJgcnPaZeZhNNwEjLvMYg5pBCx1I+LWJzDBG
ojSU6VZtlRQ7coIaMZ1nzZJWr7k/b8BADXfw8QZww3Py6XDm3nSuqq9bl79NGBCj
06WU7c7E/H91fHQ/gJ28gQQ+os6eFygHuHus6GqN9+i8hcrqUjmWEMUnshxnVYA/
jWZAe37SRjgiJcXbpfbvmNLInX53GHxRNW2+sZNMMySE0BPm/B6kwkL50aiMSDFF
kBooHb0yzC7vtpkBuN5ktsX6vRvh3esPh98hQAwlzFbzLTA70t84IId2G/HVT2tW
DVhLIatqsfDXkXji8mUhY9lMegsBdY6ixqHQSc/A8Zi8ZpicsAZ8mpAUEDq5wRTs
AkbX1CzkZqQP0fA3OBobiGuaMYtT4pk6RUXbEK9oJ8wyPG13dOp67rAIEUrCPmxs
7TqvesaIiatSYGK58JWHn8k3pB6yeIOA87BNAbOmFC9zaBP4ZSo4vogj9IsQaA7P
T/nRUXy3KWU4/UoTAbutOxAp8B4TiVFCLDkeXa9uh3ENS/wU14F0Y97uGqbY+yRF
W6mAmcgEFJ8vnGdZUImG1qaz1VhqcnS+zc4wdmdbuwB/Lu9/2007Legbvd62pVM+
cbV2XyiDCS/0yk6vcQnvZaniByQCyfOLXG057IEoR+KS5nADZiTEPrtEB7nVpr8+
vZolO8SPhogz54ujv1CxYDI0hRTay6PeZa+lmzy+O1GuVeOs1VhB5hyoTxNQ+tXe
zcnqJJlN3FWK65OkrQo7l+c/VTb1cnItDokXSDTo6Bc3PhYKSV5phpHlCSVgZySa
X+Cxxj0Q4jxfHWv7vNlo3lMiBpYwo6v+lWgeaKVTZgg+7vv6GlEUGFkA95VYhp/S
jbCWanNzxe83UChqJ6paf/rzYpy85FIH9LSU/sZmM7hiWegunT9hSB9Rft62Zi9e
LsVAsD3SpHC1WyvFw6LIXWZFa5vX+HTzTgnTkNGVsxF0Jwr9dJx2vY1hlvk1fkKO
UmuLveir9RL2lJswQ1yzjIl4N2lU168zmDhvoJNV/8lqqPizYpP9DthnH8YxvMTd
XitDlLswfiwOA5aGjYn0y57vdoqWLAJiJylH0k3m7AfV1EEBz8VQno5D9s9ffLYx
LfvA1stj1UM6SpsnyvzZGhirMadShDcq+uHwI6Vgdbep1vUFpfx4FQ+6p0uhsk4E
citD6ckKrC8r3I0G/ghcWeeU2SfiKUAkRYP9+sFh1jOaBJ8rHy8hUQx3HJJ/c1Xy
8X8PjMX/1EQbj4uoibdc7OC11cB5DdABkzxMkYHgglqpFt90S0wxiTVGSBUskXFj
4eI9At/rAUkUDdnR8t9o3vyfD6HIj2KhAaE0qsVgg2QMXpPvVXBivEmssTD2CjBw
aydJRASjMwlQkFoiBBQacXtasEHzQBu1AJxZI1c/lwM4Je8S50s8BX5hIQjZVqQ2
4lrggmb7gjzNmPErjYzp1nHjmxBsmIfKdBGJvLw+MQ+QI8TrX5Mn1Et+wZjz7gae
fUbMJOxlWWdBWRsdmi0g5lOLPQq8X4eabldbwO/gk23D+/8fT2ihXctyYxtChPTg
Jdl0SYIXdL0kvtdR6/6YYTJ+V7KbJ9RqhUtzgTmmClhcQ+qxmG/Yy57y7hsbtzzK
jE2msYRTNVxSkmSMp6gtlDhDsfCYsGgrcYDc0iFJ00Vn5hYIaZEwdbs/V7gbb3PR
wpWlGPeYqdAmkMccYCuZrAqUSWbyRFIcvr8bQNCL/vshkx6nRFzB5aKgh9iQk0dh
BaJ3wviYXfnY8uNV0HYdQWIwWAWD+eDScdSqikX75cPujF0qHs/UNmtDkvXL2CbY
HFJFVD7/iIcXd5kZdIRldKM/WpbspQZ73xI7w0i9C8e+m2Aq/ggFW2gQAzdRzskA
WOCCwkjMsGLBBVh1EDSRgVbqSccac/LNcsWwi1RqeRAhNaSwDZ+rE+Tb1NbvPLW/
CwCoJON6dV3LsQQ/Me1atLjO3rut0tn1n0pj5LnkrP9x3nGXCdggrAKN2DGzawa5
EzrDfS9VjBQzL7oW985b/stX7PiVCvi21+iVnsL6H/vxLPM6JTMZMfDcRtG0Gty7
HjqbjMKpDNIrdEeouXQeqoJL1HMaPRk3qsi7txDD6CjV5YPtdBbd6kg9AtOL5jeR
+dviqBlM3y7pJ+zLupwg9O/FfsmmazT9xHayitxskV0rhRUI9ZQjAMo3zoJsIvYC
zlIKlp0BNYKfOmy2NsaMQQ4S5bZ5/HvVKeJX4YaQxlU7kQMWFahGmSKOCEMQ1GKT
4Z0/gKdZBHWVLJvAwQdgZYKNTBrl1HtlQZOwQD1oKJ28A1fAJddtcwdmyWR+Fz5r
dIKILJYQmYk47ewwiXSKOM6doK2XbyY+oIoVF8fl+vMgy9Sz2Vo+L3xYRIRWj9qS
rPjfNYTj5XodsgVzfecxJzOQ8LyQPWghcj6elVVek9bxiiVb3r8+NOJLgPqgP1CO
rLykXTg3TIw2DeTNi7cGHIPk3zHHPwIkFAKdJabpoCLu8rGeyIUhPgWnBBWxPMgy
Fj16lIoSzTGKI+PUi8S/7Ur052JotdaiI0wPbg1lAuN2NAVBy7ZFaj9dDhbfvXHK
gEKSn0FapGyvgYfYYftTGhU87D/aqbOmuPAKkom7O09lelAmk+jTcYgaLCI2TJhA
D3/OxUd/V8J9Op9Wq9gRAvKBivAh8SSHz8uuX3wQ34waCGaP9LFBdnUY5kjLk1U8
U0E1S+3EK1JrnSwjtR+TaXKoCyTKNyDMdztcGFq/goWMMQPPPUwYNDvcn7P39Be6
l4c4OcUNamwsII4fVOxAuM6h040OKEFzniMQ0AK3kczgpj2acuAHSqrZSGkLuBiW
SIurm512zGtm14KyptylZdUXNURmbZiQroltEoTU1Edp5Rk6xD8ZY2kyBFR5dTOL
rCIDb7uST/m6lzwwKm+pwoU8i3s3/HfuFC2uEavcvdfq1+nsvF8YaiqjPPhbtJoK
MXQY9oM1ZExHYePPApFp0uyuvhiczgAYeAuX5B52ILE7wjeH5h09fqBC5pC5MWO+
VCNIDyiB3sqlM4v0ZcIQHxyvvB+D2CaP2bgo/poUP6+o5Lf8/ER2XQZkQ9B+Kzdd
FjBf4Z1kl2FmPEvaygEt/QASqGsLxJkr8Hf8VM9fqUDvXwadH5uvqMPr/gl/qiYF
WEhm6jdPdjkwQMy3CMjuUSvuXTCtHKHr/cglen5F0HZ3TV05Hxwu+PNjmKCf8qUl
KUJ9tDx7Br7F+N7RQeQT6Di8AOdrwC7hpOJlY//+FohO0nmglcaOkgsWFqH4MQ6q
9h4Tc2B5NeSqUgjikZEYdtuNt5rEsfsvQP89mhlJzdkhIhfJ/EaxiLUur8jPBWD5
CaxNV3A7iHe2BTBkWEv3P1VN91kMvq6QhWphqSTO+A9dbaMuXyNrv0VWfIkCBVMX
0WvT7NiXJxesPx+qqcH05PwI/3ujdu5bWtRwI9vna4AE2PJ/9VxgThUzULwQE7Kb
surRhAuz3OtVEjLVeAAnFQRRXs4Ere/KMQYbDdpLRxxGp49ZjpIF/txpcNlBR8JS
dyBoghbgaI9BnM1ZsUpMiq89UCZ5rHagWEagTcaXV0nA+DJdagQVAW1Ww/7qEuiA
0Jmw35+PuMnYASQsCuqp3QpwZeakrnhXdupECLxXUEPMWXN1msJRG9GplqJfnHJ7
mVuzqE900XXM/mHUeuxdwR1Bs3Js5CL5s5Du5YGnyOQguY/2NKfEmc2zjXEhqSmp
iQQ1visWrRPpLfdE3GTMe1d0bWZcD3hj3KekLeWTF8dND4ohecQWj0Ty3/xQfoFk
qDx5EiFCVgmqF7WM67erM2h+G0/DpsF7K1vxMxirivfxevYpNBoUdmRObqib0Z3U
+NTFWG08qpeIfhlQ9QVKQQDs4rc/u3yGxIte3X+Ufj7WWatninmMdG1F6Rk1qZBf
fCB+r23d7Ma4qYfUK5rF6hdwsFW8P1TUoTRzybCNhzYiTuFpTXhylc0HL2GXLEMw
jnsgltE66GlmDPp7rJa3PTlVzbMNzEt60ZSgBlq24BPltdEvX/xOKQS+vcDOzoGh
Jw9yzQh00B+we44t/5qaZn8PBbXVpG64zBm+M221/wyLb9HoNTmTeJaiTOS5p5yf
rl70P5EKnIKJSWdlxaMpcvZ1vmP2f7RgWlDZZpnv2D1klqsDLFC4HW1vRfyUJ6Fh
X66IrVCeKFm3pc4g/OIW0rlEm3C7nCTjGoLEsYRnQWJaE+UKG+IsxNxMJgbLcFzi
hcGIcmTD4B7mrqg5OQJTdWSKHV5NxaVe6sDIS3Wq+GUQnO92haRKVpQUfxgW7Bgi
CSaeuzYM6/xiXmUZ2a89lzcUQTK5GYUJRjtYz3Q9pL454kc8M/KqM5bP/bvahw8g
ONw90nPP5OIrGgtnWCfo0lyMUKy//LNRacF2zgcxvlIMf2gEWRokLTR46Xo/mM6j
Ed9Fn/nCWvQzb4AmXdLm7ooQjXVZR43GKLHX027HSrSgyhbKrgZrsZmtNc5o3hZe
T3f9ip0lzLWtsjL/haBDca8vO1v9V34+FUu8fxKW+iwMGjEBY/yQAD7AILtz7c+T
lDQLjvdi4fEWX0w5Cud4M4qxSc/3fy33NNB1qEqLutVODamBZ2GxxprdGTQfzj7G
/DKxKM+/FUmDFmnwZNleHPxp1vFTLuiHgFB1nsJzNmD6U39MjkXbw9e+onmL084y
H5Xd/NgtbMvJpovzG925lOgufsNx4pRtKQDdZUdQvgMwqbsw2rIT1Yxj9SOd+Fyz
gaBOAAfWwATXzxCEX4QNj5Vkky8KOVUgBpiqgl5BOmHf/pSvXksyXTwwHVpP+fSs
pkEFx8BHNeWgOJgq5HNrHP6J705If5+S3C3GHkXnRqxWXGVTUEgNw3NSc8MspPFW
1c9NezSSPJdsjZnfKo6jfF5cSV0CgFLtKsqo22jOp1vEtC2HJnA2wYz+o1DSuZQG
NgOvDnhVvSJMjmU8R1/WtYLuxR+PjFv8VCpHI8PQ868yYy230dd9NMrlohToWenG
a35/Ve7K3CtJoRAZySiKwzO7A/Kv8So5LQ8SVc9BrBKCoviiWoAr+JUsaW7/YPNa
MCmkO7LvH/gze7hqVTpHHjKunro0x52VK7T/crjiEEdQ0LovatPls03D6bkwX4U5
HJTWze8t4oVSJ8Bvzb8HsVKSngav0Gn2DVtkwhXMcjocFt0yi65bHQsDka2AKLnO
SzRjXD5h7aPWjTOp1q3Zca+E9JgBgRZ5f8sUdJK6K4ZpstbsKJ58yx6nDq8mZTxI
NgGhcLvi9T8njIhfm8DfV25I030ADSG7zshRu0eHmzt8fPDjIOEttbHOmym5uktv
zTlmuFJY3VUCaHdmdQc70XAAqLDd9O5poV3Ub1IRl0nSlj6LaebarV10ahXuwdk/
6iSlyanbQvpdC88reURSbEgtRFStAc5tl9OLYdW2wq6L0si0ZM4SiQ1nYjTlYRft
TQqcW2e1Ty12lPODWn/twrbns1/qsMW+nc/mei99S/LajB1x+CwQ3MHN0EBWmuU+
z3LCtQ+lxE6qa3NKyag/1b26nCq53rFQrRMYnly2FZFvHFxhIG77g15Iys2N0cf6
yIWk5mZZjNVz42sUx0SrOISRAw4O/nazC2n1hSWv/qf36Yy+3FGM1YhUZ4vVDstC
uHA54fZMbKktSZC0WAfCXF0yOAkOUQ6CKtMhwO0Ins9AJo9PdBlpxxgisuMGyNWT
Yqp1izvd/3H9FTQk9EnVg9dJ6dilgDEaiE84NreJ/i0IGJr35OZ92Pr2oT1eODMc
yokxCH/7X08yuqiF72HQs4u8JCfCbOkT/wBTnbjpZmmoU5vK/XkGZcI6NXHbhDaX
OflzCyrCPjPC01TmzgKKVSV7ivYFNbwwVagR6DKGa79Owj/t84SxcNCVx8DVapLl
yPoPeh02ogSLeFBwm77mwuD1Xnl2+wzRx8Ajiewughozwfb4X9VKex6hYmFQyMdc
rj0KQq6cjxg9X8En2sH9nPwrP4o+5BGD43g+Z1zbff4pafepS4kTJV2ZZGA9ZNya
ZXsDidnYVoc3O07I+M57iCqBQBUv+GohVG75CjUD7KvZcSMmISQr69Oq8nbC26fv
YAY35T4ixGID1wcQFtSB27tv1PPTotJ/J7ym+MPjUgauChd25PtWyTLwO35ThGUx
sGNNMNl2qKFKaxsfK82QRyBilv9toGStafvvEo6S3ANoV+66o5fPP4Je7YJyodNK
kiQkli/valoADSztMe76OD8kLi6cErgU6QjutBVvLyPGbejsUg9fdwmkRXBDMY18
xatuabQ2AHCLlt148Mn6XFRhK9KZ5hYeOHa8IJYmVz3MsNi9cEZ/UENh3fobfewx
vQuqE9f3PjkN1SMN24/Mr+EPX6q/qHCp7HoqR8pkq6HAZkJtLEsl3LEfXgbUjtn0
IH8m0iFRJMWVx8hRF+Jex1M/03oPSGNcHn9WyHDHExy+Myjo8N+PtVwQNd3c6Ksg
dH6g1DClnxcg+mwL/001o210U/3ImkSllEO6n6RmMDd1RAneheL1q9RcQU3ZM2NJ
EXS3HLBUCYMJrAKw563lqIbvB7/8+wJc65mchLTNO1iMyYQgFuYPCImMbGofn2D6
NhgqTYNmYFaGjMtkY7J9mxFa7TMMyWga333uXK+pwCQQJf4OOPTDcYL5/usXIIT7
CyFdNk4L73I1zrCB+DWTF/0xqfQhwG90QvUhQS/V+r75vSt+efbL8IOVANNJaAEI
IaCk7nseGgYoNtfQz8ioyEJIS9m3gBsu1Bayg2GgdLc+TcE8jTKzo2m+2TVse9yk
N4py7mIP6CJGWLvkAtgqv9oInre6jCDtleDaIcIYb77ln3VFx2DwsmEQm1eJGOtC
FZ+I6lfGeqwBvwtk4hYpUzKuealV+UIH6ICB07D8oon+AEp3hNci8vb9ryG+W3sq
1wjxSIJe7w7LJMOPOs1sFvnRMfmcEiPEpT24ZwwrXcgU7LwyeRtNjFCyiOXJ+lcY
uJKHBTjKnUn2TweJQ8t7RsuBBr7Ke5nsHGH86toqFGQ9lvRyo97Mu0w3nhxm5+SP
j6DOBQJxdz8pFTbPQ3L55zOgEe+11beq7lzizSs08XJxEYiwAeO6q/Rf3tOCA7xA
D5t9TmJJmDY06vIQ2jYemD2JGFMA6pNCJdOOGqlKh88cMTcx8zVA12h1sg6ogOZw
9GDatLcpRRuIhIg+u+RGpZDHvDx3gV3gywg+ryKocoRasrvDOJmv3sa/InmhACm6
mN6+31H4tA7nc2eIJ3pS64xNELPrx4WbLAReOFbVZXOu0t2tjcjRFYGnKcKAqgvF
KjCoqPPvJXss31MSEL0mSSbmeq7MxZu+9KbCI4OvdUaao8KVGgw9lxxl7l9/w2YW
bkL2ayjk9kY3RSxuWcWiON0N+9ak7XxPfL/WVWxkhOEV2RSIDMO7AjpKUZR2V4am
NrUuPcKFotms9sIsz757waFPrFeb0KQ6EUU7SAkdX+4hlUPZ3aB7UUm4x48rjwhc
TKNfYBWGH/KgoEo2W2kqzql8MYlVm7i8x7Dhg0EgQByJSDGKeTe+5rDHM3Ss8dgG
JdiFg7D6WVQP0IdxH/kDUgeJgK0mQdxVh6fu/7+N8qQZi0gTm7sEXGG570hCzk21
t44TqmjX588yx7/nz/5p4qMKDIIzttKNQ6h5tza2qXtKr8Cqfi5tO4x+scobs/mE
gmEa5yaAqlsSvGZBATBo60fhTRZT3zq7bkOoo5yq5RnkeboXpjvWtvXXu7tQpd+X
2RUJu6YcY8K5lLyvJKRfn6p0OGYmxpjUkihhAUGqWwpKzq7jq8fex5QdmiFnt3Vi
IvvJDUkV97qnuIdYom2Wihyk0a2ua/VmSZpjjf8FvPTpwsMMHs0xSkplJzzh2snL
OJoHlHT5CSnmBzq65DVoS1U8A5Sa7mkGstUThlmZIt7ITimH3cNkFKxwiISWfdn/
GlW+5nNNyqAFxW5xYko16T61apCSiIZFf/mVm2rcgF13OiBLDuz6H8PLcEa9Gtwx
mUDANldKqZxjeUpietw0TQoXw+eRSO4ZQGIF876BBX8x0fYaX3TFYPeJVyfKbdS/
aYCuJeTKpOtoRY2dzFbiNjNObc+ug193dm8NPlqUN+w9hTIkf0/yLT9cUoy2kpPM
gaVMlQdpna74Vc/Ryj5cB7syQkBwxxB9Ro1zGMqmslikl3k9Waugsl2xwLg/bUnc
IpZLxO9qDIO0OpLJDR/1ePqRQS3ZbwGilqdwOHk2g9Puxp8OzTq31BArjAYLCFWJ
+7eSt18FXyw8ryV/eMAXgdNNWFip0EwtuzEg5py/n+FZH4ZeGYyjikS06ui925oZ
QAFcvNkhfeWejuo2jLbQe0ijCfPZnD8YwxQhzQhBg5ewFocakUU7cT0S2LmRN7DO
AusMqVvzcxrGM6dFjnEuoL3LwGBoe/ZZrA/eOvvCKHIuVNZwTH7Kf7k74OKllW16
ceIMVq9Iy8JNrndC5+CNoI3xvEIpRJ+VEUXyhSrl5VWtfAIa3LKj+nlbIDnnClnn
726f79gper+TUDWiHPxMGzCHP3iZknp05kl4Ro1GXhw7yjUEEnslaedimKKe9Bqv
p/TucB5uTdpqoVV9h3ZHGEOd8zN/h1Xk7CkpMac7y8wiEglKSc+eVYyYOZTfBMEN
vUvx7WquqFTLYYmDhc7sKQxdvIdmTT9CvR+e/paNfjTSEZNDDI+L/bvMOb41TzT9
yN6EB6AYKlo21Z51jOJG46x5ajeDLDJJSqaV/FOFCupWm+MFN8NJKj3CyVvn8mIm
TFMPqmRy5yZuC1iAFCqc3RFkY9VEOHFoFh3MfxbEnMcoa0Rq4VOkAjfeFm53m876
Jw+zXu9oPPkmNoeO/CV61w13zHaxXT2THzWIJ4CTMIH31Ep7oKtDGE0iBZcETseL
VGHF6KpnpikMZpAVAtbppsYljTp+VOljcR28WeOr0Vq3beIcGDqS5GIR3havHiKP
AeHOvwnk8iTud0GO2XpgWqvxcSa1BYx9opM+e9BiW3TPWNcBYDz+uRhGi0LBjDFT
5o8duJ4FPfVMRiCRWRd4GZN1iqxq20z6jXW4e0k2J5AwzKZ62k/X1j608mHEIG0H
Zg3bNIeLRzaWh8aMSIcpr4PUx1HLgaVG5Bw/WwdtrPUIroa/WluW3kNJ0zym6V5c
Q27RuPpledPJYnKtoY4G8pDSAn7D0Z5MKUgIotTiCmUB9h0kCXahQPvV81cNB+2K
JGkuz5GBMMF/ijL1maYTFsgt+KuQHD7nN2TOL6i0bvyXUtBDXnHDP5EiMIQ8LLaU
DqKGcOTKYnNeiiIJWp/X7cgntwV5TmS+e+VFm9eCrGbCmZC1XaNmvrsy0kfjAVCC
0qqsOsr0iFirOmyzp7A1noKWysLh1EdtszaKcia9xRH0nAAY3wUTiOnGmOdU2nRD
xWUXxdcMosoK1UMF4zoef1iAWkecfE3T217TPOayh96Y/b6aO9vGxal6veUhwM30
UA9/n7DYXaJKunikzWDxJXno+VSoXbc9x9hvU87adi7zIUD+uTvm12NGVlcQNfAV
SQQzI1KK1xfgMZeVLkMZczmNNCuwJkAYo3D8GhDMA3FXhlE9UbMsiuGtOJrLehiZ
ueHdLhxiTlAkNYUjoDKRr1qa1r41BQOUgN2h/9rY/EsqksHeJuZff91O5Bw506o0
A2cbBCt9hIuB1/6QwIwZVyyEylsGIRNMpcRgpYQxzevkvPI/R4MDdstrr9rP1h2E
oogOACuwRHILUKsMi/bj54OGXflV+ZbYK59JPts0WGhCqVxkbUnJvahUybVmQ5S9
9cYACwaT6TicLgNQPV/v8sdFGhzLBB21iRsKjrLMTBYMESs6DFlCRapxeMxRQL7A
AiUTTzJ0Z0f/VSmusCqBFXx1hMlI4+t5NYmkmWT7al7erTs6EQaURbNxo6OkfpEc
qhu39fdbw4TAt94XE7q15dI7SQGPrTJFM35anNlnfiaxxzmEPihqkU33ExXosxS7
o0lVHPLQe/nwd6pl4Jwv1FmW7GOfmcS502/o2LrmMr3HX/uhpMZ1WPxC19wyXHGu
xAmPKHhbmfW1KQP4ux6WUKi9jwJ54HuzTLXY6vNXxsCT9iM2cYFnPbx7SJIncpMN
7G7eAgSl76GjgWQaiUp76hY4yZItUmYS64YV8BPHaGtDzMMqWSEwAHhIJUcePquZ
4rDaVWLTghx1mV6hnTFq/aoWL6XC9hSLX0zWUPuaHPaKANnbkr6eS99JNHLVCq+o
XxwWogv/hWIfEnbiitezrdmsaXNVZU82J3Bh2utemJ3S56j6h0EAqzwx5o5CgQXv
2nfmUBejIQuRQE2ft19v8qI5BvMRAl10YnYGsovv7uVLiAfDRw1Prf/D/rSGKI/i
hpLExSb9S/metbVMfsZENo7LaoQ9szTczv2l4QhCVHLxzZugAynPsKEcRhjpIx9r
0EkoyESecXftUOnOp5WgRW5lOJl/RF848Ety6eQnKb5je1Ad3u+B8n6JWuQEnDL6
FWkuZ6xVOBUlVTNo7awj6Fi5E38n5D2mXhqL6kCMUJoBu+ezegEgi+SaA98vxdzt
M2SUW9nq/ZvR8vFhP11kMcHu3j5zkNHs/odUrAdjsQkU/6hz0kPgBXuHROJiMcYu
zOWOXccuKI/mupQsL4rSPCWImfQPbTdKOIz56l1WTnYC36TpI+Ei2y0lBxJOvmYw
ERaynHDW1BD5DN5O4+F8dK9B5sakOQLDNPhw3/c0yA9MfxTAKDgWR75A+gMmgVnV
b7LynRURB8CwB+ZPzkjttSb/R/d2SO9MuLenA5S9QNG4Dpoy9+tHBJy6XhaSezr/
yEgkxJZp3NkkF9dxiu/8q5MDLSWuUJS8sLb+g9X4aTCMmnNHbz+yRmF2Jdl+6xkB
G29STY2kdcgUqS7QdIJRBU5rbSTBcULxT2cjTYGI5s9mnrM6fOB8DxkJy/nyCc28
0Y8XDCS09azAJj1sISVx/gx348plKMnJNkWLgoHXnl0X4UUqGcR00X8Uc5Uc16zW
pbCwBNIo4E6osWQWXxr2mam4TPbYxKGFNTIchhZXEjZ/6u+jMsjzKoRqwisodciy
nDiO7WbJ1fBRDqJsLkUgRCuuqEBBPWHVCnPanyrxdLjHDVOQ9XikEcBaT34Tq82A
ovCZDl3c8JJLdMGcy5jcZbB1ILHZqlGex6krLX23TJa9w2vmiEsZx3KzKFNDF0ud
N3QpdqY+h3P9t7nfsqahPKycqEDzw4rzKqsqBrCRVr9ls2sAidghRz13n4+5ZT62
w3RAXXaqRnSk6DqBpVTuypTIaT8VbcREux/2FwY+tv5gw4a+or1+OFUQaALS8pj7
N0lFA4PBcU/gF/txGEx/mXhLjtjiVHC7alw0wcqTvI/5XyosCPQCgTEWqn1GaUTr
Xdhrp69SJLDDoJIf0nhM2roFlFvTh/9OHgw8/Eqmt6FWCuNRDZEmyxEgxzV54nNM
p2Y/nWKKiAaYCNYtDgxeVSxs1j01SASsqY7fFzDlF2h3ecyNfIZNIh4z9gGWA6TR
1R3Uz5CWganbBbXBUXudor2e6pHw30LWlxNTEf5jx5IU9w8f+c38kmjHNIUIhpGi
C154p2EJ2g288IVupDfhNsdpbkscxwCdUC5HMiJpRb3QwkjRp8affEJevzJsXRpm
FQSmDpIkSn15W9zUkKliRFM8uJ6myO9l15JpLYmKq/7WVIXyojqPBhHHfW6PIbri
ob/4lmZU0OUuD7RHw6/3apS3iw6BNWh67ZrCxXx+iy/gnBe1OIhmIzog+6OM4NvO
Rfw22DdI31K2facc6jIbIfGEVJE0qaYFl5N9qb2022wNt+Iy/jh26TQtdzBMIHkb
0jEBoKsVM7gLEzR7jSXc3CU+etODPuyAwJEPzM4jiJdhk20Q836jioWnAuOcSuBs
qNcjy7sjDOqP8LBa8V/Tlug0mz0kFs8/fJUKQ+vN55DiJrjCRmPfufGnb4r3xQc5
Lspu9sRrWlb+dUZ2vu1lqLceXzjPG6j3K/R5/QfRval1W+DWxHhaEa5tdjx/285B
lgVNHrE/AEFkIEyr6nc8CpJu0vHDyhRNQAp4t/SOGkT/ykSnwIYx3h7R2w4FyvWA
Yco2NHS/RQ6ZgRV+bUG2jazEFbXTQtYHkQA8cxErGN9KeG7i4SGv+YwWHTcMfmcT
gkfwNkWC04l0BHSyy3CLPc5JZGm0M6dKy/z06pBn+r5CCsF/5gFxD1NbltuvsI52
PGls8pu9qmTxnS45D2DUyu4g3Wxp92dXrnR2zNoR5FtxHYg09TDjeI9ZsPnzwk7m
uyxY2CP4okSAmWeAiON8T8a/HyMvolReBkgYXF/3AFjWJ4rr3DkCcepcXWRcF+wt
VTpfxClS3ZSyrElyI7izws0A0vJho3rPA7FQtWTAsuB3lkRo1YK7rgZ1ylYkIbwf
dFJA3VhpB5vgQy99Ljr3T9Xrgr+jaZ+TJ3+Z49I9PATJ/1pcCItWww+tPRct+Epo
oOz16GAtQsasUxuIyBHww/W7WDvT/tQnJgqI/Rc7ufC7duEs89KroRgsJeV1VZzA
x6pt1bS/zSDyGOeI5w3Xrd0mIGcsjk/hv6P0jSC2iZbzToR9H8pcywzPGQqBA4vM
BM0dAk+2GQq1Lnx5ighXloZUfl3TqmkCpfw5aqoPOqs3bwQW5XFd/UyNle4vOf0g
abprwfuAIhTDUQIJNDjfKn783tTR2OFNcrwaohN0OVG7/Bja1SLN633zbNPhGnwO
NXvaO/xtn95klnLhHHRsSJQZNc7nf1m3/RGnWmEPRItpNLjwtqpdIe+5dYyrpjYr
i9//wTUqecKzEAGtYbckU+uZsRh0EA88l87c3q3qYmFrlyNQzps9jUdKZD2zx0at
p1iDGP4hEK0RAEBj2FIDm/R44N1EQD3l4rfk1BoHKGbUNpVEsLB4P9Bt7/IIjzpv
3vwbBz08bfhGrmA1RLP6K3oAXWsYko8ibX6NF6/fmqhGSQqF5E57csa4mMpoBs81
vMnmZCrMwCBwO1+A1rN8AzHaOZJ7sDDF+CMihC0g+UWrI3vY4Y6OUA3vky4mmYzp
tDo+qdA7OLKzoajscAc655hQhOqFV9O/RhDFEdPQHlw0XcujeXga6zUkTuSL2aTb
ScuCx73QUNyzNRpoZw3zv6FgLFsFqLZTMJQT7DShTAfAb9B5c80uoUL2/gkY7UTG
bPC1rGkg8kKWCUplUzojKXHNRh5MIZC7GtwKe/XKjwqvHqM3Zh4vb2GKmzFLqR7+
62NkurHPRIHU0gmFSEGsufyTsk8s3COPByPjqAj1pLVaQovs2uRxzHzgOjnPECMk
JYoXC67FJZLP7tdnnH7o/soqAw0lWTxNAuv32GDzHaZoVZVvuDfy9+Lz5mPumbzh
aLG34+hxqMnYAmwKUmJKff/aM3vFvltdfZxdADJj6IDETIMIGYr9N2jThGnzQ6Hf
IqxdBaNe9nAxibTb3gEFT71diyeySm56d0fws46UV7R+oEG7KKWhopVCpJKSo0B4
zOfezPraKSAlMfbOjL1pEueHHJojntdULOa09znp7vEB751suKuOGC+lX62/URIE
f+A2xPJky1AAzJ9T+dOSjohwFnQN+5i2BjyQjLDaArrpAzFXi6Q4XnfkpZwg4cGZ
OSk9Z4+jdF+ZJE7gKtAkuodLjRKOuohX2e1L3d3fpGXHqnhLSVxSQ7yKJO+mFkuP
gn4UbFlkw8MN5aE1dRdUekEPuR1y5V14IFjbJoPymsqf52jjtTWZNc1PAv8OausK
qhTPZ21R7VCTKU18N0i8jm0x/gtcXhj5eGWKTH9DklFJDgYbyf7n3oRpVTDyLppR
BzgNpsCvImzDBJajkxWrGTjaOvgk8aPFtJ/Dj995qUeujuiW16LTJ9QWgSBiKCd1
k0Jt4rbPf7JDMSSjVN44GNJukqihHW27/SonG1mjeuYY2U/dbK4IG1kyoKDCohp0
NxEOmbPl+AabWFvDBiaNzzRjiyUswybRpvGOgex3o9LdsykF5yVMJNQdWxKtyVjQ
cuLgdnSFBVFFcKeDQ0VH7zVWVgbT7g2dRG9Hyogosu3mt5y8zlDYvSclKhQSIu65
lROpmJsrjuaOLB0vVNMRlz+Uct2SV+jsLuBeR4jcDPiLuva3MNHKvUa+i+h6yEVq
8DMUHjAo3dJ6U2OIdDspc6ezFtc+uJvqN2O6sBDCQMKffl7A8QDm4COVhc/dlQ9I
KUM6GlcZwGiVP4hvzE2ZJ8COKGso3DQyM7TLCXOd6j8MODpujv3jyLitrITAepJL
TkGWFOXBFkgJTwDYfy3/MUUrrbRxajabG1NgEsfZgvpfwpPgCMOCNIDvx9N6ScrJ
8/OTKsyep2IGKlnYcq6UsJ+IOX3vPFy47JxeMBzSGK9WwTYm3+BglxGHgnGrItkG
3OHtsXPgmPUI/noqXVNDUHZSRPMaJSLenGP5wBAq3St4I/t1nEn/Jg5N6+f65yWn
fFNDvwFDPq5MQeI5uYzarEmFBhAu0EipxNIsAYCch86pQ9Hes9p1nCN9ObG50akj
CwdbzaZgdOd3WZIxJG2zgfXHJaXZuT0mRHg5EOh636B+8JOSuGiQuJKRsk/lFYvt
4BnE/M+h60sZYT7dDjsnFhw5/f9enFhjGu5owwif0+wnJ3/3ew7OLCoKr2e1xxzz
R/BHSdUsaY8rcpqNwCNSluDzbjRn9E9sYC7QCyJ54tjwtsPmnchphVEBy9RkTieZ
CDSEhbP88miisbx7TEwXaV6X4ro77QADB86nbnowlkFBUxTjwjYf8BSp3gryal8A
r4lHObPnJSTrZKDdIppU5Spglu17GCCEm6eD40PInwIM4ryhucVsUZOpGCtbWtIz
DHU1CX7eRjNPVHzlpP85s8ifSABjzbuiD9ZGDxCPQt0FKdi0/x3im6PsUnj4MeCI
dNoLqFYNTD/TNuDl4On4RjDE9TiNS9UEQtmm8Pe07kS8GJ1zfs3bReIkEA3vnUGk
AQ9MCP4jmCp5jTr8vm5TKiluSNJti6aL5SpzVIb1XdqkTpLVHKMd222FGP7bZBZn
649xCF5MA/pXF0fadBEWUXbOiRJNrZ2FlUXNoYIhiguBHCo9HBz3XC2SrBxMew62
oCEW5Vzul7TKjLktrI7W64xhrb8xxsqtaXcBEH6ZyGvCU8Gcx3cSCGfFcrZLFQ+j
bSntiLhOh9VWwgfLPD9uzPjBN/MmxVNwJdA0Pybq6Sb3QkTYfYWGbKGPBbID2uAa
s5GAuERYaHlINWb+O+6Lk8qf9AdB3aCxb2EKIBFzuD+O83sz7Wy7DHLC0mIcxQSG
i4nTRw4W4GXLmebJI465iSXrOqmDgvhUOrPfW0yktTw3qU2v9OKP79KzWGbyWKhI
3z9iCwhfjSdSWCIV4DHvenq/jhMhY68Zw71RiWU0Nc9vTs48jfALKW6r67q4mM/6
HpyYT2AVSjTMEC2grLR0UBSkjU51MwbI5mJdJjqR7F+PU/ReyaiY1J0ChOp13lln
aBcQxpRGs7KDfOwY+YQVwtFyOPgdJ8q+DG4eIpvn1Uf1HvMD6kzdEqbMDy6uhNd/
y4B89A9mna/1eEdu5SNupraqqKlA7HZuMUcIOQt5jJbb1l47ZSTwdsZg/sbilEOS
k34QDB+/kEzocS6MF29E1vrtLqqFBmulHKmL5dDaiaGH7qV4y26qHUez7n5BNPis
u6bktuaju87w4B02EW6gdXIcmC3SCe/J3qimwlTX5Wtyif+rNkUcEJ61GlT55h5R
GyE3rCNIGWEKbz42Wzk0wWW3okjbNGkHMPRVRuuseuRrqwM4lXI/5GpIdRbhyrSE
iEhuzTaCM/NRVgmEpOJ8Tyckw0IYXz56e0V8uD5qmIsZgzdaUMK5Ottqq7fua1nQ
gAOMF0p3oAQ1Y3F9emIAd5V5Z3ByRzJrKp1n/amExLE+KgesOjm4R+gJxrtitIMe
JWiCGXM/Izdbem4gsM0iZiUy6mUNXdN7RMhbq3gD+cJyRk4emYpIW6UN4VuSKAd2
J4eIo1RgLc2rw8j3j7665PTkv72eK0nvUsNHkUMFZYBo2Gg+zT4xQN9dJqUR6OPw
oLh+F1nUvQlkgtC9yYEzEIL4JaaPxyWP+btAFLo43pwABPYz/PSxbLuNDEx5VgkK
0JlA7XHTfwc9XFMjEX6XzlcByhn3DTSLj0s5unTubjF9EuP8exVXyHtWP3lTDXjw
LOcCJTGjuGNu/Q5cYmvVQVW6XsbjZwpoEVwaR0ulgak3XSN/b3UJOyelbvQLNX5u
wUAuvP0u2nI4SYLnUbtWPIgOjnCBGtUCtwQOIIwXabPAnpaluEfLCavOE2fZuR24
GXWFvqKkmvaP8wihtl4OkMWvTtMr+GVcf7e84RG5wKyve7JHw+rzCVJ/q97n2oJz
vxCnKQ9F/2M16bwtYLsrxGBKzLchyQh0VPUtgGjaJgaiFlnW9t0f1x/prtj42ItL
Eh3p6enB8sMloi21Cb4nXi2pdwU+uy97IkgRhs6Ayk2pwvrxMrxUsmM2koxobVgJ
idZZVN7RhYo1LLHHr4fFhkGwwyqFUXoFVGpu3lUH3khhcGyNQ7t1Dr4km24hc2c0
fQfhKH+bLvxAw9hQ5TFi24zlSk55cNsYUnl0lneaHWCpFrs0QwignCSLRvb77JJH
3Zs0LTAV5pSZX5l2PYLaN4CV7ppDFoIDwHWnZyBdiBk0Yg4eYf3nSnFst8iXORv1
0Bhwr10DtXHF9P0IBBHxvnaVF5q+14PdZviPIcQBnGoacw++XDFbX52iws3i1zis
Br+vd6OFQ9RLCwqCpdoY1GDHP6nKz7Tm/x+5AQNHsDZhAo+/VdIxLShkz0xcNE9d
Ipe7JUG4YRWLzVEKTu4dkXHB0pONwYMkchot2k+167TaSulVfFlOCkRjtqOa0j/z
Vo4/DFg6f3Looi6tvB/HYvwx+uWKUPEZxU39w2ODZGcdKbAW2UVFMwEVcW93tRiE
E1KhxGULOFLcJSH14cfEP7d0dvsW8gDcLHh5uFaNf4RS4EpL1SdxnmM2ozrp48hE
s9x1BtNTA5qNCrj86O36T/T9ymyNqRgUXWmy+UbBKch0IirmSRVadlio/PlvDzSM
ZKQ38xD26fuQFfNG4tb+fv0qPzu7qviz6ImpqRzdl/O1KEatd5AO/mTT64/r5DuI
Waf4dp5TScrQE063Tq5swFoJhQlmg2lco9V+zX5+kwNZAJTzPEkjuinEoQtSenUF
XCC9shR7W6eOzyXcQwk23dDfldHuXfRSwhGdZGy/rAEoRRqPwFud2Eh8fEDzE7fy
10uO0dU3/ASkNKSYBft2JW1Qn/OAMi8QK8RMGfTVtp5+0E+NFyz4iD0RcEV19hvB
+DPOb78NXnIA6aIoJJKXnzgBkr3Rorg7rCtZyG4XmC3byd8nBH8znecYdMRCcvgO
Rcy7jdoldd6Gs3YZvIEGxqKzGEFbIaQWUeishoVHK8dwuk6jmx6bHCa2BB7iqSSO
x0vyEUKlBAVHZCg/A4w5QR4R4HQUvVkYtQHz10649s42xAt5rqjnX4LH/kHAY7YY
M/o+My1ozvU78AhJSAtRM/GbrF5UHqA1hBSSZV7+rVGYRmTLk3PcFeheokoHelQl
6DPpMh2arMnfoVp80f0+Q7V3fP31aGnozAcI+SrFiWRDjf8FfE2xLvres4moOZ2Y
O7TR9ng93NE+eSE5zoSgEfpIG43+8KwUakdLN2en7Fw8wl71t3o2wr+m+OAXew4Z
lXZbaHmaELsGJcWQbsrRmMpnMjPZ8go03ZAmO60wPo2cOnyAl6iaHM2G0bu+CjJ8
oEyl/viR5oxbtkrSp/42xg7dAI6bVgWOZNHup6FQuMF4vdtptJB5oUiPkCFtUoz9
QNCNK1+TWgD/JomgnZekONTDFE0RUZtvvQWV+mCjy2pZW3e4F0hc7ncoQ0JwGL02
88gpt7CvxWGNC3p2sp7+tG0nMW8Kas2JEgBBHytpUo/dBjaqiK+ZFFVXljMAYODx
7Uqov2Gqnt1GbNQaUkO94ayWF3zWu1B5y/H7mQOXAo5TLuUy4Hk03Zk+wVWxa0zl
idS46jWeTK9qDxCxCQY8fuJOOIgFLPChmsLrQJaINC5dFvSfSifcYZSdp8lIawCk
q4Iyja3NHbuGGx4OgGmyXQAHXCy9kEZ62VXplx/K/EdeCVxEfNkq5NqQYLvWwjCm
AcNwEbcOoZebE112PuVmKCB/AKd8sD7ibwVjifIAIi9OKoZU+JYcX8hC5BE9iDQc
sBarli6ELyJhYK5wH67L8fnUv3xY6bK/XHIWmMrTCfTT19mmWkHe0T4FkTf2JmWE
3dywsq6lfcTrABTsQpmHSbcT9/HwyPjBj5NLKkOv3dm0/lDuMXyyj0i7WZdHOyQG
IOK+FXtxakth2FYl6IR24C7T7f5A6IIp2R2okco8ifYEXX0Hj5GOwe7J8ZM5GhSZ
WTi533KYscW8zLJM5DYqQhlD/k4x2Ff/9jUENUfYAhWHzExEuKmhrmaba0KBqd86
/duWi7ZmSOrpdFfj2JA57c6vlR7f/pcdoP/5FZWuSl4rYIfZz+/DO6D2CSSlT6kH
+tKvb2vCgsvrm122qB8SkIsh3JudMDqDP946AX0N/RWvPm/qDvrfBB+mtnnzO1Mc
WWGJ8fqJjDxTVkCA0kbLpBhYkhwzOxBZAY/S/1BslgbduAHZ0aDXMw7NHVU6Plx3
fIITObBI0qOI566YtXB2GmAyjFpbH8ZsFG7Fhm1H2HBbctnSGm2NGH5uR84blbs0
/GXPDA9krlJI1A9Bx47si0gwJFnnu1N0L3VioLS0EDL10TX3UWBXgGynfvxFc9KL
P6ZddSqgGD7TBaMEphbVPrBTvNEL/J2LkRW894qmNz6OYvHkwLOxcjf/AH+05M2Y
X/LYdKxagcJncEGQiC4zEDoMICpYVMq8iyL2Y7q7wg7rC/5HpTnUkgc+yl8CdqSH
hBfgTpug6G0vfRCFznvxKyx/8awOiCfLw1pKDy6sqVz54hnX8232vs7bjMLORMSy
s1VALalcldWHjRpE17REA+wpMngvZ1klrluAZ1MOTI7k3/Xp6WmhGThxZvnz51Ml
ZZS+TDGh2R68ePmp7VMRpLjZzIM4+ZR99lNjRQ5jIza3i26J9IeIcNz7buzquK5O
5KrCFIWqVtpmdLqfINH4l8lmfys3TGlhNSxdnA3wMwjfE5L+ickKEdu7A8anpRVF
a2H4OQYSFZGfepPTeztthfSXuD0SkIQDo9CVkIfcopGe18/yLFEkoTI53rEfOR3Z
KBymmlloOsspVvMvI9xkiLkiBq+v31nEB46H4xP6DaO13EKG0P8vB3BGKSzMMZjJ
Uw9LwPn74niaqLb9fCEr/siMW5gro+Z/MEJ+W74azphO7M9AXTkpkmXfJWPT4w0o
Gj3dutya7YUXiel7SXio9Es5vIfET+NYEgn1QCMHzTxvjNQlECIos9K8dATG9Is0
1B9GoFqZA3BWjfqUubueknr7oop0RAJ2DpAfy4+b7XRNfQnz7XXD0MmH6WIbIwwh
bOemGcWd9Phk4eC/W67IRC4uvsxOfnNIFdTdy+UW5aC6R6YZhwTuXztN1hmdIqvV
AXkzPRQCk7raXK/iqntOni/xoWlLYcq9d4hAFX/RG0JiKOyYfFqwBKICVsRZT/wK
iHs1SEYFjWv0g+9ne21jjxJjcOLV34Msa7xgOUUYMEmQAqnSRdEo/57mOOUz/pGd
JiCkkwDoLCXclvN42ygb+oHy956DFYp6WNG9CyWIs8JoiopppMzfbAo3Hq4dPEhP
rk4oT+R4tSLGQtGHU96HUNvCMbflqImzOeIB+ZGEX5G0tgooa8l1nJ059mHyCCbS
fUZBsoqX3Ccabz5ZUtIbv4YxnWkVqwKSC0kiExebnm0n3v8vf312INIYoiN6BZJH
+hnB7X5xEjJVwBvbBzAKhFjYnb99BWEVjCrHT61c0A3lWytWztMEpD9aRoVsOTbY
Eg6+Epb0YM0l/39U4VuZs+4Bnn5AnbQD5yfBBFvvjMvqJbO8cQyP72Qchi4ZN2Dj
U2/hFPjVQ5ycjBOiqDloDAv4VgB3idKEcgLssoaAmJAsFb8R+jjqyWXyH3rx3DCj
zoxSn0pSH7kdvRCtQBiZ1aGppC8bMJRwJJx6AY3G1f78bKMKaJP5mR5FhdcJX5Vm
mVMXCvmLgnf+hfpq6rzTrdsWHapC/x+pu0Wr7gcXybZ7EpAKsUvOAhrPImI0/BsJ
4rFmKWz+gNTvxMTso+L0veLXU9qMWjZn1rqZMbSzmZnqvQRt9OjfPHp0HoNpG1Ce
qAi08Tpe6nG5Obzjq6XFi8gUbp2GrxxUeyszwVbkz5DRKQYeN/0uhbpttZKV5vGm
zUfRqJePwwB5MZbbE1QsdplmtsTw7hjkzJcpUE2q/To6mj6wF+I8L5oLK3EWR0AS
e96yZ2975xCaywVIF0r21t1qMJSm2Yr/AcWHzsedpA+zymBqePZGK7CXXyZwe4NB
xvV6mvP2uvVIvBo3JV0jBMvjHtlAxHJL1VTypybJhJ32tA67pBoeXriUWb7kTSGI
0smfQHUW98g32K9kJ4fqF1ovk8O6VQYk6aPV/bkqqPPh0pzGo6DSLRg0xt6O3tWs
7f088HoIzrInswOJxfAFTj1xipQGDSQ3vzL5fMyQfFG8i4eeMwXlHKUOPp28j5qT
YpMKeNq1q5uUrQvLaH2F4a29vMsECk8hkXRCOPLa4lHf8dBxoo5U4J1DdpNtcLxm
BYSk32wRwQtN0wxhDZ6KOV1LNMLQ6UDt5HuPboaHVd9evLiaVwjyU8amOpYluBbH
nZdO6sh4WBKkstjUu+BrzwTZ9pI6sa12rJ6N6QFzxoOx4HQEgpffpY+jf8MCu32x
VgFSEAVv3bmidWLcNsTrq9LmknwKU30pR9L9zXtWTsUUzix57nmdMI1rZBEpAF5R
/oGQnAwhYiWpLRDtWRZHF8LEeGR1473WzAM/jXabhAaZ+CusZUpMzLU4eHonjoOG
jwZXMvv0oJCzDvkDoDQCu8BE6wUcOj3ZRAV3Ss8iyOdtifwfC4Foe3x9lfGcVfoy
EXCZd9033PFFa/roDcMDDqnRbG0QCpPDxaikVtcLWZo+7FwKunR/3bSVwbafQEH/
O0140AQLlzYdzvtORxJCF0C2KkcX7PL/plOQqsIBfiSMLOfJx7+Hlb/uWK3YRjEI
3n8g761DaBYMdapCpR14er9MnTswp4Uq5+YEvBtFUoVpQRd8c1jHIUsjfvxLfgeL
oA4YtIPjtS25IidrWP7CagLH54ZkQsjTMmrYoE+WACJ48haejmtCv/umjXqrgO+Y
CpT70Ke2fhX84OnmMCRDGkJ9chH5EB5KyJOuJ7aLvb1X50/DCwve16kk8ob9MJHJ
oEsJMb6vRTf3aPqnCKxx7QWg3yJr4Vdvcd2AZBINY43lhRb2MJk5ZRSjzFsm4xZT
0d+1JsCElJ7z47RjXafuDHeSDSz99OJEj94a1Jk+DuUm3uhZ9w/JVhSe0aCUywok
d+YCMqnlGtZiYEXbR/O5QMXw4QGCDi39Xs8XAqHSvN5G3Gz0L7tjv36oV5QvxzSw
J5nNhizGmkghWJGRPR7Cf8h5slciLX+WKVgCoDQouoaF4Og3yoH6eV/BEvmnix+g
E3wacBDOEQjcdMH026yRBaCdKRRw94BVHeqtJ2S5Rco6+KTq8lbl4Eq6ukqdST2a
TCdSo0X2SLb7rEB5UAq+b/VO1nYRZWMQca7slx7tVNmZz3AHCm87lWiWGq4hRWIM
1sW/JXww1bObfngAf+PeHzrxgM42CQoGKtFLcANaXHjsJvJIHWTngOZqbnDqV7tI
Su0dgTkmUvPZ7+ZKIIbU9aefqXO/LHJN197WcJ0ezC81EJGbal9GIDK57utx4mCW
T2cujZwK0QQjdxMHpGFtF5yEJFjXiT0rAxZGfGfI+sXeSnGcMllCa9tLnQRgs0jv
XxiKVGXTF6m9FHsEZFCPdVnK9mKq58ppFyrRXUDANxbKwQgk7VQholpjgoRhvXsK
wMjGk64vxgJnDELUcWXzb/Xm3t2f49Famg1QYyxcctBA5CybvcTjIDwd0kXamN6P
2eRnulUG7dEVX1rpPxEb4D2619AnoDDe99bxukkPguG6QfbNNyx11ZPUb1Kfgm5C
Pj/QVlokoOWPAn+AOtkLd5BPKkYBuOWvIARfrnXmX7LCX0gsCO2CTGOGIFHjynI3
sNCJq5ops5jizZfjDDXCBNxq2BFh2Apbiyow03+5MROBD6sJDeomQRZqwz/1sqQv
gjEeETkwRMcaQiquom9OgyOWXc5gPTU3mdoUK4sTU6+67N1Nl/XBcRcIolad9H7u
yyLF6Ga9igL0wHXmEE1RaOTvJj7PX7/e/BIsPvjBdIw+LmBdC1kxJbTKLa9INwrS
ERP8nMo0MiQxl3/t4v1o0DETAoDY/7sh0ZMxt4+ddh0dahemVXc9opLWdZX/cpOY
uzUC9eEB7u02qxOTELobCQmaHCLEkXzZywHAyWTEFBvx2OqHXtIwC+mg/M2x/Qcq
y9bsvuuSTE0+4m9iitYtBHg8USxoONzBNyoM+B4gZBIT6qMWzRnwlDnP9cyQdWEi
4yvVaJFCTsJsJeVYEnTqJ0uxcJ7RKMnlboWtK8ZtwO357I2MxB7wNqLRG8UKT0HJ
aOHONtiWVWT6prPzCzDvJXbe00apvG4daYFPF3EU/EB9wdyC7BePJjBLZYedE1o7
mpYZFTZ3e4zgFj/Ra4X/oAsBNIqsjs8vZ6Knjr5R3rr1w99ccRVzkpMjxlzj2NDB
iAG+NPMjAr0CzUatw26EV17/zGEdoPUeO2P6tvIte6c03BA0x85qRkt288a5WVTa
ekpYZCucCsBE7NTMnp8459tbJOiqSTKKNlkqXfrO8o/d9y1dIo9WMbDtRRwk2ZF6
n28eQF+tKK56eZ8I++PqVNkWSdLIdAceDIlO4pOql43uWZWqPcGOBpcgkTyp2l5A
u30eeFqntE56KRAVhOyBNRChMmipEbIUwoE/3rBwPBBNpbwClcYkfDpdnx8SzhTc
sGlaAo9AKB5M5IK+qBSPijYLn76SYmUB9Pq2QHo/A8bvt6B0vbMDKzpJYsRdu7o0
FSJ6qWjRHB1rv8pYiU7oDJ2Yy6PirWiC6PSlmOLeszXSQG7FEgk1j95+2XjFGSCB
uPQY2C+2RPgljAA6WHfGCy3b5aCHmwI5mVEH8xuc73HvIJCGNKNKicu8o6OKPgVy
/ysIIkbdbb/3hbODaqMtvZK/xCD+Xd+VGeZJSiW0MT1bAnlejgneyyvpzXnVzloq
lqlgFJHjNjj3gQi5M1HDfciz3AjTGfluiDCqtwN/OUYRkylpEdMFJr2tXAjeLeUJ
cpAQ74GK/rS9QOyrBv+S4Ui4SfTfSNor2urP4JjPghkJbVCT21CEciOe9LZJMzn/
K1TL1pUJRY41ewamjxPo79TedHAKWzt35mLFZlAfbDeHtLPY20cgg8COYLW6KFv4
FeB9GWJcENfvSMJOjiE438cSCfuHsmm2OEd+PJwqCo1EV6HB0vO91mUcpCQYVjn6
UbRUkFRdBLbqeWenY7pm9FaRTsy74ysyaUArw7ryhONBe4yfurA2lUM1XLtC0JdW
SJ5OmtkCnMFqV5FcpujtwApcbFNonZtygCKNTkfdn4l+kGEEhH/2ruWSLFnm66qo
PgL5Ym5p1vyCx3WCJ9jjnlHglEiMiuqmtU19xoblf+uX9q3tsLPqFjqJjxJcHwM7
9WnS2S2ca6Y878JVu0PUdXzevcXWwmbD33U8bbzYkRd9pqawUQZsUD3e3V0F6SwJ
SGu/CxzScYOFN301Irg9nkO62jfD+8vXasEP37m2bjmpq+k6XhN9NRmOgRRuIVK2
FPWMsiOQdjT9gMEtv5pZAfPHgKF9BH6+ji7KPy/Il57GKYrUVO6GtKb8TWpDFwOU
oDR7P4pEzIeQTzqrZEEOA0UY3/5doSNHiAwkDHwad1zydtCxWQzZQqdC0SLF5MSy
w5800MTJA5OOJAJuVWd8CX6WLbyKUhcrV4mrS7k6DIgF9N5Nh0arugViEddO11Pj
Zwn1zJt169jbHer9M6RAWk/OuTULNwaxu5nO5o1wpCzbcnwsTk5J3fxH0DovXIUf
zI6C5fFuOzCRqbtbFNeVxVUOHWWZWKkWdMeOntPqnFTYZG5DHJaIff/qEwHmymPn
qILooz+YiIJGn/Smc9yxf9WuXJ+O9wuLBGPu64WYsLGkMRDcAXOFuL8LojEMqOAf
WEkmVtRWTPrwGUHfKSnZ+oDKNAXUW+Yz/zmd+RgP/oq9d7MYjJmWWjy9Uak2+rhy
aK+ANIFOqqCILFmiGdui9T4G3uAIHNbNoLs+7vupdQY4BwJ8pttJcxKiXnroz4V5
xAo648VyF+zmlFCEKGpx5tZioZV/piuDkSbx0NQt70SfGWYA1mEzveCld7wWzRG8
lqMDml9ahu2lUHLc90rKwljBKR8/o85i2S8SzuKWbKi/9aQs42MkghjKkApsHsuc
YYwZfcXU4OHaZMMh7hFGB0r+2RTSl/HUEK46/sGDRtozDk7iMbFEN1m6+WtNCnQm
9HNxcglp/8UPTmFif2ICYYgEirVAiIUtC+h742Ha6Ch02kyDpr5oRAYXC1+h5ZWT
5CmovfTZZGX7MiYN7PrSc3ooMhq+M/5fKgOU9EAcdMskuN52toFpk9eI70NTvYTW
p93oSVyyxXEvCgaL9vw85rFOReL0mwpEm2R3EBxErQ7QOCEnenGSVbyl8Ns3an2k
cvBWpjei+P/+Pnd/743dME0G7B+18BaEpSYmS0Hsw0ULURXui4UOFmNXwLwElZjk
JbKHwgIZAmWsl6Vogx1yRBs3m6Ke//mEzYg8bQpAKMy9de5Ab/LzurEUVSq3HKeA
dqXPc0X72d6zJ6RXomyqJTdSBIcT7w5ypJUjRYdTvLbg8sBNaw+6+FE6oOLe4QA1
8u8g0RH6yc3zPlopecLT60h045mecXwfhstDkT+PCupURYT5rLw71CFv2cUwXwoZ
PRiXLE7pfd9lNm6nVj6jijV6IguiPgj0/nixnBg9M/4T9KwNU8gc20WO9bPgzh1O
E8EPn3qp9SllrkL5A9HgfUA0MhpHtG1xT5rxdVhhKIBTZHTy5UtpEfflGn37d3E8
CiIsG+7cO+ZXzvQ5dCyFJp2k35YXCI/ZZo/Is4MbGGvoDWPVY8IhsVogagQqkuN9
E/oxRVs+6g3LEpBA4jgHZCbgAuRtOmVjGKL6FsLSKD7bNkz9IySpPmGYx68F4t28
x43jQxMxpYgLwziBnl8IUAuZjM1vc/DDQKbyhjyZ8p8nsEW2XDUj4nzqDhG813BD
d+zXK0jBS69oohGFtTNFw5iaRY/vEABcwZtlK2ixaSu/BMtGRj+TUb2abD+1IKyA
ep+OfL/cXgTDav7EauMIeOb238wwuEZXKZxBioe1WXTkvyCA2K/iqKaqiSkXtg61
KMF2clZuDjQBJ3/bckDO+oBTB0vgVGh2uuffpKpn7aHUcCFKlIz40M/VTHA5uFmZ
wpx2jhvyNwZhQWNPADmi6UMaVQ5cjoVOy174qqRonB4N27Mxc1ZmSCZuB/hJhrKM
3nXFF2WbOjmOv2AZo+VnoaZnQ8NniQ149U3vGfVMyWEKIIBgeDxOTGNszEvdEDRO
qiYRI4sd+PPE/FdcD2sDZxLVt/Z8UwsYlj9GTy0+QHC23VyNmemu/aDJonPgImjD
mUCbQChqGilVwhnULXb1+30C2Cf2e2t+ULIaaogSws5s52zfvThykR1RSORBfaL0
cSxqWi56B6pmhYgQIUPAM9HwpuPRQZBr1ZR8qHyCgA9+Zi+g4fvkcM+d+fbGzCZN
1qjTFu4Z/yXS83C/bpMzzz24dLOzgeeHQXeDInt0Wz8EJznNaIsNR9Q1xlb50GXp
hIfnAcdJx+56H4Alm4rEAtcViFxDB7dnXMhRfHU0mLRfYYQOzV7Po2HWTsJooGun
Ctlu+QCqYIGdpCEgISPIcjkd8jtKkpi/koGftgHMCEqDfSqjblVJTOmmzheE1LEz
06SLP/Beg1qpdEvXt+Vdl3bY45px9vR3A2cbK3XOHfPZZg0rTGnamski8Vvd55S3
oX5fikIkRZEkc4etECZF6rmnXJpRas/xFU7Y+nwDMncw+JT+Tq9nl3RwBV6s+W1D
BMnNp4O7XsYPfyYjLIV4lE39T6/FBgOM9J5w5+qOF0m6OsrJH73HcbykFINSU0q8
H2HNf5ohkkib5jCi3GHT7aAwvxbcj2tsC9bZTen7NrUf3v2xNvBw2FwQ9zQx+/pK
ZIrYMYZLWOEB5g5ZgNmeGYFc/b+/e5JrzGXvizhLm9ySXe5yVK/1vxldGVwSSwNe
Keze193yGKw80S9+srW7cx+YbFWeL1ZcNAO7hZw2LwDOdT7lKXEUNjde1t51pVJO
OizOt5cNr9ympnyqCbdqTzfbX0wUyYmfJ6byDCyagVmAV8KAzP2mHMebEW2Gv+fy
Px3clF4cj2MXGz+4AJkOEIsS5lCqNNuAs902XA/uKxP3wcdVv/UTsQ6ORSwIh7si
xhAeR82mtnE9oJwn4XedthrvmntYwcng3Cwkh0hn+ncMa9eJCtgezLG7Mohv+vXh
NVbUYHr14kBmDEjxmEVd35tBVhyl5BIJKCTdOTxRHwYksFXJ/Toa4MjVA/K6/MA2
bOqi7V6JVPIcdLKshezc8ls1P55ydSHkEgtJX+xiPvHk45G63dfgedteQISFlXBs
suz5Wd7/z5QgoT9WRos1Cd7k8rAjMRhIOqtcGCUFi6pVI8CY5P4ZRe9nbcBad1h1
Pa7DdQDEKrrMMAum8ME96+QVa60jPQHJyvPepwVuVSFUhcn8I686PWykKvLGecxe
ssVNpJqdRDimgoDdrQ6Adr5J0R5dG8/JqXQ+hKCDVRKayXZbvwYtnwwU14jAkdLZ
QmFIlI4o1uwwUvr8voV4qah0hD6+7O9XuNswrPkCfIvFWZyO7608TuIs0Rja4Anf
PtuK0QKQ1HD62WSQfsKoEvpnjvYbYF57Pp8Absb64NUeaBouUqr4TzGFPbtOIpUS
zNS6gbGFQ8O5Vh5PhY0ApTZUA60MD4z5qzseFYqdL+7NfhxqRLK9APgdcs8NWwbr
BNVaF/R3Qv/YeTehs10YjhH9Rvj4dsERiHY7SX+rkmnZLJpy9HcLjCPlBg5ajgFO
D5B09RN7dU/1tICHPv+7oxhfa+kodZKfn2Kv9CGfM+uy6YDd3iHxOUKi1TjKNstP
qJ0wMPIZdUSoImr2vwfyIdlm3pYaOfw//ExOns2dHXFvW25pcjgXrOeL4LmfdnWX
Jaq2cGPv3qU1BeT26Mkxs890iLHhPm7PCpaUmhd6CyRHUp589U48Pz/vuMSfxCvN
kQZ2jz5wFXQ5hmaegiUZZ6xfWmVc4hCEwCxTZJA50uNwUVjySVT5N1zpqG5Vl2QY
/MGY5qF3ywQhOhXfEOtm6F4Vvxc/Hy6+Ce+Y6vOEV44ALFkO6BgkYSiVQMdnZ20x
hQ6BCRJ7eivs305+OfHxK7qR9mZSdzB7QjDJZtB8zj1rkkRihmJS/K0/RmJd9UHf
tHvdzlv7ax18BbkIMwKYEOhuVbxDmkgztxhy67Lpapgla6d7tc83Y+G6qdxzjYhe
xXnEW8GgjZWzBL3KsUckOvV0RA2MKfSYRHkJA1br+IBpGSZ17G0nLhvt5fyjmRV+
PF5xo1RMQV9HrW89QSJThGZ7oqyQJXN1JCPfRxiL1usD7DFI8FZiz8YGm7tIVh7S
HdGmC22IpvZeUvyhp84ZVkUCvf69EjgwkUGEhKbYqLndUj3dZ37abz77Juv6sgwT
ir4ZWor0BwLnsvcsWzAvxl4BapQ69BLkQT1zGPaQPhJDRNJzT990Dlyd/bDpGxCq
2vdNvYuF6VVXnN8CSwoDCkwewrW6IghkjkXKxn3QlZ2GVPhofBWS+QZtELN59HJ9
bt5mdm/QjYUuUyi41xMRofRD1ltJUPi9YHu3BMuiychXTehbLqTgC0YzeTlVdJw4
PJlvOpf9zwNdiSUEVH4Orr7p80n+GyiiNgXcJCKpW04hYBCRaKlquMzgvqRrEr1b
EpSyAO6iqWVPfYLBTH96m2UTi8gu2XvERojIoVPj/WuQOWFXUtxXLQWk3dVgZHy2
08Q+grpsPniYcUmB+wtlJhnUOpsbW8tWyfKRKbD3nWTzvE9tULsfvHsWz5MlY1gt
/thlYlTa+nOL8bTN7jLOgF0trziagMnTQBmh+yhv56ALesE1Ww3KI+KcDC8wYOsU
hmq4L9lzhNZg3c9x5miopQljbCkGcBPlwRI62Xdc5XBR96zgixA0CyO8pHE0wbDz
17vSlYGlclFK4Zr7RziTzFUkWfIvRlzRsIFJFIZpnBlRvuc3zzX9gPJRuK5k6Vbc
U37SdXXc0zPEAx1r/GEj5EFU0i1OXe6+to1A9lfoiQ81tauCC8Qf/1tbXLeS9cGL
fW/ZgCEiMhjCG7v9plOoGOS3l7K1sxDjodg9iwXjSomrVROZV7lQu8KgqBEBGLHm
nlLyTgqsSG1yqNDVkvf1H+/jz+SksxVdGlEF2nh9zWvIoLkQPnPVELjmCbtDFiDw
160YQDMu9oVH40Q69OKkVCZWohN4opADXjjBS/HoN9dpXmH087NBVZzYBrpVNVdy
TgLP65dSwUNXdEfH7gqkygQwR50SH6xDm3FTkqmMfd3pCbggG6H1VayJr2KepDIe
qsb2t6PnuiWegex+Mu9pGPJHIUO40fifYmxG0FqTYApzPZXerukInW/6664Rkl6a
wU9trWR3hjiQJ2D9B6FYNePeEdEOX3SDGSZEJFyphiYVmbv6hUfE960bQlVBEYFi
Fem5CATn1vfwg1uleoTn0cby+lw+ReY2q/KSOGHm7TYllo4ftY47RPhkx/nihnNX
ewjNQOZ2ZD6oGeF1rPEJ47/iVdCM/+LP0yZ7cck6bC6uVinr8IMVNT8c/cYDRdNY
/90FDuR+iH/12mwjt4HZmQmETxO49dtlowFirI21nFiq2A4IsbJ7+sOdR8Ovw9Oz
QrUdQ4PWSZdgUOV5+MKrJOgtjvdlD57jF8Pa/jptfdWeMKiEjqIEf9jfdEdXbhAR
UJdrPB1p4Dle3SyrvQXKd513BFD6E93fPAyLqOQczsHpW28QDm9OKCmBnEZbScIB
vwyyWJ7g+XkjRa7laC07HWVtxEw27VDJy/PyujPqZ9zxYJsEwaJCoGCnmxbRHveD
188YJwui6PGsZP8PEiT5FcIfP2LRbSrHFHCddIxDduJB3MD8xs7LpT+8T4VKatd/
KTvaS2mX0E5rEdBN3gHRq8w8pOwbv84U/Fubkdd5vK05Ghxc8Fj8CyhHpcdeEKXG
H6MuxOF5FSwg1fmDM43rE43dQpqvkxx6/iB/ev3w18pVqjVdMMHWW3xfWD430Rx6
v1UU3myewkg//xQG8usLmFrMApm02i/6o26+UrUOK/pbOpah+dnOuDZMzpcT4lkg
pDgJ3cTDPQdAZVlItUMe3ocBG8N0VqWSf5crXqWLwmJcw0WX4B+aPmqDs7UX4vWw
s2+w4u5gLQ1+ges9attHDny636ohaxX//FgbD4Cw/LF7gc3wd8OQjwx7tajQ6nBD
XIC/s8f2nNsDegKTM6GU9YL8QMkgoP6GP9wCoZbmyOJjt7BwQ3WfzpgNxDtPpK0Q
a8bajfqLaEvxm8DNIi4AUxwr75WWOVtGPx70jc4Cm2xt0L8vqBCAWKRHGxpeLYMF
4G3oQI+qwQTyvkYkM/4iIHx1/gK+BbDuTwcEp7wGiIPvXAnqJ/U2W6bnc2E2UUn1
hYUXS3cUtnDPou2qLkMwXdHcrsxLOnfhrU/PFLF4/KxQHJXc8tbkEri35hqJ/2yr
shUwjBlK7C4TNQaVMha8gMYIrpQIpPGZGlyKGsFJpLPN3WJHe1YkHDtuOlqEK6Hx
N1F6KrYy8MbytsF9TMnhGHw2JCIIvkTm/03R5E0XmOPVZjG6B14bx6/FAZGXrQDN
xNPZqccBIeVmvZl3unJPbFtXBNcHFroee6YYQcCpDU59P3w5AfGqbV8Zn9Y7l29H
uBsY8EpVMo14VrsxSzhTLUVvnr69qaGUE/5EE15gG/zBTswAEWbJH1A2fGjMGyot
sYIpfms9lAin0BSsGISaKDAh3ZzMjZa1AGokG2w4wES6Wbylyu1v18eUW6bH4cuO
//syrCkdp7rrxGG8Cnrm2HGdgwZEPxlu8Ib9i++gXsEe+D1BEr4RSjLAcVCTj5Cp
LhgsVR5FuRIOoUmFwjgmhRtROH16I+Qnodho3p99s9G5gerkcZZAuD5TF1cyfHl+
6Gx1BN481PpbB+fTXQlz2Ny2W6bso3DJx5MQCf5loRw87BqcPb4sPVRGe/aHmLhM
VPvp1XahbLb0ikSKoZ2kpB9QVjFKSGCBXZvEJvLoDXT/oRqmQa7u6yCDR+oPn5qR
VXqvI3oVnvt8e2/DT7Tils01alqlmWt2TCoS65OmXEabDreaMQJNwHRLpZDcwYrf
b/IzfwPbhMC6xkErMC8KlXrMQWnIyWDgjQ8QXsktt2ndCBMm3BvGegjLyqucASe9
orK5MNVSlJqWHo5zVg2uZpcYWyd0yv0OCN8E3E/k00Y3f44xUyZC3NUsJ8e6Oftp
tL2cJrArGt0AMEPgtqmNLo7kI4yVj3MCUP/J1OjiS3qFmxvfAxUEoaEtsYuvkmCr
HSP5YX5cA2GhudsGqt4Qw0wM33ltkgQLlAsB75Wl7enjYwt+KZOTyE96lsAOQzdc
ej6d2biJXH7gUL4BK9nE/D7nCCUiBQCvkc+w92lPX/WIuQwMRa8Ce+NbLXhe0H2b
dsVO1ee3puGsNoy51x/OjJshnWxS+3d5JwNxugbXNzVCVtOBK9xLUFPNTkY4R2tC
rUqtZxxpM0jLfyGeBlWT3Lb2lZXD2LcCzQ8AcrGAK4rQndl2O/XvfYpThQPtin/n
2CC1fqnn+FgyFF/aND1Rc5+SFdWWG4vWjaFoTvGM6M7KaKKcEX1zcDV7D4rF30DA
iP8Nt30UL/z2F0aEdgZJF0avGCW5fJcaFOLcV8346j81AZgMMavVaFvva7wC/hiB
hIHS111PWOyHfc8+zJTp1ZeJCSLxladN/dddmnFB2cYHO5CUrfQMwWOHLJ+C06By
p1g3XWOsfs+isJjj2+JkIboPcaBAb1r0LSt3zl9B+hnmi84P33w0YO/m6UlzFF8J
jEdbKoUTtjsb2GNWFzKLU2vWJ2/VizvzXjitEUa3FKk33d8Gnig06IKPOYDaP/fY
MLbYTZVhRclyYICH+fvvtNfrTgvdlGLJ3MYnCSUtrVQZMd7iK7ouPhdizhji1phT
4eGKy+wSbPyPvu7Mg5cZMwlrp2dBLVE6BIlcEJc97V/388YHcuKrpYZ9AnNO/7j6
ENyUiAp82Svoele5jyN1+AS7fBd5PzNseImuOIQN0xJ/5bx3OsZH8enWmyIN8ars
tM+hyqv7ZVtg0lDiyjekaeBYnAtqk5nGe0O8lSx1kl4/aAKicbFtnZRD+DYc6LRi
+/VwQvZ7FwYA+6Scsudqyox9FTrYCdZt2wrpVAxmSGA30OwHS9e33+l1927tNaCj
nQKKEEzsPcmsn1qLlVblU9FUFFe5Sz8Kv20fxgQ4henN53juhvsNJVEqAl0M2eEf
bjUt/XQppKwku/RpEUHgGIcV6mYAZnsRKTWc3EDZuiveRo1GZscEKVHAOofgbU8F
M/eaobSTdvwrX1EZEjsyl19ah9G7tI/HSQBZWKLK3M7lesdc7n99cuhf7kLa8UvQ
9aZmJrD7fksjGnlwwt4r1kikFaOFCeCAxSacHu+lTrUVUTnm4ZFIoS94NVoD8RRw
BdDcjJxqldgkzxmg3XExGJ6AAIl4IC3oYcUb0Q/D96GwYjTrDns0qq4ukL6bg14k
WzppzMA1+w7I/YGAJlxk7auSASBgFomo65XFNwokIiCU0mjC6HWKXYYIqnguImSX
tcTWZn3uccmXeBICuBJgff/uAkM4A1jbRhlX4l0uhiDtw5AU0gGGiuNN1dtJgN0Y
Es9yDo/ouXtcACieA0D+H3vB5D0+IXqzL4LZdT4evrJvtpMrJfBDJF5iqmUy4CIx
QDg12B4fn9UH/K5CthojFkz5EGCwXMPFrtFLsQj01NnvAozMmQQcjGVEq4yoEIpc
BhzR/0Sa9vFuCEbYmG350fInC7va1w3qYOUjxe3P4TO5IZ4ZTDtKUDE2zKPnfv48
uvoZvGekdYwGTTpzlcZtgMFW2FxMd2b7gWDu0L9TpnLZlQPb83uxMjXVbmmKlyya
irpqfYdoeWQgYDm8GMfKwmnxtpip9YIR2updS9ooKKHGVw6QuNZEtLpjhs30t5DW
PvI6tlscFVJ7hb241GVJ+taooIJERxOeIXRf9j2OXhXmgBX2ZjxGPfKQigUojwGA
G2oLLKHThptpd9Yjf819Z4sd+vGleh9DepmkX3o7XH/U+Rg6Cr232NikosJ2/+Hb
cchKokBdRAt3KGAtoF7XfAf/pgEOJB1cO2O7a6s77xTiidVXPBVNqS3ui2Gpd2NN
RPS71LbBlCpcM3r55RlN87YyCoCQJwoCOYbrj/vAYq5BP0vQunRv2zmGwO65JDoi
95yO2ZfxrNCg54dQbjgVk2Pzp5mMnPzyp/jFZjhLH1sXkvna/q0/nor6+oMhhKpw
3fRRtfKVLtZU1fWJroKX/Qm1wO5PTw/zFPltZF3BbypLl6jPeYuKvk13gSnB2+g1
VD9GTPdk/Z4S4xPyvfFFB4eXeG5CzzkYTEksUFtYAdYYnOXrccKmqOCwUBgWrueG
qx3roDK/uxK927AncWTfzOlbHqLLDBF/A6eJFxFA7FF/oQnyLAz8hJ0eW2hI4u4y
kwjmVqE96/7NcucGnkLZ9/2ML40zk074wR/LV5AH/w9A7iLtu9MsyBEZs17uL8zQ
GbDRc0JOVEqUXDUQNITFiXp/D93HBYX2WZqRP411+2gsaqlqBYI+3g/gk8xpUI07
qtU1tWQ7NYHdmOjYp397VR80/ZRQEW92L9ILqnmAFlZFBure5NniGtt+cpfvpV+c
DQmMquqG5D+YwrlzbU1hdc+fcI4GF5EUbhSfMR4G/Uhwghxj0yQ0CywPNbqhbw6+
1YZUUsWfE5ISGAQzIs2hbPjkYSGWEQjbj2vFmgqD0L53YfhtuIWmOch2jK+/4Yu8
+5elgntTDjo2k9DSI3MGMP9m4s5+nUjA3fjbBMIgROpVnqkGZPLMT4t7wpP0NSdH
D3J1Bb+ug8O6rWpqR8m8HByIaRTW5pLKAb9Xpqvxk7m3xnzLMw4g3WzZuUaFxVJJ
5fciGFEezqOAEo6nBfsNCz/J45i4i3V5ZM1QzO7T+qbTc3VyFXmJ1rWYFp6b8hZH
FLtg5x7922dCh1iBEMJAymvhyWnCRgbs96EcA4lEFUJwLoHCvflhU4Q9W9ArAo9l
eISyazdcj2jhlwQokcnSOl4D/D125qNFyLRHzCrFtMrb5BqwruqGLNTSxcDprqcG
feLtC24+GstRoY53VrWI1grOwPhkPHving8Q/MON53yk2MwMJDHMr5su2Ep/0v75
lN1F0JrmRyRRcZn8/NKlghQzro4l11FZBnjKxcOTaVH0B3qLlIQhd87EyKZS2hH/
Ce8ku2kRPu2b+HZzPNoTzFGh5BgBeZTKASdaCz/JnHHq0I2NhT2hvl26dT/XrRHU
K+xhQjjaR5eiUTtpLw9pdBs4PoRMOZ+j2ZLrpDuK5BCkTqlfXg9NW0aYyCIw+LA1
7WXlFUr+Y50Qt1yBW2gEQHFy4J20EziqOOWJ28BErHkqVgFPuMZy2hqCuzfoSAYp
MVcU5nf8uAWpcUe1vJpzd/iiMeoEIDflOxnJw5EA/lMTsAy19ykeqvon3NAwu5Bz
QUMM/lLvr0zsLTuElOUxwa7MqOgXlXijnnI+bvj8w3PHdFOBakOvC0q8PbbxecZH
Oowr8iq4cDXpdAfPocgOfbIS4CxhDha3kaVV9ZCAU8jwW7roD/KX6jFxAGyBla15
+m0U5BK2gNf57mI83eDN3yOJsGF1jXTLnCbbrjg07YTHiiqP6PP4mouuDCtrxC26
HuFG66zVBEYxpg9w3QywL6WUYXLV/hyj6d192mU3JLGBdvNxd+cSP8b9R3+qgydD
GYKgtWSDMmS/Q0eh/PD06tq2eXFrXCiP1FhYdQFt9r5DlTV8GaYUY76OE02aaId+
YE3Sjv753jlSMBbcWljYf7jd26O+u+MFNz/Y4sDhEZUFt3E8uTpYOd4r7BJQHBa0
FzFtserZtce/oOMtu7U+aQKdtH+CHswDyoySu8tgwl+hjl3opD669ilIDVCKpUvf
yfAB+TKsLYTeSEEm9VsyO6XL3rWgCKDX13Gkv1FfsLQOgr6gwi/TQBUBqUkRiFFt
JifAA4UwolhClIDv9Wbc6a2xvxvGFljLFGHmRzowcOJXWP4muvYdDoDmZYi2OuG7
cpmE0feyhG7z73HbTrq3hu/R/atqRrRHJnEYxm2CehFeHdWloZKLPV0XvPLxufFL
HZD/PET0euYHg6kDy+w9+lTAKuLMs4JIZY7GAMK2a6A/lev9gmRADiF4NIxzuTms
QRYNlr2+4dC9mSZTdgBCHPvrGQt4b9vgzlOKRHPp8nxFNGKlaGoFXnJllmFpr7tP
oGmLIqgj4H6CgMOKtgXq/nEwSH9Cr/wcfZbOi+DgiLfH4Mz5f6bhpNUtDZ/AGaYz
5W+Ycaibcc5gs9oye9mndBs3UNgqpEiW6P3yTPc7kmqngnxtNxdSNCLeRdoW/iqO
dbBkVbX2U/CxZdeEM5cfguJ+F8TkYIMxPc4MMI0WbFfD2W11cG1jRWoC7ane9b9n
+Xanw82iaanwOW3RhXHZHZP2gcINvHm8+MC+ja9jbQ1O5shjxenbLp+XCWA7Ouc1
nH9pYm/LfdM1KH+FVbVKlUqi3T688AFUmQJJs0+TNTN9ZJjDjbHRPKY3r2RzqyXl
CXfTz+uFX4B0MjeaZvKOWCwniXQRBCs3W2BeHzYABTeIMGRLjHmqCTqVVUHWH3I6
8+TNo4efvdzyZYovpdLyNpdmqol9lA9EdVaCmC47oFpT+xY/0a6nUK+zDTxcZNU8
hIUrWHC10Hni1xfueP84Hp+fZ5EpJ0y9dfBQHCRFvjttXulzqxCGmr0bsnEf2VMQ
nhWCrhVIN33CvzLcRlfx/6SdX1I2hVaCLrA6U+Oxr5/PSCT+v8yWcClQ/2RTZnQs
dnVdzGNN07tEL4vfj++trvglUP6FDqO7uDj7IYWdJZtN1UU2JHGG1jjk2+2TbFUA
QFyd16SsryGu1Aur7SsjNi76M+JBJBkUagzd54UkcTMret1CCRdMC+jg8CffLaRa
B838cLDPFOPxzKbWhGQbuld5tWqcLjRZWhJrRha3eI5fBwqpxS63uTMpwOkhVawZ
AYooJv/GNUFFfNJlysidCD0lMDqwfcLqyC8NMlQWYnfxmVRW1RVUxrr3HuDMCY7a
l7YUdxWXZJl8RW82gPhjf2E6J9d3PZN65hpU27DnZXGrPFNZo6R1HijJP9A8wEk8
kGlO8Zd/kHDFaIxY2VPzxgGphhh+PlDmVptoprZrf3HsqA3iFQ303aNqmd5pTMhb
1J+Ia6ZYsvoz1MTITPncMSfPKfdOIeg+0Kdv4AfrrTlYolRFzsZ2Phx7MQYGexaN
zaS5zzVQp8emsBj9oGxDVS27L7rfp+WoeyEnh7DVeyXLKWKlbD8a66iDyylWmcvO
5r2XZSlCP8wJSvO+iI019RMEYLhOwAO+ojvsSRJ6pX6qKfdtUYgoLySF2B+gAIR2
eIPyaIJS6FLxYz5+3HHVGv8lhn2vkJv5ei+/Z/5sMWwF3GJK02Aa1GLZTzLqVQwM
o6A2had5IHnsWJgBO8TpUJLDj2zR88jECI8LRj7YRD8RigOhNMkFEqJ62iOLsqd7
T7igSa1l5NExV/vEH6/5Cbge3xKt0hSFE08Ylh6S25uJmNH9R+BBU69BlV1PWPJ1
V3m/CZWPGRG3Wf85aqku4Oy7ORo7d9sbfqHG33r6gl5aiFds2NrJFvofopT0dBvL
2qx03SDNZ0GzzXEyAuRFrLSo4x3Hc64MzB32K2kfHi9rNuosGn2osAFQ5xv9o6qD
FV87gh5E9D5YbLoAAVYL8l3wVOYisZCotnraFfrJAORqDZwGUIpi9SrMlHCMyuE+
oRcbkD/kHPZ150d2uvfOIalG+L3KgoTB5fD1BXxJWkn4MfgcrQXSfV5ZX32nyIzR
w7yGmjA6+c9IABQTVxTBlWCsBP9mOZOhAin1LB7NlLx+M/YewngBu+BMe1cU0fHW
bu94EhiIDjRbsHQkSPRyVNfPVke3TzZ525Xv4sFdKPwnXhTdJHY1X5p+x15u1Ydv
e6xpJ41pKink+tVDc1tq7xAYYgWBnW3r43etsfnE7J0fGSPQUmchxawoWUcgSKkh
iWpEY2uw4//9KI7REarTRLu3y1yTpcGJSc8ylevMOaUFdP+rwwDCjt0wPnsXgZ2Y
gWW7Ue8Vx4V1huKMHC16+jBw9OyCjfJsXeMHUqcYyJ7tLycQMwvHc+EcK43jnSoa
CX08oCuynMyck0JL4xlCU6nG6pOgOQkZ30UwCkfB+HkFo8Q56jEkX15zuURqZQMT
DdUtwWCqHQzEBQO+EstOo3m4fAds6+AztPOUviAOans9vj2aJ5cl9d4Ghd1C02Ur
hdO+hgWCTPcKnkLwKsl9QGm47S3NxiygoBrJ14c4Bpoc56OhdApWW6UoUiS4vbXg
1VzhgcP+Y5ER1CDZB/YZ2WqgdeyBoJ45NacA0TzFMfXJcG1hTJshW+7xVZkJFxIf
G2t2DikW+JUKcnkMLQ51oJaw6s86EFqGy224tjrsPjlsP2vCw4J3d5noy82TzSN1
hC6OOqI5SfnjLP3QZ+dQVbqaKSUvYUGmOYksQe75O7wfoKYw+68ldjvGOPJVMpwy
oT0q83M596B/0nP17J+ELL5XCNtNknJNhOzaDTkWe8OuBoOkBO8nAWN7bb4mf+1U
rrx/vJFwoWhHOSJXdvPqPjerUQVsvZQmceBj/MxliV2NrvasAS5+0w6sL+ow46Iq
Wx8UmdM3F9W4A0LM1+Kp/DUxFAg4cm7Nlb7W/XvrqS7UFsuqyo48Jxl0WkqpoUDg
ZzAmVNz3Ig8GghhVMixd1SAUne9CojoK4VKnaPektGDFrc8gh4gZ5hObPDc6lp+J
Gq759pKKp/A0MI8BLXLBFIyuD2iHasMH0or//o3BojIu4sdGKOjkLGOCyXrlZOlG
NkfNzihCe+8jNi1l59EonlesWLT7elc3KzeF/5p72DS8MKURNtKKp98WBXqq+jB8
o4w0aGoCdht0+IZIDCquF4cbpws24hjA0j3o244WgjUvDDdQEAGT4k3QHSUCc79X
ZqW91LFLG9Q1Gr1jhosyVs8WFM5oIqNbgpVRztxdKf8xrlRzNu3iCWp+rmjCWAUF
FIGmGN9mtqDrPsuqoTxmAVqQH0ezEYoFOXtB99aOxvAlTvxFVQF5LoitCCafrsIk
lAg1WN/9ZZHtYsVZIZATucov1750AQKHw09T0HRg6Jac8QkbrluUaKb4loCu6LaY
CaeeFWn5vXU8QRmcBbnNVe1RHrjBNyImTm/8Dh8elvD9S46tuSGs0ufNN4EUo3gg
FMuNTc+2KCwMUFWdXUlPABILICRAYwlb6E8zaqfd/h8SYaXTy3cEOTjTGFJMwPJ6
n3XT6Vejd5Gkz+H0VHY8dhv0Ack38IzepUuOGgkwfGnsjygNtfZkta6OL/LK6uun
pckTRZkURaxQIJthNP9lYgIewGpGfbNgj9bt6AINeAF+rID6ndvcG196tDh1fXuc
KCyo0fKiSV0xbf/RYEl3VVCjIr4uylppnP2VWfLq6tE4wbi9bHmEkie/ZllBDiRL
3uLE+srVa1LvCYD9kFRmVYfBbLJL3qj4pGCLqD4ju+15MU8uwQODeiuKHhyiylUt
g/lCtRTgPKt58PtOFzueATtUqV9Z3VPeFtDzxtC69OoJOqb/CWxMFv2PAr/RTtdj
1t0KPsJFe6B/6MadfnupQDonN/cu3bF2kgqFJA49Pk0FP6Lgqs0j5gA5ca0OrB4z
CZfaKK5X3PEzktwANzuX5Eq2868COfCswhLGsqbQalPGSOMy1R2WEaC4XEu/q9So
l2yAqe8ftqFfgS5b2SP5v4Ek1q5tZhiw5YYAXZmsJf+AlshAYd7uKQr3vqY72GNL
8zBoNYDmdfsgwZawmRSXG1te6qzimw38OV//ZsuGNwtC4u7MCM1EoXiHUAiLeEl3
5RkcBoZlVjApm8ULs/syabidfFVtqXpqKbuiYk3Inn6aw3lp47pekE1JfsYP6QhZ
8bwSkllZk6DGEOnONXRqm7Rmw1uKF4GTD9D7lvtWXp9Rt6fkKtPyeBkTpV5wx0AG
RZqhJOuDCaQjC6ofgXdSeUFzIHODxDe19DCnBX9Qhi1a99cKwiTZajavNEEGwfAj
i1wgPV1U06fBLu4DPbeOvkHYc6BpZImm9TgJRq3pKtd7TkKdwnr5jqsNeluU3FWP
mYjkQcgft4BFhUanHV15NI973v2i0qNWjOGbl0XQsYa2vZY3HCUTuyDq0Dg44t2r
L4pNxyVGmLZNlqIhnJOn7QxblmlgBJvx1R2MZpU6biYn8zAXeFIoSq3HFQ6DVjWl
3v8YnS5ez2AWh2AuO4Xx/KNWZ90O/Dt3atPqN6ynhvLlD8eKLXQiB8NxSVRbUc6g
hyvhbhSq5SMWbJRRzFEQJVopDkiYrh2m0w39FBDshVWuHigGg+ePIHLIR+E/qiDk
bX/rq4l/xDOKDC3Na+jWFAXV49VRNeWiMflNl8DMhOD2Sj2z9hoaJ+fiwH+kgeEh
vQ0MOEMAPLjvZAf+eCsvgcI7ASpSooa9LGXYvF3sIL4OaaXFfSRKZ7KbLoWiDscd
6Fo7bmiR0pzs67WRs2/Zughz9tDK6f4pkx2oax6RjW2xHwH9mkMWDYlw23zD+jIV
WCCLgsZM5kWTArvk+KFkijFWcMEGrSo8cQjun6kRPSNsgEHPzCaV3UmApQFHQHuO
GNtAmVaKMR0tZtByr4xnaF2rzYCoHUYwUrKTx6noxhd/DVRSIgFkHLYmz5/P59zn
mr/xIlKcInkni2qyn1n+PXuH9FbPtxrjeVwHcsSB7ZZ9AhyEXLemj9ZZT7HZPWRY
Qj1O/83tydx6u7JzeCYZCf0bRQPxyI4rUfNcvW/AsFYM4yvSzS9vjuNvhATvVuR8
yI+H0ZARSZAzaLb7muc8jejQm8/+cfTGg4rPpesjzxAoOHiz3rnjqIPNV+KYI4Ud
pfn/zIBEeXWfuzejFfjvhrgWgsDBfZU3jaBL0CRxfdZyHagx22b1dUkjX1vvYx7H
wLXPzF7ylQS6ieBldaohNDwsV+kOJw4f2lwoG0ly+QUFQS/po9twv2J493EL8cNE
VsqxuTt2VjSgpsp1x67APRhkUN0eYVLopBd8wgjYVcRotWouMrpHbs1+d3NRPnRF
BmX+bFWycI2AfzTNdq7gHz81w8AK8BulzFvLzEL4qJnTXz/rnEwI5bj9hYscCHBK
BX1V9gxFhOvFzue/RWhsLkLilyWouX69ENJvT1e//hBb/OBHhs0l0HNvxsqUJYsV
qHQ54GKf8VngmIBbuoHiL1T0AgSEN/h4Z/KA5qkFLdrxlrrkBj3MCwWRcM7SjanV
8RXL0/HWuFrRIHiokecaNN+4Fzs5P6jRQWngdnciEZzZkC1Mc0PoFzUbx30ELYaj
DV9vY5BXDOBAoUsLK4HTQ7k3RpTcBBhEByNGLcyANxJs/UBiJqsA7jezaFDOwvKu
7P/zxBygCo4GMuOyL8UR0LuUCuV/NS58pGqoQZoe6B5OD7b4PQ5DWuBl90YOE5Kz
7bszebZmqi/ekwER9Pa69A/9IOllAmg+Of3gVc/tAvJidsLf5LHX7PSjxrOqm86A
gQpOT+X/OHe0FhLDfVkNHYpBKiBlZKJdZ4x3yG1Lk8hKgJqjlFNSl/sPmcbpweug
7Gob0pt4SO1i4JxKOGNezrxL//Q/8/Y30KzzBFOhl3g709ootjes8Lxool4agPPd
OegyHOcOG3O3qje1+8arMKZ5pvXksGVxiRQ5kzwgsEbUXYyviuvH0AKQxQh2A9dd
6cQnemMbkj26aS9i1Bahj4Fi0EXsUp8RfEyVkASRCeqM6OEc96wDNU6c4IkJOJhX
catvYaLUZdsJtFMYJ/Qu1q9ukV4aNiwSjxvMkZ8iJPDNcOHKLApMnzvYjhUmg7Ix
vfRrRwW9pVJVK19D79k38CtEQLRoPMrB5Ep9iXC3bDB3PdRYHbGJaLDQRvQmjMSW
jzXCzX3UPvjPuRQ1Wc9uwS4wlhz80HCpXUtJkf6sNiFOn8OETw8yU8ICfxE2R9yp
HaqrR+WtOmVRWKjqA629VfUXTXfHFqxw2pDvTk+I9L97mSUuWEvjQ6hllmouHqQH
kvyS8sqPUonxb80UVhU4odpfZN/Dh2d8OiNe6Mzwiae454tKDAbyMwuEMe2QI4w6
JkoWNBEtQGFkw5mtejYhXNdsUNwUPXsMjKf7op9z25mP4rvkJ1HTtq5PyMZ9rAhW
toVB++9Ofi5/pgYhBDoZrLhI23hNadKzRjJGk5qTNb7chqX+HK6tr3KEVsGrnWff
sRP6FdwxViUQL4RfRGLrPxyJpnPmgu5UC9ivDUzCbrapS1USvFMj9G+Q9KdgWnZH
4ldhFmpDUjx+Q5puBf7iQWUp9QxnizXJVEbcBX3AiMUOVEaITfETM4CkFBHlS2JA
NgvjRZugiQpo3PJhYbp2+agsV/MV6ruCqTd96717VNq3+SEcMpsxHF6KQQoWtBwa
vuEuUZdPiTB6J2o+4VE/JcuN7pKGzEaIR/sWM0dRuZlbBUUnR5Sh9j/GxrLnq6Uv
RgdxI7aMXzNrXmEEA5wEwGD2l8HLfPNhABFoC924Y5auWiNBZZbb0xWsS/cA2De+
gl5rLOoRtHYv+VVLNJbxve7nfC3XOdRXWEKUFOd/t+kzTpqFyK3vRKUWvs5J31L0
RianXxOttPoOhTZCyYsSxQsH/wQ2JPY98ll2aJiBIoBDoT9wCflHaPa0/4gNfoPP
UKq7Obwg1qfteM6Vr4dOAxCWG/rCySv5IdmJ0sPJlraXmHMlZztBuN7WAqngOxRG
2hlDzT6kWlTeOT4Ft/n9427Wyv5OqSAxZi9WapKW+y+t4mK0lHS3LqjFGBeKKB6i
cfK753bxx0aYhbx9iSbVpp2TXw4b1MSnI8MR03IZSul9b8EorEOubj6u/CC3hhiP
KAi24US4281h5ZrlsTanmNIxtsaI6s6K2Lx3hbEa9JCuwmGnRoVnTRu6Zlpk4wPr
4s880m5F7YyCbVobuLDA0eoEiKXXI9Pl99bzq0q5Aisqw2PgOjiE+KYzVML5J0G+
0XgvpVywtfmm4AlqwnxrNMK/JoxfyClg2euqPGdKD5pbA2ro3bwBYJydeKj4CFOL
OIxnMPFKFuD5FcXt4kHq6ZlcCnsRG7TpNFPEkub6Fc46JXnf/cG4PWvLgtfteKrD
wsRHLItk3QjIca0nyhAfMgvmuJGbSXgEote9oXnDbKd68rxMmus3JdzPSmTBk26C
zk7lhuN3hD4clbWF9swdSWIfw6PzfbRJnENUNMMxgL6LmEtpq1vPrt8WZsiTssDt
WA1VzRhj+9sXHAHrXWuZFKWAxuoKj7GILMq4taiup4IJM4VyhrARB4XZ2Z/HZJLW
iUQkL+lP5pCpKWkFOnb0UiKN9yvOKd3Ez7kdKMh5k1JK/wYDfOE/hP7ZGr96n1h5
TUk9EPNWmljtnN+jWRVwalKVuE2hTGEJjveauNj1vvWG6OrgPuFR7/23l2h+wwTm
k8KN+fE1Ot/X+sB1so0xIBH7184gpcWgrcHWd4WqCdiukZMf6Y634S5XJYqSqvEp
s1JEijy6AY9nT+byi+fWQnNWw8baCxZWrWX/7mVJXeNCGwAZ+lNKENyYmfwAhd7Z
SM69Zz9RpIU1NXeoHNvaF/6IGxp+cQ28gO6QS9oT6q+2KJaxXErtWVEaNjM3A0sb
sIHOUu5DJLoa0qK5D88eUhR6HiH8xZ7h8ZsKh0VHZ7RCqYh9jn3GiiuyrejDjDlW
Z/tU2uX4vQdZgoBaQKx1MbH8bVLrkxQpvD9abjI9BLfInLXALk4A6H1xegYCdnDJ
sLOdnlGoFDQTs1IPjCJqMlQkBcFD/SZAMKaBQPXYvj6hO4S9i1DIsilXJiy5Fx/y
mYW+NhsAORfXK7IfUKZPCDaOCtUEu/HqKirv58C2y9iiPEwBGTyO2aocc2XDY0f1
teLtlUOHi2guoIXj9OKL+ejjhpHqevNAe5zvE2yogaiHW3SWS70dY/VtDnRtlJ6d
j+rajdW4yWXhiy3lamLSwJyN0jOWs1MZQgp37XCuaFfNEOV/mYpbHRyjtFDRyDUq
2w5SmqqGuiA/xyoItlDW9LkbtpQxfXNWFzz7LAEQvduFtG25K6qdi4ZXCzYHFQrW
dtAS9YQwMJF99w+CTfkGsWqi0gzitawVW8hxQq3cdVkUGQIvTL5mVlEuu974EMwB
bJ4ano8p8jBbBYySXxsKcZUPw3leb6kUpf31RgDZU44bdo8Uxd96F5m9MnmQkqby
oyn/AOMUdetgD5aBiIx1Wsd5FHwEovRCKLRBXHfsZe8mD5K9Zg2g6WtV/ZWQ91r6
aTO1tAF/axV+kTrKMCv5x/KORigmYOA9h4C3IIgPjcGYXkE+tcdZ2ErsABG0yxM9
8UwAfiMVZeMbi6lObrCVJSS3sjQtg3mh+tIKsiOlyqk4p+ZBs4XsVToSq1XpKpKf
a9Yg/JQc+vNfhfPT1Mnb0qeALX2mllhf7bE6HrDw7O10//Dhx4E1CYeGk7tsCV/1
/+BZ/NBcTlmdI6ynEzTJ+nkiCxDjB4+MJimju4W8vACysU6mPtfhxIk7XSU1IAzg
J20zaR5somXvoA7AagZa2Omn7kuQCmQ2nM2H/gXkyt/ToTtGJCwwvRL2vskCFJOC
DItRSwYJ9QfzXNClvfuLYyeUzi/i9xiy7hdZxpaj5yzAT6ZssUi2GGm0bCLwoODT
2FZe8ZRSvOoPUzqT4Lbz494lvBWcEarK3lb5hQmA8iKSS9G4dyoGsgfEAegpRXE9
cXuPg2AgnXQbRVNGCXb16JhPtH+f5G5AgY9h6f3LT1Bo1DuReV/JJuISVCbUt0lR
GOIgkp9cYYjoDqRPW+otDKW8JsMmK74iVti+tYBsyxnODmxE6AQUggNUX+RhF3tw
hHZTem2RwdEKPep1XCAZaNzGD0LXhSu5IpIjSeUwlJORMeFoPR07VcjLA5IRNFl0
ScO4ZNO3zx73ZCNTmlf66SOb5/fKBnJN9gXUNVaN5M1BUnmttz+jabI39RLnQ1v+
Kn3t8AhKO73cLdzfJEroB/J2QCrjj4Vz1MB1UJBbuTweDAmvg8e00eWvPjhtR1CR
knSFiTUkdvVICadTbOMfuPatj/MBQyy0eWuQ7rN27YFIFcDtPvQVzubMu4dtGf2d
LbseAW0laraR3sPgzBxtCSL2Pr8nyqzUQDnYyZUZiP40Yl9ULb84LF/lK2rw/bn4
hkfn0U0utipE+zyLD/+guW6KmRzvCBl4cmMrgv0j0F5YThdWKgUgFufeKiabynMu
CCplQqYfs9KuKdapTb9tg6KrAsNIN70epRSeMvRxX3oi2Anw6ZohzZdsexsnMJRZ
++DnJWO+1v/tv0dTatnN4oxHM7/11aKCLut3OkmNLpgB8GaDr+WZJmkH5BlKTLxo
1qpJyZZFVJVPmvOkVCasAAdqVqwkH0SD1WRkubXZyxow0/wINS7kU1lRe8xf6+68
ZksPrd/DEwg0wpGGR6pGno2Qd/4FMmvmGKvqPIhIREEF51ntF4P+SkjqmFr45tTh
k5B0aSbbHYX9fYsXSRxph8KxVoNJ9xzCc7yY6JkxXzmyHDklpH+mIDzw2U7h/0J0
aykCthc0vYVmuhCEH1CvbJkMjGGHlMdPUp/6WVloixRL3ZUzlfoBR/tgE36QbNuu
6IfDpOAusgfnq/zG2qgxDc0eCUAuDZKLNVkDLkcctnY+e2woPpXqsoGGp4wAM+Wu
Rzadc8WemRqvUxkr649g8zz77uASdle+81VnnUx3H4zlENu9AlPwZEHLGWAZw8az
Ea7CQN4yFdVcDvPT2sMlEN2l5fyPBFNt0pSRFxRJp75m8A8usye33JNAykBa8qlo
x3Ztiew3tAljQPjWPErjIWWKDaDo+WZVP/jSsLMgRGNsc4ZbjoilEeY135MOSefE
gWdcpDWX5IHfS2YckP/+2+gqfU2SDVObgPW8UIrBb6T02opjee4mNgy+eDi8WI6Q
Gvc7Wilf0/4Iu5FhYU1XeWOsBftK6wyvSomvjcBGko0gtbcc1SdC3Ao1URp8Rp3P
Xdt0InBPSM6DWXGyQKRhwoK3biGBw3EnC1MRAWDWg1l+nVNE+xngc4d1JOaZrEnE
OyMDYeaiMdThNCiEj80v56hw672X50gLDYHK/74uBIbJtG9D85mcqPGAWxVFrTF4
6A2Jku6GGUwKOFhFug1q9nbLc4aFplnKnrmRfyL99ZbDdgsJnjzHYnc8E+OYn5AE
oSsSwkpnpjq4v3P6lfeU5ESHAzU7+87vVaEbz+dl62KhCBo5wVBIyiTqbkvoMih/
Yliy5DtCmgAgZHDCaH0wPGL4d8ED/v49B4Mw4Q81RZefZ4W35NJsLw0RK+Qm0mO9
+taYmpcIaddMK+G2DbJVGuasuuiIuyIdULLSyWzbpGRHy0bF2L1oZpHotVI3Cons
aI3zmrXsP11YZmxytgzq0LJnhUcF5Uvxfle87ByHzyZl9gMI2A78y3OFTbGUWZFH
bwMsrNmR1MX9RYd8zf8UPEP8ONJ8fxKB8xXxuU59DvPtK2A6AJwRPzm7JHEqC02j
2o1qguAwKdmbE2N9a245wqkulN4bFEELfhKbOPBNQBYqI6gkP0dp6GQVH+pVnUQt
6rdOFzeFQqnB16IWqXFQgtXu9glfOeGUUpwKjbLWfUIP0IHVNgVRjvpJL+4SD7Tq
k2rSWoQWzixumKeowoWHQl5bml0eKwIded9HMTpR1iLdg7YldcDTkRfqecqdLTWH
Jc5QASSS3u06ynkJewTNWMY9EEGrpw/54wvvm6YwZfqEpDA6nNTG96947un1732b
Bbq69dTk+FsrLou6e71xH+77Buoma3mocnoVnXl5DE+0PRoi4pFYN4Al3V9BsDaO
Ilm6aRWuTJ/Lvikx9uGanEFgPU6uF7iq+d45XjhvThqSFpsiGO/RJ8Kts1pEwYGO
kpWViwMItID4pMOTQ31m4enkyEI82ASxqVkgvXiRD1yQYhdCMA8LSI2zyb8pXQp/
kZHm35wNLG1d+72yReTa0Rnsr/iPUGzOlKlfotgfPp6GjnncgxZ2u5KSmilKl/lu
jOSUKPS4PFWfh72agtJULoXByMBop0jd8JeWPkedctN8UqVhD862OQxRH1jjAsPw
SMA2/+fwBNJGh27aJLo4WmQ3NTTe4ADRiVGt10RJRERYct6mihIfeIPN/n4i9sgg
sRlERxMhd8OfX/Cp6kZlP9ondoUJoSkgI2U+7vdpZlOjoA7AAdfanv9cKDLfwX1C
DS3bV6O8M2tDMeAl9GyufzrFeesXSbtt0gfsA4l58Yp9/3XzKbeal/jMV3Xd2uBJ
7jFjdQHZjoXbHYkbtbPeVs4Z3yRhGsdZshkLM7wpWe6jrMRTAF82HtBvVogzRhWa
fWiOFHGLUxFxqsBoVSh4OsLUQSYgfo+zLFCScoghM+u4j6pzuHkVLXSw4x6b55jL
OpoolCtjYroTu2CvrQRgyIt3fy3C1xd1196B7lNGfbkUOQhUNjHFBdfNPPXSXYxr
TPbomKBx1uQQB/XatavUBgCQcrI5MFnbnG2hl3VDux4Gg20K60DsFdAMDozmZMkt
05zCxhnSpBWlmDrp8XRY7+AIcdyofDWHDdLRpz1spAOiQ3oHn8gLx4qyXJJP0qM/
tiTt3z0GMy4EYTzDPnSRdc96WORGH/872/LS4q76SiFOwtnL1AGFF9CUX+XNOnBz
YnwiV6TgEMAhh1vaV/8pVzw+c1yIJ/WnAcUjcOc3I1CVO36bfcI+xCcsDIJtPa/g
LJVlwzHdU+ai4xSgbzndFBcwOKhCBUJgE5ZXd6BhihW98l+2/jCLb6ylgvcKqmlc
jWSCqjRI8/cIyx+QRLb4KpLBwf18XWVc7b7DTa0QPDcYH1F3EPkz8ybwgN55+Jfh
4ZfBEPaGuwirbW+9oGkCOfb4SalSjtLNi5O2jYaQlJBEzN9DF+rkZS6q4Z7YZxo1
B5kyO0Wtipsr7Cb410MVEUsEzs9A8tO5wV8Jd9WuLZqQY2479Sz09lCZvNb6FYPy
eg7NGihScdXglW9s/ig/2coAsZewY5wVEPwGDZbq1HRiJuCViU0gre3BC6GnL0Eu
v1KidtDhQIeSD2FOl1MQkkzHJUZUYRQ3hffLQC66KMcpKHgx5d1No20lrZ1Qt1vc
B0+RBUG4Xapf9UqVsx130xnvEJ3F7qPAlx4wR9fJwN350NRfYceM/FJ4N5MaZySF
Rjqpxq06GSoD1QiuBeSKIVeHz49nrmHNiue8X+Z32dXRkkD9BVYTL5sX0nnTRmoE
jW2sxxp/vudk1gmt1msLSCNz59k+1/ujDNVVzSaZ0HIpVYBoBnEHplc4m158UJby
Oxrim1gnM3gNbCkfObHySe2rfqexSbu3WwyiiDd7v06Zt4rGepbwLveJZ9DPNddB
NP9guXpYLi5lg7U2n2hPqxkik6C1XgtPX8Mi+E1tkIy3tlT8rWhgQOjaKWZpX33X
67wbBCRmq0KtF5AACCFwSqFFPzC9afYlQBWF7RyUtwx6ht0dCVCN5O8+3ABj6Bu5
0XA7k41d29G/VimXXyJcbgTiKdPxipDbVTKHzBe377ux4Desupv/06dWWHEQ3Vg8
RMNB4ZwpPMXd8kpac+7j1mvurtNHnTJ5TziL4iUNVeh0/BFgONdsC5iECCZSJt4g
FNqzbX8juX7PqzQib0mT6U2X3Ng7rcQuACCgBO3ZjMxL8rK/utDun6+mlYU9J5iW
+tUiSDqatDbyRre8MZqsZPU95wktanAo//fZEySKN9tj0emToKfwjA6uG0JWyXEr
QG7+IWADM7yMkejyjAgS+8l6djGgQZkOk30o39KHuW71Oyo0d7fTkUok59ZiwMJn
A231HC0VBYtUJfgN7+0xEvLe9lAZLojxDz5hZZw0bVo9BWIVtiriu6kHYfVUkpVL
HmSzWa97AwLzS/ijx4zXl6pWvp9WHK7vj/h73LrxIgNKuecYLQVC0ndutTTS9Rqq
+khnLmlYVZWCcj0smmsId56b/grBf7W26lOY1sFH9BAe+2nwJvuCJQK40+MjSlQy
2WJQrmmLdWqNAh7LQdIzlR+S6OVSrpLUUOA3xJ/1XjPYZFMZg8DSInitiVzAW19e
9pDBZ8FgoK1khz10ywwsYiMf5M0Gqn0rplv/rWl0uVCNmKgoGGfxP+rt1inQ9K71
VnA3ZJ1HFLEMSvHl/OjutlYMYlKbsRm1XFIPUBN80kQCGIvmSIJryc62gv5p/Fo+
7R0Vjv+Ts3IbC1yEvW4aqfXTqy75sH23YUXstmi4US0+rbD3zd/wMo1cmONzpuUc
wXFyD7FplVgfCsn/Rz40I5a1SBIGMSfXjGjuK+bJ6csfUPVJWlBJYRczAg/O/ar/
IzRYXLcM2OBDOv88NeIxTGjRPCxyGVj8kjHw4+cT1Q50D5osJ15qpKZNtuw6iCWu
bupSFrHU1vWLpp/mNb8RHgIQcS2Ue7G2T5ysHCWMwtptaFlRLFjBtqoiUzt4Xvyb
8FntaumZ7bdXye1vqXggiDt1kWDRf7dHqGUXyqdQLe+5eRfnWpZVCAOABFKv/3b2
f08j1ybhRNfw7PK9kg7jVWGz7S/ABxLNgyp5I/ZRLQvLHh4kDFHlpWqMBcPd9SI2
00iCmhXZTuN7MtSyALCLip52HASzBqqc4TRPajGfSsTOIqL6Xa0Wa1Ukb+urAI0u
zwxdJM8USkUjrrrum/VTllFa79C0JFMgCUwsbnZIxSjMrRwRK+xkDIbwD+gDTxAd
GkCAqlvUorkMWq0zqZFW0PsYdEiwgdAMn/EnMEHzDaoIGnnCGI3Wh46Jez+8KGQ/
BXVEEdxiWjgFNSxedrPy3qCh8b6PR+2xBTBD6AvwHylZ/ZwdjIvrUrSnFYnZhI+M
CP7d5B4C3rfflEvFEZx+J2FQknN0RJf3SwyOxrIqneCpmDL39PnHAvifQmqNyFAG
6kcPpEIt7XmozjoATTj/vvutAMZ747LxxfXDyn48K9EsekaR42+J3MoWPAH+Yd/7
H9z2fwEeyNMHHKWEaR/EpN91+kWgCMZm0xgBbEJ5YPyHgAVQPYIKdD843B5HFI0V
XnAKzQzejNJkTf58/U2TlddWiUAyEM6L15Z095Ft8TMECuLebOge+j9o6K3SyJD2
dEZHzjaPSeurmhYu07Gk2C9VzE43M8bi+9mRqYRtVPNCWH4aoli3pWHv8eVpKznD
w72NYmlx9SM1TS9vMePCj59P7HLUtz5LBCjTdRDFYzvK72w8xO04HolKMblzCoI8
frr8BWGPXT304AceoBf+ou7oYD2n7irQ+uO2AUOsgJxXbvwIfCCxO2RBeakhK/gA
d0pQMquYm0LsNGp/0rEa/Pss9IdUMSJ/bnMrBqHkRCSZVEvdOlnmZLuOC3kOtXVc
dO2GZQlk6x54D99k+wGdvaZqI58RxZbChv9JBL9I9rBgyiAie+MlfSLxzdVJNc0C
EN9WTQb5sgeXiEqbytgYkUBLlqC9RcAcgsi6tPxYQpRFdqZelzFABl8kx3vfpz9J
CVwSNtV0IPtGLgIj3kQ5CO9p+zcXChB6MV3gTOXtCZPubXsqvHWHRDz5K7qZA2QG
tIqCsUCvc8y2HIkwPhepD/Lb8e+Xf7VM46xvhAsLDLdSbmGtNTfiAhW27g5x8on/
oL1Af+BIox3m0L+2cqSW/NXCtenqIv6aZ2FFoCREg3HUhCmLilkJEeC0M1ONfeFY
1K+yXg8Q1QCaBiVXe/KArNOa1/+ehCgGjM6cGWTSf/JbHYeyCncdmNy9iqykXX4f
n0vYtnue6YiWjUR1q9zd+bGk8pCRmZCyU8G2P9zOLh6wd0PTBwDsvGEntK+0NGh2
i8uNSGM1Sfn9n6+oMwY9qxvLFjzwI2qF6mAPg7j7KL6lRbr7x+1RWLax2IOuy/8J
2pRffTr5+V+Jv8gPjMSxLc5qyJnkJjGhcnbu5/GB5ut1O+EwuyYkiEAJQsmDHXFt
kxoPVMbdhIeDx8spaFsV1twYvRBrcvrPwLWS0OmWfjCWREG9n7G5n/12YmeVyoYt
RfFwGmgIPMEc/ZuCNOIa3v/Eaw60JtX6Z59IvkO5WG5HoZy77sPh02qAa3CX596N
sgwunKGh5vSkz2+QBkb7FIkzAlreInllaWjmqONAUn3Mc0lZzSXpT2K6xkH88LeJ
msPUouatX4LnNFCvv+FWpz47RAs0n5ZpKj6Zxf2NuFHK4K2Vic5iC6dbYZrBTjkH
H3Yl7CcHRuBSJCUwjW4a2BO3cUyXZg/P6WbZes5Tu1PBtILJisfTSb6JAoHqyJQA
ezUxtgZ5yY5CsuX5hk0MM/LO1ygJUICMo2g1fH7/pO2S4vozO2z+oP1lH/0oZ1oB
YpOg0YWLSXnGyK4pVdYSow+sgzRMzZ405fAe+r89qcOOGDB+9xhFcJqBz/GH5U5o
q6mAmVQ55kyKk1EFDjqssXQdh2wnOvmp7Z3ucEinyQCZ71uEvGudqogRdlnanf3b
mx1LWwC0Fn65P3YPlKLhhZ0PXqgib/v1H/ISYR199T1MkBpyGTrSxzfFyhkS9D2a
9b9qVWOTyiBpx/scx5C7WpMrs4A18EGsyIcNB533y+gyeudiE5AhqohIycikGC0g
NUWlKX171WdCeQGys4DuJUc6mdVU+tMv6YepxBqvcVmZiUWKz6mpgRrWLBqHiJ8E
U6MG0IBvTRKwAiKFRHX7fOLxp99V24d5pJOj1cVcIfWdUlZKFxFO9IpSIAYTwO/f
BI9tM90hCvaQwQ7+B/aSjlB51PrfMmub6RE/KSiYKZx+aTxnr3t1xiAPdNk+YL2n
AUSSPf1uzsKf+yUa4DJ3VdL69L04yciKPH7zlA+bbHvKWPoo+7srlnVPHXood1Tt
DSVrtUoOkZ+wBKAixiJDHQ/tE1KGnLALnJ5/l2Z3434tfXMECVaU7T8gwr0sQ6Oc
ifBobOKjwQ0iOYLwAgc447pc65JbnTxQq6EMMuBQjfy/Ik8F3z4aABqSZYr+vO5K
vTXAO+Hqjl2kKBXI10mqQSCdIhI4klc+KtmNCzjnX6BJF1J6Pew80+AC23u0/Yef
8Shj2xJyMBUNvpF+/gF8YhwtlvotYeUgrnz0agFjkxLvFv9mN3VzzVV4+cYqKwOb
0t0UHvha2NPO89+7cu3f9tHugO66h7Y2LkPEgf3NzIDsNzUnXqnAmUeovQq+DdrV
A4mwY0kyQk4iAiHn9oVJP4JoE/HQ5l60Mg/SXOZBratH2/PXcMlzz6Debsu2Rn55
q/JWlU3MxDuBRMWv8d4kbqjEkx+8FrgQo1bvrvCQRpDIUWD+Sr+K5aruN1nMZlC2
UkWo47CKcmjoxMfPuA38khy1hc2E++AWRg03A0DSAM7HQjpxIYAtEwQy7YndndwX
0sbCgDyL3q+3GAewz7ajSofBND24WvYpr2Jf4YCWNiisYZoBedRF/78fatzvcuba
HDNpq+4udtKZDkhq3mgBo322ctvlE0aH/JU85KFm+SEddpIQDkm7dCygTVP5qoXh
d09iTMuE/f+WRaBPaWhnl1vTHj0wR0NJnjHWd7uxtdMWE/BZaAqu1hjU8tDWUDFe
UDUFtI8WmiCEtR5p0rnAQk7eTF6pylkS6D2Q3DjcKQ5tjFBie5EMzFIEUwLSFZv0
EfNXDoyX+CFfUr7nwTdb+um+hC5v6X7iT3KAsewSxIFWEocDEYayqv3K9fTCcnaR
wl8CULY36DTOBniubalI+dO+zxV6Kd+VYGW5/CWxOkFgS0RJQVsolISIBmLPlgVZ
9Y6/225jI7/rUUGFSGKVy7Bi06upcTsKe1ufy4H5lQApcVYZQb7vEUT8YL2DbLem
uRzB63mazilcrsjYaKC9xb/rp7qbCJ8uhXSMw9iapvoofsqcltyBV2NVmABXj6cu
yRCUAt37r9ggth8RkkM8+XuAEzdBaApMJA7S2a+zEo6Tb9YIF8lAX5Lyf9ycoguo
JUqkNZcqHaQn02/4vpIVzz2m93g+H5E/8vuZFIRGTcEugofCmdptCz609SU82GCj
WA4C6x0yElAYonVt9mavg/KOUXuWEencZIxwLA4Gk1Nq8WQ9rlNT9dTTQWYBZkpD
UxR9WWH57fghA+plTSe+orJMwWBD7heKywh7uvbQekE+G9VmuTGKZPiDNY3yqknD
Xj+H94i7qLeKHPlwci43/qS2gco3MrI0o7HXBm9cittHBYN9Uur38OJWwmiRwq22
2YhjJtvmwinxgDlIQ098jt5EB+FGr0aRlJ5cB2N8rEEKyI9lJVuAAqi/hPC01CMC
79LxOVKRgiAT9p3RUK7l3T0DTiXXi8IK4hwVLzpJdf2VYV0a7iCNRJxCSIc3V10g
/JGn4LAzwck9gemuGNY6MaCipFQ3gqGzJmqVpXKylsGmzfirEMNEL5On2z1PBTXE
Jbz7yfuSmPTyN0L2Zk/uAvpWJ/x+HtfyQNfLUM+caFJpjFDnPb/CUY9QzugzelR+
4jZvXYbHdHEGPu9MZzcWhr+OU2/TEXOK25TOOI93ydGVqep8H+pXHYFM+jfbM/rP
xveI4e+oY5QgqwUTXuZTyn9nJimXKzq50AwI2qWfxP65BYA1hoo1/iExiqf2GJJs
LT/DNRKmoue33n+B0yfDAlosPMj4eSU11ZVvhAcUbpRhTp+5v/3Q3UuJw2Gtgs7U
8F7RnEHA/PpklPDpyH7BV1xNpLevOhvRGrp2H9Vh4prbQK4Gwoogpzr4DkcPyidG
uvGseA6Hyq/4dzSGRyMAAcgFq2G2Vyv+MHOJrSAW4JdrTItmuJIGfh0M2sTKcsoi
IHt+Z63MOs81lLL8sjNTILbZ/FWpSmpEW5X+mZ5LUB5zVXINL+82L88ao5Gro/T7
VSbTtIdMx194JFHVwY1jHzG11Xv1reIie7B02vlxtfGZtn1YnX7LA9EBpzxyOIjG
8I1y5oRmElxctga0O92okG78tZuYzSO7+uZdyJvNu5x0Hmhl1rJtRuoK/B61jC7b
maR3NzaZlORuTV75ebu4dw1/39gW32t41isMeHJifnjL4s9Kn2QPKAUowV7To+Ff
/2DrwWMEh1GzMnJe9U55YpSQ0ae8qmFZ96w4GIY0HGU2FZm9KdNzleMLsPsPtdtF
Qxuycgjgz0z8iGqiwx68VeWJjSNNnBvs+0iuykc9us1sD70m0x7Ykvj1diZ9KoOW
ExvUXCuaGqVeZtgol+cF6V6oq2HiAr1R1CRr+8qgfYQXUg16FLkMs+h2exTWLTVZ
CkDb5vpahXqjeI58Oj6BjuEkCDcMirPzCmPbcU5LXWbECzkJrfpuutoI/qBeYiB3
VL7+R8VSk8jNzyFmKEjqCEnVUVuEzulxsqrInU7FwChy0Pd8PHErBOJzljCxoXLO
+5+4iJPyy3AbxtlAVqvkLOkKaW/NwZe2ddcQ/1F037Qc+NS5AEJFVZdLWW5Ih+hH
Lm36dqXJQAPqqovygAnunDhcHJefqvIOMa1PRfq6za1mh/8u8P9Q/CUyhKWDWLDw
/IONAV/RllsNAc/1rTSIDwz+/WQQqHFAVpIqycztEeE5TzV4aztHPJKZ6ewRWHwM
QqlHhhevAGDX/bu7C6E+N3BziJUa0wS0eo6NcH6xscrjDAVR6fv2sdIwNI/5HJYr
xirXq/zw+FEUbeBpBF9cF1t9Qn+L/omJczTvBlbLxzzsgQ4jnuONRwH/rk4E+2XQ
5wSvP21EVClnFBHeoxWm1zx7/nQUvoa2swhftH/Z4XLx14VtH9bYrO0D32ULsbu5
/JmOnvifMSC4vkYyZgrgfO0P1EwzBKC6YuEWamNBtaNanwz5QTlchoRLlvWivDV6
gCDKgqKrN4ciS1f39VnDR3pG1dRmCz+pQGypns93/whONKGAGfpc3ACl5Za/XyDN
bxEVrzVwiRuFmNxTg4chrnty2vR6rMBz4FYyohNMt3My1fdwpzfOcog2xJF5aImV
/H3/GpBMmU0LAPqHQUsXoR1IXYKts0r3cDMREC/SUwOCBFycmhk30VFFtBLHCs0C
S+tfPVjWDnKjZ4QIP74lUuvkznmduK0Qbmq54Cp5oVFboeKdHOpcF4ET+tkrXh1N
YrM7fR85R+440NxCZL0HQfLmQW9YqeGbZU3NH/ujyeTLvW/3AI8aZF4gUDJxO2zf
DmL681hwK1d8jH+JjXC0mI8S0vJEWeEYD8WVfffq58LEJ8SjleFNMtRJKq0IG0pr
x2GqGpz9ZeoqyaaJ4Mn2eDbIzRTdQUA1OsNEXeiBLEoF0HTNDws7j7ddIZ+3iDJ3
X08SnKdIqI8HWVyjPk/kDN0g+ycXwbjKgwTnsZZHs5hz1CDvxgdoilfiI7/n2Of9
slHQGwNZnMuTMDN/3wFJKfKl5OQJKou1PHGLuqVL8n07sPdq6bDtAmiyYxqLkmQW
J48vk0zrglK0c7Ss9M/1f+jsZf79blBJXn+0Z6a5fkkZuBsivUJ777vEIC7QIQB4
BfmCDmNQu0FHhg66n6HaVy/FcaHFIMfzeyxOb+LROcRXRY6cM22/Glohif7lf7Sz
xnnkVDPeJCUuN6MRXxFqUA5xFHfSL9pguvcMJ0AGeJVRQAu2mh72OauA2YyWo5pf
fXHCLqy1wqzhtR9xpr6BKwTubhJbb06pC8hHwGxlAwxOsMwD7+EPrMrRUs6BRrQH
HzPlIx5muNvYD6gjZZESAYXu58YomrjE/q3C2F+0YEiQ1bVadAbF+EtzJ21FSc+R
aW9DWk2AP9UjATAENZlnFneP0ikt9ylzmcevwO73GTFK/RVeWLf6kzEBONC3oq/4
+4+6gaKZkyxWfIcj9ZHsNtdn0yDZD2vGH8e8IE9w5MB4eQRhK8o8MjxqWKkLJCIY
EnXMMFtotyv3+XO4jPsvtk81+TlH3/Zruyv0EcujqFCRAG4eWTMrWIHyYVaOn5Ms
w2WN6i1/jZpI6Yd97ve6sJMysvBP5PMrjtq9nLqKVpWHGB6Os/oBWl2giruO7R9K
KbWit1EXB8+pRap8FPfVW/Z5VgPEhQwwjvpXjRwqrLA8M5peIMsfKLEIGPgeUPgd
F8EyP6l6GN98T08gUc0aDTfdLRHQjWz+ynG/3hz1t0UUZ2d/4jDrl2C/9yeyIdva
7rk6gUF3QS4q8o+E+sJxD57u920u73nSwNaKJtkeY0TzSeyGUqNHsxR0IfUyVpyV
kXyP+yprtyIcBgVQFuZ8OL1n6Hd2fvgEKNuV8NR5dulSDYZf4DD2gmyTpTUdoYiO
w0dG7ORzamtAj+jYyEUnjtNcazkbGMODJS9ssdhRwHAlgVN7n0FK8+O5UuVQRytL
Dys6Gc38YJPPQCH1X1DS4h9TwOofqeahg5KkyqZzzFi8kW7H++iwjS+7aGLa+T7y
hg6GfENz+Z4FoGZrQt+qlgc5SfyCciCORX+ivizs/XDa5i6/Yg0uYPqeNSskNB7t
Gru/oloTCBtxV8zqmHahkxc6m4WMdjj+Ga9w+d7Dmndroe/PoaiZSLAdWySI5i0P
o0CIJTGA5aeIpuQ5Mw7cxmVt3eM9jdBK6+N1+pzIrEUc5aQMIYpuc/KVfyPcLzr2
Qw4qFcvN/2LxS5kKcmy/Nc52xHqWEupoYHxs/pDRB5VVgR991Z5jOi4fStys0nMS
r8wmrQuManxO40+mFZjKsPLUeB7FRGLHzZVXw1IfTtThPFWjCtKFJoPqSxEe+9bH
qxpaCfNSjYltUn2Zkr6qYZn/NaUBSYl3y9sRyfgH6+yXny18+eBktc1swNksgXhG
ttut0YkgzuJiHPhSowa7SwjMwCnRnJCuwDgX/GDHoy8HktwFNJZ2HfT+od+XA9o2
yI8dUrpgq4yw1C22bymqeY+x1ShOikRLKZaPij5kiQQ29N6OB1AllvWXBmaOp119
g6BCwwZTbQz8ny8OyVd1cqd47x36Sm+HfV+yDT/LpdZQp1dCnHr1hgIA3DVGFGnW
wmgNiqCINXdim7HFwSonfo6CQ00BB33lBoFkManIyqMrNuPh7yq+Wns53xvZat+y
KqCvW8hhh8mXDm0BIRzTkQRm7sEpfY5fpAcf8sW055RkL/jaJqY6KhlzBnUnA6cc
fj7Wz/ZSR+dOuWYkL04Q04Tt3+QzbctKzhGYmLVn02HWXJ1BRAIoN/GhtA4m75wd
gFMTpH2bOO/RC4nVi+OpIu2U+gt6Kd9e4FAQwIHRYm3xUu8kZ7GjZaj+QFEtwYKZ
Vro0MHQSROj3XHMMvFGfRdI0Pp2ekxha/BjPSgFmLnoJxcQaaq0Tx2jsRV/DLU5e
bs1iy51FxFaojwEtY/JYuojTtObf7Qve+dMhvFue2gpufq+aOv4sLhaVojy6Qj5r
+p7EaV6zapWtFPtb9mZnPcPhidrmOSRox1kpU5QMve76mjtWowEIM4EM5KDm7RUW
6RRRCOTf+74td4Mmz9Un6wPMjleNKo1W4DDcW1ne0kiimeQ+GwWCrDP9P7OYtVaa
D0VURx7rKDU4YCqQjfoLcea27JZfhRStZkomu5k7vxNDx12QI+jEMeOWZ+Z9f9Jj
DOh+beGEZG9r/yJs2npNyed6nX3lECzMnsabkCxnGlb1hJY9uHFLrdTG7ZVmId/Z
FpOGp4288QOj39N7uSVWSZjUxOMUse+HpuykEoHddoYDJcSnNmCHe8GRPeKrvu/v
rCjvMmP5qyAS3lIICdTWsShK57i32vbixY6z2f/i/8NfQo35cfkxHg3CE7XVGIh1
3RtrRPkC3U8Hi/fd3Fl+4WFNzf7X5rC/7ZO58oTQeWeUDFoDHFYi9bl3wgGsylba
SQaOrisfug7ciiGkj1VvOWces8gLEMULc6KRqkjEVWNfSqlT2cWjXKzM+9a3OW0r
0LBmRF2KKZ1Ib+nYeX72tMLbjkSuE97uZl5Tn8si4uJPnPWD2+9rgTpCwMhAaThO
uH3gNFslp7JzTH+ecW24x5ObSQgJxzxVyVIO4Y0s3mSH2vJUsBW7aM/AlBNaLpu4
GkseviC/9BlyEHSJtDJ4y3z9U51X3wtt20yWL9nNtk/7IddvJBcWUkfKddoWdeht
mXAu1WLTiNkIPrq8Q2Do90laa9SqBTLUqRE0coRBfKeSyY9G7mVGmSE9fIN3l/+A
e1nzGPuT35G1nkzDRy5O0DlqDTvkxnux+Gi4IA79IeIjk9G7MnGTAIxrqL4e+20f
7gQ6iAyhd9w67v9WfZlxIvKNrBT2PSkQHno6u8578efKY3mOR1Vge58lVwRdphKW
2wjv8TApVOWKH/Fhe4P7lQyvrhaS9KKvISrl1UKE6yjm05a1Fl0BFUkql+draFnH
kXQeP+AVZ0cXRKDLK74vtl2ftSx6CD3860dysJnakRiShZN+yL98Y4tHTQ5BpT2N
Zv+ATmkAfzsJqQ8PzMVVu1PPtGDosCP63j4DjaOa6TG2IMkY0yNdrXv1Tt3UN+Fj
GLCOZcLWPiUBUaYocXsiWKEE/Y7OmHfn9YYB5q+JiX3x5GakfJeWPEYh3klgqNrW
Jrj7Lax06FgMRnFd6PVs5PaSodDQZkgn7C22DF65VKKX5b2gqrmHVgTmLw9Z0ubL
iyM3iKjfTqPzel86cyqvr+YS04s/0ik5S9a//ikVJW4N0HyIFEsKwNRGsLZ23S7Q
iS0FfUFpsvvmQsu3ZZar/c9Sf4xdHiCNi+XHgtsddvMrf1An57A0RtS/vqeW/LUY
AjodraX/F+FYX8i+NFbUJLWxFWzUW+TdHTe8I/7Lmi1KubF9eoHgMv3xbbtC0h/h
r9MapsWqzjY99mxSNBEcRrbKmkBnfG+lTy5+6zU2sMOcuNvLQ79xcOVykEpTBiWy
tn4mPyoFx1vihuZ+pdAZIGjq1cJDQyaXEyG3B24Sm5BG+a+1szCqQdRv9krXCKMr
wHWOCLX+mUhVVyqFk/AgOlhTYjL1+L7x6yMvpVwntY4qVjaMrsLGoqbhEdeJOAfu
xfsREFjoaMlGaa48JeJU5D/boMaSQ0PUOOxwK4FA3rViDduy/YeMw/hVsCN48dYI
plZydwqR7PBRR3Zqr0bMEeuiHk8lgQXhp1vFL8YnQlP1pRxgseVq6brROjoR2ckN
RYAgsHwBo31so7xiSjwdTIozAzFAe5wTisRHuoQnb+TP4JuIbOTYnTbu0DbQIyjc
/nTqNKO1BIJrYAAdLrYX38O+37mLW4fJwwig9X0aIFpUIbL1/4UvafORsNlHBEvI
aZCT56vBnhgslYm1l/A0lC9eUX+JBuXpWC2j+z5qViNGhVHyI+8lDLhDXlpReoAT
OkpNQ5hpk8jwOap9UQtIvXCGTyORYw33z4XcXeWFZKpTZRhvLjgp+xIHwztsP3JE
piMtQpTGsejmABl/USPhIlS3Iok0XLNINsjWfdeZuzOa+lcqD4nJcIvkmQBRx9Wp
sQ1Yy25R9kYV61QPoHT4WIbdt3J6IltXayf39dsaDqFM9pwjrLlyXAOQlDd53sRL
bWJbk7zZIL48hm1JQeyd8X34C0+JkVnUMCr2hC47MRmlh8EjZ5s13plws+D1ybH6
RiyOu+PPkD5/8PUEFTmGbdXk1bR+3gHEud4nvzfRtn3UEpDJfE7SArXBrjo+dp39
uO6X1ibfLJKUgrVomgm+aKeA809UD7SnQ9BWKoFGfPpngOIcT4nt3rYVuzhkv0Qz
bJz9HquAO4jG/YznFh4y3iVXuvCe/li5vbCdOa8+uknqACO7hF4mk4vHk8DB1rp+
DkEpPEKYbYHbtqb5d7YIcbZgQO8VwQqYfv75H1Y9MRKtFhENnY7WcgGIDneUMwj8
MWnn6ExITfUKOiIXtgDgnuOmXy5tIodl4ZE68TYPVIsMDBI5pZmay/jvOFjX1U0f
dXFwJWV8MhkVFuMzMEi0F6hvyykM4/J/Hr3Jy0Btu2tn+0d4rp65w/L0RcEGAdNz
8I/g77xUrmwtRj4wASZJWvEJxn4tcn0bhDVM8nXm1UAxEc9N37DO10HROuqMMwaj
u6rcCS+PT1gEoRJCDBWU9BPtN+nsfoGjIIrQ4pfTTg9x5OhHBYMEV6cvlFUiM6jU
Cd365dXeTnMvSepUKb125TzmJvSO1El4m5UdWMNiWzQBqehmRG1xRn5lQhVNu8gj
savALBBQTtQEu14yWbyt2PfIiAuTVUpWnawQGSFBq3za9CYXvnH/eEqjNWVLBH2p
38Tcfg4sfeiwWWp2yvGVCziiLSJ7nzK0zFEwVN+vDXyzSYeP1ON37iMCxxUgHT0s
rBzoGzoHCeJ+2lpfR4CtS+sLQXdn47IMnXjzeJGQ15a6MBf2BPPp2li52QbOop2Q
QgtKjJYWSwEnvVqB/rpKcAre+oKK7fZRbq/SRX+awYnYSydDuuOOsCYc+POX0Kfb
dUbKrBRC/IA5bZCh3L0/6qRQLf9IQw20PgFDlnXuOqTSAyWxSGfFAIUHYUa0V+vI
fV6+gKuLNKSW3R2n0knQg/AWO0x2TSkMci5N3vRRZXR8nUyK64gleOkCAXAlLlIb
rCft4yYBBrEPiEevZm4FRpnMTulAs6iI2M2W/L2ucROr6eZhtzXRe7w/+Sc09kmA
U2wyFcDcaCIF3bYRD/U6YOk+GIyvIrXDGDnlAa2Y4K2HuDJpEgEitXo/qEF0NdOj
KJ2pkl2PvHBp9en3fZuoJiUKmYJPto5FolPeNvc9CU8Pz6An7qk6FTHux1vM/My1
K4+U4xvTO/+QwMZRZ8kUEPNM/K10jKOdQ5xSmSObdzxP41c9AyJfiMY2zcvelieW
HLa+G/8OFGd8PwzKNJtO4Ud8A+M5ODH7j3JbZ+WRhMoTqiknKoL+EzJLjBnAbuUj
TE7TbZt7bbhVOpE1DTT4iwVljA7fGu2XYgWQBTFI2NnRUmQzNlakXAE8RXVJIWL9
2KgUDHPBfzlHmDuHPdW6VChYJlGf3C+zA+U4N4uezJ8lkR6z1Dfhmt6PULBuhmC9
n9n+zZSk/8d3n51X9z3xuxV2SEYjfzSWJKExLtceo2SEYbxQaX7aEhXtdESo3/Je
gbLG82HZ1lLcYs9XRT1pQlXrU+GKYSg+FfxycDj1vDLhqFmogtjpX5gvzcv7mgcu
Dk9QtRrptu1fRknjpt4oY3S9b+v4JCNp2iZEVvGKvErXrYuSM7+yyeYFTjUq6IHi
W4uTM9E2j1O9I3qZOoSs9PLjcSodkhbBUZBIn1iay4CyPNHpKj9lEX5aUiwBUJgP
c9tLZe1XgOzP9pHN5P6V9UJgthAp2d67SxfwfIShQS3irSlCyKTMSjVwkPT76CJA
7lFodaBhMEeaPGHBdzn5W7Ub2+2rnNr/L41b/gt1gIYVYn/NZw5Dv99gZwhziQ7t
uCGC6GQYbzZtRZ98CY+iOg3HA0BIRbmOiKGuOyRxgd9U2RCS2XW7bsRTwTGb1NM2
QQJG2KDwi8N5jnJhRFhXGWadJG8WNnJ1h08zFCVTpheTL/LVu3CQjLXBlUc9lqzF
utTa7AHP6GsNx3KbxTAvsGRKGcVX7A9gKIR2oAITzym1M9ogFRZRx0SQH+9UKLF/
KF+IF3HjGxJoZw7zObFrxoqgtfz5vqc8EIMbBy43xhhb+GfDRJxmMqDNS3GBQN4Y
ICNsHy3oYUH/SiZnumOLZxv9f24Yw0m2GZ+UQoW0/dqyUb/vj2oO6oB2zfnpJKtl
DRvJX1o4uB+XbiZL+vREzzkVjFwH9WSZos6zzJznwkrYclyjLhNDj23rFADskHu7
cJYqugrNANxZ7e4ZRZi9oI7kv/7Iu/+8smjVmyOljyJyrev0V+MjtqvfeQ7UE0Wq
LnBLl0AxNKVz71T7SS/F58hTdo7IrrtB/fx8XWuEKiv2o3ZzEg7DI8FgGVZcGdjA
Rt05ArnN3/aXAIvbfbDIC1pCFLiCeMaFdvbmLkV0nmZ7AkjEuc76lAdxYnmak8Kt
0zrSXo0rhlQs+W9B8GcL65h5DK4806E/5pHynj1E6tfREKFug17GJ4gbKv+jJIws
haPLRWa0/vRh3GfPOrccYciv3EJVjKMVObUzANjEA7i7ZCmkJXtEOWOCctlqmc94
VDxUI5MBsDa+j9Io7qOvXqaBRiFRR3Y7fYpkJ9OyhhpmAzbV68HcqtrCToSdU9Sz
0GQ5/ozpfBJNUHFGMz4FvRq2g+t/bRT/sDcF+gIf1dA4i+9Kmf6WydK/OlqfyZaN
aj372WUVQ+uS0cad048ChRIM4UKRFi2AjPW/SzCsw7dApOLgwVimDqQl/tT3kZng
XUKyf+xKIJx1xVPx6csD4SWPw9vNGbvnWFP9an/dLJbDozeUEPrl1eCsiVZsmJ3q
9qHlyPPu/1OR0oF6MPGCN9xq4yB38exeaU5CemcqDiw0K+V8ePxRWvpommDLzp6l
pOwCb5dVjMujgOAZZWfscGLayIPvAr+kzfuqcHVU4yuI6KZTmhac0apWzVDWSgjU
+vxFTIm4vgsn1bzdxMmuMy6eWim7QpXcGcklZQiYhs8iGZZNOR6E8S2JYNY50Z3t
o0JUQr/K1mgTNRr9EneNTBEEOAOoLl/CeE0a0tw+w/EHcCukoHKHdVIxQ7OCOq53
gzHXVFsopocKlE1Ke/VsuI8s/O0GEET7F5k5nQXUEzUH8/HxMZSL6L7CXsRNuHGT
LOLlw0JTSLgrlP+zyokm1qOsfPLSXiLjXu11oToIkE1j9DX9/SNyBFsNtpMs6Jyd
7iRKaSGCPLeyoUUij80NBRy1VbggOCUFX2FKKn9kw9GYFn5IWEhMa8XiamAK1u6m
Cr7ud+ueTUrui1O+rsTdSZUsQHoyGLZw61fZp3wIVtq4N4FGm5+XUETBd50rkizb
li3oVVmo//FGvmzi5032gm7PS5NHFyTNhy3Fdp0eEQ7X1pPlJIf6apHLho6tUrB1
8dskv7CoL+nr/N5YCJYF4aePx9S2aWdYQ4T+OhaftfD2fDsCgszDNkFcbiMARhKA
kx5w27xi+gUzSqwLJqjOqeZB3MUm2T37K49GGc+67cHcIxAx7vLiMxzy5BqFJbfJ
pTuSW9W0FkrmtxZkOp3j8p5UA3keqJb+DzP/BvYeI6ejkD2Z3lPtpF+rouiC6zM4
4LyBPUufFSfBCBydv8/VBfGy2fK+uo/nfDxxgLwzagqcIDy9Rc4+X9spHU+S8lGR
Zll6h1pjHDOBTO69Ea/T1aE6mmyRTFWU9UuYQrDMQHtsOpLxwQ47ajgRJ70bFUei
dcx8gX9HtiKivSdYzHCUeSi578+CvFt9KbSrnUd2z7O5AnHYJjd3qOKOStc+MDRz
Exvw0bkq7XfNWPoRdAIhhGyZDG+W13iMYs2fKB/tWd6UTdLGjSWTLhMXMoljp/qG
cG/JtcJNfWW7gJuokdkozotMQs3jjlnXsnBvcArdSta65bLBjIJRixPI2AlZ3COG
brJ5EpYjo1cZFCWiIDvDib/CzCfPjKnVFYQz6iOfYVRNanF+xJPYpyiqoFVlC+49
5XdQr91HCDSHKRQGxsLoW4/VAcApOiYO1raXuTYPhbuCYa6A8Wc8ojCK/dCgRPTs
4CuPLdPipLKieT4QkjGC89iehn5kqKecxYoiab/rTMMIvzfbL2qJ6ZtogHoNc5so
wsA+20HU0FBIsCXxb1TTgHcijgdwZ0v0qd+QtntlIfzUW40HUxrpSZGjyUoa9rIM
F8cpmPbBwapr86WRbUmIRSFrXaKhfJxUa2Rb1ShfxuBZUUe/6az54j9sN7cZViBh
Dqe+xsSmcNF8qyW8Jk06kXJYaFOkDQb+JVflg0nLC8qbXQ0lb3w9ok8WpWaY/Cf4
bw1ml7Kp0+k/DuNBBMnU/eVy2nkOFxFT5qYDmYZnG6Y192hNiT9Yh+4fMqx7Mnkw
8fS23Z+gYLKnMcAmif2xpFAkHio+NWvp933kUy3qYrD7lT2rnVVzgmYfG+HWPMhr
ddr7jw3OVMjBBnS0EJZxfBrciqCMLzOkkwRm8xcdBVXwTXcTxqOJZ/n+hDVsTNZx
GevZtmVURqu8zXeMFCK2SYFiiVKb16ylKPabNvBoDOTb0JnOzdqQaH8jBcHTj/8l
SCRjTKaurT053g0dLKlpn8VxNNlypUuBVoSw2GNerkkGCuPJ+iimyIuwSDyVRXYL
o/7vDMLe+Hk+HWXLsgw8iKjuAr1y/Rvb/HFeNY0R2kx5Svif7wUJBAxjFekwJUJP
RABB/WnHSoHRAzcJ8IMjoBH2gUS8chNJwQup/8uwL3UtU9nL4C0jVzrDyoRml05w
FWXhDZh5ny1+R2GDxRJv9jvskMAOws7PHoyS2pecWsnlzfN86ExU2yd68hac6iHC
AtuO8Ue7UkuSk/YhNQzGW3ub/DtdVBPyF7tQYDWDZTr0xq5DGBwLOFKiEG8dF0S4
ey+njJTCkWw6RRSPkxZuiUz2iRXaZUjtLtZhRt620SBv41aishI04nDBmqNWQlcq
ps65jOFkzCbXcr6Zze8ZrJPclyQZBHSyliLRlQSJmbiTEPyrhKLzZCEl8vqzjBvU
9APc4ba907BfhDzvOK1tjR/jXbtO0tnlPKC29vMadWVjiW4x2reNH2O8yCIW2Doq
bnzyo7UW0u1CubeBttJ88XQpxpt5ZoGGadizqjDSFx4ZPyIIyS+OjeZ8CMiBKpz4
3mxuEbh+JSW97IJ6Kg6G0mfNMkjDfNAuaus6lKawkGuUoWYKPWxH0oer4ofTfxpT
XX+ArAsynEQi2HDkVjM0N8lN2QPBDX60rUJ8lCOAznZgIcwFcDHzvZDWp2EJkUNu
n6xGAfRgMVtu05HQhZlqZOntEVnn5utYhLGKI3TXfaEbYm3snRMwMAzt4KDQ4jdy
8LTtBYNvw2o6hzGoES4GlMZftx75MaGpUAlawOGmXmEO0arMcuXVKjCiFgO0+zgg
nWOirRwT20FXF+QWWsyBHmw2yR2xhzvSux0wguxXE4yX1S6gbP5SrR25kvo7ywMs
b87I92BrnyGBENrBid32k6NvAUnrAZ0c0kjTHB91lFrjHtVvahDBM29+L/5Erm3e
ahwhjoU6M+G+F5Nbhmnm8qhvrxS4K15b2P1fuhxVY0dmoQYgcmIrYfieVJ57du1Z
xE1eJ6dRpGF9jG0MSGZGiH9Ld+FyhLKv2zkNij+umvMP+cq+OzVofI3w5e7K9Htq
Gk+L1QtUB+rrNJ3QbIAU15zxevLHb+3maZ6Un6n1RdU5oklxrKc3/ySa7vssQHm3
rdam71sBtpGxMEpnC4ocpG8IwrhQhJouPpo1MS02W6N2f/U97oPQyet+UWuMwrLD
SP/yvp9Bv155akOUfGCA9gki91jV4fGNDbo4jCuAlW+z0FjaqkvoAZJSVQyATwep
7NfO3SoNpXHr50ECcVkcgdsoFsfqKTCCL/faGPCgqRYThx72GMSu6ugw4nAZoRj2
/aNBfqPWfGO2RaFdrD5EY1ji5M+CBOawG7Lr8j6Ddr5rOPdDh8fw/faDScrAhicd
Yi82gWNPuEN8dBN/AtJ1k17fHiRiCa3rqVI5InKPotv+28nrSHbeICqttoV7H1jN
AnFPiPTang7LaEjc6u96S480phO5ridnJlxbIf0dgWrkXX7sFUT6UgqEHluGuw5y
j6IwH9X8ZjiuQUiHZlNRc/r5PlXFD7ZRyjXKUdvqt3Ciyf3SXoT0wH62X6uNJ5kB
dLNiA0Cad5HFnKY9C+5YhisR9Yh2ecI2Xp2XmcnuAMg2A5eE1/DxNEV45VymM6WB
I4B0stHjMcyLmg3TrZcF2oc90CcnAIzlzyjFoosBBdJ04XN3jAyy5fz1UkTBZslM
L41YBg+BdzNRzE2I4kqzWu8TfXWu4JSWdG1MPSaXFsqFgmJwGeRgQmSeUHr7BP1i
nfC4PATARdaXNwt6OZrpJbiZsD1YvByRMDcUDGDkmDA9iZLwuzbPoYkWlC8Q8gS3
U5z/qq8EsIdttIvrTAYViSZ6D3mASS3fh7koOAwvxyxFeZc4RzfMST0D6fpe3n07
VZwSTeWnJO7DiOqSWhLLt3NmQ0Wo4mhEzsmhHFiO7yQ2OrCmm94qv4dmZgjg4M96
vG/NJsnPg8H1Eww5SlyB+IAzUvrOHoI3lAvyUaylNfhgJcIwdKq+7eQ5rN/KAbMV
Ej5zH8bQOJDlIdEhLaCNwUuvuvdWBbbcgQLERqd5n0oL9eNXsNpkGQT3pDKTlK9/
51tsWK6nn2oDDiUjB3I5oYbYCII5JS1vrHumou8oUKgs+CmOFUKxs7loYWsFE0Er
ZrhBt4nXjA0pSRxSgQ7QJr2EfPP+i++Jg582dxvpzIt60Lckv0rmpMrg6SgaQdAV
Twf09nUFBbSLPYxI70zJUFWgc/ZMUv+MgMiimqcoSP19d1non2IJXLQ95tB4T7P0
FXugrF3yCpGwuKOZ1PobVVVkMiM5B4B/eKPIj5Wt1Hi257PSro3ZvA1gTF4alSKJ
MzOsA0yOirZXRccZmoVJaFgJaQZxXxYx8Kd0eIJZaaqVR+EU6QGPH8zUsQ2WiCs6
AtJFFGqswJbdkl8u29wmscO8r/pHItV5CUSbvTHKwUvtA75XBe8xSLg5k0+gusov
wEkVB4Pg4OKvlEIo7yhoBOpYlpGequ9SnxJBDPIa488DxkF/9tgDEa6LFKaGqwLB
NOZiyZTg9WCTM9CKYT/fMWCfqyNmw9iPIpzBx4W1t6zlQqBnJjoUGYVE2FMQ3zUb
YE9fIFVvoWmhMS3VnQ+6hxSc0FmywpWoNlgKHYy7N6GeIKfSA1q1OiysI+VlVBv7
UbYlMBtnN3SEtCrInIxHC5qh+hM9KfD9WxbDemQHmY4ysODzknzLdieP6XpImvSN
0USfzGfRyUqpygV9+SyecMui6e9cIYp/Lr2Oqvnm/I67iB8QWCZtOmhMrCXw1bIF
lf9lNA6O0sQuSmMUFJaZcD5zd1AS2VaYnNUP2xsdT31YZRKUdnYFfV1RewKIpB1M
9bhlleQPX+VzwM02HHmKO3Yo1w3eb4XsR4j3wiAy2eoCHnbiF3zZTFDEZZnA9ldP
TFB7KSll9dd6Xe7jLCtqTiDIIIhxudzIGks9kTIQQopvOUhsT5PshUtICgAGwo/f
c04rVhZgXXpBy45B6b1tpIV05SsVtsa5jSsaHkilLMNaRZZrPWLFAm4OPApKIyRZ
mqVdNcgD+j2Kf6TAtSIBujm32wjUZUEu2KKDIQ768XFuucK9MA+kVasppvOcLmEc
y8D3doT8yz6XNyDEJf3MpdDXAKIZ5BA0IRQjw9jFhl5hivH4JapISEb/aTvyzGuu
6xewT2mIJxUkDgsdvo0KKefzz7ylNrtdX8TbS1IFbG/gXST6jdld9qXge1aLBo1B
KC+G/5P+IlR3fOVR1AgaACDsrEECn8kwlNRcA536+BVGPYitftoU5pTsShxDhOdL
e+DbiXgrNeDl5iJpUGE3cdliPfexWGxRMoCSS09NjzLsQYhFfJj0rLc6rRCDjLlh
nJ84LPC9/KTM5tOf7s7r7BX0hWpADJwRmmnYPKetGx3IYkcXu1yDsRp1S9mLxgJO
K7rOmHARgnf4rY6y2hg86l7PiAvI+BNeAxFdarjptxalDcWRK1TzGFJT4Fcqx1kB
hnWrr7+v/m6YOaKbsbAvzXRFc1Tt81cSONPeTxNzyRsFBPCsfgvBaIftrG337rh5
Su66QfljMJo5+iZohmuyHTP6pFfSDPibDoA0Tiw0hvwCrWA68Cvr1k2k1pawKbZ9
E11e9s1J3i27RdFkyrVQceawCVBzl3StKdi0i5ai6WjtXrDw24SFwnWOJzwka+oW
qBA3M26G37i8+ypCweI96Wbraillo2/vBC/JNycMlVOazc/szJvv9VuWF/tqtEP5
uHZ2ThH02XLqKxviVQw+bgB4patDroVn1Cfv+chC+x6B6kAkwstpw6xUu5sgj0DL
zR+lN5MF+/dAgFMMLbY+Q2v4aubptq1rW8Rk51t3wLxoXKKz59Fig+EnN2GLtAeT
dQziBtyLxA5KUcVN4168pZXTzU3Xnlx71Eh6OOFOBfWk7jH8r4u9m691wYqjXM3x
lg8/1adzigkKs52Yazxvj1A+6j2hW3ZEmLpFvIeAQ4eLDScReVtTsGGZqpnM+3ll
1CITom2RYpjsNtc7eeRqfciLS4dNjoTEcgokX294WaXkYspVDgrCkENQuVGAzA6K
PJF78fUHhg/zSshpVMciXkxFagWelUkNxhYBCqnYxJqvNKP7ntmQ1EZfpdCDkWsU
E5Rd4L4CbNl4u7rJgsTdwuG9Nuz8beTpUsJDlJ2hU6w8M2XjN7zdonbFTV83ScUU
et9xN53XW5xcVM6d+BBwgRRt+Ppjx9h5PFDqDo7lBZ9+oRkuIGRyCf8Rjn+TPe2D
clFGwt/6+GQDGYIVhQgkZEzB8RmwxVyRBKlNpSCUMyox/ZHD3Z5/lQenqmxbWpUd
Ur7cWE1jRh7cM7C3z0o3kMdTqiAFhnKK3Of51YqcdDg7cIxLCS3phTTuKWQ3FfTp
F8IUNhgyPQ5mvqjdRD3xJcH+gOGy6clZCStO4Tv/IAuR/bNYDouVjUjadjLYEVj9
TpBJbxa0m9Cm6+jFUoVD+K58VIHST9Y00P41OADYXQHgLDRaswjvlGv5Fma/E7fO
OWikwEof8AScs/ET5k5xtLfR7VcIV96ffZgNaAlyy5aUpONZC/qJdPtfE6cucbY3
absrHxcUjHDmYY1/gt6i/syhCW0bFLdiTrsxxDaBXLt5YbH+FmmjoMOqMA33geYA
gYjY3PknBAwN1D4CoAAkDOEONvNifWoJJWCA6gWAKOT9f/oIpfdC/7najt6m0WHn
UcmHmYebai67nLijBF76IGpfH1T9KIc963hZUiM+qOU+FipgKVSGoBWT+L7U2dcI
1qOSFw8KYfD3SzgbnhiQsD7VxCxKvnT9wUdHPHZ4AtmDhb5rw2WX8N7PQBWfYsW3
21hkfUu8RMdmQ9R4ibjI6mmf0LtNhh+aYVT5N/glIjCyXD7DNDLmf0slp6mafDW7
W/r41IxaY1thtzMtfhuLYxpfT7Iy6yuTnhojhaxN0672egldbeTHRJVJ0x2Rtgp3
P5ve9jVrKCOXDM3uMJbA8I9OH5iCtUqU6w7xR8IG8/CELbnX36hxI+s8dW01xCaC
I5imxWON+fi54mPYWuXmrsLCWVOVje/xz8OWS9sdpTP7yNeTqr1y4eN2StRScmXx
UX9/1gh6V91z+IHNn690aSTzn+m9iwJ8L2SBR5zXx9bMVRlmSYRM6cmkFkrtwlfe
6aT7Vkzgxn1r/Azpw+Y9O+t2euHOUKj4mstM8nnZzM8z4mfuRa3YfKw50/deSOZt
10EPOalF78dhcR3i4FlFlVnJk3Qf/P7j0XgOrap9aArCsQOb4ybfpBVV+GO1Y0za
HxJpTw9XABEWKKGL+8rV7uEilxnsKzOFznTm6xKhv5LR3gqdHWTgXn9H3THd7GDv
0GW1dknX26RP0XcCdzq6zESVBjC+LPnxsteg6dpAYFKoRg6Le7qBEpE95u4sAat7
HW7lzyIFWlziVSr/sbMBzR58dkYvDtUCBw6fIdTH7N4w9qjtSx4pB0oy9TAiqM8S
reOq74HZGAk9URhPYoMVFYdG804eraDVXP0OCUxfc0Xn/OxUsK1PgUY09c2kKUnu
gWOyrMcHM/tqiWytiH6HaeEjbvDC6V0Vco84ZJSQnCuIyaXehjMoEE93zxX2Rryx
q5nrhpzogk/WT3XtiAt+jCWirIz5WxGhk7fJ3SfAMi9MoGrZuhzDN3gz4TF0ePj5
9Qw5DUvUtyoSYU4oh4+sgyifzDuFxz2H9ZN7ZYF4YjcjI6MQzlRShUQnwjYyJ5mF
yUJNIWsq8OG4mnfbDt2x+cjO1zecOfhfFTGz6DaGkM6lROszTIqoh7G+WD+qJtfQ
KiTPGlkm69mkZkNdn7BjshlKf93DqWoOJRZXhho4QSnsmdla0zADoZdd6dv05GbQ
KrMlNUVBy/iqywMqi/5G4+ZpP9OpB7m6bAq4qu2izNLAp6iHvo0dLXsFmwMapHOQ
qd1vEcqpOmiXu9ZfAE4el0FXZgHwDnDy//0BX4AuAwqEZ5WboFM513zrE19cUn4W
sH/X0+RDG/T4fsniq1wuaSV/8seLHWhmkFVOC2c5GDKmRIdnwA6XGV/bX4DExL9i
JzRGvMhSTAKCIQMzGD5mbqIOGEhT3EZQq7TZQWx7C8OtkVZuK86VPnF3zC1mXbU6
iguQNPP35rlEb2IZvzIy9lgYSVZr/B421zfdb/fYuiiRVbogXSLr5WKN753bFKOK
juKXd39ICbEtsjETl91KUdRiXRFMY3uMIdwG8HF+dASM7vWENYMNhbRPGziSWcmS
BbhsAdDCEInkfvhDywihVTfZPuUi8l0bd6iXtrpbNkw05FhdS0NoOV9XU+tOK3jN
FOFxY92Z3K6aRUHDZmVXH4ilf1GjHjGIign9ZTxuC8UIHhfyOZ0JOgTMKgn95nCc
qJkMJjkbR7JQh1qHgIFFepHVKhbROCCv6zm8wYHmSaEv4ZaAW0mkaWxWwGuU/Tc8
sTK1xcQZNVOJk3AUWuaGk9QUmbhgx+yA6Webxj25OydkXe+QM6vNVT+Y+GRBQzW+
p4UdFlbzwsNqcyR4X91kd60JYzLplHlZ5rprhSmMCGpMH35Vyb4TVfTXp58WrqlV
i66EzKolj7HZaY2s8wIznnnfy4YwAV6GcXtacG2pyPnQwwRP2386/N/6u1grvdn9
rA47oOwb1qpBtBBTjaYIWFqVlh6fcgtWZRrYivvaK8YWe9JLjw0QTL5G4+oGY6mu
kKbPRxRjlLCzXIchrNFET4NrYIlEYGINra9qFJBv8uFh9/Jl7NYZeaRtqIM5dq+4
dGjiR/7obNwPIQTTZC9DTZOeqTE8ncsowUKvbTQblrggEtpwJnwD/pgTKkmkpi+C
pMdDRKgYXPkHnuiTaPcc28j2v9uWTC/TyOg60yuXq1vnvMw8oEV3xY6V17A/RF43
FfRbTzs5WRhQUMi5fJTX+xTzmzC3/B/zQW2+336/16zhcbEAKF7beLe0N2nigApI
FpPVXn/Pvui4dnrgcSIQPT6+BYpXfiaU3tMryDIpUeH4tP0/niPXSiVd6ygD9wVy
u9RpCxxHqB7Gid/GfVjes/ykR9NkAH7As0B2EqYy7VHvw8GiAMOIMh6mUL/oyzsw
vhna+JfO2nnEhQYg5avU6FSsIsnDU2tOqD/0NZf6otkfj3CBz99vK/IZVxKmcuoQ
44PTUHMGXzT4uCfhcoq8oJdAcF37ZjTMZjsFUUeRXzlnwpqxaMvxfZZv7apYZXj4
kvXdcmqVIaZlHeEMolXZS01K3lnTxA9qcZQONHmTzE/7hTMWoygQtInLyoW5FxFF
8X0jfHXH7Gdu3ykBToq3plRLh1sp50kx+DTceaDY2j14MLkS7Z23ZX4lRI0Pyrxz
gPPZ9rUW2F8gdz1DTqq7gyYOylzKce7lClTvrkFo+2mpc0H9N5Dl3TQvkEK9YIgx
CerebPM38KtT/yfhx4MIF9ORhNT5cTLOi8ElMXhH95lPN1lrUzEi+l0mnk0h2+E0
Jan4ihDh3JoUkOR5imO5J4667kaSQWJkzrweeK05K+QpmQjjRJr+hlA+xq8R1guD
k7af1hp/g3y2/vEtVmYxMS1sl2DNC2SYk7xtBZWsPwNns60HGE1dBNcSTw1Dq+Z9
h4/g8hpce5LrtJJC0XOy5kMHVrVVdPzxeIqvecwZjx+PbAlJxguVQ2++9W7WJwR8
I7poYIBkKxNwNH90Yzu/aUcEVq9h77XR4UrsSEKqRKSKE5XkyUa7p/cBBABL+fB9
uJWEFefgrG1Y1wKEgxgXtIMH2hdk6gosDsZI0LV8SV5R8AEQzl3mj8fvU3m00Fzw
pQzsjKSRYmlVqr0dHmRQxRtWVKpsZCOD0VdsqkXv3WBR1LfdRhLDYVwTfUOmZdBZ
8V5eosNMMeHVinyCaEJjK2NegEOEWq/dNk0+igi2Fm7ULEZ7tL7cL6payCxmaZUJ
Rb1kjj1CkfarXWSYCUuybxu6mqx7TQ5DodpztxyfOw9BJpx/juIHyamDI9wGjpkt
8aNzPKGkT8i9QKLaLS6ShXOHQzAtScAKj3z1tTZq4Hha9N3GVaQX7MVLs+gheXAv
IJ5cqJXU3F8nZ2/vU6cf0aA0au7jP3TLIFVUx8G+R+az+tdSdMSoeW1BT+fw5CtG
JjD0XBsb0Sx2P1U6yRtz/nRx3zay3C65YiGKkkTYEgofXHkUrUSfdgMskSpBuhYD
TpLDAPdjQrfzrPbRX9HdROx5YHdvSQdBTTS6Nnq2QcFKPf3MjR73Xw2Y1W5WEfFN
zCaWd9m4yGYxA5D/BzgwdogsbLTQFU+RuxprvB4AD+zHlIX4M2+wq9Hdf62ngxeZ
IfRrwX54l/FGJPCnSLf8EoD4uIwoAMNtXE6F/AY1QcLSmbYsBXWbdkzkwatSrFFQ
pQmxuL0wMpBuASZBPqMquEVzruBsJvFl3LD8gzVpzYsq8UVNtM1Gy+sthFkMxJ1R
h1Vmu397iND6r1zTrPOiy/HOO9r5MMo2AcIynQhb+9SpOyTo14ELZhkOr/ow3YJL
4kti08OnHo/oS4HSA5ImQAol0tJXxoI2HFQN5nTiG5s3uHfDUfwqmspFYiT7JnCY
UeZSZMsyYLOfoE/TYTgCWj1CL06T40ayM45aQh9z4IiaNFTaJ4i1TWoLQB29UQeb
bJATKrGzpDoux9UqNrAR3OB9EM11oIYREU07i4t5C4yRm4jSMCDukcF5vRmgQ4es
Z1WWynfKi54BRWXSGdLyQ1jKq6GglG6AyaZRnfHfQWwgxM5oKmniHCpCTO8X6qae
KJYoMFC+jFgbkyxd1bZAe0gDKAYb7RJkV98CjmC08JWjZO6kX+U00r4w73naft1r
Lj4VPdKfczy2cjkwvRSe3vm0pAYmWc7h8f3cSsewWQVN3YBQO6Gn0vlqD5A8C9W2
XDfX3K3UfkEyh9Rzm1B0lWXNwQ06QbW+Tfxv6UM/+Pfwaj7Bj3yuG/kuE/OfmqCb
aD8IvnVbfw8XM0o06JKnSb3HF7Ybi776+jXz3ZmzgaBs0yU2DZCrkjEmxmfQTFHx
JqIylLtwzXGybaJqJNrr2RhmUaO0DHYkUWXqnXLl00F4dgBuiv/2ZPyfe0nXYgxk
3j56Sp0Z97R8vfmJ6zgjmCmRkv3Wz+H5n8wZ/w2S3vuBQiRStwML7nG+qOXfGnXk
AgYsPqY0v5sLQpY6S3SqRBfe/KTn9cmfq4Zu4Pveg9BnIbN6m8iHZ9mxWPNyqUn1
J1p76nhIkW+64CLqW2eWXuKeUe8xp695okIcLB/y59EGo5A2bAWdpD6h/vSZHEpF
QKObz59bVdMPEbutmbClAO61NVtDLAG11bJ3wkA9z7YO6SKdpOsgJNB+ppM79uE2
6mRO8zNCNm0ftUw6GYEh5eKqxl/PWy+bvxxKrsT7pjmzx11unop7l5upJRpkhsuQ
XYzOV9hls0g1IHb8WAPpriAjFvnKaajmGMQtp6bCgMU5HHlZLaJE/m9F+yA6eKZd
pRNDsfDun6Glb5j80oiVYbnJvbHxRzzU3KjKxC1DHOLCD74tW8JH1KFfzFwtpFHr
UdsmvQiwPXb+5QmPX2ATAE8+qBE0ILy8zTBG06FP11Ur6qtq3p2qOUpmX/MUl/zg
deCc9zAi4JPuQmQrm0AG9E4rgJYBCs5NsB8JcaivVQs22sh6NlP8OFJ8CFBwK56e
pVFPsxnqMQO8Y021CKbthFr2OXrkbaDUrji2bKampgETkgSWy9hR/BpapC3KRFA9
2s7CakfNJ/LtnpHMDNPNgHxTD06G1nb6+u7/xRphxT/CS7QFDBWSsnlUMjxfXKI4
bbw9dMZ33PfJrHwCc/hxPPKwPb4ZFlzA+8AyiGAeIt9PXM21sGxjFeLoxjm+oWP8
imv1jm+pFp4zy5nl0Wct1oFuwZEhHt0PDheRK5WJMTTCmc1VWRymVysutuVkBIDL
aJPsEhKt5opK+HCTpbKauUMnKD81mIdxAL5fFCyku70fMD2UjR0eyzDnIpzid+E3
pdWNNgz6DLNqfB/SV6Kq9BsxyVRhXimoJyznD0kZ1LHBhvV7zoRwadgVV2zwMBIQ
yzmszRhNFySyhBbytPLZ/+IyIiiTorBTQuea1+0dC4igh3E4IHcwaZeH6IszB8/+
Gp2Tea3POHavjvY61IhTOngknSAAf0+IiSA4I5o1UKT3LTjwm1HXKi9Acm5xDy9X
CPSQ5bGCz9CFMXeZUrGN8fBY9r+GGN76WB9GtPM1lSq2SsAUuwkObWYwcnd+8ITB
7DYoQKOX3Buar9fdZrhDHNcduLvmuGU4T7cnFlUfvHuCpbHo2KURlwEHD/yaflB2
xrLs+YBbvmSb/PDb3bhlohlZ3MAkpnGVFbi28ki3vbdWZ4AQdMOPLPyRTohx2GlI
NBMSF/UOXBKPs8jArLQt9qmMuFLT2vKTPxj5yLT4qLoiBlpETTTGvE0PDRtsetiB
efQ7JKWNcDfvIJoXEZdU8E1ONitGyhFHq9JTxNchXVyUIgJCVTtPxFA9Lkax6wf4
BiE+786AwU0h8pOil3pnwE2WrXDqkUwR5MSmWVmh9zuNmLCI8K5oUwMDX3HE7yAe
7WlKxIhBhWHOSvbnsmT9mwejfX2DrR4p8gYY4nK6sgPWFXlWPY3g/e5y1dLTV7P9
8BNcUsTn7iU02W1PkvKmGN/3PFePvhKPyX0J6PhmakozlWNcTaTkUmdSnBKUiEXv
mf8UhisK8NNPbFvlaLSnFluq4pa6LyHRjdjDmUMDzpwCoithYGBHHtUxKwBOf15D
gaOCp3Yg8wunCcg9dNDQwbLlVVa8b7IfQIobD/E96kueZYHlNnoGDHqXCqh6IbYU
z0NC+eeYtaK5An4dcTGU4vrgi4qI+0K0lIaCs9I52E3rdDVJKNOwx6LbYGid6XZN
VQ6BUHrmznR5+QjRoyeJk/+Nbq/2PFNUyyhKzaiWHoKHeuAF9X6MfpPmdDIZtqng
BTfhH/svSG5KRquthRPrlGIxPs0VW1dehru31/YmX2jbC+jT2zrD5M3zNDjBoOmD
FrCaZbkoLi5rosN/xXWspm7Ksdjt3R+oVnaSm+Ep9TXy8lhp9JeZFuo037sngOg3
B1r3lx7NzRC3q4PDZn6ihJf/gQcwgldRfn4/ZpHRqcxVKZEBaf9aigJSUIEOUKDE
6HK9nxvce4IEGVsbHO6u/1FFc1OIRDMTc6BrLV+wBpcY4NospiPvGG7xihqT4oZE
qzGTMBucFtrO2t21f6HL6UuPr42BcE88Hj8kYJokTmaG6lSHK2+AAG9GE8Hcab9J
fB2tnita4LOciu4CoJFa0AQQvbaqHtYRSIajPcY/G0ypHm9iAbuU7SMZnORIdW9g
85XcPXn63C0IyJIRU6btGxowUGVWNCtvXtA6V6md2qXrBr0ItQ4p3hp5UGqAfhHD
ByXoWmY4J2R1SGaiOEvrK36guHgniMosKl11Z+vOKcfPslzkLOGaIJSQYEVBKmSW
4xGaC57Fjve12M7JGd8CODr4+NEUbx6phwGZF1abhUXlMqujf7TGvZSqtrqBDY6y
amiSyDvNib1hStSUm8YmXVb9cb6TGBo9371e8Pk+WSCVcmSILAypvYlU5n7VILoP
Ir7nbyKrubKJz/8m2o+ljoq+tOykqtuGO+D1cVUDxionTRIusamXdx6QhdUnMGjn
7nvQemVJS3ucqUcbdAWOtOwtAcIN/EaX7uCUCHpU4ql9V4aMMWzysnL+MahJoDW3
iLHCemS3/UfEjEbqvoh03cA95LpeVWtRKWfAfKjkczUyQOIxUALIhyiPEV8gu7nC
mBDHvR0+wI9Ql8UaA0W1H+SWNzyJRCSQ5ZPEqI66PTyLYztUBH0FrZGRZ2F9CqVz
iaXNc/0bVykXRzojBoMe1dg1Y0MzuoqOJtBZWT0OSpG5Gg+F9N9MyJaZh8GKo0jM
6JnpAHokSjvH3P2yWgSTyUHKX4xlGFzz9nnNxcHpXCtdqjaK9hrRIYXKzTSsoiJN
zfBHXaLODEp18ZbZ6+o8mRj5jBuW+dmtzB0fv5hy/AWfXNCmElbROr+oTTd+UqQq
vJzF9r7c7g+MmM67c4ilGg++6JjmOaN/1uMMBAbrgOBNMjZF6LDjYsftv2RfSX3y
DqqdmntssE20jvYvMYIMGBXQDXmiyaIKyZEYdy/Q8wWXxdI8Wt/lCSLtRdGjZFB/
WBL+kNFslKL2gHOdrL5xO0KAi3NnGboZui01n8h6U+JRHf0dQO4ME6mEzweRDohT
QgOgKngM0qVaVMGiJDGNgPP9Uz3SZsYqpeVwUsMiaxv5roJDxfeeNjisiUd7qN7T
IAkj8OPFLHnR40v7oqMRJ7+ieCrR1h3ZfSIjB7XXGg5U8p3AgHRKKX747/sVG5mZ
7fbS0KlbSRE9O4bICgfHhIq8x+xiqztGZQdblF+/ML3hDxSxryEGOGNXqhyoKNa/
ywoVnGgpMCNaulbLOE50RtQOHh0MB2qnZuEcb5xM/7eoJFS6r6wFPt5zJjT5IR52
XiY0peiczrReiInYFsCFH+1h2a/5GP7kYwsC7BY130PF5lUCWLMOkArpogxJyEoM
EjkCiqWISRWx1S3T7y7HVrcwrE2Sk4oksjxGxb3hRijlhkFucPh41vIx6aAFEm5T
vJTDvtzY8YZxr6pWBxFI64t3wnAUNn9YNMVbgLXUWjsNdFfWu2dIo4wdQz7JwAGR
+AXNXrG7jkh089yLDs4j86apn7864vUCNGE8zkZ0/AS5HPrFfPeW1bn+hywgRjgj
2xn80NSL+zsTIMydDZGvWJZFgY8zWmuaRyu4LXw7rEP5on1ssCMgXP0/6uNDfHAG
IWdZHbtQAhAQgyFY5PBrkyXPhgSs9apU1LiNrCzI/PdVudfQ1pzl/9u5hPsqOs3i
LdxAlTMZyOvG4qVK10znrhPokwoWE+WrIBFkStfKQn9sH3TfEAVa470lJcltNi/M
sfYY2gxDY0b4PZ7ckCMrZP85W4Sc+hPD9QZBtIYHOxk2p62jU32DpZWuZFKKZvbU
CEJGPevjrxLAzD9aA+VHcNUtQVk4e8IYnqIOy/9BzgQNmBImMxY1sWDWGAbB23xO
2DecrH/5/82Yw1sSNXjksQueyNtiX/EoookNLAYzYAPrIKVA6uxbTnBLEnBuYfo/
AKXYDp2FFzoWJI2aV729CRhmbJKxJ4giNMGbTHOoymVvJkbTwqm86tpq6rWpaBoJ
oGl3GB2aAYEePcEkdodO5quBi7LeiMNnYTu+iaXv3SgCHMnBvLZTStHuwbGKPyd8
9Y2ZREzeHE1byMLSKPmwbu+iUNE/fiWfR7SMY2jzPviV0EsK4Vh18GElIRGan041
6oAQv2zFuPNnySTDNqSzoCE21cYgDrrfalb9Xw30XYvZhaLPCt1m+H8azmRXns9L
MPIdSnW7n7bocjDreTX3pFWPAHiBNHLQcYREeixWpdMQ2nB0MUKKAyk3DvcqfPXU
x3FWKYOeXQbHjmhIMutKaaKkdPiIsjsz7HGHVnj1MWx8aSOoS0M6iLY5PzcrQ+zR
hD6CfYPYSN1cd0N6jw33w1DNG40HAbtI14LbubCHZnHfxhhopB5O0CXIN0A9Qtt+
x3ZYTVnBIK/1YRO96pVrKKTF+zC7RMxpFYqTjmElLwDv66WnMWu20pBZMG7d2/wW
t7E/FsKUlV2nFiCluU1j1cH1m6R1zkFhlROz2iaaQSzdXSn9QLSra6wc+odUuhul
IKMvjc/C2iXH/iwsFqqHl+t6Qc1uwV9UwMtD3cJbKI1QpcbxQHr3vKcFjmgjw568
`pragma protect end_protected
