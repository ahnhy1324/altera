��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O�k}.Ż���"�����x�u!
�*�*����K�f��\ �<��nFɚ��f�.&V3�t�_z����RZ �UP'���I"���U�ϓЯK�݁/�G�5��#
/���R�|�1{���_����,$Gn���G�M�J]^e��Zd~;Rb��N>@���O:G��o�)��A�ڄN����z=$��TD|d�c"v �y��qBL�����f+O��Hr�u���?�\�������s�it�Ư�9h�dI��D���H&��=�8/�i��x�pD>�่3��8l�Y�#�`�ώQ��oE�h�V�2a=�|�WB(L鵈�?{+N�ؔl��YI��iQ�8#�j��ӗ��\�1�Y�Dhv����@��Şc�Z�\b�v���I�j�q���V< ���Hc�3��(��~����J��Td(�Ɗ��}�C	�"�y}�}x�r�E�/Ƿ�  �]�#u�ş�N~0�|p(�D/�s���~�xnೢ%5�.
HA�j鮦���z��!���U۔���0?���m�Pf<ht]fވ�ly��8��7� ��3�0���!0�`�=�|�Nzb$���I�q sK���%K�Ƅ�U]��]�sF�޽{_���+u�� m���?P�@V�I5#�A&n����U@a�#o�#8,�����B��7"�����V�m.��w�*W)=����p����C��3ߟ=�E�Z<�쵃�QFT�<�0�.jj�ckr}b�?�ʣ��J
G�4�2r�I4��C�{gE�NJ�M��I��[k�a��#\O�{1� s��Tx�3YүTBM
]׆DOe�@S|����%t�}VD}c<�Z���#�&L�1y��P=�1C��9���`2{`&�hթ+!�/�x��)��5��M�,Y��[��Օ�����#��kb-2	N�D�$jT`1 �j��1+E�����
܁'�oC]ڪ�R�]��_.�uR�����_��#��I�I��8����p��g�����b< k[����1��'����{���O�`����n)YO� q�PK!0�
��8)44�(�5O�i��QE���)%_����+����%�Ƹ��o��5�d2�9,|� P�ͩuKL1��	}1��}��om]�%_��]\p�b���j3%��	Vx�92����1�$��lYC��Jd����y���fy6yx�O�ʣ�� E9gG�I_�[��g#&C�P?�h���6m�s�%p%q|i����D��DpwZ�o�Q�����Gb�&��_����$��%��������A�픅�+�Y�Bb��y8p�#��^���O��E�z��7��?!4���aE�E0�]���7Z�J�N��Q��SL�Q)%z��=�L[̽�G��F��A���9�د���Z@�m�����^��V+��Vip+����.�"�E�D�v���k��꤁�]WC:�[VSA��Wo����n��:��3ļ�'K너`g<�Q���{�c�Z�I��䏲ѭ")u��#W��>�� 46��)Qb�U���!If���'�����y���4ݍ�c��x��!�г��h�E�&x4m����}�FJ9� �2q3�����775�x�"*�B\s�&�J�S�4r�;�zdk�l[�2��i% �k)G�'ɾEJ�Tº���7�w���@9*���Nn��6؈��+�<=�6C�1+�S�9�.���!0P.Ia��׾t�),�g�Z@]���?H����A*
�4��;�"6o�Q1hnFd��SX�A@e�G�o�	Jq���}�1���gl'�~C�l���.�Ӧ�� �� }~�H��I���	Y�M�H�7N�GaG��ỢSo~��:���c����B���);�����m �[�C'���.i�'���'V�ېVg��r��}O�wXh���(�S�Q#��;��T��`�N���=Tƒ��fe�T���]��8����?ҫρ��<�EZ��d�Ȣ 2td�����"��t�R��м��Q4��
�����Az,�'��D�E���ڇ�q�o �`��U`��}�ȓ"��7f�+�f���N(
	���[�m�'�JpXzU��
���j�:�G�=�i4d�[q��޴�&U�K�أ^�⟾�+J$�Ez��Ҟ�-��#���K)���y񷲁�Ѽ�.Wnv�xj���#�!�9#_���]�{�������a��uݔ�k�:ݚ~V�$m���g��9���g?�<��p$��{i֧K�����V�:�2y��rZ;҈Xo����w�N���X�����:�x_{"Bg����}���B��0��;A��i%R�t�B�5�}�*J9����Dk�=Ⱦ5H�7)�!���S�D���]%Σ�Q�����'��w>�b�BI�d�>_,��(��9K��A��Ź�>�4
�z|�_���nI�{`-ug��K�Z�?�cR��3��Xqd�qC�⯼|t����m�;Ҕ�?��e�0\�!��^��J*����ein~�:�-��x� .;�v�O�{p�]�UL��iǙpÀ�"��G�WH6�V�G����������>p�r*4��=Q� ����w1����&Z����{<�L\�6�b�2J@	t�[� =n�Ͳ�UFa�������T�@w��B��j)͜��Ҧ�Ý}��z���l�_��ï�D�q؊�i*�#H�(i���4]GReϴ
	��� �3��%�G�`�Ӯ��Z��r���Vlg�!�ӚH��Q�|
�;�ה�j�C?���������+'���r�L�������5�G�*V</�u�`ѣE�ky�* ܱ�tu��:��j�Ob������|eX~Q̹����֕���!��_�ҁ��E�W�9R}�}an��w!$j0_�(��`�kc�����B)]%���q�fT�^�d��5�����_�S�"���h����������A���a�E���B�~L���p̡l����7)V-Y|՞�n���
��]��H�pT:���*W#j�����ڇ�b�r�	����?c��P[˓>8a*[筝�^��*6�M��n�K&"�U#�Ϣ����;ܪmf���S���}б*�ō���8!R�R6���#���jx�H����w��8�jg��	���	9�u�Z>K�����N�Y�@=B�	M$��TI,��z�Ln2���eM�v��yH��|�ݵn����r�iΰ�F�W��|F��jlFJ�(b�i�/V��V�~u�5}���}�	�Ac��)��~��L�u���%�'�x����c���.�cX���/�BL��:����-:�����=^L� ����E�>�z��E-�G��C��<��(�h��p���J��W�w�A�i�yN��7Ԟ�*�bᨍU{����!64�y��rQD�A/~���[���Y�$$���Qt<��',�d��8�2V�;�x�`8��U��N���Y)��}Y�<,`��0�UL��y���p�PŸ"}��5ä�	�p�u�[�����=!p�GU��=��#���?	p�'�{�ÚyWbO1��9��fR�g��·����O(�Ta_���Q>e�^=�".���\'��~���J(K�[�,<����qE)S�R����G���Bo�0g��p�� �8k�f0�6[��i�6�v:���Î_g��2�}PR���C���<�SG�M[�^t����2���e�)]j�ꋋ���M�4�4+A��� ԭ�H�W�F�9eM��=�D%]kd�,s��T`RUjȈ8�W�@wz1��G��ͺ��pS��� ���?��&�攢	=*ǌ�P�6굓�E�}�{���X��r��^hj�yv��(]�whz�,��ϯ�0��B��Ϡ�������:��ni���̫�.�E�[�6�Bd���#��=�x�D�����?�������<�����5F�۞�a��PF�	V��@���j��e4�~W0�_�Y����zqӆF����Wc������0H�l�e��BZ0�K�.��"�T�۫��O��l9��ha���gg����:y_9�T���M��0��乧ݭv"h#�����[5
 �}���V��B�mh�8�	�����w0#�о���H�RJkw	fڸ��2�D|^�?��Z�J��?�%��v)�;B�|�>�3�B��ժ)��(�*H��`Ox凅��ux�e��D���L!gy {�� �,�����~��W�s�%����_���鰯���F�8%�7�o[�tJ� �E���V<`�0��?MoAV���Mf/� ֚�7/E�h}�c�ʝ����GXq��|^��� ��R�l}�@��C������1�|��u��m�(?+��(��E��B"�
z/�}�+>`D�'+4��zvJ�B�q�b��O
>�h��5Sb�*�PѝP�!E��ĝS��o}�z��\Rdv��%2Oފ
����*���kH��hԁɄ�EIOv�$�*`�>���#$���Nɨ"� ��hl"��c��~!��ێ�#����6���|p�sE���3uĭ��1��Y�������(G�!���/F?X�n����n��b��c�4P! �U�m�U���U��(��<i����Lh�;������@k3rsk綧8-������-�����9!xXS�ܵ�7�W���rlK��t�w�{��U�9$xҕ\�-��u�A���;�E� ��� T�*�s�u2r��	�	3{��X��-�\:ӌlN�k��%��+U��ݱ�Z-��s�_<L�jÊ��{�h�c��r
�u	j�m\� |~n9�_���Ȃ��XN���-!|n�@�Ģ́�z��@�	�J�W� ؅i��&ܖ������/k��)�!���T���z+��Q��������Ǧ����C�0��ަՔ��&���AD�����C�DMs9лi�'47�7������w��|�ԧ�O�}w�v�(�}F��<��c����C�"� "�Y��������f李�)G���+K��/���>ח�ǡCGE��f1V0�w��ޅ< �Rb���S��
<��]*��rE����|[�|v���f:�$��(%C�D������ҡ�%�J���to�����ɲ��hv�/�JdM�Y:�?➷�M��*QA�>��f�>]��I�Dv�	�  v�K��q�]���b�ϰ L��NlT�u*v?�v�H÷��6rٶp�vs\Ph���m�l@2���'��:<������$kX/�K
!2&.Z��{@hǛC�5��49.�#�lj��ۋb��9�0�α]�V�k�O�g 8������tL��4M�c	����򰆨�L��sҫ�������טd	���S!+�x?ӵr��q~�rn�~����aʸ'�H�����!ua�%�d!3	��޹{�5�}��'0���YC�	A��s�J���}�jnR�%�z˸�>Q+go��:�����9p���	
�ů?���ý��܌�AF�ga�ݴ ��Z���&����s`~=k�2����^�|8�6&Z�T�c6�a����!�Q��~>cP�ޗ�Ri; �VP�}R�7V�:4���/�_�0E -'�[�����?jD��]��j�!��\nrB9�D|��ÜUX!��q�(����s�z�� ��p��A5�ިjrT��!�h�Q]eױ��!�5��~����U�'��-����~ok\g��#6F�;�9�4	*�HD�MowU�]ӳ��}�C��w~]")&P�%�X�Zm���A�M�Km^���������2�Kj_N�j�G�9�~����q�u���V�A��Yv�C������N����fҞ5`���35&�F�D=�,���C�%��sj�F�i�Xp�>�����!����?�b�����[����ƭ�TW�>�M��^_�}��9\�s�`������ҘuX#Z����Y��g�.����6w2����sw4&\�r*}Q��6��W4x�Tȸ�G�8�B:\Kb�6��۸
��sh����կ�G3^��A�~�H�x�W��ܮ�ǦD�����1�q'�S����Mwq*ov��\%���z�n���BY�B�0��qc%3̂�ن�@r�C~)!���7Mx���8>7C��[�](�At��� }�X
W��m����*���X���Hi����A "�&:i�A5�,×n���G�i��zG|;�L�����5��و�RvD������d2�THf!6���/�_D�t؏R&��ړ�.��^�e���@�5O��ɧ_�cC+��5�A_}���ŗ?��yn'uj�#w��lO=�B�OK�l�Љ[�T��nVu�ɍRUد�M��bzKjL�ݎ1�d���;3�GLm���k?n�����O�k	 �z+�W<���[����Ib}���/�9��X\�{F8�ua��^O	����@��P5E�oE�5ƞ���SH�k�ٓ|��f���Tx�?v���7!��<_['@��)OR	f���Kw�~K-�#�[�/ue���)J���ӥ'����I?�ǐ&��
J@7�ա�.͖��
�k�w)�������
,��*�ԍ�ݥ?�-@�?&��4�[BM8�3���s�ۿA�b�W �ߟ[w"r��2�4͇ܕ��'Ǯ�U1���Q���])T�5��q�(�����Њ����~!7����s��<G���a�0T٥�^��A�+a�k���ϡP|��4?�%���:I���{�q
!t�?�		y)B�Г!c.��У�Ż�S�>��jW�hQ4`���Z���kv�����A�YL��Çғk���/�h���A���=Z�G��$�A'�FPOe}�	���F`��xcɋD���D>%�.f�O��(%��<,˯�8���5�T(��������0�t1l2?#N{v:��O���c�`E�?�BзҢI��Ú�u�f�.[ƨ"+EA��� U�DV�*��n��H�ɣ3�@7�\��0Z��؜��hU�E�˷&݉Y.M�F_�DיU�)0I�T�b� �Qf����oQ�ht�)���vlF��L��x�kuX�U22�a��=�����0?������:E!���þw�O^F�>�QO)�yL�P|i�Q1;��u\C4�B��t|�
�)Ч�z��]nݐ8;�9W��u�{��	)H�'��N��y�w��� �i�K���?� -�b��m}$1�^���swQQw6(!�G~e<��-�H�B�� �@�OI�7�D_c�$Hg���%]#��*�i��Л�Bh�m��(��y�7,���*��B�T 
���XI�N)�4�n3�R�X�CrH�"I�ֲ]o.3���q4�c�����%�.�;���2L?� ��^莏[�*��9����u�M�!C�� �g	���Wg��g�D��	_ޘ'�f�ب�C�V�#�(xD1��gia�`L��V`
�N��'���Z�E<�˹��IV3���|�b�����*I0�w�
���e~���a�1�[<��y	{���x}�au��v��H9f���Cn-�D���%_�jV��O������G��Hxq�nU���Jo��IVKR�&�.Yx��/H�Q�S���Q��J��A��7���6)����	��m���h�5�K��j�v�ݶ~�������^�.����Ph�.R�y@ƭ��p!��ްu�B^�lF�Q}Ħ�¦K�>���*���D1�kC��n���T	��&q'��kl�0MD),�O��v��'�)���~Z���'uHw��-6�?�\�ow��Р��Xcj���'~cPչ�1�)���*����b�v�%��ã�_3�M�IQX8���G��Z�Bj������̒A�M����"+�_�|:��*���_�G�}T"�'��uO�l���0q�r_�d1��ML�g��?Տt5����5'n�Uzl+ZapZپ�G�P����S���M�%k<���#&�ಢI��]�Jy���7���