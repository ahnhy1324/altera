library verilog;
use verilog.vl_types.all;
entity smul_vlg_vec_tst is
end smul_vlg_vec_tst;
