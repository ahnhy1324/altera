// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UGc5+bl2jXWunip+t4tKr6CKvxzdf8UajqPZ/LNStYxvVRjTKV1+h5+V8Q2DfPRu
JnXT/JSFoAXDLEt/muOn/O7YfOZYnsP4OaiyFIuziZpCVpw8RSOqKOkgaICY7P8E
hgnko20OUmFQvd+YBHb/rgCfcvTGjRhzo27GUDUI6ZY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9008)
yQtRsjRsNFucUhIl27KCAOiKTTIc712QVyLe1qeql0NOV1OOH1rkicJpaA12yBem
tkNeLk56BoKhgwOvhnbdehzTUvXlOI7CTw0QednQI6Cb/5mZ4UZ3R3snwDiPkDOU
JM4yTlDVhsMLGzqgjnvexBku8gMtVk7MRvfuE89Tgg5mBeSi37McU8d77XOlu2Q5
P3p9Tq4HMQujfHGqjS3Ueg1xVQwLKFxpJO1PclJIqKbmnvR05ExSLT8e2U6FepLH
AUrIQsoKrfmOaMcLfZQ/n1hbZ2pakNR/Eq2YtA8GsutLlbts9zhNOupWJ4tO0pdI
dUolyjzOtzBzoH1kBFMtTYHCLfCNHxMqQ0+M3tdeGil5WDMnBURw/ShTWpluFRX3
8QVlsojyTdqCSv/YDNun6nvmVkpgRuafiJFIG6fGOG1ZyQhp2Qg9rEt2EUf1a9vm
GU7ZzHc3PTgS24LBD8gs4OQyyl5Hfm0eYohBw7Zh4lVyAAmTZtY4yq/BEfmJhFuz
06DqG1LTdYLkeT2NzzXoc9tlLQ9yCVtQZf8lDC7Sg5F5Svp2iH5n7/trd/Pe1Qts
ZIvfLZCLIxE02yhijBQbfyaRK2Z02rmM2ZTvj3aQuETXDfv09hYFJF5vMk3iTOSt
1aCeAlNlvda8mLZ5XqatBDteLTYx/7PkzbjRpBRqJhEs8Qt2iXO5a2VvcSBivKvh
vWHbRdBwHlnUJZb0T9LHTIjjqGDVSsmgU3ENo40E7jLZ2wuf8Bx6Ty5oa+VP2Ety
/L4NHrqAUScdY34LqWzVyP2GTczYsUBeRIqxOyHaeitaP0Q21dL7DHpE7vw7XHbY
cLM8j+OFKQioXEvZ03IJ7PidAZHdaRkBM8d+vOiLNNRW0BralPiKCjwFXRofQ9Ky
y2jIHNe4pc1gbfodh8bjlDDhGgzOKfsB/i1CNzcqQYnhwEKq5vxcZSVohYSy385t
7CJVKKP70KZxPaUJZNMO6Q7tRPWIrd1GswQiBfb5QDI/n+tN16i0hGhTQmqM+H3n
hW4wXiHUm4r/SyWOz43BGUM/wTPP+OZWCkrqet0g0J6qYoyDR56B5frp9PdXVHfp
67411s0e5nCa6nkjAy70mQxnJPBvud/lKT7qp+Cr1AN++Qt1fshhYFNBzeSILT8I
k6nv++zmy3L3HDZkOL3EV5uJGGqIYZzvgvRhdBPfjuxK4ae/rpp2ZTiZAJSJNZB7
DN0AxH1Kts7Qn4RazVRBUWD5wR0Hahzc5rMJKcpNYg4JcPda4b6sMLOKhpiP39UO
zleogNhMabCa0PfaLCm8T8Z5cFz/b8lrbBL1+cuy0ow1ZTf3b03svWFq4X3yYJ2D
/KPyV3rfqn1Wn2jFuqS1BR5qHQS2+yN4TU/sAEIi8XJzkUoNrKrr0aEN7mwY4qWD
PLE8WjZkab0O4nzM/IeXCi3vAHNQxFaaMzXYKiVAGPPsED/JDG2pQ2eAg8NVo+91
kwJyNdS8zsThs96hSFCmObYb+rHNkRF2PWTdwj0aKkVGeqPOm7q0Mw8G33uE2dRZ
LAOMJyDhouR3azuYIa15Xd3gJW54+KmCpY3EitT1APGK4o9+t5Xgh4DDcZzwevsX
6kgCQYZuQev+QY2rYhj7jTuA2jRWPOkdKGDbCZL7V8nhMKd4fAMe/gowClJLyDu1
g0Z+EPXdTwL2KPS/1L7JoXB12QLcVlJTEyEYLYwNeSTVGcpt1zD4PID5FKIT/tbC
cYLmSrNisSd+aKWF+0+xV/YtsA5dUSNV8BgAzKkesCpdCTliMOujQJSeJ/k0bawK
hGWI3DqkuIqVOv/u2fbGtXk40f4SUOiSMb2/zCgUnTCDNoRQSaujszKTEB0lnVEU
qoD7NndsFRuYUjRZp9u5VbLNaFWkeALwwecvCh55mzXue1qq4138GQBBRLL+X2nl
GX5fJ0UM3RtF1TvV4zkKOLALSjftm1q2Yik92YD4j7cu35SHjqp7fKULTflQ64Kw
m7n/1Kz39/K2XmRiamQBlSRE+3VOIYH9gpoEzf3/JYFVxN2m69w55MAt9VdJoGUg
A3LEiHhCZDVVHUqidcZGn7+plYc1I8geHumM6nWekXm6X2RXPC0wJhOzw7k3t0w4
LGUZ9NNYT6b7JuU+flENzhv7VmCBCm+ni1V79Y3jmTQPqKZXdt7JZrW7L3ZAfRDj
KjN3OrHKz98bWJZkbeJxahkfHWnS9055DeFxgl4qbnDWGuuaCQJjArXWMq7D0jlg
vIm2WYnRne9N7lzkBCv193Gupb/UZKt8HDYpe/wly8qInB3JaEMjMxwvvZaZkBjk
QTnCHFNfwC40rhhzRLvFX8YWH6X+0EQ6jeE2bE77K3iarLnTv05v/9eSi8tqqx5n
k4rVReeZAukHZSsqS4L1AO6hkMVzyChBZ/yrXxtL5QikOzNE6aEckVuDZRuIk/os
MC8g4sAoHER1Z/LKSrnY+FnDGX649rVoyZOwPAwnfRph4H2q7yrok8YOdyuJpjbF
3Cd94C1A80Uf18emWDgxKFve7DLNXTqxVhUIww6BhrKN7IBs1gxOXNcrFU3OEzvp
AcdvYi+AF/VtICAswAaoCFMagnMTKYx6Rnsm7zpDnRXaWgAjy+x/RSSLR0U81Fry
5efohko4uYAu8t0ebLt308kYOsfzDAK7kKPtemRpFtu9UPEELx51pyc4aRnJfr8b
D06e5dL/kSArAMjOLg/lKRMytGbPxPEhg5X8j/E0kYhjTGqNBm+cQHOy3WgFSPRd
RQIaHqQmSvDPymRI6l/h1DXvfKGGjF95EieXzFG63AhpkzbrGE4sVJod/Ovand6w
LJ8r7AMbRuoTU8oJXkXf2kI3ZmzMzvhd5lubJPlUAC4j7c+1LjbJGUrioiqBbVXf
6LcYiBR/ACsBKbCI4FpigQX9x+06TzXMzKB0xTC2RmaUJXICGNtlnJsfu92B36BT
SsKRyb2b1pv3B+LSsfPlXZO3otu76oe7L++CQSdS5EY05HqLgEqk0fVHeGoQj/H2
+cHqvy078c1yo0ZPoPCTkIXxG7lbucODuZ52rfxaOfe6t94WLbaPMksImakN31r2
zuQGAtCpXGx3xkcE+n/H2ExGBFUUF4981hVgf6DAO2AL5hOaWsDzjcnt2/d9vBFb
XdPHB/1ttAFVVrWJVu0XfiKBJnsdQlYJLhxbJd0VfpD1zEyhU5mnOQYWoHTgidf5
2DM+uqcyaN4xI7U0kx9YXoIy+dRuodv6coGW3RkGA6jGDihbXxJIhJzNfM3lxExb
Iffu2g6lokWR76pIA3bVJgO4QCxxBz7MUtgjLrh2XfTz6dzfVvG7tcEPZTk2T/mi
4kzQXSCRdEArVbuill9PllpWGhYxm6UJzfxRCU4nCZiSZ9IS1q1b4pYUEmznqNKS
ifWhWylAcnKdC4FwwVUE3P36WBNU4q4rSCQrB+FYhM8X+8PFfk/4qxOYBov5NkUS
mx34US0O2CHY5a34vN7M7qjaSCaE2CK3FbDViVEmrPe1YQZuZiG1YrRIXuMnmgXi
ON9SSASV0pOHYyqjNKEgo6N4x5hzjKFE8Wk0qij2spYSKgkBcvNVEL81PWEf5Jpc
WVNplS7SXeQiBQusnwxRYW6111iGXn5WyY4dN+4P8NuMbhpLh5SWGq8WcoEcBCEG
KHk+EDmgTyf586Kw8cyQlpPZ90dyCLxeXYd+8cJg69jWnLJ739yVTTdrzlZ+52IG
Mhv5K0GsuWaP1LzpRpEC51eD5a7GunFgVSn9pbJYO/zcwH78hnfFcOHcRusi+9qr
Nn7My0ZrY2+++881lymEhJ9/1YmtDn6HKqrDG+WbgO5N/LjetbRaTWA6iaDLtK+8
wHssDEe+R5Oz1rlH7RjPeoLGwfGxAPsYT3I99JMJA0HBtVuWUYa+AHE/OENvfc98
fhj4OFlxNvD3dQPIOrxIbSDQVpgO2GOWHFyr0P8oJkIq8M9sy+rEpo8vau/DRRug
SX22jttsLgMHZ2pnZdpaGeH8M0k4kyo1ffVC3DxJUXU8Pap1TlN4cReKMoAbPQDW
snUooJR0CfMdAgZeBbiPYuQq/M/u5JVzNnXYpyc+8jeMN0Lrw4zk6pZbQtnQBNzB
BWnyPDSBBy8QrcbU/Hl/MskwcLONBNwJZuv8vhK4M2qMV1cqQmqZYmXxF7OzhjAj
BCcXaufL7iKoOp18UyaDb4VylyhOb8ppZZr1BBTMCJEzutOlE8kFLd2tMyhj9caQ
A08+cE3af3RHdO9Y8TSvruSD9nQ8XZ9s+qshu1igjwxR2Me+MIor5ux4HHA6YKZf
ENhNSt/oWzTXc4bCYK2krk+M25JGzMeGXX9wk28nBwO4g5v7p6lgsl3GFKgBL6t2
BDFFCaXjZyuTga//pNfnpaxh8mSiKSLZg+9ZxnSKIEzuCyP+ktil6CCTtl963xqZ
aUZagJA+pG3WIgyuZFarjBnrszQfjIwmiDkT/g5++MnVGen5k+l0txV2CEJQ8HoM
Z/KIi79yTz7KdahixgfSa5pSI7v4/1a3jzzwdrTGbKJKCnGBqNhWaXa/3CJS4O5U
5XWsoiQkKWZFDhfx0e5KdRkSjTuOFOJw6k3yAVumb1PYmnmNBxpM5jb3ZHUqunSx
gcEaHLx2ZbcV+P+Sj0UAdu87YTmzXO1LU5gvPdisxcR1Se2/Lq8gN9yfuYQz50Ef
Qw986z8ptVeyqydg7ZTxjkwQWD9ndvjiKh/qWHdypaF5UkAW92cZcTNJPNp9AScp
ZERbZImZe8qK9QrgC+Tvo7YKXuNeQ2oBMbt/P3lz0rhbxmzgB65CWzAIZhqMmJyM
vIjpAVUbIoyXbFXPkK8YTo+AEfQCih9/zMFBJKZ5PxI9Hv2k+eNf5wuwpvd9tVnC
48OOOkE7BWswzzx+mxnQUlycyP+rL7JGBgNdP9LzD/O1mAjP2EPBIJ7Ba2Rw1Hra
vxkPErSrwhM7AqsEls/nEY+LZ1zVJfpRs0+30+t1Dv5VFfFmHYdjVkhbJvsRhw3F
Ar1kOYy/cBI4/L9Qspprx/1M3OrYdDCcIxEYNI9UhYl3znBCs/0koBdWyeyPuN9+
cyI0NQp4QtOsbZNB9AoLUCLeUHbkBsSPKWnJxRa7ZUVP+lVBtAtQUofEyGxZqRF2
17YK/lNP1qgTaAJNVsP3+Al7UlymneEpKJLu8Fri41z6jiX4Ejxa9SykQaC0V2NM
otMpNd4x8ldnlMoDkdtnnZVsjA4pjotI4wmiW/Eqj6CiPx+PEsuiCZPvnXSF9QHm
L/Nuyiv9cGQjI5QJ9WfBTvQgXIHI2a/yVCotsecG4v/O5ozz7FYNoXJqexr8dV+Q
sy2/Q1AWCJZ+Fg8BDeLOPjqVOf2llBvqSUY/ySJWeYNLCDWMnJeI17Gc/QT447hK
liZ0rFZBT9eCl1PEDQN4VOBXk3Whn1PFHg767gXEoq2TM3GrzbK7MmyrFz6vcgWG
qqpwbItPxwO3+6dRHEK3QLrMKLwntEy/G5yItDlZMc20Xc8UvEpv3ccjQ1jJZ4z4
PEJ3LDCaSCZtuBnKNORwv+mHWCYLuAXf8JmJQLYmc7cU9rRVvnYxQvp2XnwE3Q9z
HorbHS7w8P87yYsVZqecg+YwATpEuf2MbtQ53Pd8BVaGXf8FMggr+jtE3daNbGCz
7SlS7B7wwmgpWUTh6qi8csta24QKxokasVMKFpAYIl+tUdNEJvlMYTsBYdQFqssK
9db+Qbs84zu2YAkze7Kcw78MxkzJeTbAdC4wUN4F4kM1/UKsWhfKTD5Pi+R5rODq
f5LEf/jh4WWbGFUODTTkMtA7g6orAZw7GPB1PeCJQxY1v1m21mSpdlxRtSku+Ul7
bwDcXaTBiwYdQBs/VgzV838AXmCUkeiktX8TvqqD/8I7fJkjyy08S056BBR1W9qf
6DwHVes6sMXGgdKvRUacnkuUMZKlCDvhQ+RC3wBU/1AqGzGD9VSXigJQdLrdU4KD
vm4F3yXiIaMyO4cYu8AxEuF4jS+VIggj7xcARYcoYbra6MCKbF8bC1u4NWRvUoZx
YXDaw73+zLb4ZCTtpzLNheNtsQJuco+4tKTyTU4x586AASvBflGRQHL0tDDKMtI7
iFMuFzKMm8MlppcPpTHDfyB1v7x+ZDwmYiSn63X7IXREWIqhd/vHBIVZEmC6cYjq
o/KS15iBQv7pAlDPVwzzExYL5Ngm/dyc6C6lwjwu5vZmHQ0HPfvwbyMnoTc1O2p9
ohyrXVIEAUZo2IClWUxB+LP3MEzCPKMMPqbFc7+iQo2RspwrsIzagD8AlQcrzJT2
5kzK7DHf6jVdFUYweaV58b0CTBAR09ubglaf2ORxuwYfsuG/57kYVtuOwhIAhvAC
njaiyCjiLGTfo6DhERd/kct7wzoGkY+fVVdrYC38H28RMg/uYe6vHxUoAPMN3twz
TmGK2NK/z9yOjWYlJEP+pS1SHhs7iyuHHtY4wXn8RU3oFsBvqsyGBm0/s96ZauRP
ailagDiXkocroEEuL9cPWLrg8bWyc2RSPl6A6ai3o4RIyRHheyyxZ8ikdIESMM1a
lrR6NLGKiJs6Xq2yNTpgoJJqfaUPgTiRdt29OMz8KE4qLXYcHDz2PbRvDkV5eCmF
ZQcus7s2Xlm8Ez5umdR9Ed9mkma9dpuQv0ZoRLthQUc92y+kDCxsndI4mcOh643n
tyBfyQSVcRO60H3N4dRheAp91x3H7ONyn3Koxh0rX/crA7CgQf5/Ccu2rPY5Qike
XFc6jQLfF9jP3iMQwUcUcf3g4zW/MuqzMTXGD0pBzbeHOUu8I7huV/wtkhYtUU/E
j00k2GZuHDHgKdEKIrGjswGy070wHi11UkO37xGAFPsmWJcOuxoLbenpUV+briG2
vHvR/JRGIWAW5D/x1TnHadZH65oZLqX3QvWteHzXbM1HcE6bwuftFBvE/VeCQUrV
s2+PnqsvEDyJ26hcYvUzbJI6mAFlyDa3twfjpDA7ZuXt9oTdUrmjYk7NmnTShrcW
c/rQsN5kWrEZap6MY3MSEmnNST2GCZihr4Nnq7QbqiZ8wOtA+eOmftG6mvnZNGHg
4oDT2Us+HG86ICOcEsKPfScmZoX5Vid7Yet9F9mQaH6UShV3+74ZGaXKfiAUP4Ow
D+y0mynJ2Uqg/kYlfoq02GWuismZJusLGj+Nzwaa0S3lUwZydSc0GBof2h5a74Sf
asjiF8Mme2v777lZPepSj3NNmJpPdnrGFDQmCZRbwbUjNzvSI30cbMAiFXemXHdZ
iJTjGchI2atmD5FpH82ASmPi0RDfU2xAC86gri98xZDr0Vz0cXE/v/5OiMTuxnoS
kAbIfgD/UhBde/paOwR9jVTQZmpHzxVXzvN8mSOemFuEJDqhQTkfy6R3UeFF8Jnf
H9eKMXLErEaImGhWdjA0gsyMe2/coMCNlPCeCyDh4bRosFecAQnDZKzl/xGv43ln
dRGfppCSALCo70VhaMr7wpJ4UzzgRH3wV4JcYVw/Tgdp2jIEK021CLROaplok2I5
ZVw4WVgrFK5uWaDhMXDjVx2Wm5WUP46vaMEeVFsEguOzr7qUoEYLvwa8xBXGFrKe
Go3QRdL4hFt0Ppf8zYbc/LYYolIGtD8m/Gy7pn3F82TTOQAQ6z4cS+Sg2tyqNZuA
qGpcARgJRpURTT0JYW/by+MoSgdfGw09pET/oJHOif3h0Jj1iJwgbcVOb1QebY53
aABFcLEDAzMmjFomMOMPaUBWvgGZZkWO4M1GhojqeSv09jejl2IomCt+j/DE/Rhf
0FZdzFx1GwvV56+zUxs2/z8w93gVLDTi46A+MlZveynmN5PAHlen0simavZwIUOJ
C5CPplsfd2grJmIeXCIRJG7HxJgj5ahYc7BF4dmn4LbYHX4FYmLZ6AIOKnHq6kHA
4y14Ja5LUda9yGOWBpLMoIRrnL/9s4R/cOdpUS5weIPMM6BJQ3JfLPWrbS2+Vayc
/wog9a/3jLnCpCdb8v15WfcOw7jMv+iUHTHcUHmxLSp3X6BEAHPBkmupwOPMayiu
yEV/P7SrQgZ/plAI04b/aA4/MXkM3z5EkVp1ITUcBjbCdpYzF2vP7LsXnJFvu5xC
oiGgOajVAun+lggeqbWFGkOzXOTRCd3qyU0RnFn8VkKnvqs4s2qqjMWmCEtVouUX
rMU0I2SbHos8kMZxAVN1DB/ovxyEIi8g6LfELq4n+YIg53t+CYcR3PDVd21NFImT
zH4EOLnloMz31/TNrrROSTyrE2P1FKRl5pdUdxlBnAG5l3yGRkzjNwLHFKiO7yci
eF2uvDhL4NURpAPOhwMqNK+cL+mbcYu2GTeaAeeO7FK5sOh4HcuW84nT5iVjehi/
pbCi6wOuEd1feNteWpG19JzoPO2roecWiGS44wiPzV8aILL/C3fGosItiVFxTqgM
NCpSLY0RuVJN4JUOVBLU+OBf3NcFrsl7KM5Ig1i/PAAFEeNpFACaCudajcAkzBth
y/nIoSIiuVQyFp3UwjPDBUsQZEyD4vIC1QaloXSUaKmSsfmeZhqeHNs5jDk3n9Ie
q4Ee9fboetoofoXfYOB1vaN1B24MmijHIhA1CzzHwYJSFzMeWWY2KWSk6AR+taQi
9sKphszPxaSzkZcZMgMOml03h1VakqkQBGzTfxD1Rv8Mbi5YK5VRWkmWhkCsdeJ3
OqGmfjW8nfhCo6gGGwJgdWjL41uMOyZrfNKxyyBsM19AfxFB5dx/OsunK+eCa474
a6PyXICPst4nSzVU+tXv2x6pn+dcOnAF589GSQu87APOJei9f9UhNNLxjv4QbH8F
/0f7Dx5Wx4cZPFvfJ5J6uLJTZeS5d/VkDFFDbSESf9Xp5cRk7/xLlVxLjeYRZtAA
GP8PhN+hX4BiE5+kihncds7AXUmvI2JjfEwN/Inxr3E9A1NMdYqZE52wS+yLKIKZ
EKC20fDRX4IkPq2rPBz3nbTvb0IMsF9RVOhASYXebcIOAPn5pUdmvzvxW7b7rQX5
H9I+61QKwlD+FzN7ty2XwC9kVVPdjA0LjM6IFE4ZnoW5u3hbFCAawW+xL7a/pSDT
OiNgG+iXbPJLEJOSv30+Zf1VWFS8ud4UOoMYvcYlpRaBzR34jZ+/kRzWUvyz6FLM
jlfsnp9U8e7vDEJ9VGrxBl5lR60R/G1zk2UTS2wj7TzADl8eCDLv6KuekCR6VKgD
UAAuBl8j2Qf37L8oVP9a9nBaGyejN7VYQQ+0Av4LHh3UQBFAFGGBTm8A4wOI6Oxj
X3A2SbnuHcUVWVI0habtKCX9Uyq1YnYYHfeD/vsqXaa2FlF56v2ahaMV2LDN1txC
1rpKpi76rzDjznAcsxLOODsAvmRxp8XAgHzjQ2bxivUgVZglCBj7Nk8L/0pVZNYy
6nafb39oxvA21levKfa7p0N1SCADkKROVmnmIoDqZelVZiVlQqI7WsqGOAyv+mWh
UsjDXiYDCDayug3k1J0CUmVWo+e8YaR7OdDZOIW16vHlw8kj3iF/A2IWbpKVzscJ
y9ql7KwCT/e20l+rpV1vOzxnwuIjNTZmw7W0XhgCPrFo9/VYw7CgS6yfGtGVlHnx
6ub3ybZ6kai2AVdT1JP/2nSO8sSsxqPFZnDZN8va+21dggv//BbC2+V7mj6e96ip
z3F4uYO92WP7nmZIeV3wV000UojV2Pn7E584SVHUUNdMF6URrto8meFK8Il3TCpj
hzNjS/VieXwuT4tnzp0s33XflEVQ3oJN9hI1CKPalVioA78bDrrODmvjO/53/RAk
aRVigNcyJKW6ByRwGsUWUG347PXw4yFz6v5qKrpZpDCo7OA4XrySKOXwbY/vEieg
uKbYskwdr/CrNl8UJt38DJJoSx0hKPxDTQy6KQ9eWZuH5GlqPzOK9YF/7Arrj72y
zSRJ/oHfFR6UhdiHzUYOq0wS+QRfLtlLCqxUsFQq08FmdGINi2AQrVhVUSkAa75d
JF521UBEJVwe/O2C1ewpruwBplWHYZaldsaXqculmj90r63v3t/em916wB4RNgkv
6+G5ZEKWmyjqaBSzrdJPE27TJ30Ken+GSqcRxxlKOPC3lS98pm1WX0dLVfxVaCxp
RW5eUVuw4SVLuzkNHOelpl2jVieaG3KIuHDSiAp76FM2/RGj6RTBO6kxVAnC2M0i
I826BC1hVUm70DKq9f51DishQ0xrirvT2kz1sMd0qe2HgCJMMPb0qxzlpeRj1vCE
bqDLiCQ8ZIAZbpWpL1DX1y1rxe7IC8G4CCc9/yMBsxX2IdG68jkQdIMj/TI42ynb
OZrZAMq1CnNmKuYkD7+sOVQaCi+mXMxI31c3KmcaV1kQpF8eNHK9kEjrd4qoSINm
PGV19KuBF6MyjiEiw6LX6WG1pstUh+EwVPTIHh2OS8eDPB7cZEaABjKbGR8W3Pmi
D5jB+u9ndoFjdBzBtoLjaiWd9BXCX7rfemiNOd6zPP2H2R5fF7Dw4QKPjaELoQxd
S9EdrvAYToYI/wPFbmZsUcFUEjY7Q7SOw+CYhIsLKHpa94+MEbQntEXFtB3DNZZ7
rft8WoU9OFS8Lvdo3UY6pflymjGGK6NZTlPfLVHobi3yKKLM7tEfvx4sI9mn+woH
pixYG4XyuQc2A4rjKTShX08HQhRP3ioNzLlgBhdPEZ7YgkD7kwkxXtxOOA7GoI+/
2hJmHtq76/qh7pwUqZrxLNBgccuahziQkBlCSd1r7mHX9m6BmsWXM4xwrkat1NYE
qk1JOKp+UYvgiRO2oCyatm1DtHuuFu9Hul+R4QexRlgUOmhRP3jj2sLPddX8sl40
1unZKNCBwc2g2ouZ1uzrf8htEc6B8AUpv3myDosZSaCfjHr1rA3FU7cMEPal05EY
m0+kD8mIxYmwCQnEyJX8ZXMHeAPZ3ZNtAt7evVNcAy37W/a6GArq9j9XnMe4xBKj
DhfTbvyMKo7y0T7/rSsL+vrF1Fr9vEqC6ridvz6/M7YRnwBlV1GhiplY7p21jgq+
3pZBKJHlyWekC4A1+k3fj0TNUjmMZU/EJDHOqhRCt8oTc2VNWrjhEwFGTcDcR0kB
wtCpnBIRUQyWBSarJUFAVua4HDiydzXNKkWp6Zhn41XkHxX7dSyWs7oOv1OjMiSN
ZBjBNIBu7LxbaE8/gfBkXBQqZOKCFtbFpbwA2bbNFt+fBzUV0060WBvG5p6L4E8v
cFsEbY1IP92B1HmEloAJ6X2116FFkQA082gZXrFzG0fLjbVYGDTXbmLjzfb24OLx
GI330jrNp1C9FNJ6pmiJK76PMz5+NL0hoIR0sIqraZ4xrZ2UeOyvFNY5KFJ71pFK
OwRxGVi4AXiqe8Rk3xnusrvld5VlcY6sDAZnpIGylq+dV/yZ9gD40P3BnGnoEoBk
UTljzNRQnjGcK/rDSO/cznNTULwuWKgdlgqQwxEVeLjS2Rlx1yvTUZLVxqI/pXuN
TEiaHg6+Ylxmh6aScFMr0QX1HJutKSPrFtlb4+84mc/Xsnisamv2Te2aWgEEuYFQ
ojUOyklumB95+m8BjYZf0XXP2Nsq1NFWbkxa9oT8CoIgIKNHajLkCRcQFhqNf8AR
QYYFN6Ru4z7Tc4j3ct6se0db0rhlpUhqRMjIbTn7lr6hK0nx5H9SW/FbUttSGHr6
uJj8wDN/pgtnBqPKPAWlISBugEgrVTQpL3EG/Qa29wTYtWF98QORAmnzsuN8KEni
Rb5nPUnvlfdQoiT0EdnxWKQrmtbB1uPjs5EYg9sqcqBqpl69W8UmEg6tb/em5BrK
d1sCH4nkoqWtmUaaj+E9WZQ3mZN+EYM3JexoRaYi28/qthsAVnmCNsNCbSdBKedx
ift1Qvw9wmBRloujEfS80B31lL8mTOt/qX+JPXf2LGIhAIE87SMY6D1A44+kNdbT
EUMMu+yxPsgAcu8L+Md6OibaRcRVy+tONEyctwFRfUiLTzs5rrHbqaGo6hCKHIOo
tztVurN9KIhPAmP7vuHt/nGdlLYYxm9r+q8ODo3m62abcrMVbfnYdplOHaWePo5G
eliJnP0HXEzMC1nwJvi/oz0bZDOecUOri9sBjbMR96Y=
`pragma protect end_protected
