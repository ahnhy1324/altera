// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
YSnjFWgut2tI4MX7Ol0Z3wtUpqr7t4MhgWlYdPDmk0Utm1Jra4Xt3tAuhIH8A4ObOONCA7i+yz0H
jT328G6yQGWjHCDq9rMYT6/X+K6RNxMXeWx+lU/VSSd7XXJ/BmsUBMVGCh1cRkBIVqKBWGOyM/YI
ghHwpTxCULJYQK5t//hXqYXfE4QKTZywy2SNO+PhKfaw2EEdFmGsJ0OPcvOPeJ5n4npesWCt4kX/
xTp/AEtjVhDiWIBOWSUxmJ97jzwEms/G9iMNLaFcaMAlz1eGM6VN8e81geoNONQeDWu7MsqNhpMu
3GHiL/z7smbXKAsPmzHZx9kC2pNeCN712buEpA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
hpWmL2ADzzNxEXK99BlgNu19UfsjK/bFVpSJeiRvnJpbkaawf15omk0HvNOwoXMaccNI5D4TPBQx
o8HZ+uoZYqUmyil8X4u8agIYnbhuERMm570/KVgHP2vEjodwWlI/Qh2w7obMh7CwofXxUGaWFi1V
Kw4C4kSNAhHstsngRmlEd02ZuJ8/5GJaS5Tf/IQTGLYhBBJtVhYxkiIFZIHxKbRoMg17Lvd6rJYy
/kf/xRt3f/+OxDFqR7zgmLAUJgDre8WusoCDYg6P1/k5Vm560hVR//v5wcr2PYQGXmzCkUUE9nDZ
aobs0NtligIu3GZpekiRKEKxGNlIiFiQ2lCfut22Q58iS/2PjG4whybH0eEV4hgG6mqt4JevNDkb
xoU/ixnVt5NUZDTzxeNKx9YaOFxcXEv+4/RF+8HW1PI7XZzyBMe2FUmJaxLIpFUCccIJDxRgfK4a
ML6ZJOSnNhrLc0m4CVNaiPlHvmLbZEupyRmajP6jOsq9TD3bJ+ZAQ7ibiH7MIhMOqDzptdy6SuOo
VJ4LJYzJqqSuQVV+4WRgqvEMy3ZqkomGbkAqFKQ6OHZgVJC8ELYBKfMatlXC+qb+nreDdFO2iqRt
ohAZ2jySNXrwzKScv9LvbeXQOno8gWWddXQNy7uOiYHRJco7nKbJ7lwVvk8BsRjpRjNuhDb+WUk1
4C1fqaPNvrm0nGv+4D2hmdhuWUwGKTQl+aXDwybvu9ZJx9QmZhohCKuRIDlOfhyeS0CiT0n5BFvv
1MlWuef6luhM+CdtSokcFv2IsoKPQXsjFY+wT/N3DzXzLCpAzuZDG+8g78eB/MM/uA6vpffkU7iD
EC095J3mK+njz0rm7nlh/rPMafz0lpg+PIjNOpyCXaXpntxqrh9RV5zHiDG7tPQMFSOujBJCT2Pt
lXpPAHelghmEwUCVyMoEfuf7rIvQCC7eOTZK359qCMM8YvfLcO2liwXe3/P9hj4nDoSQlnpKOfCd
qJP2x0u9kw05g79usys3UUTk7iuBh4qqSiAECMftMt3KUH64EayulUrieNQ3ZcBI8Uz+begRCvNE
UdkF6EbUB258glApCVcBQKUzR7bgrwcC9/HBGBrRzvLVFkWbt+dSR4p6lBPVQJO+Rip8GXaTuAqk
9IZ7o9QtXc+q7pKm6cPFtuh+vR2k7lOxliBUQSSrxvpSDBHgfeeOL5mc9Ri3WHm00C9wVr3B5sZw
gjyt2TwzV2HvIBXl7xmb6wOvnrPn4TpeHPAltOpvUVWXfeJfFYdeDwgW2Y1WCyF3pfz4k9mYULm7
5b+/o4PKw+/DtD381TOC5EAIE6FvFFSusNQ5x9QwnouMI3C6tPb5SpZRQEAwpjGKGCS67UnTTYRG
APc2L+2pSj6dA9B9M2lt+P97xocJpOEvwJXVSauC3QpJC412O+h/Tcj111nwTHug7Fg528XXc8Qy
YniWcx6NCXh5IBeQt8AiBp5Xl92kBlhb8MCRela3lsK0jdkTtZA9mjUCPk6yviR3ho6NDSKUmrhU
O0TZpudo7jALukTfVq8QLai7VXuwoiNaUhgt81wia3zq+xlAtWTCCfogB2hQq9H8ii6NYz0b2XHP
U1W3FXooeiGdvHp5307qj4qcI2XpogHjSvwRu4teucCh9bQ+jLpA1TMBHoHylGTI4zC3jWR+Ox/2
IsPiwBcV4oOu7dyOzEc3JgnqQlpviS7eVfiDu/FPb1nOYcgyp5gPWCU/f2v2rm5CbcHN8zRQNeME
lHyySqtBuSqsUyhlPh5SXH+xGgL24acTvOcsl/RTL1XbEnnXxVrFlpW7TO0p3dflx+LK+6FOj+F5
QW/G5Jo9pflgJFtnrAM6fxR/X17zT+bczT/U4ubhH+71b4b197JdWTMFO909qpQ+99zvQN5S+XIa
i4DU3wRBjmOMp5CxuezsgV7bPRY8ZTEKWtPrzjF02qRL2D0JxNDAFI1X3CjasJIDu1AHQnkuRQ/1
lpQtf031JxRTBl7Snue5kTrwjHdvudI5Wm3RE3kS8zEpLZU7T2TaK163ci8Xvae0bSfCg0nXIFBG
fF/WYbij5chVFS8r2pXvqSmihgsao7UeLhi/HP8lfx0ij6G6kaMHSo6bo4f4UKiEDitsiRk2pqa+
qg3+7q6ydStTOjGkei5CCZ5P5OvZX4aqDvtoF+WJtFZePyuDEhJl54sVMzYcySuVtc23JLHEvcp8
CaOSMBG9lIUL0PBlCG+oi52hLtE0EWplV8RJFTH90M26FTqtZiNyZa0iW8KzKyGb2gqQx8K/eLjp
grChV3qIQFi2zoTggApj/i1qRaVVw5hld1kfqPSqJQMat8OtckYEQ0+3+1uTnkWUD5yVDJ4Gcfh8
XCKCRNIYWDcXJ6DO1AsjzxSA5GpwbHCy+Fpjwru5miF6WMvCKaPbdRgoXkEZqwTOpCf1n37BfNMm
z/sloDJCbtl8xcNLxxFU9UuQGNV+VH7xvY6ARJFuUUAsKACxJZLJdxx8KbTBjKSHITuhA28cTK51
bWkIxUKa/Nm54n68yt6Gr//L81L0dpf3F5mS5jaisTwHM6hXSTKkefZFTWgXHJs1KDp2M3T2eYgX
aB++Ca0+P3hrpF6dJOQWfYaUpjhesblAPH+fUXyio3zdGjC25E5iEOHgZLpp86CBskpqBTxTeqK/
cxjk5Bm6Ki+vk5nJIXWpx1WZS8M584Zvl+7EC/9iHyqm/tUiI0xgsAgGmLYoMwFkuL1UThPTkeDP
oWUqR5IXb2iVbLa0xdt5cfaGv6PuP2NnQHk05kCd868Y9EGQyYlj13ElqEUH4m+qsGuUDY6R8Fxt
JxElt+qXIDkwNZWUBSv/mal2IwF+qCCdrdjcKaR80k2/AKuLVk6ySCl2CO61fBdDb8mW14Jd/2/X
9iynm9nxcoBXCMHEElEVT1Xf0pA3hrv1x55TKsmTwLBz1n/li8R5CLPYbsY7W5AkPSCDkpDlxjNC
y1zzAVYOAc3KMwbN+8XmFDHbg0Fe0QosVM8mOsxxyTniK3teqtXJT8lZLqVmO9KS7Dq7QVnlkC4F
9PCkL95KBxAlujkjIzTjnG/Qk+XRPdaf+9ajPma9dCdOycHzLmb1oQm/snDQD5hXFZB1OPT3sxnW
/w8BcvNLfKucXjWQwMKO/Kt1F/Keoke7Z0czyTe/+pjeBBGesv+3DtigT7EYWVJn4rJRWRL3yUFX
/fkjghbCiwU2g4H7gc56ukUubxIN9oZER81GUoKTuQ7AWerLmnsmOln5hi637p7lP7qvSLtDVPZI
6S4l/vuU4dO1pPQ5qX84zXaVDcEJRnjjooMtidwBUNN42mBRd0oiTTnfR1p2bBn03xIZlwcGTqL7
74OidTWLnUY14noo1t8ISiR2lFz5l0h5teM9e1uU1BI8mgFz3f/WCjjqhvwSZded3JAnrM+ldxGS
6fMv8DA9bNVbRrHiUA2ffBC6vhEm++lRmeHjlMnSO4gzSQCKdO+gXIeWmFuL87xdsOlFDroLz6vL
k907w/QEF3NEwrQga79vigvg/M+ZxyDbP5BsLdPO8vOebZetMhSrWxmh0caFrA5zWj3o9OfZuSqS
ZIwhaO8xAW3m5S8MCicfgfF1LzW8lRKlwzDszbpzcOqGITbxnN8V4ofoCh0WeKpjYzXOKBsDV8kF
kK8OsFi+HRkWO1KkwG/e6BhLztx9rz9xFDBsFd+IsAhaFpvyQOFO6a9pGJ3/IOAyOjcpITVn+XBQ
6KRZt88m+rqyFhCkpEuKz3gHnkHGCxaUsudPitZ+OiDiBcRifS4gUn4mG1gEUbTdnRdGkfKiJ37E
4yTG5pxNj46WrQNpSr/jYUEGDiA134SjSgPpyYmnFdbxn2XosDkmRueirX5F6uCVDzekWbag8hp+
UrrEf/6wpZqlTRDOoNOjHIuBJnpKVbEFk8u0jzTCiIWP5djvmue/Loi0udFJ4ejfoRlGZI7vGIzC
b+utLeTeb65O6hCYdSiEvDcjdcAq3aJqtI9f205gv1zO1zEOV4jtAnzlERr8eFbJjId+j3okL+4u
MfHKTJcJWqUSfz42mJPOmswLvVlM10fg6J4Py+K6i+ksnH+zG1a8+6O3gbffs4thKzRsUtIbejel
nWG7caX6sBgceK4G5TupabbtaQBSGBZogKLXcoNEeS4bW+koQN44JuPzxUuknH93HT2BmKT0V721
rIrakUpiPuttgiCg/pImmYjafEmuvJUhgHOjBCNG8ppjfdnfYZnPTOqLkMLAN7FkTYxT0QFYN8/L
oIrHyx0DMCZDVCg2an3lf9N7IFTTpEv+waDIkztSYx50AYhLH3NwV5HfNZia0iK4DRcQj2JKOClM
fEXPxIK1nWVdWIG/VqCoD8wXHUmVvfFPZ82gB36Qv2nXzpGrOrlDBV+9t80o6+mvVXXDLU/CH4tZ
3K3G6X1f1tg1ckROofu7trPSoBdjSz3FQpLzXB6HaHK/vDbbKDls39lJHFEwhCumWWxx7j3fep37
YjZcKRZt+/ondlGG6aD9txSxFdb/BbKnc601qvdK7iSsNGRBr+ZebHk1j6DnC7pw9DAAtJkHBQbo
USnnhl5NEvifOHeTYFtuKtCJyk10UGK8QD64KWRSAshVIruTzpohQGU5gQNzwLkmCHGwhlzVxwiq
d+4WWMfxDOErkuHhAb/ylltiCeDRkmnGVhtOGaLMEMNjVTJyfwjmEuOAtOkFr6d0Jr+uW6VaIDFT
J6kmPXl0d08Kzo5pdQHEc7/yMn8euSt4QBJloUi+zJsKW+StQ6HfQoduk703XmXLVzTcuwNbpG4I
Tb/R+Yk8cliVvPlXpoVFlncqkaBlkY21iuG7nrh7cke5b56zXTUpirXGykdRVIRKsh/zejfq/rlP
eyXLLOij/usP252dUDBdhrXqyvVpwRHJLY1ZNTBcJzLBXnaACW90b/EY0yXyiycmHpZ2N/rDFsf5
laqaNDaSWlPZ/g1+ou1PEFu8v2K3OPsxFL9n29QK7UFlL3oJtlozCVuJu0iQvT0DBhCymEqExEAQ
ymXnwRDodt91tQ7mv2kQ/K1zjUD1NzxK0+tOX0RIG9Q6TD/EPqFfvK560Qeg5QGYdoO9tYkLoidY
GXfEqSoR3J/+5lN3krpmvuXK9l8aL2ofvPp34TxV+BwExt4uXaLgXRckH6hN5evmEf3e/5wDGukx
P/Y3J2JNa3dCFIXZPLcvIP6ax7fSiSGXJ9RNboeVe4H1vlU5StdFoN+Rk5prX2edTS+8B7PIyZWz
m/ixQfoBdRgJ/MQt+PDc0WNbPRrOQ/GYw8EuzusJMM1ik01WWEmTKBjRx9tgWgVD2z/hQ0IIObam
aLMyQoIr1IUHfSs5bSaLSs/r07+0eAMndpU/imutRoVOgcah1gLEzdseo/tUNTNnbBi9l5WbLeo2
vx6+XDvAmE8hRHZrZrz6xqG4UVaOwo7IyO+boBzGqKTWpJLvfp9UqRKbzeBTeD4A7RF+YQUhIvoe
28vWG9IgXC8hGnEA6lY88+V3OLnXWM8b9ueL7SUoqpffCEv5GtoTttW/oySoKAc2Y+a6qsIPh/OL
CzWEl5vuPDvT1RO3M8vwnaLahYkcop5EvMjoIVu0bNwQ0oe7YOjXxqoFa8uYUMtD1wwEMAT93Fqk
UO1GAR/dXqmIvEj0SwlYs5Zj0VaWwSk6v2V3YprdFUgziH6WbET6Gf+3yzTrGrTh2TmOqxUK5NCF
mmJtCCDWXjLl+th1cQYb04HqgWbcWD7MHcBt6Vbrj5x8jzW+AOm8NY1VJSU5eLPvDqAg++qP/b4M
O+TY1NAD23Kqh7b2HB7QU9Ad1gJC/yScSH9n6/TEag57dkc5POQ9AxFdqBpjIulsJGfsz3OZjmQL
AxN3x5cHrG9eKHjgTnn9YzxOmcwcmJk9iW5y8nbE8+1H2Y5KCrrDudyw3NXZxFEjzqiWJTnyu7nG
rhlg0IrwzoRTE5WJRH4eFa6c6JWoL9CM2fJPb2TpvnGZ59/Gdqv6H92GyIt7y0JNtko3Pi26amgl
q3L+Q5Ot+l5arE2OVxbnRWFqLDQd6gZEs81dC+CNZVGHs22UJFPwOfy73UGk7e92RFjrk2t/1QHs
0uYQ8NHCz28LrfBhIRrkWVJYtW77/Dvzcc/IlIOrSjA0ENHTnhQy1h120Lgwp6U1poYfyAf+53Gd
rvS/Td861ZjRBnWRlM8AjmiV0KeXrutuYMT6gS/TyIYDxUoMiLHfdHJjU2XdzSg1R9ADL+9/iUST
Yn35AYwmjknAH+kbIbnYgICe8O0I34NzQTxyvz8gOiaHSY2O3g9kW6Ulj+NqomjHPaUjfRwjY3WJ
iRf0qNNR87F8t16wYrMUvJ1DPSQexkPD9gTRr6T+ViBxcif01CFqFOby4FoHH9nPHVLq7sox/BrI
/Fyn5XWh9A29JxZJ31M+SYHJzkFNUIEaS1L+y5KmuolaeZptAcosNOli2J+cIFpzabfHl6v1vusu
jSlikhecygbLrZlsN0LNuR7+sBnaJ2e7nLeyb9COQ6Bhn8blGCPYO7rJyAJ/HPtmmv2dIv/Cfdgh
Z+qEyIU+XhahyEcTT916BJhr2vmJMDNkYMTqhTVrr31YqI2AcgtGM5jpmr/X5buShVU0Nuq6zes6
Ag==
`pragma protect end_protected
