��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O�k}.Ż���"�����x�u!
�*�*����K�f��\ �<��nFɚ��f�.&V3�t�_z����RZ �UP'���I"���U�ϓЯK�݁/�G�5��#
/���R�|�1{���_����,$Gn���G�M�J]^e��Zd~;Rb��N>@���O:G��o�)��A�ڄN����z=$��TD|d�c")��8��|�N��BK��1
i.6ME����˹k�9�ʎW�3���<�?	�}�K��q�� �ٖ^�O�݃�g2h�nO`�=�Xw�Qn��x�";��%j�ʅ��d>ފ����`9r� S�·�����x����҈QT���tZ����-D�]y7@1W���㿛m�����E���v�	�7[���ga�՚O��0�L��o����4sA=ߪ��a�uD*�E�����ŐIb���HGK���;��Y�J����<1%w�,W�E�.`�z%s-�T=��Z�ȱeԉ}?��E�9��Pa�t��T��*ޟm����̀�z�P��`�8Q���V�5�P�R?�R<o�X�Ď���c;T�c���Z5m�t��Q �w���n䇒���S������,H!�k�g��`��
1ӑ�f��X��BC}]���5&��֗�[�|��|�Q�48^��w\_��̦�'�	������W�n�u:��R:f��R
u?"��TsD� �]P
�:��=˼�r����7�Hq�c��B�J��|=��ֲ�s�~)N���I3����?�x�X���Sz���[N��)e��j�$���@¦V�nz|F-��6���F׉n-:��A��Ï�Tҟ��J0�+?b��t<��]s}/G�^̈PȴN���l�����~��19����q]�����4&"[ḫi7L:��G��Q�IYzQ�G�	i(!x�yLI�>P�ҽ����M�|�8��k�s]5����Q�!��R[IȾ��}�jl���3�v�Ѕ��e������U2e�C��fkg���B�b���y�[��u�"r"�nP��*R�>M� ����E���_���1��+3B"�(J]e�  ��7�M'Q�S�I�Us��*]O���u|)E�5mx�f����J_�P;�?�ސ��u��@�/�벷�(�Now�ћ����N�DUE�kO����r��4�zo��~9���u����y&�lGt�̺7��� ��$�E�wWe	��^m�0��	ł��t˒X�Axw�Vg�n�Zm]�O>�NS�T��^J��2E�E;M����Dp�e*�K�72>��,�u��X&�CP3�,H��U�U�D�T��'�z^ZM��[�G*ڊt�&N��ܐ9L��/QA��l�hʖb��<��
BCŅ�w"9U�}~�&�$��J)%?R�� �Kw	�|�<a�<�n�����y���t�+ɉ�ut��2�+^��[+z���#�w+�tQS�)BHM�����_r�� %bZ9�o:|�O�Z�1������T
���Y�18W�[�@e��%�������,X�Py��#<�O��d�r�O�SUi`G��jc���kld�P��n�S�X �&�ȻK���������F7ؿ�%�� ��)��R���,��b�穉Y��i@�\��?�%[X�!ӝ�(_>0�W��[*���B�*/{�Xs��mA5��8��Ѹy�{1�%�_v�L;�9S�;懲&5�� ��������k���*�J`��,���a.n^�)ݲ74�6�B�vzt�@:�@\�؍�R󪽷�;J��h��R2`/}/�m`ct��B�#��%Un��5���nR�3/���0t��}���G(��1�a���w$a���)ķ�O@cc�T��wC�+���(��_aD��C8�t�R��|�Ջ%2v��$�]�9��V��<9���sj� �R(Fٲ�'��*��Hudo%���aL����3����Q�<Nd��f�8o=Y?;.���c��[�g!�)�K��B\b��o5�J�5��j���BDVՆ��y�M�����w�BIJ����-�>���DE�X�
c��gDL�N�}��Db����ر#���y�sru"��9�w�/O7�*f ��`Cq���j�7��{b���������3�6�����>�nc�G.�u&��w�qJy�du���#����.�7Y�`k�U���œ"����ұO�/�����K\]J�{?&z"��C�}��G�~e��d,�u����� 9��t��OF7�
>K$/-L��e���:�{�VE�쇠,Nǫw
�Xj�%�qg/�[x�����TK��Ua�қ�5��_�����1\�bn�W�g�ιs�M^��d�M�0�k�������&�ZP�	�ܓ.n�3U7_��	����^��D����nc��Le�LV9������#le������m͋]�þ&��d����ʫ,S:���G���<WR�(��U(�!�2�B-j�K���hR� Vx,�j��/5����Z��!��x�I(q���_���<z5"���,�}'���t0�❝u@ǌ8�e��k�$�Ғ����M)WM��,hZSt�F�2#�z��'.
�/�����_M:B˩=���9r�s��W��C7gK�/��O�1@�ȷb/�uo �Te��<�g ;zX����J������p>xqf2�&�Y��	MB�@�W�f*�-���g��n�NK��[r�JhFes%~���չ��ǖ�e�^�J��6���c�]�9��kp�w�%����Jׁ�p�dxKxD��W�|�L'�����Z�Y�B���JAB�7\#8D�u�aJ��I�#;��u�������45�ڋb���c���u��ܮ��e�=X>�Ï�u"�e<�:��Օ��LnE�.�Y�hHx��5�O$��,k��%�BX^���l1�&n� ��Xa���܅�j%7�H��G#�~���O����	Q���q��r�}:Gԑ������9��vuU̓f�Fo؃� r y>�͝�y��4�h�ؕ�Hr]�$��ׁ:���=u���)H~�	h�:V��遄��P����Ѵ����a+��d���gkb;�O	��6�[XMn>��Zt�'�+��!��O�C͟6�&�o�߭?�;j��-b�Y!d��)�X
F<�Ih���:��@S��υ�p�ֻ2ʼ専�M&���x�X���K|��:�Jи� �Q�B��(5���{�b�Q���,��W�m�^����t` ��uLx"�ALR�]Y�W�&+�o�X�dk�ԕ�58X��y����>Y��:�"�X)�p��Ds���SS��}3"��?�؞zDP�p�θ�{Hyu�)5%� �FwE3M��utؗ^��Z���|ޫ5�I����G�1+f3ョ����ÈB���<Fp�i����٪؈*�X��_\��CI��H�&�N�|��ѫ;=��N��+Y��׿5%kR	$A=kR}������Hz�Y��W�UA8��ܰ%��%����؀<��qt��F��T��&�:�W��b�@� �Vฃ{n��������ׁz_��;>-��NVit���cP���H뉂�C����:W�pv�]�w����u�Z!�l�I��	:�ۂ���̟�b_w��"�Q�_��+�=sy��4��|��X*��i��NK0\O��,��ɮl̼����>��eNsy����^}Z���R�g����H�8=%G��nCB줲,��.6��'S�-ek4�ڭ^�^l�$q�)�wM����Û	��u�*v�+x���_�\/}v1��|����=\�s<�Pwn�a]���tײ����aY"��;O���N�$ե�e�����SK���n�|j(�W����4�Qsq���-u�&[ ��V�$4g퐑8����G�c�t��S��Xl⯎��Հ<��5�{�]嬩�X����X�ãy���V`�D��-�.*O�������/N ����	�o�FD�|�`���ߜ�:��>��&q�}�����$���绔׺z��S��F������� �_) �~ū���g�ge��ecuƭ�7��v�5�jJ��~#����ۓ���5�13;.��/�����y@3��㰼%�VKn���hdsd���xH�r�S��qs�;�����<��t+����������B&�)�7q³z���V��$��Fj����p�,�)�.���{�pF;r�Z�P�ߓF�9{l�ܼ��� "�&���ƃpqDL�D�SW@��|Y2�dd�q��f��TcZ���K���'J�c~��T�VB��3l�$�6?a�hi�C~Å�����~^h��� �EiDf]y��5�Y���a"|+��;[B���g�C�����0�s��f��� �e��ȕ\�_�>d�Ϩ���ccj*�h��	��a�be��n����ڦ�Ug�C������D#���A3@�.ة�A��jw��UZ<6�p�0�?DZW	��C��O�F
0��"LȠ@�U�ák�[H�]�}�#n�7���w$X}SL(u��1u�Si��v�.��j�n4*a686�����+x&���ɕ����Q�ĉ��b9 �O���1�
�q�G��ޗi6y��ռے޵j�v��� ���p�n*���j��gB��#8�t������5�"*S��<�D�r���M�ǹo��y�Vj���M��t7�!ݑi��K5�B��R�I1鐗���c��7Ӕ�'�P廗P/��h|@*.Z�O��N�S��B#�ø�~�M/�O�����8фϖ�"U�˦�Lc���kP��v����9��)�?����]�l=��s���~��-�j��@\�f�АQ\aɊ�ǖb�sF��E1�^n�➮�F�=Q�͆��!����u�6~��h�v�6�vz�T3����r/�."F^�ߗ��%D�)6aJU����a��w��|M�`R4��<�u���X�)����&��L���i8����HM�>[T�-��?��p+�++r��$B
3
:��u�>�)>�Ja�� ���0!��lRm�m�+�rf�j"M��b{���K�l����"Q(;�zN��/�����d��OɈ�@���	��Cf��Џ��쫥�.�����e��o��� h�Q��*��Fb�L���%� �b����'L�,_P0��[��"8!s�+W��+U���M���:�E�~����_�E�V�$�>a��$���+R�Z��}$��ř�fn��_$׼Ă]�q�`����*:���2����(�Kgї"mb����:k��o?�j��5���O#Ε�Bp���ch��4��9rI��B��"ɆClS�ccb4��?�R�B��$l�0�(LĆ��**��� 9i�2�+(�S>DmHZ�I��>�^A�"?��&X��~+��;
�����~�����F�t���
.t�pwJk�!=�zz�WW*p>��6(��Z�ě&��+D��dq��@�`;�m�1��s����̦���ag�OFi_��%Ɔ�|R��kB��ޔc�$���n��sk�6*��@�DY42y%��77�X�P��8c�R|��@�e�z@��h.
�RD�>m+� ����0��Ln���ua\�_j�[��)D���H�z��f�&ͭKW
�8�Ηc��V�[&'��X#O�@�fLk,^s�^kv�J�@��V�q���8o� �l�/YWJұ�S�d��l���]O�?ی����x�q|�����B���(�Ƚ�s���	�@5_��\�ٔ�$S�����\���hJ�F�6����ˑ����ȎO�	>T��D�h~r��Į�����q��αf��C�o��3�K#��D]=���o��\2"�+.�J��Q8��t
e��� >�I�FÔ���va�Sٴ�t���z6 z�a<?t��BT�k��9��I����&j)4��c�^�Wn�/��x������ P��r|d�(���-TF-���S[ٿ��O�"�眄j��'�2G�fE\�9��<�9��)���0`�<�t�)�Ǵ�l��W}�ث� 5�]�߻tzm�;4d�7C�Pqze^n~�����NOwl���4� ������J������~�'�K]^�m���`���i4TaR�x.�p�zn���p�'� ����֒��s��ǭYU����mP+ǌ��r��abYh�j���0���X� �U_�
�R�֣�����.�-�Č�j�pu�\L(մ�您H��j�v�9E�X�Ar�[B�ta��ߪI��_�+`��RR�K���������������xG-C<��>[���R�����osX��GRѯ���7��f�l,k��:�R���v���I�����@cQp�#�׶u8,����a�}�$J��{n���A/i��2���b�'�_ӗ��Sl�e�H�q�������t�ty�B��?d�7M��k9�ٸo��%h8.��qE�JT�ICB�3����Q�B4��� -����>������gr��s�[��s�~&��K}��9��Ts��@����f�ӹ��!�����G3uv�F&p�)]zYn�y{�U�U~"8�n5`S5a�}����{�o]0'
q�[���������;�v\���I�+_�N��({G9YԂ�ba��3"`L���=�f�74�O9T��B�^A�xg+�D�.��C7��J�=��Z����,g�Ԉ�B���<~�S����s~8D:�IR�j��9O��6Ow{u���J�$��eˆ�<K�d�lIƋL"F�վ4t"`�쏮i_�#.�yrR�������/X����<�ǳ��`LF��b�f�ˠ�s��Y������\� 0UB�b��T���j���	6lP����9���{�B�)�p��9[���Quގ��$���Ҽ^,Zj*w�g����)�t@� �����-ZT�Op�Wo�^.��tX��f�T�L�+�(��ʤ��=�ҏ�tm;���	�z�Rc�ͭG��㥝�i>�=�X�,�j�8�E2³E#;$;���<����p&�ds�@U�X &�c9Y�B��+Z�c--]Swt<��d+�dA�_�F/�s ��^>���E5�Kh'�Hi��3��[?휷�Ͻ�������!a�Z�m�v/$X��8{F��q���Q��cEo.�DYhg+�$;�U�\<��F�({x��b�c�݌�ZB�u
��C�a�ג-F!g���ȸ�r�4/Z��إIͱ�	�QɃe�-�MÁN�.�������*?����!w��_���$��u5��x��YݱP��,]m	s6������^�]�O��~T�c=u;!��M��Z ���Y -}:�h9kEh��i�R�vij��~S]t��ڻ�J�>��%%�,K}������� |=Y�G^Bjr��0|�i7���6a�����'Mu�<���l/�r��̩���&�;3ٗ�JN�Dj����a���� Z~��I]=�d�q�>�_�G�&��ڨ�'�p.� o�X�9�����:+=*��Z�?F�εpW�0%�s��>})�����D)�>;�KT���P��a)�?�����̸T��Wi
�g8���fn�@&�lW�0�/�+55 ���ȇo�����R����*�z9&���1�r�b��w>�t��v���û_�.�b����%��Y�P^0�J�G�(٠o.@���?�4�1B�[5ޑ�rQqw�͈*��>X��é�'hf�e�\����gߝ���(���(�� �W6�Rr�)��F��e9���|<c� 	<� }Q���ˤ�KN5���܄P��l��^������ġ?&l�Ѭ�}ŵ��)q��V�+��`}������Dk�;�U�w�8D��[��҆��/�
��m��j52���z_YE�d�#����2�)ӣ�Ν�Z��I�u�""��ښF�j�)�b
I;�mOA,�r���ro�˰� ������ۋc<7r�3�|�}`^��S:FL�m���V!��aw���H��HZ��ٜ
�r��eNSRz!OV��p�Tcѯn_�-��c��V��@X҃����DByk���D�q<J7�����ξX�u��[�sbU�H-P���1`�Yzy����ˤ�Sm���t�24��]��7���p��:O�pb�@��$��b)f/�9�)�_��0܂
¾9�<�|����u�T��A��gp��F�&p|�dw躺okPC͡��������7���O�S��*�f	�����ru������ZV���Q
�vq��_��X���><!���R�o6����ѻ� ��U�bq�5����p7T\��/!�q�?$�����FǾd*��tL���|8[�Ep��7��\�"n����쑹��(ߤE�&�Dx��:Kx$< 与�̅������ܝ��l���;1��E(B-�����\�M�JY��Z_9m��䗭��$��x���ǚ|���0R|Ǽ����f�\%� W ��� >������;�+��F�S&0�0�n%w]':xѬ�$�^+��a�b���D3����8	J݈��O��n��>�q�|s�;��/���$�� J]��v��װ�I�-�����p�Uh��De�XE�K����>I���4V���Th��η��yV<���Y4�LU���dGS�1,+K��\K�,�e�m?U��7�U�h�嘟�>*�@ⓚ9Y~��,s�@�RD����_�=CR�*`��AdB��u��}��B�5���b�I�Q͝@��u����5�HW��������D����	X�"�<�'�׺��:�N��'oW�K���|����i ��Q����=��?=	�A��h��}nH�?��I��I�p��p;���H��� �-V'V�i��S�kݪ���\���_�쫦u&k�\T��R�դ�K��6Mg���H�2��֫�w�	���5�4��5\'y���/1[1������dG�SU�_zofE�Nn`��o�H��v�|��� ���`��e��T��#Y�	�#���-V�A-�X֪��5u��8|��CK��e8=@2���o�u����jȢ� 2'��yn����߽�T��K��
��Z��d�.J�R��0xDR��Kik!F��'��忮c�ɋ�<2����/$�h�L���ޕ%BR?+$Ł�#���t_�Q�ݦ��m� �:i�}FV�$!{����k���\��&u�Á������z; jii��Pq�5�r9YvWQ���sG̀셷� ���2��H�o�x����iӻL\{YM�4�K�����5�hʉ�I�R�!P��^~����h���D�s�J@���i��9�G=�^�;��(��K�;��p�q��!�\a�q�R|dO������^�`3s�b�ג0[����<��c��>����3*7�4��<�]�Q�*���|#zϮ��:�s#7�x/8#�ۘ���o����ۨHޒ�#�0�E��fʦ�?�$�V'LtSѷ�s=y$�i��j_�:N[��Sj��o���a��?ǣ��=���:_�-���m��ie#������}�K?h�+J�wn+��E��=CJ��&�QK�A��,n��T������}��7�G�?�ފ���þ��-�o"�T�RX���M:��9.��y3(��K]���W�M�[(1�nYҩ4�>ع9
���GyV��EG�kXu��J�1#ؼ"ER���'b��0b�aQ|?���@�Ɔɜ�0�0xÈ����(�h�����*xY)��m��]�[�r4�h)7B�*ň'��pZ����ًr����#�o>�(o�y��-��W�S�� �S���^ަ�kz����F7�M�.�[|��Zs���3;^�V�G�ס�\8_2%[����r3�~h!S��D��5^��a�����\�m��m�m����P_�v}��a&˳/�c � ��0M��Z�ϫY�˩���e���tQ*!�2�3�%�yU��~>m H�{.:��k{0�dU�U6$��4�����vD����?�����u�o���\��w%��4c*`̡�H��]�j�~���4��է*��X���岙~���U��"���_LimԱ�|���D���> Pȏ��t�ڤ�]֢��-��k:������/�tU��J������K���OI 渁�����Q� ��5g�a�|'�ƌ���" i��(3���.#
6���FL�؝������2��ݒn�5z����Nt��t�S [�����/M��}����N`0�F��3-�+L3��A��>��ps�U׳�d��EqO���&��e:'5 ���+���qD�;i���$'Q>ޞ���US�PD��lY��Q/��;:P�pZo7eJA���(��,����+���p,u��� P����y|S ���g�
�c�%�c��zA��4�4�`���z���F5ꅻp\�Gh��k'L��K��n�ɟi�0��ŷ���Vko��M<詳 �z	��I,����%�m5%HrO��0���Q{M����4-���<��^�]7�a^Έ�+�M�S�5�`�ygV!ń�m���A�o�n�<�-��:�hu�t�Gm�x�8"v�������>����mOQ�A\O�F/9� �˾�-p#��o���Ƞ6�B#y�.&��zH�k��j��P�����"�2�6�514�'��ÈỜ�'zA�1$��˺3b~��h24(����lOK��70-�ҝ�uNB�\/7HT�)-sOM�P<�\�<`P#��Hΰ�e��7/c�p$~T&�ft���������)_��q��9� ���9p��U�f�QsUkP��.�q��1}������W��3�9N$*��*�	xy
g?�})���[�L��^��AuIpy*FY� 8�V!}�����cˈ��[�_�_�KQ ,Hy��014>֮e֋ V��	1*�fI@?g�Bg�l��B��DgH�R��ȨtL\Sa ��YN�y��H�P�n�����D����x>'n��W\E����6��Zo���IԽ����"��|�?!�=��d�֣g��Z_�����l��%�p(�a�Y�+��]?R�5:�7�*F�^�t���ʔb��c�!�(8�� �W�����8�*𽼦���a�)~F4uō����Eۊ�����ˌ�q�E쒆s�:+40ܥ[6�X��Y/{�2��'�7G�'���:̺#�WƂ���C�T���f���p����w��@�Ӂ��9b���)��V5BK���|X �tU��X*o��눈(GB2LbEt�b|T�b����	B�y���Vѡ7�Gq�V�b�`�Wտ-�J!��Q%��8�_�i�����Zix�|E�k�~;A"pA
1�8��z`�qc�Ż�]��(���ȟx��I�x��eut�*D6�9)�_�W{<D�R7�G��B�oyq���A�ց�bԙ������������I�~вq�'xؓ2���~�bp��YbPa�NJz�w�J_d��s��ڔ�/6:%�.��ӄ��ԚN�k�Ѫ7w^��L���7��`��u,R����m����uK]������(W�$ �{��Meb�:'r�$x>�B�j؂���	�:ND9��}��dݛ���D|e�ֵ��m}���#�,.#�Ac/�@�X��s��D/�]#|e�~�妍«�h"�3_���~o,T3v3��j��H`�P��vM�W�X�O���wi?�@��C(R@��m1�#�Mm��?"J���ٹ0��[İc��n��h��ەL��:K%��GP,M0)��RO���x:Ǔ>ӽ��f�՜���{D噴��؀y͕�ѺKCx��z�n��Ѭ7����� FI\V	z\��(�:���BB�"�_[���g����U:p:zE4
-2k�ØF׊4�v�� +�g�]��UR�byy�ζ��p���_2��p�����;L����5|S������5��`V�4f�k�f��3q��ckn?�73P��~J��2�����gJ�1���ԇ�W���b�v2�p�|Q_�Φ���ٚ��)���ۇE1?�s\Ύh9���^���?�]�t����5��,<�l1~��5�A�S�9E�2$���#=kDrHTYUB�w�k�/�.��E��T{�5q%u������y��U�fu	vzWY�-ڧV:��f?>��7�s"���nlU�V��*ޏ�\�_[K�t
m�'{�c��;�,:�4C��:���,U�m���d��g�<#<��9�.����r��s�;����� ubV���P��t��|K������¼�4�Ԯ]y�%��� ݯ(���A~���ICl�5Vò�]ǻ���FN(B{s���H��z�k���sp{FVKf[�@τ0 �!0�D��N�ǉS�����q(��qq;�����gB�"��Կ��  �?�K�|tp��
bL��e���\���W���V	�[v�=]
������'u?Ӽ�܏�$��_�R��`JL`���v�#�e*Zb���8�0�K�����Y�{}����̾'_9a~B�<�Q���	��ŏ�Tl"��8����u"*��c��!,�|��V�኿�c�O����4<z�3�P#���Ov�H؋�ls�o�޷�b��Pn��^�[��[%�2��ۤ���It�1n��<Jo����H�f����w�f��;��0�{e��t���t]���)��l������S�V�'������"�k�6|�x�w1�'���7^�� �-4�͐6j�p/��9���n���)˩���Edq�5������g:!�������2Y�{,��c.�:S�x�F$ʮ�tK��1v}�;��4�і)���m�W;C��9��D!H���s"W���#����R�-즩o�㾉�$����4[�^�Vr9:�g�P�k3t��6�8笹�n��.�mjX|��v;���b?�Xe�읧�2��z���.�?î���DN;5|4kon,�����Bh����n��<��Qt�����p5�u��G~ɴ�d�CG�M*rEI�~ꤎ���)�R�{ 
��>�_HR�Y�2§��Gv�w��[_�ڿ?z��gz|�g�+�����uf��i��ߙ��u��>Z����<�4��^~��:=J�/�V�Z)f�r���Ε�'U�J��K�+��S�C�XC!]�c��oX��m���So�-���J�Y�\%G	Na�S���g5�tb�ׇKV����M�2/�#�ͣ!~�@�8D`�jr��A,�m
�\E,c��������qr-���t�{/Zr:�)��7a-{R��I��ki�fU큀d%��
���d�Xx=Wr�����s�_Cf��$}��L�;+��nN!�/�SL7������>�����]�xb^�HkJ���ӭ�ef3tӹq��=M�Z瘜��Y.��G�`�*���P�R�
��Lw�a�d;t-^�#�]������]��4�jL�.�����j�G,_e���A�� �l�pj2_��Ժ��k�v,�6񎴚���>#X �t�L
��H[�!�b��!��
T�Ѫ%��t���
:Q׶�Ey��%��aS���
�A�<ݠ�g*P�����?h*v�)\���[&t�J$�pc2���u}
A�O�t{�J�!#W����vBT�]�f�ŏ�1	�1�̆�eV����n��c.��b���f/����޽4X�FR@�f�P|)�rG"��:�F�Q>I��Ļs�0���:��?�p�Y�B���l�7g0��=�0O�ͬS�e�B������	�"��lS��3:c��!��< +�`ŲS���Va�P0��AR 	j��P�U��cc��In��I$�Et0g�~�Y� �YȲ{(�,Y��d���(3�͛ 8��1�W�\[91БМ�{)�=Wsn�c���F�=�XƗ�^Ӂx���у��]�G����Zm�uW�^���Y�)?x�E<�n%��~;1��)q�4���� ?$C3F�v3�ɵ��	O�����]�%<֜f��;*ډ�#�_)��Z�4�C6�$Mݽ'k���t�+e�%N9S	�	��	2.�d�| �k�v_�:�5o�ډ��xM~��Jm�f �5*��A/�\�r�j���O�Iy�-)��L�[��0��Ţ{$Q|Sf7�}�-������4ip+6������}��:]��s'�-�<z���VV��J����l&���m��ToF�쥽���-�/�=�U޻����}�����Jl�4��Kʍ�1�y��@���_�\���2�;+�u��{��//�Xd2#=y4�7�V��>��£�ߩ�"�W��w�ۈ�m��Gfé��`Hh��`�_�?Q���j�Dc�"��2>'��َkc�N���"��l���8���ȸ���/͑r��j�)�2�k��e��?�)���PI.�b����|����j��D|G: 
��?99Z���ݓ�6#�ڵ�fM��(z44gӎl�V�勺�rK��԰�Ƽ�߽E�|8d�d{G�+f��{�*����k�C@6œ�%���[�~���+����4�Ub���ר��
0�[�$^��jvyb{�m~�\��Ǜ���+����G�>lR�nK_�6�`�cC��5,���@$��B9� �Xqx�
���\�ʍ�����]���+n�4�Ӻ�ϳh��C2�x�=^ *.c�.=V9��l<-��Q�(��y�lyd��n���<����>:{p� ѐ���çI�=؊�����W���V5�5y�7�1��'=;��r��8}8y�o��HBխ��_���Y��#�L��#(��%˫wA_��Z�\��BV�NJ�aEb/,��+`�:�~OG8Dވn��4��&�x�`x�@�!�t�ژR�K�6,j% ��f����K��%P"F��o��6
���~�P�S��g��h�1a���&=�wfqƜ�ty��T�z�jB�6n��=�����]=�CnF[�uZ-�E}��5(��)y���׹m�(�}%,�u���G�p��Z��ۏ,��~CF����!JC�O�:�%UG���U��"���Ţ��9Z��į(��xŨ�jaۈ
�ɀeM�T�6ߺ l�>Pg>�7�����u������r
�X�ɻ�lw��p�G�R7�Ec��T�#����D^~����#�>-���a}�6��a'�F �$-�dڙ�|k�����D��Ɇ�q^A�P�鄴�ؔ�f��I��ݢ����� ��o�ٓWU��v߀��S�L��}��}w�ت&e����	�p=&K��}���!#�:���iw�7����Q���,#`\�A��2�b�+q��,�U^�) �p���ݛ4�,���.:�����2�ڡ���Cu\J�!~�1ড়�Uѯ���`XL_S]����X���2Y�Y�d�� ^�d���㰤�^�lD��V&�Z=˅{4�J���)��V5�J1��5~�x�LN`_�e���R�s!!��-?�HhB�۫㧝�x�161���L�P	��1�$Ed7:uϮCj坠~O��߄��v~�;Ec�F�W����QjLU>�^��>uݵ��BG�>Q)��6�۫���^\��	�ݳѢߵD��y��]�/m�fHh&���� h�:O���ۏ�nՑ?���j�e��Ցaz��[�9P�|F'���4��c��s�&+��yl�d�����5��7��V�R�����~���\"X���V�V�ű6~m����)�y5�J6-K1�������/�x�>�(B�ؗ���]Iᙤ�&���5=���R#�Q  u���e��O��f1���x���ݙUm7x5�A�X��6#��;k�\4���]%3E�׸x�,b+	 A�d6��7x`��Ai�Qͨ5s��A�u6�#����v��1��y�6������<ʋ�yn[)�����,B�pi�Y
�ֲ������Ӷ:ģ幦��x�Bʫc�,��V?��C���R`��I�Zت>n~<��y/8J�wc6������rR���Ci'��k� ����E�Q$\0�T�w���Y�� ��%Ô�Y�?�}i����o��z�&�ĺ��aE)oyԿ;��c1*�s^��\C��6���Wl��e+;����J�I�������.�����}%=>�t/C	}F9ɇ���0�9���E�M���l�ҥ�틫�T�$�9��랲-֓�T1�M�-�s��&���-�T�سJ8|s��X��l�}�id��.R���T�����-i�����S�}tW��/�\�i9�d�-@��]Op�]Ԃ�<�/�)��m �VPk�'`�a`�x靜�
ѹ|AJp���0j?UN$���HG����"���wI&zj�f<�Q)��ĩW?�EXF.5��;��������T�Ѡc3o��a	��-���5�+�{�A�5zG� rć��uy3�#��#M'�gm����fgL�1��f0�����������qE����[]RI`_n�gKX�9K״��Nt>Z�#�E�r��][��-#9�v��v�������z���x��2�#�$M�I	�֌f+�8O��Z��p��*4
ȟ��H-�*/.O�}v��]/hM"�⋴�J��F�+�t���9�,���
5Y�$�-]�nl����-Wi��Bc����� �ոR�ٴ����۷u�"�	�*e ��%t:0�6�`\n����N����=���yLn*�-�0!д�M�*��ߡ���{r�/X=rE�/���=O����(ץ�~5%'t����p��Ii�%ᐶw�� PT��P2���X�h�e\���(�:C��[?c��v֗�;��޳�
ۜ6��͸[
�� ���+���3�1�n�u^�Qu���m�D�;DWr�GL��o�Ñ���X{T�P�v�]BƼL��ɇU��4-ׅ�ޓ����	.%����J�B��6�O(3�����V׹8�(������u�M�eY���1]0���v�I����՟���l�|̨�g�a�9�$�J��Ked�6�,�0l���~�up���­�]��a�1�m�~o��l�2ښ�K�f%�M�:?cN���)�����b���د��gj��o�8
 �Biʽ�eJ9XQ[Ǉp�Q�v��tjE�!p@EHy�i^�4��6G�8��vyM�6�}�����Fk�
K�ݶ�'����l^��Gɿ"�dYB쓋�)%�ÙH��«b�i��)2%2~�g�����v9oY��F�7���-����+��a�Z=����J��DgYP��0G�N��qu�y;��s�_�����ᾥ�+e�N���!kt��i�o�t�du}��ck�p��ƥ�7�5�uxX7�m5�M
v�'vy��̇�ه^�&?;�$�®�P��>^=mÕ����fգPp�w٬p����3�"w�=��	��a�\�4u�$��p��
��yG���L�TҤ�V`�j�q��j����I`w����yWͪ�)R`Ί9/�	������ͧ�/MR�Ş����c�}>��%A�>ZG+�M
*k��j��0�M�;���D#31@��9���V�d�������u��C�v\�'��-)�����y�6�fZ7'��Ԭ]��B���r����xh�q�ÿ�I�d������&z-\6sRw+��� ���d�@��~�7KfeNVn�de���ʖ�����]q!"!��x�\�3i�V/���qv\ٽ3;��5�:F�<
���y=�<�����T8C�h�}B&:�۸l⏭����hf1Z�i�G6�N_��y�B6�L���4t��.���37xh�NX�V����(�̿F��'��Ó�h�@�@�1��}��?i�k�51��-%�Տ$˴�.%�(���)h��"Y��f�+���w9 dQ���}vс@If5!i�xO�U�T\�����x˞@K�+0�]�uk�3��c�X��V� RɂC��g�D�����O(�[Ps��MÆJ�������dボ���MϦ�Kg�'���^B���{�)� ���1���|F�k$�ۧ���p���Q2j����M��;�>B�1���X�u���W�Q�&�[4�ApI���@#�zx2�@y�[�T���0��$t^`���~;��Y��B��~���?B_���W��GIIC�S	8^W@��.���%�7�i�'5ezB2�����S�NTi�Ff�����h ^W�͆�=��pD]�i]{$��gi�����AA��AkGg�o�9U��]��T���u���o�2Qb����<�8�� >��6����m�Ҟ�ZIT�.��[���xyj$rm��/�b�`MH���P���|:KQ�X�᎐����lZ<m5ư[�,T_oQ�\ `�g���@d*.b��rQ`������:r���!���	5k=6�
i����cb����ܑ�}��0�WY���5a�EX���2�29�i_�`{�t���w �݅�_�;�u�ʝ�x!�T���w�Y��~~����u�=r\uʮ�q?�|Y�*�:�E��bk�>��u����L��n��+���sע��ǌ�'�h�"��q���U����`b�!��?t��<t��=�����{��HLC���Rn�-��m},�,��������C�	�"���aD�B�����8��0z
���J�ި��,�4rZi��YV{�`�.�����Π�� |0�䩋�x����jX6�M�_D��X>h�E%���h� QJ?=��_������M=V� �˧g���Ix���[m�E%
��.��!w�l���JS�<�)f|�|�^߬��nF�O)-�P���B��L;�8��d��x��O8j�ƳI,NH}%�����G��ق��pq������[_���`����K3W�3*n-���+w��)Ǒ	$e�7�EV`;��sK�I(?�`tt�:�ne+)������1��e`r���+w�w�Gt��U0�!�$INT� b��H�w]�"vP�9_���5*���}�E��
W��ˀ����Vi�� L?���ϒu?	��}���V���sݎ��u�%���d_�����y�eu�O4�L�g�5���I:d�T�橞�(`�G�T��������1��{��V�|�O�"�oU�������ˁ_��B�ҿxSg�������/��K�`�b��*��G��vf)�L�أl1�G;9�Z"8���""��K�J�I�a����E;�����X���-L:�|�`� �>���	~�����Bf4��-�غ1�[d�΃D��������K��e�� �a��SX�ֆ��n�r嚤x�a`Ϊ���JI|�F3����y��� ��KNNT
�]_s|��ا69����R=�9ѵ�Q�,8�3U\U�9��5��j̕C�^_��m3�m��R��~V�f�c�3o���\X����/�P6����0��4ਦ_~�JB�wz�1g�����ZS	^d~ݎ�'s#�J.2w�U�wλ���W��n��>
l���^��!p7�:V����R���x�'+�/お�y��0SU�r�ͼK��٬EQ�khgD%�=��86�Pʑ���u��7�d�M�#J�į������H[�I���鎙�����a�W�q|�k���=3�[�4x��� 
��{_2�3�oe�{��R:�e�s m�W��xt�7a��P�?@���YpJ�Jf4�Iً,��=�M~�/�#@I3^W�|����5/}qW�;;���C���]�6���+'�8YM]�!/��lx���C�q�RA�фA�o�x�P.|~�hj��\a� [|�A�7��'I!%j޿��B�V<���e9j�x�������a�����6qH��Ct����*X��*�q��E��Rl���p77w�˩}���<^�: �@��p�G� �'y�le��dmt6�����#6#��^2��h�_�ۄ�X󍦭@�`��ѣ�1�_4�t 4���e~�%�>�� �W����i�{��Zl��B�͆f���txĬs���ݡ4��v2|����A����`o'��w4pt0�.��~�K�b��J�9�8~������7
��i�d#�1�#��B��)�g��0�ø`X����aQ����g	Ӆ��C�ܶ��aKP0�Y�����;�t�*7�D��>즘��b$_�ש��&/�~_0ژb�VSc)ǟd��%����6\<�(���M�MW��0�Qg�m׭$���|c��FWD���ׅwR#�^>���a}�1�����hĂ��F5?��? I�!6��(0!��iz��nb�2]!�����:ڰ|o4Flt�f��5C��x���A�Ci���HQ`���NZ�o|w/�p�ɯ����|`���ݟn��;e:�e�1e���q	�ԍ)u+	�+)6E{�� K����WO	���s򡭿��xo�|������+9���� ����*>˛����Ĕ	��ԭ>��6|H�<^����y�q܄������]lw�5�u7A��'�K**/�����)LT��2����g�L��^�>�\4��F�%�n�h#�V�W��{I�L�W�!��τu��R�,��GLs���� zţ�.eտF>��7�X��D5i��ܺ�f0�3<���T�g=�b�v��&�4y�Z­bӃ<���YG]K|s�Ww1�9�%�����|��R��U�1+z��^��=;x��o��eE=_!5��Ϥ��^�rKWB18������u�c%�%�-iI4�I�A�ԩe�+�@F����ئR��&�(A</N���ϡ����n -x9Z�Y����Q���Ǌ�l���z��O��q���dϝ*�S?Ck���XR߻꒬v�J��{%.��h�W��8�X��D;�ĝ|�c�z�qa��E��m�������U�ț_:#ʰ0�_J�����K��^�l���И	���VI�M�>�@���1Zo��XM�y'ܰ�0ˁ��߮�څ�,5�<)I�͹_q*#���;���r���L�܃�kє�s�r��!�GH0n�޸�jRw��V�;��rfz;��Ör�����l����)���"���J�zH8���]?e VMK��!:.U�"��e�2�J��^~�I���P��˧�V2���r:��7_����6;����X^$8�rގX�*��VPL�w�t��e:�ep�3֗?eL�Q�k�Fۓ�v6�PB`=�5��������ө��*�5y��&�Ȕ����uT��3����.ǹef��]b[{7ӝ�-a5#~��	�=ԺՊ��m ��:|sϿ�m���W��m��4G+-ᠡZ���f�iY�i�t�?��}�'���*�C�2�7�'��ɮy���G��O��u��;9������:B�v�! ��:����	�R
b�) 7���������?ۺ?/X\W����D��~�B�5��v�QJ.�;{$'(�IL���xh�A.��Bz%q~���}�>�b]a��6�&ȣ@������R�����2Zd�l����*�k;��ߘ�l�P��������Ro��@DHs��'{�Tt�'9Y8��Ov�6|�������
L$�6���Gb?x嬣o��ƃo�������b1� F!Q�Z�׎�"~�\N���ͯ^oa�+޽�����d�/8�����}�j:p~��
S��&ƅ��8t=� {���E
���F�0\�禮F��T�1�P��K�9.Cո(0������_<�?�3�q2���0��Ƀ�X\k"��/�Q�Şi���D!!�I`��e7?�����_������Vut���wG�Еl�(]({��aᅚt��&wԳ�/�D؇������!^�!̿�'/E�QbD�"3�(�aN���'~��i������i��:������1���	`}p
��%�[pu`�|��"a[η�p^$�:��:N�ې@��i��}�e]�q�;�����[��$⳱�t!O�_[2��?1���
UF�yl�����|������){�rd��V#Ms`��^I��?�\�	l�Tr�<Ii���v8��q*�]!j�7]�h��v�z8*���Xm����(���N���p�y���H�����S-ӏ��0a93��4�ށJ��>W��v7*,�)�;�8E�2pP�E���G��څti�J�B�"�MӍ�m�6�[�@�M5��e�\:}��0���19*��gj:�'�	N�0���ShT��t����2�+L���y����܇&02)H��^�:�'5��}�9X�2eT��/@'P���%eZ�+jr{�g%�8�?��k@���(V��W���Kw	+��oWv����i��Ā��1z�U�������?<?����O���v��)3�m� [��ƾ��>%�߁�%6��#�S�}S�J��*�G�5I�u�OV��׫~$�{\�g�rU*g�j���.}���z�yOZw_^�c�yg�F}�w:~�CH�KV�j�oJ���n`�'��	`J]__�NX��k0�/��������u����vk��Gά=v�G��
��ߌ��7kl�AF�|��_ݰ�FvVIQF�s���7¶[��B@�� �>/�,�KxDʟ� `�kb�yQĤ:�@�G�P�\����������T���^$T)��bك@���^WWC�!yDA���˲@���
�v'l�h\���M3�L����ݠ���LÖh�5�֛�(ًKE��\Mޓ3�`/������^�>!4��	៟�G>�k~n�;���͌Bh2II8�`t!z}�\
�\�,�{�4���W/<�	9�S;y���=���A�D�!�{��ƃ~z��"��!��8�lĦ6	@gd�; �tY1i�b���m�ĭ�P�&/1��7�Zz�ސ�O�vQE�˫�)4��-ͪ��q������d�\��œCj 5V6O�����R�1���&!QQ��Ji�b=J��"�p��8A�i�Mn'|���}z�}������Z���?·>!��/7+U�ȫ�_[�M6Х���A�����G�ŹF ��!F��*fV�\�ו���O*�|	�G����Z�|<��]�ҁ���Z�g����0�Ħ�Z�gU�?�-�K��5K�ACIV� dp�F�=t�F����Ȁ쥜��}A��`�g�Z�6f֮<�ƔnQ{dT��V�{
��i$M �УZb�`��ץ�����ӱ�.�.��@]��R�|�vt9�u(�������3o3>ZPDN��9�n��ѡ  -�f�E���}��L;�lH��6�3ʿ�?ڮ�u�̢�9�U(<r���ɤ��#��k�,\'s/Sn����$�V�i6QPr#�K�6	Xu;/kO�rs&�0�]�b�,Q��ޟ�p^���rX�~���a�"�Q?*�[�˔�� <�ka���L��j�v�_N~ 9w��JlW�Ė�+��*�v�'�h�����3&��q�"p^Uo�F�������e�j3E����d���ze@D�;;���!�}����$W0�|�Q�2&H�Rdvm��!���n~������q�Z��y����yЬ��{�K.�t҃Z�|f�)jJQ�����a���"�+s��Y*Z�!�󄑰�zG�B��B��6��JN���S�\�����0M^E;ݩ4������q�r�w1_0	�@q��7��<a�8�I�)�gz0#���W!J[�����7���Ċ\�􀲕(���}�I1a&������	���q�[�F�~�Jn�V�fU?=-SB�v^ة�����C�6�vw�wC��Y�.L��FN4K�@����k�㟤%�Q�}���ƜG��%=��Q��O��pHZE�l9�<�������Õ�N=�u�Y�1�"�KB@%��[�q�^���#!�z+��2�'P�:7 o*�;�7� X����壔��9؀����ܜn�uӧ�d2��'�Y͠ ��f���!M�?Ԋ^oFT��d��-��Òm�;�񑦊�`���P
�{n�˂^Z�ٝP-�_t�RcG*7��B!6�j�[��!�HӤ��,n�L�+^fG���>r��Ϧ Ч&e���V�����>�j���+�C}y	����7v�~��[Cq�Hs�6���bk���S>�w+�L��7w��9��U��A\��{AH(��&��8�Oi�3-X��5����{�Tri�j<���S�ƣ��%������$���[�髿��y|����M��s�q��e��_(�F'E8�J+�%�mIY���W�ܕ���]�"������`�
�Hğp=�Ds|l��'43䦊�t�ݏ�����ЧQ��Y
��1#�\������o*�����`ߌ+ƭ�7�u7�0��D`�sK���uZI�T��o��3������P_�.}d��G�=a*��M|�Sf�Ք1�>�K{߂m]�مFW	�Z�@LJ��ɠrFE!��O	@��;B�M��r����&���_��2-d���c�������?���qg��L��zd�.T���/f���-E�؆?�hCN�I~:���y'BJ�������K��j�ki�1ज़X��t�� `J�r�(R�joo�6���h��˓v���@� u����/��?W�*�\ ��d$:���X�������}����ٟiA#qfO���t*�����TDX4a�OoѠ}�w`O�T����]�᠓��]�_�hbB ���y�z&ʔM҉�Bۡ{�<d��+nż���8(�P�_��a�-�0�d=�7&�Ӛ8\�$����O�Q���v���)��"e0��(�;��5"��?���h�BK�I��)�0�r#J����Ccm�΋pe6a�K�Zsd���Ѓ�`�~����ҁ�����֥ \ �ŵ��]���2*tLFy�ˎh�����_b��Ao���n�v'�C�R?�OV�X�{N���(�8ΫgT���ap�QS\>�x��Kv���1OG	�ξ�ѮA��>n��6$��t3b3������,���%_��i˩�`�vQf�V6p�W�\إ��9�h����ݫ7��)(*Wt��s: �[�b.!��ܬ��&&(��(S�A�v�"&��ލ�)d�9Sn�):@����X�mG=b�'" ��pr
���k<?&�B����V+�
#u���mxgn����uK�VںS��	5�Pr�O�;���^hj���K�Ю����}���`�3O���m'7�@�a����ں�ƀ�O�3ˮ�޷�}��kK�ϳ���j�[v�,�᭰q�B��68�Ȣ�0��#{a��0ㇱRN��5�.Y�Imq�$i���P�`X����k�v���i�� ��A���*)Wu�]��b��-�Ǆ�I�w��P�J"��8=��� �f4��$�'�q�?�4شۗ�Կ��b���z�m
��o� 1�;��U�e��`�\eK���}@W��a&D&���v�~�ҩ���/%���t!7G�d31���������>H��<��:@7>ED��V0-�>>��Z��&����/��#��������?H<��K9��r)��us���ySrI���*�}����f霵�9e��S�,�����'��.���|�.��}U��`�T*������ ��^p|iF|_�?]�mM�S]���0>Uy��(\��D���ʁ_��v�ܶޒ\� ���n��.��5�J�՚��wA�n�S1�U=Ty˵jjj�ݞ��{�K#���x�7pb�\lUY���䤒��5��f֪��\��v��+Xl�x�wt0%A�8�yv(	nyΓ��lVx8���ZV�Սp�	V^�i�܉���
��q0.�ޙ��}�Ke�>d����u�`z(���>л��w�^�|��6�8WRhS��D�H5'�tөi���+&F����v�l6@�v�o�;|']�\�#�n�`���(K0����)O�Y��|w��Z9�h��#[°=�K
����h�|<!�c�
�]�}��Zԩ��	�)�Y���p�jm����y�n���UEF{�Z[��6�T�E�3�y��~�������H��� �n�-I���W G6=�c&�Uio�U[�q����>`5tܚR-e�͗w[������bX��R�eM��iB)Ӌ����$�1��Ck�Z8���-�g�D��PE&�W8I�/F�L��dWV�q%ьۺ�:k;��������$_�����������PMu��I����
�4a���BI�Ⱥ��ui%�m����$bu]��W�"�|�}���G�
�;p�l`W�7R)	r.�Z���PkO�R�������=�w
��iޝI�&����	_��oH��	|�\⍝���Q`x ���J�s����s���V��7��?�9�\c\���X����xc�����L�:��l��iԝV�9��uW��YK0�03R���Q�j��e��7q�R���-���1��r+�>���*�X,�#͆���9���,""U�֙�e}l�|R�Ly4�ZƖ�n�B�����/�2��d7QҥQB�F~�I���LP�H��Z�r~�2\\F���k��Y�CW|.��8���Z����|֡/���O��ߜ0����K�C��h<I�wq�U+Ï�KX��0��Vw{���CBtAxy�q�6n}�q�죬��"��X��a;�4�֭�3p�Y� ͪ���W����P�빹�e��$�.D���j����,Ք>�eQXxhlc��L��F3��Y�%��{��G�=�����\����2��s��l��NB�$K��cA����V�`�Ѧ;��l_���1x�IY��@�o��?��������I%�wa���MHE[;ˍ��FL!�^{N���QE��a>�*g�ԓ5�pNP��D����#´O�J@�A�Z�wZ~�ķd* �,�	AhE%�/�r5��*�vs�E�]���K	��<t$(�1Sƶ�?2O6g�
��Q��$@DЉ�gj���*˴�"TM�O@
�"-�.���$!y�5~ܤ��æg��v���PPw
�xq�Ѧ�[�I�zaT��.*S3�Gz	Sn[��!٠[��>ۥ������):�\��y$y�D�OW���)��2&,x�����h�,���%���e�E�o��ܶPzrF�y�Zq�f<[�W�|��7~��^2~�R�jD��΍׍ƕ�(�����x�9�~4!�I��@9��Ǘ;��v��|(���Q��0�_��x�oz����(C%��k�,���ɫ>��Zh�����ټ��.tQ~N籵��Dԍwl�a�z�R�ޚ>��4�St܊{v��2N�f��*�r!�OY����s
m^7lx�]���;y���5]�xG}��3;�4�C�(���������s��{�*!��~{�yF�H,��%خA�:���ٺ�kXU h/V�����G���6%)8�mz���;����dmmA��b9=9t�<+��h��e'��\�B�原O�S���	q+3 m���Y�t�<�������1l:P�C��{7�󼁣�g�� ���N�<��_#�����p�����n���w�]hc��&�Go����(l��'���J���s�����)R]J��J�8&:�.��r���W�G\�5)\�6��|r�(Ԇݟ�H� ��&�VLS�xѼ�d���g,*���l��`Y�@vUC$���ϴ�9�=9����(���B
�@�.�R�aM�䦮��g���Ϸ�H�������L��޿H�(��moo�ni߈=6Ny;;7m[5�W��.p���	"����}��pAiW+E!�q~�Ż���]]h�X��p��;�VS�&��ڳ�:@�[�k'���xDwg9����,t�x1U�$��g8S>� ���Qu�2Z��{r�E�t�=�=󩈮
�ͯ>�q,F�P��G�*,��[;FL�_!�����d��UBk�2�I|��p�$[_>�zk^Fq8�`� C�����N$B�6�S�P��S�p��Ç�=D���&2��r�u*{���LY�=K���%kP����ϙ*$*2.DJ:����\�Z�L��j/*i��H����]�=�~Bf���&��l�H�r^��K���Y��M�i~�q��X0����x�-A�>6w��T���,���o�=�X�� �B�l|����?l�" D��	һ� ��ȋ� wG<�`{4Ob-�﮽fF
-��d�4Q�3� (r/��؜�]S⟱ه���RUx�=Ҳ���v�o�������UP��9�PFsWƶ�����!�-�Nqɸ{��B�g��ɐ����gj�Ċ���0U	%B"jJ���t�]���\�BT�rU���|5���݀E
��i%L��6��>i���e�Tk�$��3�" �q*ˍ?t|?~���3�&A. � ��8󸳃����90H�I�*�j�/�& &͡��a�9��յ6�4�����D����oº���pV.?q.�U�8p&�]�b ®��9�-:[� w]b�)���%�B���v��EM�M�IZ ��G�K���:xx,=0�,�"�.n�c%X8�D:3>���ٱ�t>;�B>13��������29wB��ۺ9?&G�	��_��]�ȚTf\&��H���K=�sxy�Sx�4�4�1䢲:E�J�:��	�Z�l?Ao9ک���Xƞ	_�D�ö���0R�*�f ���������|U�r�X������a?��4�Rr����2�-��l���v��.��lz�p�A�s��x�������y�g*
�.q,U�b1���]�XA5V
{_����'N	�]���pz>�����x��$�P��&:�.܎=s����B:\@b�hp�0�:ݓm�W�j0�5�U����<ʒ���-9����n1"J/��Jvk��Lѵ���������kh�f�����le.�+]jF�t��U�uJ��?�~r#m�HL����ZT��m�oa��ƙE�R��yȳC�fx$�m��=�3��"��/�Cn�w"E�}r���g�=4�s���'[���w^��KD+�}�?Ԁ�0<YڦP�v���~孜R��F�2�y�{���d�Hϲ���b\AEU�����*�"��F�����j�7e��C����cn!;A�k�[U[��Nj��[j^*�\�l�e`;B���m��ꆜ��=DF�Ӯ.9���ÆtB�20�E0�:����Lg/��DҎR�� #E��z@�E���-bO�}�D�smj�HY6*v,�If��u�m̂R��O:Y�B}��	9�y���m/���9��6��/�2W����̳΂3V��{�Mb�JʯNL"D	�#r�'���]��Ä���K+�����6��ʔ�n	�4A������5v��G���V [�r����i8�mA��KS�#�E���::�X�p��M���t�f��BFC*0bl*�;�.��H�҃.�ξ�U�!��P9A���B�s��I�Bo*r�l	�~:��>����+q���L�Q����H�ӳ5�ʦ�#��T;�!�4� q��r�O�u�t�A��_�Ѝ�y���J@��0~�ZN���)G�q��9	��������qwu�G)�<��H��+\� >l��`( �I
cW�40p��ԃ��$��.I$I`�`��gC������ృ,�*&*��}�%�᪊Iv�+��l���}wd�B���Y��c�\�p��r@��r��T�����贍}I���ǿ���߭�9��V:�%Z�J���}R�1��0�1qQ�r�k��+~�"F���Cde��`�K;�.�n�2���B	g.Q�X��RQ��f���N��[T�*�E)��n�o��⡨} M
��~��e�B�7?�N�V\�i*})~�T�T��r���cMN�q�g�SF�q�h��MƳ���_�N�<��Gp�(�ԅ�
N���Aw�%l�1�7��Խ�������%�z�a� QQ��;�	�*|�k�,9��1����Z�����i�2nb1m��v�v��U�HH�����������<�T���>K(˫A�1F��T��5vNm���	������ip�
N *��0�h�H��v����������/���:~�qI9���v��S��ۀ ��Kd� �X9�-���}�]T��r#��4�I�.IG=�-�!�u���6�|��N[^�n,��>M��y�����Dq3�n��+�DZ����:"��� 9
���T�ȸYaÿw�$�A�$�����d/HNk��p!�� !�wO*�*ؠ����^�WRV$�su(BI|P�Y��:�R�[K����}�.˃�	��dF��W �������+ }��~QT�5��e��SB6#�����Y��uݷᘄ��@���Ӳ�4D8m%��U�os�tҪI3K�J<Zn��CS�/`���ߏ�8�^���ل�=C��`����靹�q-�U�
r��������������J�>iǷ'�5�-��oe;s�$�d�Zk�7H$?!��񒚮`d�T�A&��1�f>Ua�����f9��*�M�,쉻́K�d@O5��pm֮�U��@f�Kư�.���D�\�b<�?!iu�b5ct�>�$h%܉�W�٥?����i:�+꫻��Se�8�vʑ���B��1�=��S�¸mu����o`w�����V'R�9�n�3��]���L��=X��UU�����q�
L~��8�Z0ݼ-�)��Byڔ�{x�~jI<�(������=�q��)|��WG� �����~�|�',�4�7̶��4e�+v	r�Iq������N}��KHT�P��9 ґ?o��x{_������>��48zy	��� �(h��w��v[)*8&8�����V���!~L{�>R$��fs�+Dv͚�_f#�?�3I���B]ڇjZ�N����w�0'�G�~���E�u^�Z�ߍ�����Xy� %�jZd�+�WZO�� &�>��[��X�Sb�8`P���Y��`��O< G�0�)����|�LS�)O\*Pc���A��c��x��pz��|���BZ�_3uP�6��e��줤$��	�� (�7�d�9�p��Eш��
�D�P���&hxO1�ǌ� �d�ĪH#�L\�5����J���L���F?�:fl���y�Ӷ������rb2�J�y�	�C3�{M���Z��6�z�?{C��=ss�ٳ�1̶D����̴��{5�Q���qK�"Ch���U/Ls�[���{j��E�p\*�����F@�����\y�;e�m���m�+���d��6{��Y�tM�O�rr�D3��w����æJ�\�;{���")�?�@�|,U����*3�� �dF�J�-��;j��Zt��}0�E:Hz_`w8����sW:�c��뜦�R�k��Iˣ�w���6"[��uX�0�Vo��*�&�{���Ԡ@%����M W<�J�M��퓗��\��:;�s��k7@�RG�MJ��4�!��G�f�ᅭ*_)�#�qӗ8�n��15rwK0��u�6�/^}�.��xٹ�5:dׯt���1I^`�G+o�G�5 �S6�G�)kuh�?�g)�"�*��E���C���v���jt+�X��U3yF���b��(#+�Pr�!�/_�ݾ�M�7l���d a��!j��8�LD�5��P8��7r���Mv�<�v<�a$�7��F
�M!�D�&w����Ķ���A���\��|���F8Ր�?��G���]�[��d�7�7(�N��*?e��2�g��̟�f�Ďo����Dy����	"���Yٓ�ʎ�9X7$��`+q�>�1.wI	��I��rG���ȋ��`����ʙ�l�!`ic��TT&^d����
��`}S��� V���V�W��Ɋ��s̾i� :χT��K� ��\�~��k��x�0�+>~)FPGz�6�����P�+&�ۯFN���a썂��8�ث��!����S֏x�ݱ�Ԙ�n�$���"vJ��\O��)vQjI�FF,��i5Y�s����6&b��#0&Oၔ�R�#���KQ|u����F�=f¤^���K��Q�AW�'����Ul�ASu\�g�6mv�Q8��j��eF��0�FͿf�A�9�w�|����U�T�$��{N���S�p
x����Ѫ��3'��Nt�/��%xxOF�^J����Z�>a�hP,��p"��V6z7��_���>!�� 9��q1y*6�q>0b�1E:ƚ�䣌R��,O���(n��3��Dm�mA05�WP��Dd����ҭ�M���(�fZٓt�"`�^O�CY����[6�]���
�g���vL�j^���_��x9��Օ|�Cc�l�Y��]�j�L�>?K��Q^7l�u������$U��e;ͯu=��b�Q
a,CYϼ5/����5v\ѯ�[o}���/^=�����~��h4 ��5X�-�-��
�xnuۊ�uB���	����5,��;���\ٴ���i}=' �<�ׂ-f64�ؕ�GV�ORP� � d��'�M̛��'�5�8BR��3r��	RL�:�c��l/G�te�b���F��б0�q��O�λ�s=�3
���+��с�����Nn��ڷ쩁j�o�"�O�ӻ���uӠ�^�4������!���E��v��p��QB�|w����M�<.�x�׆5����kQ �q�(?-�����}��<U��;m�������ȃZM^Aq����D�B�Ӯ�B��=��Z�Q�=#�f� ��Q�艐�d3~au^Qx�Ɯ�����dQ����Cy-�(���|%b`�xd�k�F���<�ҜS�R��fe�o��B�cp
���)�ܶi�i�CuN���e�tD�@p��M�r�6W,	]�ן3���x@�n�$�q�kX�г�q��_ �e��Iaߟ���E�Ϲ��v����b�QV������Q��)=R�vʙd�K���bݹ?.�o7&۪v����&@�;�#���ᾭ�AF�x�lS�|	�x����vM��7�~c/���Q~�-�+�\�y����,z[�Y��zW4���<�k|zkI;�qW�#�/�^"g�CUt􄕂C����/S:�mɈ�c���#A�ĻK�l��	�ۿ�6!�ƽ rW�iy���w�n�*7Ӟ�8i�ݞ�s����H]�i*��m[�B=��P�1��B��v�� ��r���},�����U�[��e�̨,}~���a���Q>�lGB�l͓����q'�T@�kVu#�I�v��{iS~�,�Y{�8���A�����*W������Լ���v��!V���rAK��|Ӣ��Vc ʜ4�k�Y��.���g������5g��̼D�Jdg�{�Z���,�� lFOFl">�<��>x�hT�ٺ[����%G�:<��$uTZ���,���u��k�<]l��q_C�֔DTdB�l/����T�-;�u7��#�Q�L|n\�m'�HiH#�-u�uJ;���*F�VMH�<y��Iǥ�����D���Lh����H������.��=g�Љ�����,.�\��T��b&��e,�ye����T _��+���*�&�N|�0��sa�z\Ȋ�ܛ��R'v����K{y�����1*�ے)iAJk��q9�G�dp����)۱�5����3�_{������5�3�]��)޲�ё����3�PwO�+���)��,©�B9���h�����L�vs�7�f�wZ�l�qT`��ܱk4/����7Y���4�@�ɰ�,�:t
�W���H]��%�	ݨx�޼��JP�-��b�\�w]^���h������?������Ρ������%F�[�>�k���,�릛�$��V̞Γ����4�FϜ�l��p׻t�H>n���J�*�C"���I�i:�V����Y�ϝ�1k��@���B'����=q�tR�v���f|�w�?џ0�K`^(�A�.����D�1E!�p�峢@�� ²�2c_'Զ����c�w|�{"IMlAp?����Ǯ�1$cx9��36ߪ��p �,�rxɖ7=��J]�L�F���u��+	���]��:�F>�`t����t�N�^����j7̤!�hI�)~K�9y:�	H(�3�s�2�d����њ"�g�=�0si^���8U�������U���L6ve�zh�mP1�H)��X5扈�{�s�'J=c���̦�[I�R�	�x;�/�|��<�T��/�{4^M�}IaۥB�eI�$J��#=/fҾ-��:/dù��=g�D�P�zuf����4����)���ش�v���z�u�RZ�t/��%,�08�zʙ�{|�c��������	�.sw@�"�-E/���0���J����V��I|�52�zN۽�p��������g�7>s�Sz诡�.�a��TMO��Q٭���e͇f��f�/��1�CP����QEiHc���u)�r��l`�*ioY�y������d���LN6�8��6[�^-̄r��ڽާ�$k���dXEJ��;E���%s�wm����҇�B�^������)5����q-�Ũ�� &Xܞ���Rv�Igթ�>�G�o�x��`�r�����,,<w�J'F"s��<�Іa����_�D��O7p�H�:��L��A�r��O���U�u.j��L@j0�h�T�V�/{��@q���*#(���f�ȼ2� >�!SG��<��hrw�����/3���e�E#�����C�VK̼TJD��	]YC��r4�n�lEO_�8��rZ3� L���2�MY�����=:%8��E֛�u~�XhmH{�H�7~_Xo�>��XK��>����(�l�12��{'w���������K���p(�_�I\����04��60h�26SzOx�f�����54g:�Ö��d�<�'�H��0`2��/�RtKIM\���Z5F,��s�#�{sf��9��l?�ݏ���`Iv9Ջ�}���cg�W���S�j�#U�TV��k0�1��F��.��@�GN@@z��P�}����'E<����`���tE��H����GĂ��i����={�>���j`$f~� Ejި���l��3S�Z�`��EK13f���/��Z��P����$^������~������f#?b 0[�'O��y\�,g��:B�ޚ�pd�GS��s�v�� ؕg��|@�e�U`�-G[���qem�$Ö�z���zK�B�uC!z�f�h46���W�>��Fl������G�E,-�������@@�EVf�ߎ�'�;Cn�a,Ԧ�p�G(�c*��EE̓*w
Vu�\�͎[�kK}�2l����V|�xf�9�F#�尿.�LS�����w"נ�c��e��|&PH.G)��_�����$����}�Cy���<��)y��&�zw��	<Y��S}9�]?��:�9IL��/j��h�%����a �W"�p�PKH���{鏊|TY��&1`�d���g����'���I<�u�ei7. x�Al=gA�}󢏴�6�D{7;h�7,q~��K��{�F�#(Ҫ\����X�|r�~������A�H�h�������~/͈]���`�� �{v��U�` `(�v�
�z �S����Z]�MB�30"%v�>L)�)����C|�V?7����F!u ��as�lF��2m��_�gwF��I��A��"̤�@�۟f�?�L�?�*-(��@/���� ɟ����� ��G�y ���Yc��4d�xh=�UN=4�_`�1#�����ҵ)Ui�
1hx�H�3�H��_@�V/i�J�����0�^꾋1���S�o���x��᳇y�T)	�m�,=�/�)@��[�P��;�C5H`]�����)k�54?��"~��_0Q���!t���K�+%Rh���U0bC7����O�*�}�Y�
?���pn��@3^�������u��2؞���T�������a6!�nA��2�?7M)h��S���󉛷$�2�/���
߿L�i��g��[�b�g�X=�ܯ6ǿXr/Eu`���)�&	]KH�dZ��p�\�g@�E���^�p5`�D����?�=�`�Q1P�(@&��I�5��d�@#�p������G1,��Wv��w���!��M�5Dtt���a)ÿ�ׯc�nj����%�^(g�#ݝٰ�"A��誹j1#���;�z�%�J�bA���$?���T�X]�j6b�($��?|]�a��Ï���`�3�3a�b~1�� ��<�oJ`e��Œ^�fƜ���9`íL���@�նoX��/ȧv�I`�V�qr'7���upȲٚG�c鎯n��Ti��tʱ�k��).�
E,��kH����9���i�����>@OIE�2 �mu$KS	�|�&��n�'���I ���Ձ6�b@���jA���g�@��O<�xv�RD��;҉8q��V?pg+��&n+G�-��'����wx0]��s1�f[�S��I`���^1��A��ɉ�C6��gx��aش~�S�o&�i�1٢� �Ow"�/a���N
ˀH���7vU5���D����~,7P����b;�|o��˔a�6o#~j�rE�;$n��H�>�;~�'�Oڪ)�����A	�,�}��d�J��tV���#E_F�c�}��@xmL y�UA� �$8+�zzT}"�+tk���%��CX�#��a�f�n�~}C.!��|�c��#F�����Ԭq����So	���pX�(<�0�PMAh���-�\�lVv*��4ġ������Nd�)f[�h3/g�/4�����_���L@�0M�
=.�J�������F%;Pƽq�u���sÐ��+_���OlHdr��q��&ji�yg{������Eq����+1�q�\�H��r�i�1b�`õ��=��`�mnf0���ۈ~n�m���V������tn�{b��gWS�M�3t失��X�&M�&b��ĩ�ұiVոĒ����LI%�̹oa0��H��:�!!�<���Y�	.��م �Y	BV;�̈��JB�A�s��y0[݊��x|�
{�e�)eXeg�J���y�{qɱ���T!�
&Nze��<e�ӱH�(�X+�UH��^__��z�y^�)�	k�J�Pk ��5�2tI���<��&x@P�\mSD\OB��16�<�Il��p9o���D�NN&��s3�2y�7��)M�2Է7���D�Ƃ�!�2r����ÖU��#7>��9j�;`@�b�T��f+��_af��?��n�x���Q�"��C�.��|��D���u��sPB��G�j��l�`��b�g2���&�rnK��8���[��՚�+2�����q������*N>mO���Ζ��ֿ/�/�j�F��@�L�I?m~s4���p�Kn���i{] ��\L~�N�R�N%U� �V�,H���O�;J�_x(w-�_�u�#~
sAI�OE���b]��ٝM[�E�æA�Es�܎�	�
��M��
�lMf
(O,��_Ik���}A���\_�c�LX������S�����c	�֒~����5-��j��������-?M{��zQI�̏���nv�u��l>�\�4iV<*~��ڸ�7��'}��⟊����I:6h�(�� ���x��A@�S���|�
#K'�]c���փE���ttcTO�Kn������"g���:����j̭[�l�a��%G�ˁ��z8�v}�%3��\���Z}�X-�Ѧ��,Y)#?.E�-��P�&��Г�!XB�>]��̈́��$����-�5�j����b���0�q��l�63E�9�kO�R�&w������vm�	��?��t�/��
C9�E/���n.�[�{K�M�V�h@�+!ٿ��E��*��̥:"xѺ�[E(t��)0AJU0bUP�Ÿ��<&ôc QC�S �tPR��
�7�T�Q(�n�	�ߙ�tW��!3�`��lG(������$͚��M���۸��V�)�UaV'�
�K	���,5B��u �9g1���q�+$.z8�`�t;��#��k���#��~��l.���-Pg�4LG<̼o��;6��!0Rg�j���?��o�i]j|/Og��������s������">�Y���*�,]��g��o��7�%��V�K��=�22������3N��s�X>�H��F�8�G�-���w;�����&}������v��]�C��gû>&>u3�F�9�⛧s4�R��`!��9Y�i��a�i?d��?쎼�RZ��!��J{Hk��q]z�8 ۏ%:��T,���C�����D���+g��&��]M���k����y�C�3ʬ��%�e���u����y[!��w���x�e���	�N�!���	�R�7����r����+sF�l�$x��C��vH�v/�'%�}{���(ua&�]���gMݬ)��kW��o��?���Y����Û�)vob��H��J���R�z�G:�V8�U�������<���M�M���F����y���ڌ>i�e��>�;�A+=3��x�0+� k��m��e�'~jĻ���_�'q�d%T�YK-�<q���(���l��v�^�W�=��5��F�	_��?�a���]!�FH\�4.����X��TG�(�޳o�,�ۗs��o��q�0� �~gr��]���-�9�s�В@���}Fe�[����u�����~���ub��������;�yV�ڇ��O�?S�Z]GLr��L;-!��xo[�XQu��%�=/%��I��W��L��� jN��4Y��;�kaM��2�Ga�:��į�Uw7�v��RY��ul���׺�He8�B����!���G�]�Y��ϧ�m�I�
��ѽ͎�<���;�ơU�$[���I[l>��)y��������:�FaN���|>|*U��q<r������b,���Lק�0A�[���;5��ّ\����w���Qe͏��L�� #U�߂�ƻ<����P�����`C�T׭����it[5��#��;O���NAoܗ�;��+BA����L\��uq]<zi5R�ceS�w �V�Z��@=�f0H�p�ս=��:��ۿ�so%�0G=��J�
x��{{Fuݳ�� V�4E,��wx'�Z"́����u&�ʼ;j�N	3��<벾�g!��8��V�F ��Y�3�j��Z>M?O��bSIVkS� b���B�߳���;���=��ܲ�4=�rmŢ�fJp�)?[��cUf��}��2W%���)���T�߁�g�#L����4j�Bsc�!B�4���b�ߠˁ��x2�,��P�a��b��^����G�M����;0�E¹�]����U<��J�����Km���m��H������2���#r�=t-W��аJ��S��eq�O�|�]�0I��͆�G�&�ŃV�YM�n>�5��_X��?I�)�	E��{�H8�Y��$�Gz�˳�%�ZeD�f/�`vk
�!]�j@ �`�R[�´F����ޣk;�q���`y"�ĭ$����Aݣ�ֲ�����c$�=�]��~���۵�׷N��.VI�9�� ����Q�ʫ���r��7��Zp�����D��!�'Q4D�ՐV{T��y�}1�=6�8]��r $�N2i�{@
�;�\���\羡�K����:���K�Ҵ8Ą�i�B��\:N~�������x�#л�N��h����t��L�tI(pc(�� DQ_/���.�R�L�[W]W�$04��ٔ��h�o|� �2-fTV��p��Y��ג�X�:A�V.s�Tg�-g�mu�6�� V�hfc�r=c��9�Fu���9��<����Z̆>���؀z�P��~���l1�JW�&���NH����q�5�dC(���L���R"w�d�g��Sn6?a,F2p�e�Ï�j���
�11cj���3tgme�w�V�I2笒��R��V�p�x�[���@��K	P�[�LPm;}regi�5�]}t{?����38�8�k��A���t�Y���1���?�8�q��2�X�Y-D���ŕ�1����p%�[9�Z�s���s��\4G\���Oe���sP�J��x�qpA��=����h�Ocsi���=��ż4Hy�׷�,0�M����C{5���ᘖSX`��/��3hU�г�:ˏ�n$��`�D� Y\a�^F�����qXz�mhv�new��$ _��R�%�*S�@�����܊��V'�f5�P��j��b�/�Mu�2{+b;��5WJVĽ�ׅZ(z (ʑ�|Q�	#v� s�1lJ@�uˢ�(	%���D��s9gݭ		P%W�Q�&q�<���f/�u�au���`v�����_��xAe�=:��5 ��2��V�L��k��.�D�h�� �z���O�P��Vu~��q�"�i�{�����y�lJ���wV�N��(>B�i��ʸ��b���	K�"��{���N`�H`�Ԓ�0�12lY��=p5W�"���� ��U*qGQ-�8�PD�ً��ֳx����@�
�32v�|4Vv��g�6y|I�2���F1��+��U�i������j,!zЭ�P*\umZ���]�F������0a��s������}���ց+ ����c�L�H���*��
�1�}�}�"���-+�T�Im�4]��g�^͹��4��5K"'�=��r|���W"`�_w�y*�u�����6w@�*�w ��~����?U�Z��Zv��%;���o._ҹ��&�@�{)[���F���$,�m<w���
��?ݡI&��=����� ��R-tRj��
�"J�ȿz(�j�%�r.�~��"xu(�A��`�1�rr�٥��!�j�K��y��X�F�����|ӊ�j��1�0E������mD:��q����uQT��w��>�ֻX�r>pU`�ݼ����u��<o����lg���3�Ǿ���F���T�ٚ��QԉS�E-�� Q����0�����H���g�Jb�k$=S�zR���#r4SJ��5�w곧�Lq3����+	�T{�N��Q«�Ae�1<�.��]8ˀ�\��ݏ���;�a$@M=�s��~��>��(��Cޅ؝W,�� 2Η�Q�ͭ�U��؛a�o���R"�w�4�؇�`��U�iRSy��>��BH?+�e�	�Ӽ����r=��������z{a��SF�onk�",>"⷏��W�(i���)�K�f��Ͻ��>iꙃ���m��b����O���bx�]�mB��;�4uN_�,�vT�!9ٙ���Tb~e;H����-}GJ�Q�N���Y ����C��#=���!E��4r!�p�Q���G���e3w}��2��'g�m݅j1{DaW�H=�q�qC��R�嶓xk��%�OR��x+���P��g�G�2C���|-P%�#��w�����#�D�݆U��'���A��LS0�)�JXd�_M����M���uH�n��7��-�R�q��ܽ�I�ʺ��O��x���
u�odMo��(=�/F�*?��;�^�x��8��S�1�;J�o�qȖ�$�cz�e����e��~n�x�[$խ~Ҷ8F�?���0��]JZ�q<�:��1�ж�h��=��!C�n!ݰ��K���^c����D���A�1��ԙ Ӵ�lm�L�WE(���%�SSW8���S(M���%$6h�ڜNCQTezSZ�I���B�b��y�z,tr` �*$�`zI��z\���/4�P^O���(�.DM)��-(lڏn�i� ��j�j��pm�B\�4KPe��n"*�X�6g��H�_�7AO�1	�a���8:S��^ef^_���YL;��>����HLW)xW�q�C�����hd��(��L͂�"I��X�T �y�o�=]����p2p��=�$ͥf��*�t��`E�<'��^_? 2v ���{�W�g�y�/F�<��#�)b��F�Y2C�`P���u8��t��$��|�7JT�P��u���)��{MI��]�(�߉E��5���ifߴ�;�S��L��0��3δl)�t��QKP1�(0'*�o��>��A�&��-�Ց�#07IwQ����#2�,�E�u�(��r�d���������O�8��:�x�`,)K�<B�~�8��U� ��+�g��w�i����!!V�ɑ�)�� �oZ�����u^�#���k��9��j�o�f
���k���څM����˶�z3�jOF?���`�a�iT�C�Ԧ�+
ub�2oϺ����A�Вb�5\b^oٖ0���
��JJ�X�5�2f�&�GOk�'�k}s�[���'X�b���A��5wg�y2_p�ػe�]1�܉� ���w.�Cm�����>ERQ�0_9�*����)7���������i�^��΂���̎�,S�sk�M(�2��\-�7d����I`��gK��ԑ��=�
D����:|�8/��;��;��J-Xd$��{)(�H��W6je{\o:a]�V�V3k)�o!X�A��9{ Hm��+l����-��F4\��)�Vb�;σ�A�NT�Wg���1
lP%���j ���.)l��D�F��8�X.-�����G�/jO/�x��.\�\=�rMȓ�|����f�����=}c}*�P���\$�e��'᥎v�/������-!��(Xa馝�4�C6a��_(�L(��{i��AKW&=��k`�m�mk�u?�؃�"�B N(�r��t����{ۋ��h�]���c�9�
�*�N�m=� H��R�V�DX�
-����]T���%asa�T��*�����h�ce�+�r7�K�&$ ������l:���3�0Mh�q�-��oM�m�ʽ�&�/E�����V��G���[ݕ �a��Z[���,i#�q\�F$IXS_��{�\u5�c�iu��l���f��)��?W?���*ha��o2�������L�����e#����4�S�g��OY;`�y�W�d'hp�|$����*��7�,�C�0V��{����1$�7`�|�����!��B� k��f��KYW���_�ق�Y�L@U�
�&V��gj����m�"���8fY}&[>-Z�$��8͌��V)%�s�V�5��=�w��[�`K׮η~����nGVFU�B$�֎&f
��V$���ɑ,F�+g� ���F�`]�_���?�]��K��YhW��a9�߱�����hL��WAT1{��ra�<�@��m���L����?�,ཌྷ����b��P����C�B����?�eg�K����9�V6�6,��%�Ȥ��_�c��5�,�'��a�3U"J���/k�&��ќ�A�	�J2�l���O"i,'�ͼ`|ѫ�ӛre�lȶ'#o��>"Z\gҡ§���r��I �s��2���f[{���)������z���GT3����_�ͪo>l�����J�;%��P��$laV�5�h�������\!�7�^9�Xwď�wv����j��Ye�������Y�̈)00^�ӻYaLY��Q˕Cv�ൕW< vO��rȵ`���Y�-*���MeBd<�ތ9�<�sﺁ0�]�-[m�%ҫ���Ϋ�z�ϴ�:E!�*|�Y(n^ᄜ�"6�[rna?��Z~ޤxD]�w����������S\T�#�=C�~�4�>��Y�	�zW�4��:��Ę��2�֗��9��Wf�&}pb:!{e���; �2�0Bdݏ^
'����"x����ef�L��ᙛOw��,��L[Cs������a� �h�ׄ�Xor@��R�	���٠r�].�U̼��L�)呀��c���1�G�f�_{�Xc��`�n��z��!#����*}�y $�z2�頕Ѫ=�9n~3q_���Fdr�`�����
U���Nkb��\z$p�lL��Rي��r���H�f��J�g�KS�n���3���Lː���1�ڃԠ=9��/9�X@�mh�
�8��(���ro�ۅ������*���R�H��	����h�v6�e�Wzoc'�#'J�g}&�ў
�����%c�?`��ۼd��GC��,AKz`��r�w�"�ϖ��8�d�@0��l?|e�<ޡL`�p z^�դJ�D����j_O2hH&�o��V�tS��<��� ��ط:��H^��:b8'�85�Ґ+��?��X,�����P�vA�F'0_���!50��ڥ��u�W48a���aՕr)�	�߱��=J���۳]��Es����j
����fi�7|��ÑvUC��0yGO�<i�{;�������<��|��y�n5?q蒽�!���g{-��ȭԂ��V�zZ/����&^m�)fZ�K:B�/����.��<#ɋ�i�Y�/M���`t����Iw��w�r}p'Z�JBa ��{�\��";i����a�s:ݟ����5�$�7��aje��u[�Mp��6_ׄ��D�"�<�D0�8�dY�K�(�:D3�t8h�2����}|M>��u}��g��J�Y��a�.`�lΔ*}�(Y��gw�k�����6��gI�B�y��Lv�%��s���L�p�o�dc�b|��R1������J� ��ш.^�}���p�R�t��֖��\���qb�Y%�!L�-Tb�^���~@���J�2���_��з�%Y�� �(1d%�WEIɌ��7�J_k[X��Ms:�<Ly�n-�j�2��>�����C�43әg�<��i��?���aN�2#�	EL{N���#��Y�����a!]sF���?r���r8�S�9�5H@��0zP�|e�
����*���%�n���mV~�ګY[ ;�3`�0� �89*3Q�3��x��+�*�M�K����P���jC��d���ے�-4�p�4ڄ�gx�
���'�R֯	��71B{r��H2}}|)1��j���4O?8��9�˥�̽�}?����^^S���O�{jz!ŝ�6������oMdb%Q��PF5�=n�i��7�R'�x��[��e6�꠽�2�i���l��ER�MyB29D��U7�͖
��ʋ{v�8
��з�l<�oY��8�B��|	�,�NK�&�Md�g�)����w@x���:���M�����!��è~zΖ-s"L��pZ#��~hc�Ы�5��,WL��{�ł��A?s")�-0e���� 9���/]�م<X��M�/e���9�{c��"���
��
Կ�'��q��M`[Y��q�Z	qK�~�lk�}�WC�͠��p����H�����Q�F7�H����n�p��'m���.C'���:��(��].�?�%JW}4�Ҽ{��Go�� k����-�ib9���sC����Xy�#��@/_ �lS�:�-��")i¹ۧh-�ic�!f? �U���H� �}� �a�g]���&�a$d�x��*�m17/Ѻ�#}��k����oB���`h|�S^�3ӍN5���y"񤺜�)�_A��٤ݪ����\����C��z���6ɫJ�)a&f�����b~<-;��� �M��8��Q��g�LtP�'E^�'�	�?l��+h2��O�ۥ����EMȭ��e��BY��3L�w�;�U4p
��v#f�]C��r�%���eZ0�`g�t���y=�I��cr��7���l"��4F������.���}��*�_����s��R������G�"=Q'|s���T�r�c�j��1o����,L�K�:1�;�^��C��F���2y3�Q�=i�I`K?)�^_���q�w�<���fe}\�~�)Z�2'�r�B_sy��֊b�ŋ��onH�<�%�fqpb�$c�d��|L)V�#�:w=����@�%5"3��)ùaC'�﫞���g�Wg��"%l� ���d�Z+Ӏ�QNX�?Z�TYmǟJ5��v{�$b1�m�9i��M؉COMҐ<����-�Q;w���Z.V<��(��ƉBh
i�������g���c��6j,n��lӭxm��[�f�1B�U:gf!�`��xY�]-��?e��$�QV]��oŸ���\$���}���B���V8\�N�)^���|(e>�5�B~<�k�40�uc���AOKz���d�t=*v��{DI9�|�_<&S%�8��5��=��.F�ia#s�=����?i-�T�ϵ��^�A:k��%2ea'u���W�Ӊ5��/(��L���t�1����v�b�O�z�;G�ϐ��/{��C,�ӄ�dβlW���O�W����*��ab�S#b��eas�8�d�d���	�2{�_��3	��|�1	�?)=�'�e.;��dr?��7�iJ�M��ۻ
ׄf�K�[��<5b^Θ�L�KR��ߴ9��V���vd)Q�x��9�l�y�er4�r�����"7 �g�J*��s�M`2�V��#W{����;t��'T�LM��:P�������-�]�8Մ\ʎd���R�YΎ���8�|��@�>3LDRo-�0J�eU� 3�Ym�O���x���-6+-+:RܹU�F���qœW���.��m���[�ӂ�G
#b~�UoO��n��m���o�wY�9����-M��ەI̹㮨���>�3�`9�^Ǵ��������-��߳Ժ�v�	:<��3�D��;qĚP�+ +h[��iL������2�pw��K�Ӹ��N%�(��~��Ҥ1�� %X	�zM���]�O�6�X�ꡌ�kCo@��Ek�ݻk������i�alrӔS��I�'1�S����!@�8��h&��".��W;��2��_{>��7|@$�j�sd`��j�J�
��SUBa�MwG��2���	Bx9��y�v!�K����"��~�&�z̰ǉ�.�EH��\�ǂ��Y/*X�u�Wv!�&�`PK�%�e�k���8Oў嘜v�,,;%�϶��ce>��-��$GEa:�5��� D綬��ν'T�5i��y���h��0,���	�*�]��	�G�P�v���@�`}��|�ם�FϚ1��i»]I-F���{Ewʊ�B��ݖAoh�5��..��R�a�
*Bp��M⹩���u�t�۷�*�u���]7_�P��rRc�?Z1�|M�Y��ӧ��?@�ϕ6�nQ�FYm1Ԁj>�(�Bݘ����4\��Z���/�@Q���o��!����
9&�~�y�}��o�_Q�v�7�s��hF���6ؾ�0@f[G+��nG�,(
P��@7WML��}.��/�<m�>�t([�}�t)c̒>걧ho�`��pW�v�g�)�2֧�g=��	���+Z���!"��Ev3o�IjM�C����r �̃���H�!/��(�M�X9��"(�����~s
���z9m���
6�H^~���^Q�a�sf˯���񄒛u*~����aa|����Iآz�kp?}��Q����'�2���}V��l��2�G ���f��3ڳ�6��x�����S@)X���K�U"�f��Bq3\�A��j?bç�%jU���W.�9�7ℍ���o!_�X��q��g�n��I2�$�O�]��m^��;�g:sU�͗ߚ�~�"(��:6�[Z),��(Yʹ�H��H�
�kg�`"������Fl���g����D�g�C�`�B3_D�`�z|��[f>�}��tp]Vw���0�{�n���z{ު����B�iveJگߑ<l[i�S�?4O�<�������h�`�K��n��ջ��6ô�MC��e!t�� {�#b�f��Q�E�,���C}��.d��+*�Qg�Yi!��Uo�#��&UOb9=O[o|�(�������j,��{��Vk�(��|��eF��fv^A����i����vG��~���g�v�=D����i��;`"Zn(��7����ż�.�L	יT\4�9Eke*��	��@���J�Xg�Di��Ze�������qC�_��-� �̱�(}��e��X_�꘲���F��ZusOhg�"2�C׮�}����K��c�~f��!@`/�Tj��Ȑ��m�S�1n����#�\�Br k�Ke'PS̰#W2m�'"-����/��]��x͙���8�Cl�)u*~�N�0�t���>m�� k��Xߤ_-`�rX�;`ݲL�V���"\�hD蚈۝��9IspL� ��6D����~�#�4�\�-L.��gB&��n%���u�yƆ}+ĩ��0+�أي�{<�Ъ�'�&���V~M�Śe��P�1��Mr��c���X{6�Y|�;0VR�8Y\ut
g���W:��۶wz�k$�k��$��1ݽgک��u`��+%#j�j���ҟ��դ.3z�@�bP;Qv�$x�T�F�y�֔7&�pi͝r�-�!��W,�N{Z1k}�[j����0�5O��o�T���`ü3�i�7��� ���t�S�B���[k?���}ᣬ"l��U��YXiU�-��'D�=��������L�2�L��0��st�����Ϥp���`*�=;;�%���h���,q�^	����sO0�;D�,H����ō.��v~,���Ȕ�@:�-Ũ���q���&�]��z�e��A��A����?F_,[��le#.8 �*kK�} ����[��t5*1�"��-�s[1��u�	�7KT΢��)v'{K�,����ag����ךN0oR�3�������x�L��q������PKv�b���u=/P�5�!.�|y
����(�~��\�ZST�0a\��D�1o�	G�[�_6*������f�KW^�)4�nd4C>ZJ��Z��6�^��&�~m*�Rn�c�J0l���o����ٵ��mk-&k8�����Ҏ���q��Q�]
j�6Ͻt�A�)`gu��]tZ�BS�'^��]f�:���Dk�����n��z"D�9>�6���f�Ė���Tm��}��dl�J�g�G�� �����o��O���ú����W^{ ����=��ѯy����
��"�@���	�Vk/׋N4"�u��T�x��Ö��6SF���ss��=��C�KT�'�O�v`�r��|�b?4�����-�2��zK�,�۝���CՂ��i��ŉ�z)L����eq��E�TN��_@}����7Jbnf���P+�?�<ݮ^�3���D �`�
�"��q/yS���(�:�\{�Z3JDa���c�-���m�Ĥ�s�
J�����ώk �K��QS* ��)�k���	��S�������q繅�^,I�Z���}H���J7\�؀��_�L9�r�74�ڃK�8���X�Y�{��Ȝ��%����=+�p�h��飙���"�/��3�Έ��z���Z�5�e _[�҉�gL��vfV��\B��e��]���W�:T�[t�O+tYbkV��*�k����?�;��b]ޣ���3x%����X[�T���t+eS����f(�z�pt����	v?��l��Yy��>cmd�����>���y#R�M���v��Sb>?���7�M������k,���2�0�F���ӕ#i<̩�Bߤ����T��FP�6I�TdG��2_%b�8IH-IJ+Q���7v�f�3V\J$�>8V��	t�T�D�`th��ş'�&���@���E�������2�[*���q�ݡ���{�v�	ۨ��cK�t�!����j?�~�t���7��ܟ�r��,f�ZH�j�Z'��==��[�O'��<���W��(�� o�ƌ�h�����k��6���h"�acaX\t�w���mՍ��Rkf�A�dJa^-�W��:9��֙���2��W}��:=�j_@�L��\���Q�*Bp"7ӹ��~e̔57=�d榪2d�]8	A���k/��$�ߐ[�z+Wu�k��JLn�M����s��"@����>`1` ��t���׬�����x��̢���O�9�&Pٛ�O��-Rvz|�ʊ$��v9���*4�l�9�AD��J�$;�'��Ӊ�#ᡔe�D?t�m����i�* ʻ}�l�!x�,H��@�w	�S���Ud�t�h^��C�k/c������f�bP�T]X�O<�Q�Tn7��B�/�]b��{��|�x<��<ł���N��ih7ݗJ�_�x�w)���v��'R#mj��ş��"u:K/e�>y��p'�"��W��
dT7��=��A��8T�E��tT��4jEР/*4-`�,�
���ߝ�):�/����&�P��>��2+�H��l�h��a.�+��u,Y�{��6���a�"d�wd�ù�烪��3�H#^Y+���7�gb�|��Ou�[L�B���C����g>{�}^ARe�̿ܾk�β���hɮ>]luc����r8��
r7�g��}u�����#5k�e*�H��(��g�����`�*A�TdFx_!tr]����+mA�FO�%�I���Z�֞t�U���@+9'��M�fwl)��J�[MGϹ�VO?���X5(�X�Q�-5�LqJ֦�7K�e�5f��o�)�|����O�+x!��0;!����|mJ��ǰE�������H^��!�_!�~� \v�/\��CÚN�
��D�*G��0Y>���m;]�}���3ҡ��G���<BN#�[L���%Ϩ��L�A���еۆ�ˈ-喪��I�Q"Կ
��\���O��?���[���z��@B.����'= ��(��%�W��	���t�~j�qFn�ʧ&sO�ZX����NTS(�;��>\G��#����Ǵs���h.H^[@�VQ��� ��ӡr<���WKz��I"�>�{]��P �%�RX�9�m�d2�H�:+��l�ʵ��j۬�l��<�k<C޴Y`#8�.W�ܗ�Cpj诓ӖtZ�����!By���%����gj�|w�l:��B�)U�'�u%��'B�:����[ߺmtNk��z���O&���39��S4Q�4�6�uۑ__\xɢ��(h�*t�2������BN$aԔ@Ok��a18h�nƔ�2�u�J�ۮ(f0�NIl��̔L�(Ό���"Vz9?�u�Ui�y�@P����"4�>+�!y���M�El������a�zѭ0�S��H����/�;ԇl?K����Q�4�FL$�S�4�������)�!��
�"�Q�-�#��p!S:�6����y$,���y�ӡ�wڙ�;�j�ڞ���e�IEF(Li��4!1�&`�{���U.hA`(?^%ݕ!
��1�/"`�3�jG�6'�P �8�5}��{��̩�Cҝ-�H;A�č��A���& P⌡���Mꎰ$��$���D"���u�d2���28θ�� ���$�A&�FZ!i�2�8B��]�X�f����(_�"��~����Æ'�72 "�mks�R鳵�cT�v#�Ć-�&�x�#��a��`�W���ϊ��H]:8T�HKՊ���S��I!ݲ;��&tY3S?G��]��7H�_�߮M7}ѧ ��v����:��tIg$fus��פ���NN`��7tm�zW�J��@��-�l�A��3�K�n��!^�%	tO������GU��*�E�N̯!��U�yP
�g-p��e�0nv��A�b4���o_O��ȃb�֡��4����u�K�aH�2[0��3+��Zo�`A;��w4�d*��d�ٺ���/�#'�ÈVl�2Lr����)!n�q���';�B��=���9�����a�vm��(���������4=PM�_}��#�Ł�힇!)��d.5՚Հ��1l})c3���7Jı`ۋW���h4����;�kx����0���#!Jh�o1�Nľ��o��?�\Xh�f���2-:Lc���('P5eN��q�3�H��e���+ȼ��I�ե���̍۱�|��d�\�d���?�190�_�:!H�������=��v�բ��<��&=�@֚_����	~����E�f\!�EȐi���-��B�������!"aa/V[P��Ȧ�C�L��������г�ց`f#����J[��,r˻�!<�m�4>�4Xu�򐩫7�2�$�n�3���J�1���Ү��up�d^��Y5�j�zD��T+$�0�0�͈Z��UaǳI�ҋ��Bp�i�b��Eot��~	�/;^��֏?s��-��zq��T��Y�V��xk	pQ�#���	�(s������e֛���A_ՒG m�R�����)s��G��.����%6Z�XS�j1�z�-���ޒ��}� �ad]���h�NIqi2P�2f���IBDI6�q��M�@+
���ȭ���!+�8ش��@	�6W��U��q� OI���T��$�P�I�U�6�˕6�z��"����4��=��v]���쯫Ƨ���F��LE��/�8���A�"��pa[�^w�'�tO+�l��h��O�v��э���k!Z��^<"�#/FFY!���W�P��:�7���!�邈��D��e&�3��ʚ�1�r
�*h��{T`f����Hq�/�~���S��$vX�(��+Rz��Lq��?�,k�C�e�/�d;��iRb�d&k���@���F�@�~A���|5��е����Pڹx>Q-E(���Y��e�\w�8��A�4Hf�9v~%�"�뢨�t<�1[�*bn�3�%�Qm�B�Q�Α����4Y�N����y��a���� �i�kP�/�L=4����ó�2�:\|a�a�s�v�ތ�"<m��]�}���x��?&�����&?C�s\���Ps'GX>"&�����QK��p�t8�=�r��dJ�L�� �qgf�5#T�Ha�f�6�7 (��EW�v�*O��8��u��*kt���rE�n�}4�U����^v�^qpq�_}5Vl����T��g�K>I�S!�M���+�|��D��3w�@�Y�@E��Q���n��I#i5�ί�����#�j���'e�RY�����G�NǮ�XK&�:U�Y�X�p�P����� ��xt_�����wKv}���^o�<�$xG��}YM��"�Ae���c
�5.n��%��^�U�^�-^Z���,,~��v}�P���rk})��h[n}�������%ع� ��p8ޚZ��ؕ�\������=2�`�=i��ω�� �4=fg$�kd��`�`��H�a�"���ho\��� ��[�|�ɐ���hn<����Cv��D���U���ٱJF��*E4�QV+�Rk�2*�:�!t7X�.�S�N���?���>���]�����<
�_>u�<c���!_fDb�A�4f�E�D�;���|��	��Ѕ��[K���U��2�����=�
��ۈNj��?��c_�w����+A����^�����sJs�Ml��f�	�T�E(�Q��e��{�̒��Z���]�4��Ty˟�fT�".�n��x��Y���RU ��N0*f_cwM����Cr�ϴP[�|&�_��v���NW���T�U���)��{ײ6�en�{���<���<)�d�B8�t9b��;n�;�1�93f�d����*I��;t$w�>���۞�v�;5x�����Ab��$|^/�$�_{C!E �3Λ�eRV�*M��{R�.��pH#�!�m��s������<'���:��)��z<��lp��w}����r�"���γ�<����+Ň���J���� ���L�a�:����ƙ!����/��ѨT�>-Fa�	��	�掼�0��i(IQG���MW��̴h��w���pYAٴ�ig�EX��j�	*����U�����1.!G���S�W�hQy��z��͠�B:[�Ԁ�9naG5�T��Z�M9Y�;C�l_(� �E�i��v�x�Wc�v�P��q�LUh"����7��#��m'�HѿRF �IA!M�	���{��ӛ*�㕕\�������X:��?��x��<v9w��+�!���1�y�p�K��4�(�;��sEqy\��{p8��"�j��mL��A��4�X&g���)w�S}c��K�tY�l��Y/R�5�
��P�L��J��	 C���w���Z�nѿܩ
���=2�x�I�o����q�϶��D�hE�(j�ye��1*�h�����g$�,f�{ݹ7pT�97aq;vb|]�u%;4\e�7f��#�,o��H���(v��>�|�Я�>�|����Y�\�'��f�|�@i���6�`k���n[�}�`����h�M�������}�qU��V̽�<ȃ:��DL�E#�38:E/����q��0�`?�l�xb�O�S@�H��c.�ە�Co(`e|*�n�1�)�j����Ֆϻ+��7��ԣ�d��&zA 2��ni1��`w�-��`۽P=)E{0��qsdM2��_1*�6GE�`�B~�t�M�Sƻ��%0K}���#`�@F���q�T�9�Tg�NB�.��  	��x�%Y��`��������N�b��̰Tt�X"s�I/|��f��D����jͮϘ�.���	���J܋�� �]�����	U98)���OP}$f��E��ʟ#��F'��?V�3�+���`f$S��ᑶ��7
B���޿�d�H'5D:�|g�]��[A��*�㬐d�ʯ�Wa`8.j��R��_*����Fؒ�_�%��c�eB��_� �����8I�oK���3��}���3>"_�������؆�ֳ�̓3�0xυ���Z�����
˾�]�LK�Һ�sx˅X�Ʀb�����gi��5�Ճ4�2yr*t�X��JZ
d���F�c#?JG1}��G�q�Me��8 �������:�h�]�+l,��d�fc���Fȴ��VcT��7f��l�w
�;d]��T� �ʏ����d���ktq�w�UF�~��-A=�a����V	���S�f7�>ľQ	���>�4^!�ڣxOx��B�o��I4�x�h������,ο=
��T�@��<si�����a�)@p��8f<VI�o[�ua�"ZQ�؇���!
��!�Г1M8}1����
�ϡ�����)(��Ze�V<��lf|��T�?�69����7	��P|��r9�7��D��	�
t��p2��N��:B�����l��ֆ�ˁ�3Q�&���m:=��g�_m`��~�%*�"Rk�q!���2�&�n�p������uoq`f��UC1�s
u?�bt�B&	�\�aKV����P��,x7����%���J@���o=v��e�V�W�$$v�Gd�BA��H��*�_d��6����;$B�	9 ��Ǐ�{0pvi ���o��`I����F����֥�@Lr��/a��䉘�a�f��ޭ���od���L2R/v �e`L�@0���`=杨4;�gǬ�m�|�y��<+/Cj����1I��}h�+x��!
���ؕ��/��YS�C�z)`M6+�]y�ρq�Q��mN��������s�-���}�[3��C8����0h�B�2ہ�H�������*�,���].�e8pm[0�=���焙��+���.��R�g��-,�~����9j��W���H�6:����B���AK�J��޹�2~^���"���XYKN�ȝ�H3I&��I��+wh%��7p�*��`^#c'���?��Q����{:�D�У�D��R��yQ�Q��%�r�I)e�x̵�+�m)y1�χ��_��<�XX�`5HϤ�
���D�Z�P�e����4z�|���f`;-�UI/�8��\��Jc��EP���¨W�����d�Ow�[��\��O��Q-��?��{*/�0L�r_W^:�Y��J�.����=������3��ɫJ>��4B��Y]ԙ��o3�2+�����B!z�w��|� %)��ȧ�܋MQ�;!��))���O�����Ӈѵ�>?G�x���;S܏�̆��pe̺͂�1L�N��p؂��rYh�����[[�ᬜ(�K�G��t���4�ԧ�����B�h�j�v�5ٟ+�!<���:ٴj6�<_~���avɈ�v�0�:���ʊ�é�L6*�A��߷I�X*A?n��,{��Wÿ�%Ί>�1��,R�X�v�w�R(Ҙ>�>���&�\m8�r����f������t�{B�u	>s]Lif²[*�|]�NEE��'�'	�Ii��þ;Mu�3vH��;^B�P�>�6H�������#�3����ia�<����:�)<��U!�j�Y��u��?����rO�������Q<��9���C���He.�m&�F3'W�U���(�E�k�W�o7�
%H�{��S�?k3ꔡ� 1|���U��Z_-_�!o��J��Ӎ&�zW;*�z�iG6�H�n�y��4���Q�A[�}���+�'XK���M�8
v�'E�aj�㫉)�CfAF~�8�����`�+��@t��	큖 S#�Np�~���o瀆q�d�!���Ճ��1,W<����b����8F�A�J�4_Q��iR���2�e��}A��s���+;�;r��9�1�E��S`_��	�v�lC�ȁ�tG�ęd;|X�MH$���%���@[�5@���L���+jl?0ֿ|���-�4^��	������z�iz$v����i�^�!ho��X>�W�{����'�������y��-��~��M0uEiz�פL����Q@�x�{�ª�D�k���b�����دY�V�c����B�V�Y�(ԉ�A��V��"++Ow!�f����\�[�40���t��|*����/������B�c���S��s��PZ��\����l���g̈́�2y�չ
{;���q�s��gڗ+��֔�6>O�C�2�!�"y�S���[~�9��2�bGӦ���_��� iD.�5�zF�x"�-�#~�詽�	��O���;6��;�j����=�$Ά7�p��V&|"� z�G�N�.�Ҵ�.�L���]��QV�<�'�%Tו˓�%��0I��J��uI�J�'�M�ȘxUɛ�G��jO<@aN�1�b�9�p��Ci6�\t�dѾ���H�(9f�?&�u��Z�c����|�"9)�)8)�]�v9�絖��Y�,\��1�H{�d�P�@�9gF &`��������UR*��Q61@<BF4�����>��+ڵ ����ց7�f:^ ��͉<�c.l�z�X"�ړ)X�aƄU�=J%Y7TJ\�?j�,�d'�H.qe��4��^����d��m�D���j�x�=��{��>����v�d��қ.��ҳ���9��D@��E����:`�I�P���JiLaK��uȪY�"��%q�M��NlN8�*��U�� �	��7�`�������V��A1@�,�s_��V�jȘٽh�_�r���(9��e�b;,�._5Q�������_۩��gt�^����<��=�z��L����cSjr��+d��m�[n�-�2>	���^�FZ�[��JJoՖ���(r�7�%V7Y�=U^_()�s�)/0Ce��*��8�r���yHs�4��6uY�{G39Ҁjjp�|K�r�<ԅ[�9MN���E&��o��ŉ��zyx[���]���4��g�D\A����PJ���R�X����ҹ�f��8��aH,a�XEo�j�f7�v��WH+�ͤ��*�I,�?�g�kCZ��^E�?*r�i�í�����+Ϋ��3�G���A&���l%�.EKH�\t_�ѯ̔UQ62P]8w^��:rNr�̘\7�����O�=�z��NOg���Y���3���&M���5��ŏ�++X������N.R�P��dc��!�G>>&�&�}/`��^B���v�d*�����{/�t�`�J�`��~��Y3��W�q*)>��2F�`�$����=�����Ռ�~.Y����RF�d���U�ښ�"��1�l%aic�E�Ħ�q�7��xТ(!򪸖 Ս��	�	M������7�^4�j����D�έuߥF��(�Pc��8s��O]�w7@���KR�6�ݍ���M+kQ^⁍�,
o`8�UT�d�G��u!���y�s�y�U�������t��]���iq���&/�֛�)���_ݦ�Ȗ���{Y<MSq�;�����J��R��柲9������`t�B�\�
�	�Eq�<���a�Ⱥ`"�zm�i���y��N�/�fbD�$n�㴵=��]�x��S����骩�~�;�ы!K���R�
	�68��(�V_�J>����o?��Mi��Υ	���q��ÃU�}���Bp��u��B�Q�^���?��v4��hў�f�9&G����n��w��A|�Z�M֐���ѕШtP��=�U���%2�s��2�#[:A�X�! M����R{�{$�l��x�t�r4��_��E�[�P���Yh�0P��l3�U�1ѲyS�^~�:�5X:Zz�92d�c%����#���14�e�3�~]�\��d~cf��(�I�?�{g�FZ��#�Қ�=ȴ�T�>)T0�7\%>?�r���R}&��7
��\��|�p�����9�'VX �PX9���~�Mc�^r��̰���>M+e��`ta�c�4��`|�1Aςn��\�+��Ѯ.��֡���/JB/����Ry ����I��}T���	p��4�h5�Ƭ�|�K$����'(��v�ALVX�����:F�/��ɪ��^�_�B�iF++_6����o����wT�x��tb6Yw�G�%������b���-}g[�9�G�����p��o�]�ue�� ��	 ��:�fT\컱�j�>���v�f�@혈<	5���o2o��G��G�~Y�	~懶i��*�C)	�ɚ�����D�%��U�j��9o@<��,äjb��gf� Df�8ӯw��od;$��xᵛ���<�aF��%�suD&T]a�f����;�u�ȳ��,�J��TO�����:�c���sϡ$(����xZk]��=G��_<"yOȫ�Z����u��Y2��3tP�
�y`�;t꼙=B#�$������UUp�jM����V6E�@n��4�j�tYe$�C[t���	=%����XV�qj�u")��lk����;ϰ7ש)(��M௿c�Ĩ�2k����<ٮ4�_(�Cһ�K�H-����lQ�z��+7Kr��f�Gh�,yJ^��@�f�)L4�qq�jx�6�mxٞ[�(��.A�6T�'س��M��D0m�1/�	kD�%�&��o�]�>?�#��_"fq&��(�i2EX�wx򀊄��z~#[b�i�YC�F�,���C�}O(�h蜪ت�雃�ŀ�����:Cms@zC�qHS�iLd:��5%}��k_I���;���e�fK�gf�`┒���t)-��9ڣS��1&�l�dX��N���oݖ�h)�s*��}��S��|N��)Z�G���N��Z��Q4��h ��l��0Dp�Fy�4vv��<H&m���h��*g�^Zmf�+� ������6i���u��_�rM��Yju̦N�d�c'6��fm�h]Jݱ6nP̘�|G�ò�+�6�ty���v6=Y򱒒�c��mj�#j�o�CS2�*O)���������Km��쾷MW�oa����f�WU�B��z ��g&#)e{|1�hU����S�v�Xi���E�lR��4sv)�5%|�l��̯,ƈ��6�O��ts��I�`$~��Ĉ�Cݤl���d����0�ώh�u�eB����i�@~UѤrs� �m;|��1#��*~	�s��i��Er8����;nm�	َ�ai�W�G��}���g�/�iQ~#S�۳J1��k�׽�ntY�j̟�e��4lv�)��R���1_��_R��)
����������G�m��dD��_��~i�9]};j����b�Օj�Ec������j����z�.�z��IΖ[��d�cC2{J���O�~Q�ڹ�`K�6�8��9/\S�� ,e�.ac���	6@V�T��}}�����2뱐l	i5Z#�D��T�7#Pq6�ضI����v_�6�w�U�o��o[��h�Gu(|�6GW4��DN�q��=jn�͌&�	�g<��E�Z8�1��8��re݋��g�-�ָ.\O���{٨��Xp�Y"3��PQtѺ6۞�\��\KL������85�3:���<�� ��B�q��/���Hm�q���u��ۼ��pT���!�V�: �X�l>m��R�D���Kbf������[�#��{���bc�	�$���X��(�>�r[���gdiԺ�����]�n��:UtT�H��:�'U��@8~�P�/��0��[(�G�e�4�1���je�E:��=t�ٲޔ�X6���I�(�r	3/Q�C��?^��J�]<) -���V�^�cr�Ʀ�%F�$h^MPH7Q��n��Ȼɑz�+p6G8 a2�U��m�g��RǷ�u����2���{��D�Y|�ɠ����$�,�"��'��|.�b�ᖽ�$���g��%�Ǌ�!��B �[8N��Y�9��'3��]	��#-(��)Kk�E���F�syF�,������f�u~�t#�>`��p*� k��y���ut���G-�+ԉ�7�-��PbX֋w!O�WC��bu������d&�p]����m[(Ȓ��	�Z�#�S�߫9?��	�+��a^���7��k9ز��K�nH�	q���eV�|�hs
Gb�핆�^���i��F���+��#����N���&�/e�hl7�����\t�V�KNC�3� � ==w�z~�7@�ñN�w�P	�o�t�J������0��Κ�	��R��1�z��[1Ѯ�iL�籊�7���}��('PZNHfq�GM�d �v�������/q�_b�J�k�M7��zz�J�q0���{��O� �	�т�RUk��/�n4(U6�#��[��s��$����Fe(Ų�kU*N��lW�N�{Zc�z ��tP!5�^pQ��`j�4k	w#�{�-ܞY��$�W^��0%R��*�����>�O���%O�	�MZ�����J!0�N8OL�Y"d	3v�L�B4�Y#�;��_�?o�=~���O�,��Y�����aʺ
۩V�R�N���"`�c���E����2�H-p2�������*�Lܟk颷�[�"�3`rK��`K�׸��
�M�`��XS@���-.L�=v�ׯC(8�]�1K�Ko����i�PE��
8a�c��<�����ͺ�2��j3f������� �vg�*�^�N���nh��	���`^�P����@Q��Ρ���?T��(?)�!���&�8߀21g�j���Ꮢ^�s���YZ6cW��185q����w�SOF�/�bq$�>C/V���Q���C��8Gv�H���%5�S��m�'K�Γ�sR�~�I�͑�����Ok�>�����?4���h�m.F�T;�՘��ln�&�_�ڲ�kϞv�s��/K<�O����o����~���l�G�/9�qyϱe?&#�*�K,NP�����B�D�|G~�U�P��[��
����<+�k��~�L|hB���Dj�����`#t�@����UEW���%��'" �w����O?8^��N�-Z>��D�����K����I���r�"2'{��I��c*'_2|�<+ZO����o_��m��y#F��@
�y�ǰU�~{^��-����c�:��W�v��i��d���]2"I��%� �G����|�OQX�1�����������F�5ݍ[�!}٦�M,� Xt��A1f�x}�^���'�0z]|8��˖��`�&�h{��Mje��a��0�Xr���ę K�0B��y�i[�>B�WJS�h�R=���=�h�+����פ�����M<)��ցB���x���G$ׄ�H�)"g<���)����ʠ��}�E�#G �$\a�2WL�R�"CʳK#T] �4u��k�w~��h ј­��U2�Hy�%,1��k�~���1j���]�>�QQy�x�R��̚���\����~�'�m�u�L�3����JO鲞QLI�ǩѯMK�C���/�%M]:��V���^�haK-m���(�����f~18�Nzܵǌ�.� ��
}�O��{-�˄���S���2����?X��g�%'�*�w���E�����PO'�g�^Ȗ�[w���0��	f	Q�j��~��;�=b$�!��1�x�4T�
'�G�� ?�4iY\�#u��I{2���A�J/M�ְ�q�9�Cs��R�!^ �Z�A�I�/��Dƌ�fg��H�y���5�x�=6;)C��As�}j�6��hǶf��ڵ2�Wg���}����凣:�4<���(e�w��o+d2����1����+�Ѭ�>���4�Q	� ya�O�Q�����ױ!]=\:�'<���Uq��cc����`	5Mˑ�]�X����'��l2���
,���f��Gb=c����EذE��	a�A�b+��/_�S
��@Ѷj�l���ւQ�E���6|��
@���[<�y��dc3%{�/�ѧ�P�a�0�V{�K �5ɰ�xp�&9���gw{�_�쑐wt��"�Ý*П��z
�M\|z	�y�����;���N�����fO�Չ=$�j`eGY����I�h\�[���;0�濂\|C����8�@�EU�m���ɰQ��~ڍT��&�\�֜v�^S����n��N8�}���%1�Q����ޢ �)��xQk������͜$�D��-�H]�d*̲o�7�����a_�������Oz��V�%m3 �|m�9�Z���W?N���fͣ�;0��3%�7ΨtD�b\&�z(s86$�Y�&G58'���>�u�jB���3ϵ��b��ֹU|����7�޼��ыg]����!������G�$��U3@鮠��ռ��"n�Y����:QS����F�p��� ��P��֡�l#�"<�y���UE�����_Y��g0��r)�.�̅1�`��y�T'$`�� ����-���{`��AY�ɯ]���v�yX�)X���=0ۍ�v�~��#Um,�-�]�K�]�E[�.�5�tJ.G_[Z�;И<��*���=�Oh�8���m|d}Ɠ{Fb�^��"�k/i�^���+.��eS�h}��H�D�~��������ͥw��IR�}�����������4��]LZ���>2���a�]��lQ�\�w�f��fN��2|�&kM�?T7~K���j����H�����#��1�&�V�O�
��~s!w?1���>@=���ٛ�잰��|�ڕ]8��b�`qӺ�W�9U4g�Wo��y̸"X���ɥآ�3�D�Q�:�я�&L����#��dnY	ܽ셢ύ�����		�!�C8� z�l{$ b #�#��L��X���%,y,�V�Kީ��~���
�}�T���� ������*+iS[e�P��|��a�\���Ũߤ��/�F�#�pYĒ����'1����Y2�����.W�a-���GΞ��?a;��{�C�34�B�v��8����	���E1�z9�@�����+�n*M���bz�ݨ��,�Gem�E|�>�*��\R�3y�4����W���� �lr�)b����@�o�e�g��	�u��Tׁ$nt-;��3�!�Y���FSGiUC�-8nx͈j!7���}����T(tH���d����\�5]ծ,M�R�@�fMwTQ^z����Xs>؜0����|b�u��t�C��:`��.�������;�0��RT�.O�-��XD�=��%�\�w���V�
f����oF�:�! ��e{��5�lo�J3��vc�7�_�:���b!��Y+3��0l��F�[�4%MOPx�D�8��_]�̻q���2?�_0G���+�F�>e縰8��#l	�����C�R�k%7��h�]3��VD�DR��>$��\����D���>{Z���C`�D?F˚�?�v$�c;#QB���Uc��$;ٚm�nc:��iN��l\X)�[߉�:D�s�Nq�)�k���l���F�Azj#�d��Ԏ�T}㙷��%�4a�;��:�t�jR�yzp�ˈ��|������Q���X�+��gZ�H
�������*&q3��
�-ƈ���9���M�Զ�����[~�x�,�E�K���q������<uߟX��H��7��ځ��)��4��^qD���#K~��FG0pUSU�[<�(}�è��CT�c;gs�Z�f:}�s5w�����U��*?�+?KZ�vM��Z���IK�'߱]R��^�4"s�a�2�dZj��i��[��і]��Vc�$
W5P�e`m���'a���8���*2֟���{ �K#R�!�i��)_/�\��Y�C� +]�XW��8�r)�iOD?���ʖ���߿�Bod-��8�������@P'�����&L"��\IL�e�%gי��IJT�i���m��C\\e���DS�f��U��u�d�5Aab�(ʹ��t�A���:l�x�,�̚7T#>��8����p40���|�k&G��c�M��֥}W�s: "�{dA�o��F�r���,1�m�X�o�(��g����F�t�bt�-U�X�$�}~RQv�����HJ�2v�gX�&6��a`�4;5�W�-ߦs�D8r��`�IV�
�����ě�WI��?���е�Hb5��Xu�jvs�B�?~���热W��#i�N�P��ךZ�?�;C�F��s�% ^\Ə%���x�@�K��DDs�M���.di*�0��z�z�I����z�MQ�������*�����+ 6����?@�VB���r�l��I��R�{����"�n!j�M�KW0��8����ڕ���L�'�(��X�>0��<#&<�?}x�]{�GX�eQё~��-�t<Ϥ�����#��䚃����B���?�_v���jc��'��M�u��:����E�[���rN:p$Z�e*ft�
S�@1���ꪠ���� ����Bܾ�u�i~RP�-R���a�������v������;��<����I���i���5�+������>J�*w�z�] ڢ��^�+ѳ_7N2�{��������YSm�M��j������{/�|�:��f��j�c��Yg�l����W`k[��aɁ0���`�:ꭳ9xs�1�Z*c��E�[�(fJW.����T<��p1wi4Õ��7����}��&s9�l�<I����F�� �T3�3�S�F|hr����ؿV�j�.��̃E9��k�z�XB��5Am�i�-M[f���؀eS���,ᵉ���o.�x�.G'��M��F1Y���\7_�ޏ��6�`���ȯ2�U����Yv����ل�s,_�\s��_��Z���&�zk�)������J��ư�����k�8�Fu��fy����u;_�l�t�Y���e	�WTɝ?����@	�O[���t�R�S;Ξ|�CЄ5Z���!��dӔ<��掴���1� ~���mU�h� �UG���?�yY)��,��{�'3�/P/� �nZ2h�Ri#i�r��*W>iY�Z��7	�׹/�:*����	�ნ�e��x�2��T=�a�6 a���QG���z7� dg�=[CX�H�DcZkU�+\��8�m��$-������]~����Bkd֐�{
��U�r��ӛ}��L�çY�R?����U���[L0� 4pU�f�����%��'�L=a!���<B���������?��e��s�^��|h#̫�i��8;�07��t��M���׎���������	����������k}Al!��O
�Qa���?u��GyZ�>ճG�d
>�����~�8�0Dm:�E)�����yo�wo�{Dc"6�`�=�rj��uX6j�vQ��sk㶢]��������܋E8K���GO,"��i@��V6�L���7@R�3��	�F�G����u�����](Qj�7�3t��8�X�Ru�ko����O ��d,"�?K-�ҳ���͚���_y����O��u1���
S�zg.�sP9�E��$8Er{�8XSɭR�.���M�D͵�����[9��)��=2
���I����h�ã���ߧK�� '�>J�����8Z�nU4sǡ]݄�(�,�����$�@˧�~k#�g0��u��K�x��}t��h�LhR;d�ar�N����y�T��?�o���&��N����v2����|KA"I�Q�B��x�����y�����"DX��xL\-��t��<���F�2o�{�Z�O��7��`��8E:�KI>>礜5`���>���oZjN\���XEUZҭ�M�p	�<~�<(�׍*���z=��Sz�J���?{%̹�vx���/�����Vq��f7h\����+�x�䟸.�c����^�!��r����^��l�uۃ)�q
��ՠ�sGɮ���ra������s�m�'�4���<��b�Pٕ�	VG��!'Kr�����}��_L�f"b=F��>�Ar�JZn�4un�)�
�Ԧ���p��H���q񧩫r���Mm���C��I��QnI�����ю�����M�	׋�F1��_����NA$���l+�^4T���é./@|3�j3AE�m.7�������c*���͍Y�ʹ�����F�Ї���!��]��������N�V�AU~�2.=<;��
��I=XP\�0�S��H��lH��t��Q��89��R��?v=( ��O� I�-J�41�=�\�s��H�FԹ���c���	:Xc| �wq�N\:=ڲ�H�V42��N������vrV����O�X���D+㰥�g��YW�Ӹ�O�tkm������E�!b���E���c	��7�q�xU�
g3K]<��F,�d��H��kS�Q���ʊf�hp��u�)dۺ�[٣��`�MH��-���$#�uT��3R�a�K~8f�@���!�&`Gy�Ǔهrz�r1EE7�g���-��vC��v�b������3D�$p� �N�B��I֫������	y�{(4lpU�l?�m�l�H�!�����Y��9G�����01pbN�g@���X����V�*��g��k���'j���`怲�a�0�G�)��^�����N�y=CX%� �%�E�g1+�v��=��F�����\֛[k�U!�Qz��KLw�3Z�:�� �qTL,jzc�����ٓ��G[�0�U�3�`T�����܎v!;�:���E<�^X�La�k���ŭ�WH�0	l��b�]S�%E~�h�'�ǥ@�m0�)��M��s��@�˺ca����&g��K�__��ٽ��A����-�>x?�.�/�$��F�}�^��q k�S��ZK3��TL���j'��|7�%h�C&	̦���� H����X�+:1%.��ů2�j���;�d��տҮ�`8Զ��~��Ԗ����
m�Z�^���hq�U`p��2�I���[%�f��!H[F7�t��,�o���(*�N�w$׌�������M���VH�"�Z�^��L�+d�k���Y�E#g�V�����=]��o��^w�9��_�#+��KK�k�Ѫ� Âz�]*���.i������Q��4a'�:#%˥�NaH��#�\{�/�ĝ�E�/�%�r{�`{h��fD&�'Ә�y�g��K����i̓A�Ƙ\���~����2+�/)I��ڏX�Y�x?�5�$�O8���v#�S�<>)��D���'�`p��3f@�TUJ9�p��i��Y����g�mo9���sз&�Q@]�X`5�v���U�b��kh%�re�͊&G�a 
�����K�Oh(���?㽯p�@3�ǉ�6��o��ܻ��U���>�+�+�~����e��9�I�~�f�Z$u��:K`(we��}w4;�F����\�z��!�6b쐧�����mD�!f"�A�un.�,�ѹ�<h
%�"3
b�W��cGp�����t�q8P����g$BP�h�w��*c���"��\X��5�z��H�Ɂ~���{n,Ֆ�&����Q�6!�3ԅ�<F�/�#����L*���6R��ɐ������k�yX��+/.1^-��up�m�����Y�K�i���gw1�G����	w�#A��+{��QT��3��U�<�oM&�#����[	���W(UJ�n�p�����,{���%IV�d� �SJK�sO��d!\Li�WŧQSq�����4���cl�)�Y`�u�F}p5��<4���|u��AyԱ�sv��4���oi1�]^���-'O���4�[G� ����j�`u�R��/5\3�M�`U^��*�`�Z� ���e�b_j6��������x��Y�R��<�59�˛�LT�D��E�
���d*�7��s�z�(,��F���N�u�<�ڲl��~�L�M���e?�3F"QB-�����A^?W��2p˰Ci� �)�q��/ɭ� ��
����Z����`C�C�h��Ч��j;*٢,$HI�[����x������k50������"�R_q$nj=o=)�8A�����_�Ӎ2���Jz	$^~�W�9vB�`z����d� ��+����΋�X	=,pH5Xoݣ&m�kF��<����a,� ������v�����0Pu�$�*6TN~O.9���8��>���;��b�Ie�ǐ~XC�ku��ڢ�(��_�� ���@�#���������+��>��a�x������f��2����D�!^56=Nq[��ar�ѐ�	j�\�L�.����C�ɇ��ҥ�䯽��{\/�5���_w�FuB�1�K�32G��*��%��nhz�U��<��/�Z������ytJ�*~��`�j�bYp2� 1(`��lb�RD����2�[��V�əϗ;�D��>���}c,E*�=8u���G�3�A8U�T�:Q:1�E�sP�m)�q��t�(b�=�qI>~�\�q�E2'���M�pM��!������W0H^t�w����qD��X}k8��l�����?�`���x�/��L���������9�~��F	;���&�,���Slv-�����R�#��_0��,��Όz�II^0{�T�>���,�ﴹ_���F��S.ǖ�Z�L
�w�o�^�O���ȭ܊K�a`K�kT0���lt�=k7�3���T\
���5��sq s��{�n42�⥧WόT������~5^��p7,-�
�W[C=�<H�)^?]��?�*9>\�;gf֏y�d�����Y6�,�-����lG�����@y<
+�q�=|�7T�8*�VaqrKec�J�
&@<��>4G !�a�J�k�W.�r�H�ݣl�y�T\����;Z��(y$G��vW)1M.�\�$T>'*�C�e}�=C4~�!�(
��cۨ�)w��DPw����Ͱ@v`��2�_�|�����*p�~�����c�;&0p��������K�	aM�Y�� w5[@=H�@��%c�ltҺ:	[�<~��"��գHz�# )�^�-��˜�	��a?ʐ��|��$��L>�v����I�?�.��j�[q�mw�r�Ă�#م�B3D�H�T65��"�je��ݜ����Mu^�7g�e2��d7*/��W))�p?��S�2�ȃ7]Ɵ�o�%b���i����T���Q��X���>묨���$�z�Q|$e	N����0Y�l]��0wfAJ�H��q��U���3�Y��� Zu`��!����Sd��$E�RZ��?2Q6P�ҁ�u-�I���5|t� PA(�X�����?z��Q'���п���ZZN'��9C6O��S�/<���gze�(�AVn��ٸ�����VK]r���1�a���[��٘Si�䜧��1�p��KJQ"�׾>ќ`�MQ���,ˏ{��M�磆o�c͉T��h��q�r?�N:�1�m��K޺�WT�=5��6 @Xژ+�!�w���qV��a�������.ڔ��,K�3\�xRc��!���,����b���N�3I�t��oI��9��x�]�7oe׿���Rq��1��^a*_��hO$���R't�QN��[��`΅���)#U��̟�����_�[R�7�$��?[��7�T���U��}�r�|�=�:�Ād�aX�wC1^�mH�+1i8$4��Y�H���/�b[��L�0zK>̈�����k��ݐ\�ò9g�|d�eq�f7�qP�����c�Y ���\����%ŵ���S�n*r��e�=	�+b�4��E� �ݕ���z��FS��Ɛ	��'k�c�M��\B��>ɗ���#����Z��Η@\���A$
�	�lX��  �+�3�A!��#� 
¶X�8L��3Ux����P)	�bPmDٌcr
˅�1k�CC��%������?�h��R�@k�vjA.��� C٠�>����N�����h^!�e,�<M��du��c��sܻ$��^U�'�^."��-rlS�D��bU��)յW��Q�7�078���u�$������w���H�z�R\�Yfb�u���(A�0*��vz|{�ZO���ι����a�n��a�OHD 46�S
�(N)�F :"\��=9��Je+b�(c��eؿr��=�e���'���?���xBj�	.�M�fP��:��f�d��6��Ahh �u�2�|ĖגcGbP$K��@7�x�J롡��,��M(��QN 4U2$�/Y�㲶�����)'��x[���Jt�>�̬Q��J���n�mU��Ua�� ��n}y�=��f����1,Hl>�Y~B��)T7$A�A��Y	��4c�R�x�!��)a�b�ir���y�ͅ��mi	����ː�j�i�֘��@��9���%7<�l�����NI����kǈ�y4-�H߭��zvo��Y��� ˏ�V�b�����q<[����Oנh��(%�d8�+��K6l)ܰ�����b�wD��6\�jm����=�R��5ig�uP<�}A��IkW��?���M��04C�����]vb���e�\�8�ꥢ����Т� v;bY�jiF��H	ǭ�l}�o��y ���py��죁�v�Z��`�����&�N��Ԇ(�Q�NV0y�o�a���Y|Uk����d�$���	gsQ�0��#�J�i�o!���h��F�{ƛ|��}����>!��L����fup)pk�	�Jw��q���y��Z2�!.�vR�~����y�/�M�T1L���N쬆+�`�ٽ6�Trn�"B���]�I���8� ���e���;W)���@�����3�8��LY1��l�}r�F��o �6�}�@�H����/�<s�.cS�a�N�ٚ��k*,�C��w{oc���'$����'r�W�[�׭3ͯV-���5��,�6|âA
mX��*A$�0<�,;��2hp��I��9-ӡ��H���ሉ�b�-��o�]p���,�f��D�)���XQ����)l(.@*��u��lU�Ǽ��W��^޶xȝ�c~�mo�qh�=lg9�j�ؚ/$�����t�j%O���c�q�DH� ��ɓ�$'$*`�`R���X'C�i���
m�_����1ۈ-��$�"{p������J-�a�d
#�8NV-�?�lG�����3��;���E����8��&�p�5!�¥�Vq1��ۜ!C�4&�K��~�RK��k�?��SdM�%��5��p��oֵ!��TԻ�>??Wif�X}	�Z��W�7�a���.E�]x�&P	��s=L.aL�bqe+D��L��!���81xѸ�,�n੕tB�W!���6lWCR 4=S�f����nU�QȦ�i�ؼc����_�/�A)��S>k�K��z�|F���`k̵��p'�λײ�Fٓ��황99k�n����h��8�煰.�2�`�	r(2[(���ҁ��d�K��1��)v���9�{$K����&�`�"1������z��QR�c�6A%��lV|+8r�oZ�f?�ę��i</Ύd? G|r�Q-R�;����f
����LI�|�t"T�T+�Ñ?@m׈2��l=�$���3���\�a�]��I ���ng�WB���4�h�d�+F��)��A</�Z�R�����V�"fsY߰2�1u@�P^��K���=~���u�&Ъ�!�^Wڧ�6|L�d�B�j�C/L:L� ��.���k|_3d�ެ2�_�)=��q$B��SH/� q��u{c�W�\ⱁ/Ъd��,�U�m�2�s�U�-X�Ы�8�&�S�������Z����� 6W`�$b|����𓍽���@�q*e�Y�����vz��2��r�����.��B�bCٌ̟WP��#���ů!�VW���A`6�u�a@y�Z;\�K��nw҃J�4��ͽ)����4V㦭H��S>������U`^z������͂�RN� 4�g�;��ؿ�@�r�]7�����O�w�!��$)�|ʨ�x����I��4��F4I5�n���!��]���}O��e�0�H/���Yv"A�:��Q�Q�gΠ�N�!�} �%+HQ��5c��V��",�q��H��>��7��b���������u#<`b�m�8�������blṂ=������Nz_��v���Z�!�a�u�	f���!:�xc���Ȳ(�rʽ�Sg�}8y|�e��m����c��<�3/�'jI\�ݜ%�ب|,�am��5��F�!=UH���f�-WlmBK$l�%�i2Q���j]/H�_ǥ��8ه�*] 3����{W61��\�٥�hلӬP"l%2�:����f�挨�=�ݼ�8�nܙ���m��_�G�LX�~#�&{���܅����@����/�4D����;��i ��U���5\���a2��b{n_�<H�_�Gg�Xֳ F5�2Zf�(�c�M���Ӊ2o�Gkw��w����[��3������M5��`ߦ�]��
�0oO��>�5���'��ʎ�ދ�.���+�� 9&��&!�D��H-+)��0�Ԟ��m�����imB�̑s*��/���e�砬n�1�;��C��<t��0�T��J~�6�2��7bҋ��g��t��UE8�[�G!j̤o,%��R�Ǭ<qޑ���U���Ժt	�` K����pr���G��It� ݯg��HR!���Mӄ���IqW�/�ʴ��/�.���9�Q.�w�G����3_'TE��߆5�nnL���33�K�r00d�����^UY��\c����.1Y���",/F-�o�$"r5*����=����td/�����Ғ���(����q ���8Ă�Y��<mq�	?v�ɷ��z���n"���b=#ƢQ!�x�	�F"�A�t��2��5�?=nY7�X����)=�����e�۰���OL�C�Zm|�Y��f̈�DФ��z�o�\��א@���p?���Q��p�W�޻;ؕ�
!��Y�dT��(L�,�Ko2:��,�w�\T�F
�%��ͦ@���@4�?�����#��{x�lCR��iTw�}��E��9��{_������-pP4u;�
,��Υ�r�yW+�u�;b.v�$���1�,�@�;�Do��r��?d##w������p����ϰ_�
�b�²��>q�_;��N0!�^i,����ܽ�PC;	y�/�^�z���g��1�c��>�s�7]���L(��p�w�����񝇉���^K�M����~x�
A�to��>	����*\ZY\�P{� ��l�w�R��`j?`����SW�mB��I�D���X���M<O���@ݞ�C��q*O�4	�
w0w�X,�)��Ϩe�̽S�,�.t�$4��Qf�1NS�_jO���_B�D����ݓ� ��a��-�"�,�T��d��^�=����Z�>௦�0��c�`���C���^�$�Y��w�3��0�i�IЫ�!+*~H���N#�UƩg�z_+HX0��ב�t��#��)m���iܝV���-����@������Ic��3��'#H-�.�.!�~�g��*둎^�iݨ{���g��!�R4�[Tg+������9do���p}7�i�{y5��f�|,�[2�� !2�r/H""�7�ȣ� 4e�f��Fn��M��#Q^�J5֏".b)�^� B0@�;u��BO=�a,RDn���U�s@!�[��9^�s�V�gZ���p*ᙎ�w#7»�3��뺽lU��X�j�]f�uQ/�i�L?8��b���� ���Q�Q����`v�,8�ն+�����BU(|�*a\�5X�ĝ��on2�/l����0���5�W�,3�F�6�17�
��h��9Ť�0Ć�C�9s�m�?�xaĀ�'�b����f��=��f�֟��j�\D�3���oebl���Ԥ�4��� ��ϋ��% aws8jH�+O�1�۹nxn�gߩq���j���O�܌���=v��*3���`M{�3�����C�ܧ]h2�x��0@��%/��0gMJ�� La��U�k\9B������x��s�]�f�������C�B7��B`��顑��N�ێ�>��_a:XV6��e�P��u�*�QS�X����f5��?-jȒ$QX@`�p��������l�Qz
���6<bZ���`&@9�y���	_t��9#�Եe?�f5n����@�2�3��clw�ߔZAVl�W%ۻ0xw`�����������j�ߓ�ﹺUZT̔�d�^��K�˄��?�'�
��h";��0�)�n�k� @ N��"!�K��#�LMZ����SM>��X�FŘ{��L�r�����B��|V��U���\�z�4�UHU|�ɿ8MC���El�@�_���D�ٽ�56�
l5y8ɴ�Y�x4|����NGɅ%*\�t�p�N�bh�K2�夬q�UQҌ�f<���"e���q���Of����3�ă�f��rQyw
v�pGUޘO��q�$��L�v�1�k)a@���g��-y�]�F�3A~ۙ��:ڋ��)��O��nE��/1;������\8�������$��^W�X�o�f$%��o=��t9G7���H�k��ON;֝;��vO��i6���f�H'#>�/m>J��ז�ײl]�p��Y�'*q�ƃ�p�*��}8hT¹���Q�$LF�G��W�7�Ux �� ��ƈF7e/*F%��p��ucg���_6Q���Q���t����X�ۗ��"8�P�����:,ӽ��;�x�9�Eܪa�+�-혷�?�ئ�(��Am�X�t��P�n='6��r�,GRU&Q.�s	3��	�Q,�B㧁��PA,�@�n���˧�P϶d)s������*��~Ȝ����D�|�4ڲ�d�\��\m��ܑ��9T��H�G͆������F�ƞ�J�I1A����ۃ�$���?;��;�lj��%k�|���]�E�'�JJ���Om�.j3%�T�i�����x���%�ƺG��-�v�o�����L¨�D
*)�;�V< M�E`�6gH��	_�R�<�/��ϔ�m�`=7���B�"���O�S��� Q�h@�֋�u�N��0\k�rJU�5V����׎y�]��1���TMk���f��K���mS��k�"�KP����Y���%��o�	Ffć�!�lۀ��D+�Փ����uϟ֛�t�=v� �u��򑲡���`7t�z��v,t��!���������q��(w����;��B��T$xD���WcW=y��5���e��S�g��)\j� �!Q+W�V����јC ��Oh��Z�g���K�w+�E[쇺P���\O2�
p�ծ)Q��eZ���gf|k]�z�ß)r��x����fO<b1z;���W!��ۺ�-�?'�D@��o�s�]I��bz��	�ڡ(�l友�uVL�o����M�'�U�&�k�����@�� 1�j��$���"��D��"ԬkУA-��n�D����?���Տ�;M�@bAg��-� �hr�%t��
J�z��FU��D�y��H�Ú��Ȧ`�n'�.+}Q�1*�u��T�$|���E3�Y�,�-�/��z�F��
���0"V�	g���
.�Z}9���@]��3^�S�1�UX_����R���%2�}pe�g��,�Y��&��0}�yȍS`��r�~O�ɛ�Y�?v9ZV�]����*�΍#�[��RޮU�̐�,�~z*$<Z��c�Uv!ax�Ԙ��zmh�F���B�Xu�� 2�$�R�|�R�*���k�A�&��f%�̖� ������ >�2��8J+K�� >/P�G�[d���d��(��)��n&��>����M��2e6o�d�f�+0T�����Y���%z�D&0�b��!�<|�3���؋��[�z���]{쒱2�X��M?h2� �p`���~~HbL_�s�ٖȘ���^'9�Y��e��p�K���R0���^^ ��@���<�ޯ,O��8��ɣsK�&$�+ƨ���Z�v�xg��u�s�"\�1����g)��~k�2Z�ג�h��y�"$ h����e��"$�D
�Y�ǭZ>1�W'���}�ކP ^�U��4sl[{V^ p�כ��8el�u=��QV��|��6�+�&LĬDBF_���ϋm�yN<�m��m[�׭�x2?�\^�G׈��`����H�\��ZPG���,�Iha���?�z�ȴw������`����<l��u��<5���?�����Z+�#c/��[��Yo�K�<�[R����<QW�H�m����-h\ѱ����vC�pȤ�g�G��e�Mwo*J�)�ӏ��ߵ��&eK|R_:�ts��u���o��|�7�+m��^\gn[�����_��qb�̦#u���^\rр�Tʭ�M2�R��!�'�����Z�ܗ�$D�w��O&��&ı��ͱlz�'d>�V�T Vm�$�� ���; 9���e�ګ��"�������8�ŵ`Y�s5(�)�ƈ�m<�#�K�a@��.X�_�)OcU�%��NБx�C�l��t���1c�Ĝ]���j �W-�����Ls���}Z8�uU2a�z�3��[�j=�9Ō��8�;V�H�ˑ�~�)Ο��:�U���ԑ�~�x�Fg���n���%��Q�x���r�WE5�(�;A�?/n���4u��1N�O6��O��=����)��;큷�?��NZ_�ʆ�̀�R6FN.R�c��yES����b�1ȏ--z$`���qGнoCȅkt �y�9V���4)Z��젰�}����J�"�|nW.����t��8��{�f�=pGoE������/O���ɯh����;���)=�6 ���> �{q �h��C/�z?<?{V���裟��^1��5}m*�牄�5����薌ӛ�ϣc<i��M�����Y+���Z	VE1���/�qw�k�"�#�ظL4s�F�ZjX�(��ğBֳ0``�k�ӱ{��=�1��"���G����������0͌�U�������b�)�1��bV���xz���o�v�m�ި�jWi@�B�LP�=����Q����M��� �PC��ou9ݕ��y*�<�`� ��f"��� +�v�%([�9��&���Zn��A�u�� �"j2�)�%��e#r��Ǘ��Z,Y�1�Է4��gp���d�uL�g�	���~�����1�2٦xn�1�==�TY�p��a��O��F��7"���;"��Sbpg�-�JC�fކ�+�G8�@�n�ϴ�L��&�{��$�&<E��K1�4���/f����a���7ۊ���,ЍՐ�P�|��Ʋp�����@z�zs`��y����7nz��N�t�|ƅ0�E��
�n�*���X�H�"{Y5�d��R$!��{O�cW��Zqe�t�̔\���Q�`܂��[�ଽ -��0�x�^���JNlʒ�6\+k��Jhʎsn����9#��a��F4|�*y��)G��;u����ڧ��Хf���>M	�m�>����!�Ͽ���pK�B,{uDĺeQ��M��.���Q������؞7����%-��J
-�FKS���0u���?�;�6��h��Sv���Iɰ�Ek��~�=!*r#ZT�+���+7(���o�G�Qw�>΁۝�%�u2�xr�gȧkߩ��'�#��Y��.,uŜ<�LD�����m�'�|��#N���Q"�������i�F�{���tb+mC)��ڃ4��S,J��
�j��L��Jiܤ2$�s0`��e�a�U�%a�j�rc��+�Oiej��Q������?qC�d5>��R.9�b���  ��>�.%�g���n�$ǒVC����&Jy�1�v`�����o����?�ǟ�
U�R\Vr�q'
Gd+������ơ��|��0J�ަ��	��6�p�������ӫ�2�H^�9������"oXa��HJ��>C�sC�b�*�  +0����7�{j���)���'���2���ul[���f�I�Ǟ���0��1��~v	m��T���z 䋣u�FxX߽y"�,9�ȶ��n�[�V���L��I=;s��O>��7�מ��T���*�SV9��h�8fd�˧Nrfդ���&�>c�o��{4�1�ް�9���0���ǲ&I�3J�gOB.ى���ai����bF�=l*:�4VoI�;�^�����_t�M�Ӡpʑ���ZX��8u�2ߵ�3�%Ob�����Q�|sg�Z7P;�fA8��f�e���&��&�\��0�􀑞X�hj���<�H�5Q��.�vz��pw������|T.q��iyI-Gh/�/�#����Sxq$>�$������KK�P���0�z��&�ф�A�}��~�z����0�)�$M&J�V Ŷ�fw�:�
i"o�u�rm���$���3N�d��Cc��0��<C��@���@�^����|��L�zO���U�J����\��GX�$�9���]��J����-�Mv*�4(�n�p��b�%��G�T�BO����<�\�kՖ^z��9	m)G�P\��4[���]����.H��[�'/��;�l�u_e�mT}w��A���a�=[��&�0GY��ᩣ�b��t"}J��deX2g�����Ǵ8���D)�Q���c2���X��V��_�+A�~���sQ���΋F93�۠�������j�nJ�v��h��G���q\�F��"��|@�(k�ss�m��{8�;�x\v�x�K$۝��SM3ᾀ��I���>���\Wa�5V�R3���w��L�7t��gN����<_]�7椄_H�߻#� ���Ū�~3����"��>JT�*Վ�x��9���	ɭVh��[�p�ġõUZ��^��[�/���r���K��J��a}����d�E�tX8�!w�,�,�0w�i�v�?#h!P(�J�3%s����������	p
���J��oh�%� K�����m�A�4 =�+�O&�s�ΰ�{����!�:��|#�	/Ƅh��>��7��|X�L�)�m�O3z:�G�f1\Pi6����k���޿�޵-;)A4DpR�ݝr��Ă�G<q!$�T��>vf�� ��`y���35/�ش�_΂]9v�bP@���
=��!*�o/ڵ�h�P�uN5R��7Aj�Z'?h(�Rs	-���#��,�a�m��4Bz6�W�����xs����UKK����JdF�$�P�%)� p�څ��@�q��,���V�R܈��o>Ɵ��ec����X�����ʢkX�j��n�� ,�_f��p�w�.�ś@QV䣀�:
d�wjIN�j%l�i#���G�{���'m��|ea�?eQ�Kv�p�Ԏ��5�'���	� T�Zς?EV4`��t[c�L#�k�6�B�}�nX��C��(e�,[*B9rG�q���NW�q�'��*�80ߔ�-G%��k��>b3�P�$��4����̆��4�}f ��Z�q[��=-1����M,GQ:�?TU ��&x����[�U�¬�<�������P"K�x)��,@�Ɍ?��0�>�L
�<�/�����n?lѡ�@C�@A!W�۳�gR�y�q5�`=�G{�\�6���r �/d� ���P�E�U���n��|��'v/P/3C��B~�缮"��z��&��=Y�>��V�ވЄsj�h�<���Bz�n�o�	��h�{�&�~�fc3�/Ƽ����q=M���-�9�#my+�>���`A�-2�}#堊l��v0�d�u]��Po�P��S��r�9��9e����/e�5�Tl-�:�_?�=b����+�EBf��X��)A��o�C��"��yx�wi,l�@8����|�(�_�����{B�����B��P1>}nv�i�l�����% �����6�e�U�* <�j�N�υE����J�1'��Ug8����1�#\X��cpu�l6���Ɯ��R���<NW95�q��>_k�B�������UI=k|��c�F���+��!��.݌A�VǮ�	(��oF��F��'�r�T4a����`�f�;�(�}S�a�d"b����i����QR]�|�� �Q~!{�k+/�*���\�9���D��ut�
>�V�^b<^c|u�����g+�j�C���\�|F���J�0�o-�#u3�����<�̫��'x��6Hԙh-�G}Lǭ*#��ge����<ըLf�����ptS���3����<L���ް���������.��Y�RD�Z�/	`df�����V�q���[{��-��l�U�
�m��H�r���-q����1O�$�Q�yW ���	�n�R?��bF�_�����9&�����L�L���84�i��z��d���8"T�"�n�+7��2�^���EW��b�p����:���V�;��S�~n�մ�FjT&�g�UR��:���,�^�(~:�����PA�����Z�N)ߓy;�G�~k�M�Ò?d�uF�T��N`���x�L��u{w�~`z�HnZ[�&��jӎt�RM�8�b��/��9���f�j �j�	|�F�[���]?�5��!:&��T����h}�˺�B�O)f-�s��	x��o��R��/z��]GG����2�P�|��´��6�ɪu�28��zE��)`��
��6�Z@M�N��h8����b�jOM�ߠ	���1�gl�rq4�M>|1�x��
��PڝEA�"4��js��y
����u�\ZX��O���b~����B��qz6�DV�_������"7�3�͑u��2x��T�ޓ�4`��I�\��g����:�ֈ�1P����K�KU=����1��]H�
�ɬ�6��c�:mH��FZ���b	�}�۝-\2g$����h�H�G��e�<�(P*�w�Hy�� #j?�[Fp���W �BU[:�7o�(�Ĝ& ����V�r��K�QTO�����AG^:"1馦��Ml%����U��"U��dB��X��gv&����倢m%�ǧ_���*y9(�^$m�0�Z��U%/�d*�2����N��zL������Q��}<�D�M�k�1R>d"%A"z�����7��Q���PJ� Z/�A�!�i�M>K�T���)?�m��5M���+�b;�=w���N�+��_�	OI��`��	�3Y�;&��� !�7�J5 m��.T!�@ qufbh6�|p�Lj��zUJU��p��y ��Kd<	Fn���S�7��q����]�+Xx?F(#d h���]h�8�1�x�43E_��R$�G�_�eA���܌<*�ŷ� �pSlg�*�ݔ�R��ڵ`Bx���izy� 2p�	��E@��4�OIk�����^'R������~Q�5�ͻC�.jAT��� Kr�ũK(�k��-�T� y������(�`�
)�4���Q���/���Vk��ݖ�3���v8de����9&�^�;��#X��AIz�Ay�D��٢�Q�R����lQ6��Aܨ�n�7�RM�"}�������=H-T ��ٸ��li%��С�́ț`11�U*Ó��3����ZuM-Y�B��}�oP�>sv��5`�׆��|���A����d�>�琍�0����z�z�Y�1��m���]*�4�_���VyyM�N�ʫ�Jb��P���¼�ƾw3�xzy8�qc�i�#^�>���m|�|aEs}sʙ�s�2	3�(#ma�q�'�{s��J*��i��|Xu�~[�J���s�t�1��E[�%�SVϫ�'�@q��5t��`�6�W\FϮ�h�"��_Yv�.�Ib�7�[$XD�fȵ��&!3����3�g�D��D:̮����ws�qP�|��]���Uֽ-ؒk(�FŅ� �Fk���!WX��f	a�����"
z�5y�mR�r��",�����pj�+"tU(�Α,6�;g�d�-��y�pt�#�H'+<�X	��\��'y�3��o��"|���� ��FkE�h��d��e����p!�KA6��*�`�εs5���{KA�=��V� ��h�����̺ ն=�
zvC� ��Yf�kR�u�RC��Y�6�u{� w/��mtn���31��^"k�p���y.�?��E.�/���O�4�Q�E��&�"�H�^�_L�R�[)Bա����X?Ͷ薡�X,���o�Fj3p4��4��)F�hO� X��S�D��y�P�PC�=N9�aa3�H3B�< �[{�|S����2_��M62� ���<p�y�{�Ĥ�{k�2wJ.`RcebV�wY��P8�f�u���K|,��eၨ��L*��f�#��GQ�?WA��#�1� �5k�*VL�YH �[ `k�z��a��3,@�b�����=�:�_�����dT���eq4Gp 9d�>������Mf�n�=���_;i9��w���o�[���恮j=����C���~��B�9<
S�hS�ȶ���.�����0�#�B��k%��9e��?�晻Vl�m���$�Mʹ��'IavB��b �
쓕:�� h7?,�_� j�Ƶ�1ٛk8�K>�t�g��=fֲTc�
Y�de�����d����pU��)�g)n��P}��J�Ѷ�[X	Ay�p�����l���d�{�_k<%���s�N�X}�}3O�.n�dR] -����n#�Sb��I���⻨��܌�3yK��4��Q=�_��Թb��zĀJ�rH�@	2B&�j`|TԚ���o ��_�'��bR�! �����O��h���ooS nJXH]9���h�=���E�,ԕ�ጧ�A��_aH���
;��"B.f�갗S^{��I��ż�`����t܋5b�^�	���L�a�o�?����͡�,�}� j#cT�D�	�+�;Q�p�V��	��H;"� �pd4Nl��j�xDQ>nK�lܺ���2,���a���;�DEk"
/�ɐ/�>�����:�3.)�~���)t0�ǀ�R��GN��{���v۰M�l[+M���+�k)]��g ��`�cj�8�JF�F�ǝ+!��p�Y.����J�T�=�V[���7͂��_�-�D���N������
D0%��~8�MM>܄#l�O9�k�ɲ�=m[�Mk"bv�|O�r��߮�-������jf�ȸ.][`jnw~���d_Ĕ5�دPw,��s��T�D����Jp�f�����4lE�#��?��L7���Xoa@>��E��>>{y���{�փ��ðWW�����yo����QuAL��hn��DT�&Wq�?��#K��X��P����i�[c.�mo���-����GY?������U����1�&�^�K*���E��2���O��+�!(�@��2p)z�����&����F$��ܹ�ًP@d�5�h��J�����6?�K�R[}����J��pRî�9DQz��q?��:�����������γE(��>�F+��~��͉Lp�s��I��*k���ȼ�/����qʸ�K)Q�`RD���/�36}����-�H��`H�A5�=����p��F