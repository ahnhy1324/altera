// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
PWpobWEgKnRulPsU4AD6ZwuwZbRnP+8/rxmh6o2flfR3hW/flqbEhAg8sG0X/3nZG5GxBk3BQQvQ
w+V9AdvohN7zp3ur4w6240RdkSWxkZQX2azy8pywUesdedqgZZSXcxp5LG+NhnZJ3ub36IT8k7/t
Gu5ZsKFXdwMUSLr1U6WZXYeMK7AdC2gciAn3Ijph+2Tk8ZZ6CDt7HGIxzVXTAAyfXAvFKSfWgJtw
hUfJz9wu3q86sL3lIwDUCG6WFUnAA5gHbUVcgrheaeZgIc30Y8Fcep49q7fWtAGdvtEF7DT8LGLb
c1x5GuMMtK+Dwz4fbt9GJfBcfvcOq5iQC1nezg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
477W2oyAAu/fR7669BCR2E81zmuGhIo9TkQmauclKb47Xl6HH2g2Iu9yDBycd7dLLxInT7l+DXDw
Vunz9iiZneN8/fk9kgj4XAnRdRcvUDXhJyc/qe9ln3YDJCBF/DkrGuWL/wQ1GTpNdknz/4pqPLZG
Rt6WiKiaibjqzTVVcBa4wZDm79/IsvtoOiLljGANMHvPuWFYEGsqmvCwlz7ug8hQf2GjGKdr7hCP
ToTiIELNtWRsSx3OIakYvD2ZsSpmFHyTuG3hPbR1zIy1J44OSaVvbyulXhZL21wiwEjvf1gnRE8q
IbdACQbB0rE27u/XUnN9zj6hb1ShPOEk5b+260TAESrL/iPvwg8ulGmy3FXFmByyAAY0asP9abcf
5B76UOiUyqXc9lXYJ7ps+VgpMBkw/e9KijirLsb79Bixs1ccuMhftjnoufFwJ2AyCBpijUd3TeI7
WKDpmLd2kx6rFBc1z4akUIdalfB/vzeYBctKZsi/J9F82XGUj9RP3hydRVl3yBevSk3iNlQOAKgw
3Nf6nY1s2jYoApE6bR8R/4e6mEDoVste+XtEU8cJoTPgI9r3ESbBPlpVtin5pjG9951MbBzJvr0Z
sJD1006gD+WGYuXScJSdQAG1mE8IQCW568WkGUHzKPOad4SnyHdbxYIF/Rk7XK3wTBDifLPkoUGB
vVeDSwyFtt1XOKgiuY9LdPTSX0rZWkPRINw48rzG8z/98KL6LwfK9LfvQuONhUoMHEtWb6qzmmUc
FVPwHvm68mQl2CiXIuT9TolOKoRk5nwHwDK8tZBIwAVrZeQqpplsRUqP6omPgL3LMSYFCHu8hQ1B
L6xX74HGiRj3fmsLxcAyXVRqpm9q7BazIgxEGNk5+rsEetOrykWTASoOUHMi01N6Xmehj2N4zqa5
uN7lIWad68HwB6wlSjLFzk9FQIaEHZc86KMBt7uNyZlAs66wLXMzFzSWXUHWJ0yLK6kn+ZcwLGd4
2m5bH3lK21XS/e6vMjQF39Y38RBR1ONVHXIE4W82zzEs17pUbh8PDMn/+qi2zJ9rapn3W3mWg80T
qoQolT0oor3M/uO+NXGv08bkOh3Ne8zkRc2KgBk0JIxEoy8G5QB8c48rls+dnUhSja9lz40auSiT
6X7m6faTTuguT+LKSUwi6FjisOUitDr6RzYN2WdPiilejTao854SOO4Hq4ir9aRttu2a6cc9hsUs
mXJ73RxpUXH3Nr58d+8htQhMIvwAvc09XV6epFrOz3lpq/aWu2Wd27BEJpBSv3UTy6Uj8W1cXlLM
b4+hFxDrWiiEMmerJMyknwrnYzkkwmVjATibVaVok2kQIwcufqxF5IbKFHnIxZGmG1vNsUFAM0fn
zgRyaY3mk+WCDNtzi1epI9Mq8FC/Y9Xw2vpVnPRpHPHQkJlwQKwr+he+Tm3lEI0c7mOHfUvy3WmD
WHQg18fdtv8KVNKAqJYMdWPGzwrF2GQ8ier+Z3vWEfEWStpz6+DY2YUyxMq4J8U8LGc8pbMkZwPa
0Zz8cXHaUH9QbGnoMzyIGxxszoG9xSVooAYcQMIvABoxi95BV1hoQDdHzQfKb6TGMIUTOBgD/2fa
LiB27wvyt3yssmrJlfIwBltqaOkQOK9FtRqWEChR25hSsQer3LQyLaR4bUohJKkPGT2nzgwtJ7Sl
+nzOOsfxk9DHzI83dDdNPeGIXlG5WjmOL7apTiIV/ZW2IpSwjaQLpawAUo6xbl7oUoiymrssNvoK
BolGot14s6GODjIR7hjurRjLJ6+i3FKV9fjC0bn9ffq8Y+D/KfDmDIcozdFy/bqbPb7QH8cEjIff
es2Ue9r7YFKslPmAl6o8kgPzZVoNONdr7++es9z8zkoILE9j7niou5zBUrexinWqaHA0QWtUNDnq
Vz3GTYUyjNDfOtqhi2v53jOBHl1ArF7yV0pOmszdnTc5wSsm+OeGrCXet15ws14NZzdJp/umiLWv
Mo6NPg6eubiqIlO2ogCCiuaJ3GkV5BxfiOAvhkIPQkRVE/NCFZGbFRjURkvXHfhujbb/Ks5DhkCC
VKDIx77YzNYbGfBhZeRSeJVs084Lx/xeWJrcGgIxfSvaL3ue8ifONPJEbgACfxmxOtc97d2Wpox6
hNFWlMWt8xLjBsCHSd77bBDlbhnyantT+v1acv2Bk9ZpVDkGb5xSyhEcLSFSTleyCB30F13sZGhZ
hH/NWOic36R2iYZhWjwyrAN0g+e7t5qkPKmeWWklf8df88lqjFVhxjEGbtMxey7ewHFPcAbO+AJE
adhbgnl5tcz3dBpjW2fWVYWCRWnquDG8093Vx8Z8Gg+h96mduwocWp2pbTCdEXwxKZLuRfAiOxkg
TuM+P04H6ITdGSZsQ1iEr7uUi9AGL+p8YrqI2m+sM7vIYjDGgkh/zseElqyyhCwzfNEwGEzmDPhM
1lbfU65FIHfgn+EMdAgFJ0URE/jNLrWyNhgaIS50+8JrWcMZXjUV5whNfKcyWUoM0YVWByMTbFVe
yCuFhXNoKydOU0Sm2jL0Cx07Zebq3LYPJihIZDhXNI2qk/D+F6jLijbWE6L23FuyzMvhuSi+qFHb
4c2Xdmv3Qp1ZMgiQHbybhBCSobqYp3yw9qN96FV8CyQB7nttM+cP7Vle0godh+haqt+ottf2yEMx
cd+rIqa/LA2Z6g/wCNPaV+sWQU3HuigNpR2EQTzZ6kx9+Fx9esyrxWRsMSSzuNSUDWn+c/RzcbkD
TFbhjQpOpd1i8TIjUYX2p+C+Wy3uGCDDf5Lk9fd4juUo/JhvpDUnSOSaZyMxeU9SwGHmgpyxVen3
QxRaZmd8mTMJ18yzWJ1t/ULm4bVJ/X/nBiHqm+61ePrfvpgOj1aFCmFbRbEL4fsFT09OQ5bsItf0
r0vzaa4X4WpDY7S/BJFmkMus8KF0AcX7WYM4rg7JsSKgzgubkSsj0edOSKO7zEk6X7FmRqq6vItV
aULEqK26u7HGhq/ChmhjewV3rbleFmp5armY6bAmvQa5TJc9AsXgZ47w5D51j1xDHAyLoPoKRrEs
/ZMycXsaDnYy6y/xqSGH4+jdBkhOCeT4eabYSmpmKpf0nI0ycujYr6Gf4X2Gtj6hvVBi+5/MQ/xu
6m0z5gVfD2UQw9uicVDVcZhZoLsO5Wg4tRlIQkfhZ7pcCBwD78goZkDJTx/j3QKAIN4eyNtRdieM
f8z4avlrkpVqR3XlmfQUO6JQuJFmIr9yoHUgPQZiReSyVDEsj3DMk3uLbX2L1B5XWDQXvoGz9+hf
N5XTI7mkGWqCBi1dyxM2dtODHohETd468x6Z/Hn/J40mpEMg7AVzhsLW9zUIYYnRZsT/D9HIzCc8
mbjHiHVGC7ebmSVFo9APUohstDaH4KWuVKruBNDt0st56s8Hfw6W6LqKUbqd1eTV384O9TJ3YUfi
vVA/iXxWe5V1nIOLNtTtCT8xp4aKtCJIlf3laltbTp2TqvBy63/7s0m59civJ1jGIaXmgcR4jJZH
bK4dPLPCDI/cxsovmjgZ9kKXWrpLnzAlMwjd8g2AuPTqbQREvIcONyhWxQpq1l/9TmCCIvRV1GsT
N3u9GGBkb6ZhRusr7OFy8INd0mRg8/EXJnknv3tlsKJmmQH6nu+rkoTSjyKV7B9TxTHmbR5SUsuE
rFX4NpPRLsFtGXvZY0asPRFwrEbPyzNxqIFAFF8+v+pIAiiTXUkWDy0SYwgmoENKFI1Wa7NE0yu6
Tl9mKhDwodIJn6mydbWCJNOq8gAw8yyYOXMeNhmKycs8p55orX8MKamx5CNMqDu/K+giMT8G+cc2
cQw9atnmMNB+4vZDINcDCbTxnlI74098nrnohaXnCSKAbzcPwixRpckxMBdRexiZ7FxMHbjcz78h
3ySOBuucXOVJj+nh5tj8FtaQQLUjxBYZoUTtBE3/HSxc7WxcEVeDj94UbVeCoIY4jhrdvGbd5GZc
gjHLp5hWfJZQjUKtiCXI+uiUEQnz4Gkiyoav6XRN4s0Yo/lHw20huWcdIyhrSxu1FtR2mMIhdnlR
GAQ9JEESl4bDmKndSdjjo45w8/oiVjH7786u3BfYe7qQaVvRxeUSQ7Dkl4n/5DlVPcbGupqruk3i
mw8/1XBRLd0A3rt4qjUyv5zp+SLLdxyAMq3sZiV+qpkw5jjPnINdInqzXkKKeM1gOp60kaefYUgV
/UG7IIBj3MvytWvFHeRPzlF5qpL5Xu7VpYu2uUW6E/5C8T0OBYBOFECXXfyZEUhI2UZGdirkmX61
9uH2KRl+LRBSRsBbkbYjcdd9bdt+8QS5LbdpS0bNTLBFNpOh7imYOaBDW2xs8zuGFuQiU0PsWfpl
gXBlVn5Mt4K4Lij1iuxQauPMbE2Ttn/0tYhFYqdtD5Vd981BfkbGoP5AImgxuxA36IHIG3jorjuc
w1M4NcJR8PCUqVMPECwy+bXtTGGBaO/mwJ/nXHo5RIFt1qFHRGmPdBSCNRzwPwyqszZJ8pLur5Jh
yTMaVIF3tOWuG+E8J7ZSQ3YqOf5FwkfmYxf2reh1zKjCQ58wRtACalFfmOAJME+d5E40liWCGMb7
8vFFsayJ6DeetzOQSsfG+z62UPvTdA5JFjn+9HW/582dEWI7xRzQkgk8bm/V0ze66LWSA99YVBeu
1RPod6YCDzGB68ZDlA353BfsVzgENbFDv8WQEfWhRCL2OeaoR9kTSV+yFU+w2GmNSzlsfTQgSWDB
ZrLMZldKLhIoXkdC4hvo1wrXRrz2KgPFZqDk/fE5bt4OmOmRgwG/SE2SD+eQFBBxdy9NzTcwB3PB
XPdU0Qr4k0KnjLhXDgy0LKT8jZ2cbJ8of2hOSISXRqBSixK+eYuroCoWoFm1UHUXCIN8AAGuD5/C
FuiUDoYqY0NPQTY6nzZz9sGRm8Ntz7kz0xWJaRAvLwVQpolxmtMgJJC1S/lVELt3vNXBasO8cDi+
AUc/x7mgGwG1Sv0ITCqNS4oHoumlu+pV7Wz5C4jfYVuoOHzdFvmZHF1wm99cpDi0Mibkez7BuBbk
ZQdahtD7nbOk3a3/z0EmTQ24fgmDHAV+1LtTEC1zQypj5KukLjKpH7QWrZSlZ0V34OgSLOof/7fv
g85Y5yLPdiQKzukHDWLSgFaWqIQop4jEO73YWI9Y/Nh7lF0XSCd3jJs4JrAR4nBTtC5i/yVA9OSt
0TtsoFs3r77mK+2pzowR2ilHltZyDaLICltQRKZ13M2whEueSXx7Edwu3EKo3G0UnGSlzTZX+xmV
btQne1Ard1mobZYtQKjz641NGLnfknwO+KhyEoAGW4dgoQadzO11j59yLY9Sue6CuKr1QPYD2sHD
i0yKLr00p10HX8iarSxl+94bCZjUfRI45aXLSdzGWgg1B0AkbPFpPNIcUIhLi83JAWzvBofTYWPG
8YaJZaJN5E4UGzaSdgdWwKxjDfgmIhuWN1lafRDKp/sMOdvBw9Qa8JUj7d974k3emMtsQiLJZbxx
jLpWmC4VLHcsul3XYW+MALugtgA7PDxDNNedot/uD7Jl9wKDqZrZboSdZwNkm8slar1ANRtKvL3Q
M5I231Ysc+7G+6QBZwhj/mbBiWIWa24eu/lz3Hlo/OXr2NpDYUws6Tw+M6EAleWpj+mQwF7XwbFF
SleAm+W40KDWYdndWobOZX+xdPPIQOBeIW04mJJCTPwzkN/XvN3R7fBdml1iIfPAFgvdLIIEODHV
uqps1Pm6cabE4zIEiOorLJmoyDu3vkSDCPfgYMEzPWhloPRaTFOX6Ac4m7lbAWagMyPfz1ZJwin1
hWcyU3nNj60GOkAJOgXg0n5Smj8rDgAR8jqgQaeJ6hhZJC/aJ5lPKlectXjOc0OPyDEikSds4/KC
q8qIjUws9mQyWlFP6ZYM3QoNKQaFghs4jc/94DxZ07gJtJ9wKuqm9FqSmqeU5VV5s0ukk14OHWhW
fowz5W+5/zlVu5tUDFjS8E977ITPx99oH6l4yilfuSdwx2keIz79Vv3POD6Axok2cpVVVwBxavDX
IHF811YOxOBvHNm7ySqYJ8zLLseRvB1argYHwZ+E8mE4eMvz+jbLHHaUcoE3urTUypD1zk2yM1cb
mbPSviBJC8xoSdrEqNeHXmwuRc6lpGH/t5C1E4kE06AR9Siy69R2Qd7zbW4FtFtd2FRDYTSeSCJa
F7HSaShZuyAx8SpRhS7FX0HWzHWDd7l88Sr+zZfYNeUtEDO7fu6ZUSMK7psCti26EkeTrIcS6FH9
hsHAgxAeTMsXX+TueDCrsnnywzZrXDLfkzd7PeNoY1E5hnY5c/a4+CqJDS+MXRmIafD5mSNvLqxP
tKwcI4vBhSjb7tSbuRn3PZ9knRHDmvL/WLqqDW87ewcYKWzHscNWTESpJaJrVJFs3ddgLe8WVz3k
gO3kPV9nqHAYC67zeCBG8N4RBHjLQHGdA5lR6bFvFftCEkPficqE0co2gISWvJCKpFonUzR1YRxF
JqKtVJcyucSgohn0Jmg+MGFDd2saA0fJmAMudaAKae9JFRd6VCNkOJUfRQYsuX+XtPW0+FlXNYu/
JAd49G3zenisy3wYrssrLLvjrFkc+t46MOwPaZT27VM2zfT6ZQSWyaJWgjB7Vmt9vSrqVcDbur46
7aHrIqL5BNVn6EDj/Apo/lpySJHQHf4LyVgnG4Ich+Mi0ZKnZbZIf7XWC+5remEGztZnb/yiexL9
BCklf/gv/EKC4qmZApKxHOQPeqi27rQSZtbYjj71qG73JDjmXz7mXnrzEXtWVqqw2jNPxgl1O33P
4djkcS/PRA/B1vRjeqAvJHrQFa1xqYeezW//M8w8b7+yHgIlCBjezsMdIZpwJxbu9wqRvnCGqmYs
yW++9Db4pdfTy61XzYyz4xhOi0KTFJAtsqm3MJmnlSOtSCiQxnfPnQEeSsUWIfDlTkQD4UHQfyEF
s9euWHC9CpNiBfWzIMT6s7ybr8X7A6dUy/3YJs2YRbeaqtUDJLqiKwfAGBJMqwjFYw0SAT+lfwS+
CqFktRBCD6SFhJEzATZKJU0SxUWxBEHivnWOCXDrX/4/M7uQcqOc3hgHvMQ5W2rjoc6Y/bDmp6BW
atcehweYiNDJTBr3GelaEjsEqgbTXgm7qjMeMVyaGqIeBXPoGLRFW4gv34sYL6Rtc1ckdmyc4FC8
IyUD9k6gIScbx6SxAxrNSv4T4pC4/HatJH/eyN3tgsD+6tIt6CArGdHnE/sFWxT4/0CcYl1NJj5D
lKKFmy8LrD+97dNfU7q5va6f4LML5yb0h4FfMuAFwNzHT9OU4PfhbucsGkbjsqEuwSHqAZ1yH2Tn
vwoSrR7AOkuNzUsw9YVNum1kzrrPZxQF2+1Kpy4ogcNM2zYsvHrMsF548BYDMk6BRYFsZroAwahQ
rzW079YuM1dlcb8+4DqOyyGc9SMw1nxKrW0tu/CckZMaK2gxWCwNzMre3ue6PrWKGa1WdQxGkaRv
ygkHC8IKqBXo3ygG9PyjTrGv432TCJDggUGRR0xq160xBD65UyVOM2OwAe0lTjxfHZpNuA4pZR3E
YEcVz3aDBrMzklSgeIr3a41L0Z3F2QqdV9xfJz34MDT/L8UqQXtnnKdCroMd0Z1JdVpR0cU+t0wJ
0lg29s/2By7S+Km4b0dQxHTDytx12ut6BzY35AvpUH6Y0zrLVbF95dM2SIwvjwX5/S2Bg0669UJ1
ZePel0XtbZYlyJatFCw7/NQ7zj6J2pOMKhNbCy+aHHMyUB7eP0Udq/Z41/GhH+P0q9BI5/cZf3cQ
aqmTVbsWwZ3BANv63A39be6Yi8/N2OHUulU2jk3MlgQMs10OZmUSItoC5f5gUlN+JKWWnYNroqeQ
Wza7uJYGpuEpOj+2f4dclAb80nkfrhDvzNgOm3aQh7v6dSutErie/XMRPOUdCLUh9vT1eNPOsZ7P
gX9SGsy5STKfa20n76q6J4nAU5CSFLqG0NeCyAbN1Ai+0IDGC8B/TiBQMestf3/HnjJceCrg0Zi/
5rZHk8DNHua8oQdKV1X0HjnpsjzKETFRQxNVJIYeJZu4l7ouaKADxtIdGi7c9H+gZlUIBNsX9Nqj
410SwfwkW2CjRpUIP3xYiSkt0NFSWOAHy13ZQis8O5F2Nlyvgjp6mJPybZt/6z0TGB+tm3ezpRoD
wcSYYc2bWxgCBjU849DXwaLoELz1bJxHqLfz7UxGB1q8zW+Nz1uvmwn1OjoxvYlA69KoFwqq27g5
WGJdWoIMES8UTotBqV34d6NM1mv9j8L37nFalZB9FP8XXXzOijenLdvVhXJZOhDErJCW+kVLsQBy
ZESuwT85SqBEAX5+jXpkVKak/yzHwTVCJG+fpPzpGYGWkI7qQJjkZpbxjmr9t02/EFYOMvYKQqDa
IGhxcqpggriS1A0v43p9plbyW8Sn8IvxINrdw1SUmrGPkPhHfiGl1mlY5ZynhVrfysinD8IEnPWJ
meIOUiFxOhWW140z75QIEvrSILyM8x5eV/PpY/Wc8aOnRzcAGrPOXzAVN5PEcqf3Xn7Rz3yLKrgH
6OldZ9ckZTQpMZNhhUqSyw96PUCe3NACPtu6rBH0CnXydrZkMIHP7FommQ6hByHGCvQOf1RtQW8C
SooT5f4UbzQAAmR1lqq9ui0Io5nrxoqZwFUSQDQaF4NlqWBGNAM+KqQmrPEtHLGTTOOO1lpbXVOK
0FfPCpRJJBSk3821Ynftqmj9JVU0bon77VkhYmAMSxUOp20jn3DtximxtT+hQFqQwZZlP8AgZjP+
SWSdQKSBSOwEg0ON2Y7R3PE2RIbAD1UbjoryhFIS02a6VtXfcd4tV1rtlLU7gqIYaLCyOiG0FYGo
UGnPzmb7fIPYI81sfaJzEtRkRRfwyP5d2IubGIy9W4YE3BRWpW9yt/vOSvUGCx6v/HJVQMAY7LyB
SDwk37suAzW7aJRIQMdW8YKk5oQY7gOgDhnLqy/Ci3JFKvuWKf52Ni3uSJM9TmndcD/eQORB1dAz
cmp7SWBXviZwL+mc/SbHoRfRfZa/Ng34sSyEAPmeOIeScW0MQBOgDZQTsU5G7gAsu0tlxHpxxzLO
G+1dUKAvOPVuNeJ+LRmdl+v/+ZZ+9UVrWvdmDthnmUiJV07R1PC7ly/GP1+1CHVCFN840zLdbgsV
KI/WMQGf+sJKcmv3pEIYH4o1zDFQM6uYnLKzxw0kdsRtp6SpfvEHuwmiwf7thjL9j3cdwKvLnLIn
zn8uOZlLROkVPIEhYRFeeRWrPynLcYlhPLmD+z/cOUY24kokBH7BU9S8yM3rk7Oe9HXhjeujjRtp
0pxKoubwyKpGVZftyvoCxj6rZBdOnY6t6rmSPSLxZFmUYjkf6HogZYET5EqnRMWHT7ge/RUksQA2
aTeQaKrRZl9yAdtJeZrbMhRswraOWxHhiEx4VLzuyJODo/I7cGrPdfxNSjgJOlsuXiYrIx7bvC1N
+cW6wSugl64+SCPpicCBGmYk9gHyA72UTNHhAe06lDmjAHkGjUqiGMrSa6zrlgcnqeHuGRcHUoy1
Na4bj/A3Jy11CCtKVJe+JIdYr8QPZYt4KG/ob4eNiWeax+aGqXHbDfP0Ix4QOrjzjHcl0WekUWjB
ML7OzQRNb+TMk78yrfyUrEO6aA8OVcebw7GpsUInop5rC+8JBsqObLUfKK5YzyNdzfFP0Fqg1+Cr
kePWcpIM6k1C8V254IJDFPtFUyry5ypbBLQg0dtzeIi0YuhOxAd859JBAe1uDrIS9bldIgiD5B58
r2R4sBMBuAnaWUYs4IZ9BLUZuL0TxYATsyIrFYk+d/nVcFtBoc0pD1mGXg3hv5rU6ofq+wIm/pe9
kDff+12OZFw9youKhNQ/wD8oc1T9lmcawhRLUInb+0+F65S/D1/c1WxPTfjkqTBogMliX/K7sPXC
mXi8MeIgpdcVAnAMPeT25BOY2Mbr/L6sISWrTuB1SaKnau3Z51EZGt5WIg26rAXPgxr+aodfK6sp
upsaFsT8XKd0QpzeQPQ/Rm/vbgnAxuRPmgcsPEXb0NxRLfBwNtjsq3PkLGbp6/klOTgXalVa7kIE
v4zVrMDM58FaIyqC2ZfYZp19U3EeUnj8IgDCwa5387/E3Z1IDxlRj+w0ZdAQ/cgCQX6mr3wa+MYO
Yie9XPQ4ro3CV2GkM1SHQy4y50njBtFgmYCIbhsbbNyISg3mDL9IP9ijdYDshSiyUmggf0s2ekX4
+SuWkTnQPlxfVEvlHyK9Pa1EjS1ITc3EPlwZV4L1FzB7sYMHIHfMMb/GKMoPHiJ/yx+/mp3bICVi
zDae/hTgJjvrrHbfDFL+MFipm+sZ/dpfpnlFLOQW4s5IEJH9WwQiJffx5BBU/YLspREAWhpU21+S
rAtUDX/OKFK3bEM5FDokKZ4CdYCUeo9G3/e2QuUQ+GlKyG+QJZRAmfAvsQbQKNSZq6XhGhBquEKc
mdQhU5CBLOv46m9gEvmfqxQAUqROx3CZfWSOD8hf6QdTX8HPwUW6McY8GhIyZrpVvwAHy5dxsDPj
oDzrpUG2wKPu2QcV26RslVOL+s6SRVbo7/zbRP/Bbk44JpBKq7Wrc/mAX+L0TqJenLRb0htWAKvT
O8icHPfp1SAMLaqfmHRoFmkkI+kl+agkmd12bU8pu9GHo5Jg30UCpRusXzXfxNWRthjDyuMLnhzb
GSx8GNFpqZPnTGA9BfywdpgZnRlqKKe7boXmPoqPfZ5Udvix2Gu70lJpnt9uY/MSAlMpB2If857w
HtVi3Ncqc5FX9KlgqCM+H9U2JQRBn+gHNN/g30eggnb8P4xvnArbG88w/WQfVt4v9VYefn3mJMsj
wTWOZRUDiMvmDEosUYh014mCrLNf7y4uAsl7IGi/rPJzDCbvQulqeBX3jnKFFL3JPb9MnSGmXt6P
IDF9s++BRRO6YwHHWTPTHHeNSLzSJCyqfvK37OV/xBWNC5J5tsnec/JyMEu3QO87UOnpnXuGsptp
rzPBzq3z1/b0T/q2zIVmZV1SnOLEllEQQbBV5IQapxJeGHkpMAgOMVOnvCBaGM5wNfrPDb2Xos+A
QGXnTpI/TyAyGdRheWbVydqND8s5j9kzuuwoj+loml3gJXjXfMzS58Hoy+cdsvFNQ1uNXuJJ1w==
`pragma protect end_protected
