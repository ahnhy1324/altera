// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
s5NMfYSfBbpHbOkVvV5K8lktbr/RTfG+HHccvEEhTJoHzT8VMAZIrESy7OxtCNqvztf4P75GkR9s
H/P2PLOztp82U+BXyMd+Qv4AYgubklQcLm3MaSTudWUKa6ekckhgqNdedH9kO03woVy8l5Y8fSX6
t/zcOJmArWKbJFYg8tDYVkQN+88zOBlsfOd5/nkKtImug7Iadr5Z6Hcc77sBMCkxmbGYuHDnKQG+
6jp+Ddzar/jXd+Nh15fjfb00gxvYLwlDm2is6VPs71WP0SML6eMEO08xRLiSlccHljNE7xpAPjUv
Sd1VKTVYLe7x9/Y5vOwy4b8UGW6tLHrVJu7D4Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
zEcDPnnRcTp8QIdbXqCkGPGiuAm+rvD4PGma1XMnPNg1OlcJm6fRxtTyw20Uhb7ICwXlhhNE3kWC
cebtWFL7nINk+K7LsA5cdbGVU//1OTFrNRfh4uN1XecQFpFW7syAwoRDk0e//uEgO3tZU/XrigNh
HCs/E+zVwjYEosaPbl9kH3BHcT2ci4hQHdObg+k8ZXZJPWoK0UfV110VjrXNjFCHiTwDv32zd5WO
9398nV1xE2sOJ68kZcicsGJZx9DgNPpq1KtCdLQ1PeLUFewQQW4o0IsUExI8RfGe1xNPHwi0nsq5
UcCK3u+vq/gRR2/G59KUeHT7bIC2JA69rcdoRSYUVnYmMuCrk9Kpg0iYRHpFmKTwi9gFuvOya3O6
JHPNzMF5LFYzISO6sQyqg+U0f7cAQ61hzZuHs5ynCjBd+k0IFeFRlJdez7zeyg+evvi2It4SBeq3
8GuVOWvQKdytCAyF6LIH4GrDRcKgLyGSqS/9vBZzzqQi3xRCpGrNTgxGgh/kCbfYZi5OS1wByKkK
KkhYx+0FNbWW6BTKO9g+BAWTxxvEuxu+a/UWhHTZikPntW/HmlyBUTioqM2W4Cok7cbnXTQCyVzH
mRizMTaPEbS/2O/L6jPKnDDErt1i3xLWl7Qtdj7UJNWMGWgc0bWAhzRphU2EjLCj88cGoRfvWDzY
w4o9wK3plDacmnULTwHDp8EKfVk9hXQWlQQybTp3MfqdTN74HzBwYjjm6r1S5MCTugYV0iou0ieX
Q5iYaVSBE/4/vYFMuFSkVata23kZRFgYXHRZWDOeTKsyfohqP2xbS9ZSN8y6H1qQdtvHFhmmJm06
OPOfMujUQiAiE2vB75kaPP25raj5k1h6+DoqHYVAZ9VePBCR0RUOhj2MWFALC44crj5/4i8KhDw6
C9v6u/X05pqoI6a1KIue/9r4INE3K1hk1dhHnN8Jf2ivtnOcyYDga/iS7e2MM+eFLXp+0W3x7YEY
alwj2GhmO/TgomMxuiAEMjKSN/dIwN47h9QRi3iwx9b7lS1rEodjeK0p3j/+Hxi7g8RGPbMX8ZWw
Tk8Bje3nxwgCf4cjGVpngbshZkCvPPRLFWrsBW0zaq8Dr2CmSt1bYr1pOLH+25nF0MsuFbHbNqV2
fCtnCAB5YO4GWCdpcc2WFJShq5UPZgeTkr8VfQfDFdRvLaUBA57ttCv/5J5tQ+AaDVuFpp+Zunma
s+/w9aunfXY4npI5cY27BsrwBwqGnZd8MXS+c6fEI9P5DRAeVY1Ey/Cr5NPlvQwjrM8JRSUly9tH
yKoghDosaE5fG0CKeZFxS85E6Hp3S2cP+vJLp/Uhg/izI3bnhekND3wVGL2XNxvTPlicII0GNSOk
EKbIP3MxrWy8jSn7nNdmWDD28Z03kyN9ZOsUIU2piyTNWAw8lPC2PtYkOwOlofcw2Izxb9kIIqWh
N689PZFmhTkpk6dBAzzNAQxcORJJawUgofp2iCINXaREQTkfU4zETeKMgdJQuzoQwCZndDCeKdMt
ptpkOmjAyKT5Z/1Day3GAydI65CmFswAQCSM+mVrqJ4AF8xQKOEG6SDXQYJfyZB4/OFOeUjxG1bv
7MkIHEXXofsBglxkjF9L0ZrPBVtM+vStxAmWm03IlgZHTYiqCJS4kYRgRePhybUM/0ayWC16hq9W
GuFEfGYSU1K3kcFYvPe1Fz3gwRiWh79H8NIuUAfr1hvx+TtpcUm9gbnPMLiM4lHET8/lESG2znni
yBl307MdxbiMwVDHN8JeHBLlPmEMPcHlpGfQC11TWAxrQSE7d2mRClRGSB0ssvsVqEswTTD8VsZA
qV6x0iFt0SKMurxpLHgW6gjsVdj8ZXIBID1lpjQYpbmYrynK8qRavARInVALO8D0hCMEY2ytPWmG
aBIX6gjAb4ajjon2AoPKadMcU87eHfQ9Vi/1Ejn/bIXxled0dMKJbKqRIUSbVsex25QRrkGWSFcj
unAQtu1Bb3XG56AZg/5mjMO1O4C+wBq/pOzUdptvg9eUyExE8c7tubOdnqWvquLnquqfjTYIDc/g
aVViLszCLtB0DEelTv8zDf+sz6xONvoWx8KBm4NECPvZmtTOZ7tOWG/KfCVFBVLj+rlSWRAXlhJ8
iibHnGcZnHtOpDawIqEEmG6UxhXnh+I/VCBRkBaS4ZJauyrbfeYPtjn9+tPiZxRLVnx5N6uSvbdq
eIbtAA4TlvsdRQ97MewEDNGbbmZkneQQt/xNvz4AuPMrjAq1AbhW1OjRgLa3o5fGagNtSaxLFBJx
OAfJCYOdEX+ZutTN5ym/5vgl/20cOAU6DDkKRr09vER7OcXb8zwsbbydgD1RC8sgEYXd+LOsbV2M
txFnsCHW68Z9D63HbYvvogmyIsxCGnY/Lx2W7E202ltgydZdHrZaIgjSzlMjgX8M65t9m5bzZvqM
VpmutpzmUdGUWe87QR2t69pZvJyYmAYCNuxFqevy8VDqEsQ8RAUP4ms7DyTHnhXJJLwcKhGSP1SU
gkBMF1nODeTkT/yWcCv5fnb85OQpf8ekoiNqjY/7p7K8TY8+F5gLLBEctuE1ryYKL3EiTo8s8nDh
OU7ea8dsSeFsKMNoq5+hH+Z7SBquXbpIjnIs6Xr/AZkWwvJ1LPbu1mrD2+PPreCSJW3z+XtazlcN
o45TNlvB9bH3V/MKz0qlkqUbhMKWSyHNmCOHo6kIXG+rDqMUoD2juq4LyIpOeDHmJFYIPvF625pd
HsU45g2lfZzGK9cyL+JfFeYjGtVFlx5QFaKA1CjaAoD6o0i7wT8rABrNUCZclnqFVM630gYrqmUZ
dNIesNTdEXRsH5yBR7J5LknXCLqdhbkak2XI8abkK70hnbRYRwxCAfJDJmNz/04xlfoLfMGByDJN
yOFGCeT3CbWt0spiITVZNZPzjBEFwqrIKDHV2beQ9eiB7YD/jrAIpK5/czu0G3VEAUbFHQMKGdZj
Sm9/dye+w9dhK60xrzcxL/ZgCjOPsSiUzkDKLTJbRCztVvc8tT3l1W95NmajybWU0MwsdHfFF9zz
RwnVAweXNWHU1NYgMOSrV13cvdiJ9a+sGkN4/yKalJboKuf5noaxOqy8rd0IRR0VhMKnbVNw0hVn
SsW1873ifgS1kKLfcMzfweiSK7Gqn9M2roSZflWG5VAuUqrIyR/ka9iEF/75UZ6dQnSBiZjTHOTA
mrAVtBeoIFwLOtdIMQWaYN+OVvHt5oGTsrNQ5KrNgD77omX2POYBFqbkFHTInf+C5g/itBPUbCsa
TnYwjVzkAzVDjzT0uhw4P0buCjLwtRC+R5WBmI01oF0pa74xWKQ2NkLlyJyNB4gtpiBCevzRVKsR
e7DPFVvhy3gMly12PINZoaHY7yZ8fvMl5Y43UCryhcUDArq+E6yVBgRHNQXwGoUGtm82fm4CsJ0F
Pz7Gc3uS5WMMn/mRDyTAAyyzZ3XZpWvDqn7t8ANTIzN1yR81+pZYrzq7/cXxLlq1/SxiMyERXXT6
YJsTJK5UAPx+lB58fSAHLjwRyReWKQ5CMm4Kq3M6aH5VVmA+LDD8OFm37A/7nXmvevSn1W5c52W3
wiaprBMJBKDMbHjhUzxRtzqqq5Z/VO9xK5u415LB6N3Mf7Q/mivseQ6rrwsYd4tK9LqgrGwzwvJT
MqJaRBG5GdPeHeltOcUtBY/6sKQgWGFPk6ILLw8n/XfHQ0KrvfJgBppv/tydOP9TTTAnhabhGRi2
eYboY88n6JEISZ3EdrD96AcrAPv0p7a2T+0Q33oyw7DwlLQ8qNhcFhOZRGmcq+OSIWsvZ/PEElep
O/9fZOr/kL6Sj9U4KhM4jM7uRaoRfig2FkIw4KUr6Cug6GTyZx0wnAsTKpY4BmPELqQL52E6YaDG
l0O7mvEEvWl/wTEOCNApDUBwQjPMt0uV9weVm/Bp71MvHx4AQ3sg4mcpXIljp4XEiGbFp0xXIIsy
AJELy3ibfVk0qqmu0ZUEOHE8Wec1vVYlmun3UhNzu23CUXSBDXfhAmypZR3/Azn4X9vZnQo5jvDY
TACsAPIKDzdgOIQzncJ96J3R3I5Lt6wLAFlvfBXMEo+pMydehw9fEHzBwldWuC+6QyiX8qGgm5fr
swJ67gdSmLBp51HcXymAJqMGpQ1IR51mr1/z/94vgsOAWLIj6/hZYQbbtHxkMhIt2k0Udr6U0H0G
Y4geJBVy3b0Mo9AbwzH2B1iWVDPO3cpXaRPbr9OhhzdQkEVpVg+97U+rdrQ2D5u79TK6kREJKsVC
8MYV5FolZbzBDmf2G/SPuyTQDREGcPsh3/6r4CdbufouA1j6rVzW1pI6rG58Zv377VKQRHr6p2ja
vVo7BkHZ5L9EZVAQ40KcxEoirumTpTdTL7N30H5TJzV9tRV70SitWs5PSjduRWP8btq0xibITYmd
cOcaBmVCcHYCQKP+p92g48N3aSlM/Q7fc6fbeUH8h08QCynqmXeQpgs117FrvbKLMNZMvdj5frRb
C1wxPolCyuGB5PHUXgOzh1sR1iTsek/Jr56IhD2GUxoWOXdHtmZt4tQUNn5cync/Ik4JSrLg0p+K
79MYxe+O1NfGBYPlXdqP9hYAPpXKSfMVMpKkybbRKeyA/Pjpa14wjmfBqJBMwk7IS2CkuWpZYteq
iIKrx3EQb1V2USMUuaUyb5iROybqx0LHWHCav63wZjNjzXelYF9t4W6C2mZKBmhL/bK8kO0y8c3b
8IgfcNC/PPHtxCosziO8ttY+7UuRhQ693FWdGpSg1kCDD27/KuV8fJ8LLSM0yPj5ZsE1XgJdatBC
++onC4I7sVY4lOQE4MPtB8TIQ5STPYnGpuJIgorpO1u6/yXuF6FZsfdCOmDUdkB9YtLqJOX5HXn3
e/XabDOujNh5iVUz1S2pkjD4VgywgY4+RY/tC8SBubatiF5ytLUpoK+OI8X5wmM9qNmhHfwiIGMF
f1a7vV4QqKRrRKpzE2AFoVtySDTQ3BYFMGS3nthNfSrx3u3jlMqfkJzshBMhnGXbzRHH+rKmqivv
AhnCtjU8CujO3l8jwzgY/emQfeSYOi0wlB116zZoGWggVd49Qj2HhcJKFf+n6tqwHk4p4Gt0TMXO
xZphhzDnmgknVbYJ+/cwOIFEfTJ9ZHflNE9xO9/1cU4RYQl7Laab3It4WEvNqMCB2QmrXRupxIf1
vrO8JFxxmXeM7tnT4q2kKKh2iMTqx2MMvts0mJHJDa75rDStinZtkyVnKodIlU+HEbfEEehgkwXL
QllDbwY0rytx+ZJo0SBCR1T39R2VZoqTaVQNIXNT5P2tht6ZOt2mSWwunL3ZL9Hy2AnkuROYeEaj
zHqnGx9lNhxgJwx61m/RWXwx0uZ8XuQ0lDq4LRWpp7dHXcltjW6OwMweQuewVTyocL7Bm/+Ft9Bh
kQ0qBo+trMOyk0DVi4er2EPA+JKVSrrDMxH36PSKdfIKdgd4YDDsgHkkY/InORv5Nx/eRuM3jYMC
+vA8CRWnDkqq7a6y/K4wLavn6SfIwtS+cl6b4/EbYpUvzyogy4bB/pD7coP3vjinwYEn+xWLNIZT
2EE5WwNfJzpC4zsTGX43CLnebSnrSqhqjvocj7iq/7PQNMYNvEHw6P5wutaUotBI42LSCgzY2o+s
xf8hP3pvjXaOadJOT4tnjPI74xkx+VUs8VN/0XvDAFoYwfxh2cT9MZBDmauR5f6wEOhsaaA+psj+
dqyWl79CnMhHtrW7BPlH2ate/wydorvoMPa3LTndKpQCpBm95KO0sSX6JmEqaLnohPpF5F7qb/y9
eowII06oOfj8DFCqAUWigBUirzfFC4LgTkXkgWI6ZICNNaeM6ySaIami/RfIv19t9ct2APTctIA1
zerOx9aybeIYU/y4BnUptmNhrGEaEXd3vWC7wF08KAUUSuKcZouVhdc5DXGBhBgAEeJlsOX2BVGF
3EMXKaYgIqmuXzy5BFSh+eVPb+OT1nTxSBAqoU0SMpHSITH8W3qnAE07eTizQxqT6P7T9oEybi3L
qhtpR8ucp3ZlTKNTJHj6DKnNeRciRC7qeNU29omDqSVmYN0f5/1qcvH2GRnxEYXBDZZueXIjpvhs
hFxmji9DALJuabksaJqEkxSfrcF7Z/t1xkuaugbtQI0mqBmjSKKNQHIx+5bQPtuio6izvn4rJrZj
h+WtxOjMZKwEbr6Hl0H/lIW8LKqReOwoUgc8lCj0TRZPqGUqop4OC0amwXsEqnjaXCyBcozr0mGk
5KZRdQdHyW1rMEGZapltdj4jR0BHHhQyXTxDshdQGN6V/9vSi7e8fHUJN23bF0EdYxxh0xtsVLx1
mAjtgN0uCnnO4jewc6aXuoOmxRVsztQTUqqctNm9GIXJTSYHPiZVMdYWd61SncB9fn73dQOjEigq
VSyCRr4EG5HjbxOBCqQZySsSUeldr4CPOSI3ZaVPHD4GlWntXngC35GyzQSdfo3OroSxwOr4pONK
KGlQAZ12WAOoLaARSzCtEWRoZE/RMiztB3J3wHsOkFJwBuAauZmMP3u/Yd+pm0drIndkCfRHu4gn
pKNwwwysxIG3sT+TMSvrhs2rFH32H/psDGPy1uMsSRU7oIn38CcsL1i+HYHtcQtKcmsxGHAd5iEs
Az/pZxNhTM4sy1EmKZr+t2wSaTDHuLGUiRICpmHFLA1pO4i1i2dUKmJpPqlK3D8TKvLIJhvLK9Zt
lphQDsZtEtMMPaixKdr3Rx+WLDoXEEQyjaXMedom5bldYDivfnNM+fmsC/iQ0MXnGTORZxB/sFAy
zSwzqUOrzgQIXr8EI6kpOflUqux5IxDdxt0+PBzzJ5iSmOTid97A1gophBsZGIem0rGkv/qPaYlb
27isbU3/DzpjVEwxIaofFcsxJA3lMwx+N5IwwC8Ux0DkHeREzJGtocP2mGVmoP/GnCZZVvDZsG3p
8FKrG0KaH788vMUylcB4jD1MDWqpnBe/Xy9pspnTILHJiGwQs1BqbTWP+DjKT43jzDPimf+wHt4G
rJGXYUwZAhPHZnRPG6hEBJv97S5ZjAXMFhDa6GzfPany8gd9EZET70Cd/6OvftNYL7R3HrI6qpZx
trBmuAORiL/8xKwod7WKVt/3sDTRUgeUf0yFcdkUIFotS5460LZnOx/d5T+buVAiaJHXr5VZ89oS
rxNlQ2pEHzvS617GdW8xu+DpFNlrMJZCTymmrCpYW7J0NkHSiEqAuCnWsys2DNBvmxUQkd+Jy1IV
ehq2AKM8kJD8Ggi93s+tTRrzDRdkTlUXWzPc30cJ9G3P1BfFI/q+DN9HDvnVmURX4QmAZSc8hO0k
PE/QBVtPUPLNW0sXOXH1t6Q02c2DSUW1xw6Sj7xjBTrZSovGoPAAh6YdM0M0cX+bqHVHQ1mVzGg2
a0osob50fc50PrarEj10ngnMaJM25B8+6AQdP1WR77ZQrCLv8n8hYhe+vD2T5FPlUNmBdvzqB9h+
d8UkIK/e5vjjVkH3UjN2Blf/3vrG0JkJ+oWIuia0EKpQNiRL0oz8K9VJt8brltnWZpbUpG2lEo1r
hYuBr3U9uq9x7uaBDYsOkQ4fNAWXoT0p66BTXUCPPJYJRYERPE089OStnYd4TKx0fa+7TYQFImhL
WokhLONnDJWzK5jWpgYepD4wfWR2sIClFPSU+zLNgQfSLLRV1R6QdUU7r4a/S1dNDrQk1Ea0TZZf
qV+HL5aMxrDDWeMsKARyi2ccElS7EGxNW3uSFAIjDMch8GSBKP38sOzBJ2QnxLwbK0/gzLnVUjUi
dnur4a84WXihQvsCyoD+f/1oCNXqkRC7ud+TWMUFZf4lpBe8heMEfdq2uTxqvzta+1ysG8/MxLtg
/3aoekSOrQxrVtNaaCqc5sBxL1KEbzbAuy7uVpHZV51C7EQsKIXTYny4eufEymj/xsNvE27jkpmn
X4b0073UUqNKOEvdqU2CvDpKN9bjkW5tuQzPW6n6nEpwOAes3ulCiJ3n5ydJQY27zuRewtAlMEbs
NSZJ/50W3rq5gJk3+PfHfnqpK3oH5qq+IG0GwWd0GNWBG0HqYwI2arD3G53wugtf4Ofx0+3aXZZd
PekmMdIboQo/cCPSFP8Ikw5Oc6vwNhnbhasB4OCvXSMskyN7bV/pBI7RRhqJHQzBa0+nKWU2rE/r
BSBrLDoGNRYX9rBVEjjh/4PTz501yQ0U4ftmiGuXVr5wK0gcAvL8m9k6k2GfX5Elnv1LiTzQGjfw
Op17mAmZhFEw/harkzx5D/ZhmcTtP3Lr+IrvRzG+PrIHf/Ci4CeUGdY2zVkPhiClpOwHTeOLTAkg
AFs2X/WhomkWzv+6/u82wBjrbkYdHgEhasy7vLq14nVSgonkWwVwLd75N4lkTAq7WGx6Xr6mhOoa
iZdU7mESft+VejWMzp6FjnP+ExR/nqemIGuBnUSaI/coN3KlRkTj4YKnDQk1Ywege9fLDfRNc8vl
9ozESOW5b+zWAY67Pq60o5GnWizYabxVQKRLMIYRqVu7e1goCksw0wg8KrtJvfwXv9J3UDuiBI0i
zDAeJmMwcIbqOMYlbw+TFqe8cxdx5KLMRDMCxKRcIt2VDDDnBttGCb/frFT8rurtL2+3XLyGzrr4
GMZZH7ZXpVrDdtP+d258UaSyUdVAQQjLImHLQkWbWXkJPqjTDXATVMtujAwGloSz+1civ2Ff6Aql
DIXNmXbxnKjdzlvrKq0fV5czd3U0fR3VU36K5ApLCiCZM8y0Iwm29AyyyUj9J/xpG5gL/eeWKbYr
S4qo+rmUlgoc8KhIm2/3izV3gOc5I5cBJ6kVvwfxuY5tyfnmn4MEBsI7BsgUPZ+8jAPnqmohNc4C
zky59EaeP9NS0XIBVjn5bOEBC54lLC9uJ1iPWpe8ULM1SlcDG+XyU/81LYGqWx8VZEdFESJwNGLP
1/XAnupdQK2A1EE0qoJiDLl3JUwXh+O0b/0ytoLS6nfreL9AsSfzVS73PoXxzyT+CrZCpJW9wI6V
/Uyg5KPQSSvYE2Tkc2wyTMDX6vD7pz0dMF1uE0IWRqujfeSiO9DPQTVoTp5xgFBAZMhJpSYJ9fB7
CeMJrqXk7jnUgvQrN9MdAoqTvxmCdaFmq32v/H05ZglQFVgJhBzVbh7KDYS4T4H09dozXdUHtq2K
Ko0Ey3mzvDzKTZl1cC+BcUqX0ylDjp/Jbeykbv7sp1kktAlSH4F4SGWq65XTNwIiDm+Y4kDsXZ5I
ipdlx4i9dw6LjynJ3A9mWwjyBo9rRp4DdUjO6tZhVUNSzCCcGoA/EBBUc274od3sCuAPS6eZhAVb
9YKET3+idl8NqBxcnU8lEIwBdbk4YFW+hdNL32OrtYT04PRSrPLnvo0WusYVuHAl9YltyOx62Buk
G7x37Zrfx4/XWUv7Y3ii/3sipBz6wpXAw82OftlPOfli81/I1NZjfgnKR5i3F5LsCZL3wS+Wucti
ZDBzHB0iYeZz2DFIPdS7wG5NX2LrJ7a3wEY/U3JVk2TT0UHqKllq9Un12B5mATLwN5QvmniLk9u2
9tXsyBgCrK1/g4x1XVPpfm+xbV5U0T1fnzGggQDGI3XHL4npnIpGH6RVqrbFVGGEqQxfipVVYtUZ
UVvFBcC9teR0rrF+zfogBWP+dV2Fxx4a+if0yeiT9RtBXBvXiDkMEDwAzgzT7Tf1nFPJJHnlFL0y
wJAhJWPRdOcPe43e3+baBaxfQv7UptH74nj1zA2PbapV+xFIG+VHSsGLxmhnKhPoLm7O3RFvVNOB
x9uA39/1G0li49Tpe8lDZvqf0uIfcrrtTe60/WUxbSObcgdQGs4htDt/qEXbu9BUQebHaCaybhdK
wCWJcSjzmeNm7p/qqvbkD5vX5zdvZQ/8Yj/9XnB27fke1zXEWPJau7LcxFyNR4JV6LqGhdn4Q4kP
LwAlV/4w4t1TTWCEh2MHby1Fc6OqAWXrJmK4f3imHSoiBtShL1hmiFfaEK7mgVG+9NzFO3x47Hpw
tCZolj50mFAXkgpb5Kw+WeIh/PU6v7mSGFGUOvu+4G0m6DMTYkeVIv35fPdtxxXH3vbGeN7ZRDsA
lMXm2YXsQIuyXmgk9pB00HiZIy0aZuSzxFBphRfHXWtkT4hErXA4MJdIQaqkXI1wMjE73u0SPs3G
EOMwkRApLl2RdC7xt82m5P25xfx6Q6Pp5tfwVpv8EfMBDbqqH5A+fQGgHhjxda1xagmoAAZpviP3
Og9SM5XZfFi+8VNzFPBmhbrJCC0Pjwl8BxevckCNYAuPQHMPqP9srvAjc9CWExiDqmFIgtexB8mY
FPLx3wMvNVm5hKIWwfqZYE7lKde9NnrSXJ76WATEIHzGhOXatRBfU/q4RmTPsw9fv1Gg/+NMPTjU
QAFCramJ0IpsCxxYcS6bZoDS31mzNKnNTgapG7KdYF5CW96kJJpg+woR+4JMRmQEHvBBBsOHpIW5
wU6BfFyXK61j+xKCLqe7yZRUcbuv3vTTqG59Y0637LPGgHxPESZ+wuqIyLZGrTSStKHu0Key6WjS
MsgMygOqIUY7xQP9h86GmQhJ8U8643WHVUziVH7sR4oNE4RO/CWjZF/UvRbIZ3QWjU3Gxzw/EK1l
Y4qav2jWkV4/Gpevc40E/AZuhD/4r++flw66h9pW6P/QRkFfnNbyWoMt9v6wBr2sAD+uPwc+nINX
NNm3FcHCP/NFOuYScNJ2kaiMZ4FQrF4+Kd5k17ey+87l9ZzA4AzbShuCFg7nWpRsPbylY2zFAL5j
n/luuNdTP9L4qxDi9x2PD1S/BQFbA9HG1I4cATNzgyp0SICsfsSyD5Avhs3nQgWxOy5CXnF5km8R
sqI91ZWYP1YwQvCnEnLSP6Exf7BLj/2B3FBxGDeiv3atYAwW3najCjkLEfqqHWnD0rAq00ZLHW4r
xHTNI8vCp9CNao5567lUHcAghsp5F9FLNMtlVOY24KNVIEg0mZAVp0WfPpj89IE+/8vJeaRhBLhQ
hFZpe/KU3HQ+8eXxEfbqbMSI/+yRW8L9lwR7wn4ZwNKccGEY4eUfGtZykiVI45r+qwNlmP7Ah4kK
E71ighxSqvE2mWeWHd/d0NGLSjqhXcSPcUdD1AK5XAtbulCEbJQExhxnY33gb5gwur4rk9CXNQor
AcNJIh3Rn+dNjDu/QH27osenNvLIXmjSqyI53usovg+hlmO0xzOePTgNi3qNKXj5pO+OXwcrr3LP
0LgXi+riITUNR7so0c4g1TK5RQKCdHrZKPnmG+vj/pSAHpymScLoGxOy8YaA1Wy/SDerAZHsnWh5
dVj5wxPa1yiOL9eKjwdBCejhqldT5+gp7Sw+1C16/Gw5NmVlEMCDJ9wgj57VOnqiMXyv2J9Nyg/W
DSa9MuBfk2MwaAecANDoRnNVF9eVK0nE2iUBHFt6peR9q9uRrBWVMEY9wiqga9/srYh8hFSFd0uN
WW/9ygrl1SMOqbm0M8FNV2oHjCXaqAxcOObYUIlZt1ZcemWT2WpzujJJ7sNCvV63JtiLyFB8nbB+
ALm1XI22kXTRRYW8HyeLKkGJ+Sz6CBP8KEWy/RJ2QVZLtsjMrDSdJVfqh70myAMO1TX+3nSxxHqd
k/abucOn8G8EjvUDwFWH43SWEqMdLSP+kf9uSvJGD7ifEOUcChNuqPFfGwGdvXuegF+sg1fxk0J1
ugcF/G5Cky4he+9q71Ra7DA6B44PCinKydK4zzoWqNsgt50++HUlOAKhzx4qDSxRSX2Y/Gpw8CHc
Y88G2DeIJEaZVGlTgBwmz9zt4BBuCBi6xlKako9nXbTJdvSm0vrITv91K1/7oQdeMrSTIgR7gDLF
h4R038kBIp/2EF6oTKpa9Nt2g5Skfa7w6Z0E4LKX2lT1kDDDc3PvsgRno/4itRpDgIhkm1vKFtIe
YgB1rYKVPnwF//EYSH66baaeuy43HsVCkA1yZHAJAZPmoS0YnS7dvsh01UYB6rA86bmEwpzfNJzc
IPaSetMQsnSIQ5+hXFxDlW9W7HjuGclMSe1zSuwFZvH13UbGhNItp5wy1D8X1aHnFz86tvMsJZN6
BocSNdgMgzVSsIHr55qn4kaT98EcyZoZBd3AGaV01YFOEX09nKipvTG88Q8wZR6phx4=
`pragma protect end_protected
