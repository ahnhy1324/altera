// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
L5mAopeKfjCZgY2A5JhqUAIIynjzu+V3sUbZEtxsipRgHhobWedPgvisoADkPiNaF23GVPivwFQo
mOObF+3PhGrDNX86QKehA8JksQEoZjR2nRzivhD6b9sdUqE4yMueu1LjPWF/xYt6JP9yMGMbAg0P
nTiCE+Fo689melptMpr+XGXMaTuPY8dWhDB3g4WYZXyq6HdRUg7H07Sb7+ZbnW7onaXkjja1zDFM
f5vQxhtsBdx3doIRYzlbzqpQSJf/8RwsixGugcvNxbMJJm6pk/QoZiRR8EkKW5lZ4Dn1T8wES0s3
y/toCqn6IR4x9XsTL37q3g+M+bt0t6+7Joto7w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
2c497e00R8MouCxLUSa+EdO0ceGfsrpG0yYJdqeDKCys1QWV2Zw9udpsKyrEb2Zml2pXxNznJCtu
JT6YO/4/CWhs02TyuFGWDHbc15T2YM2qnxJUEGAuctHLIv1vutppAzwg8WFfvsom07leyL2NreyO
eAyI0lkaiffIqkliXJuGz0tIqlrZ/KidH9hXSBqXsMl+AqLQQXlaczFT3CvdjHfC2IhAnK/BFUi6
J3K9xA4ffPzNiJaqTMuLxN+pb/QhG/yBjQmVk2pEfu/ZQP4R4schmOT0yt4889ZVjBIbkLMHNcYz
4FCmanfSXkeaIkjm+J3zCmX7Op2fwZZ6iGVIWDfTvbA0Mh0QCOpuUNsmSRB31J+hoCL8t9r3nq5L
fTBDEe2u+A65yZhTGN2THyJ0bwI9lPVFtX/LkCS78aesBbOniMKlNl3wcPsku2ovloRLg3TUJzJB
hnA9IK/QVNeqwZxQvcPB4yyUbpKduWQJnTQOzmE5b4v39TVRCbZExI4BmhRBoml1pvwGeOjh6D4o
4yBbwdF+Kddr7xceXmtO1cAnxbcEaA7k2XrFaoSpRKIkPuWm29cP47i/hbzCye2Vv8cQmd0DPbXn
I66HNHKE0kAj8kHTjZ5vLHTNdumjdiqHmIQbp6VWIYT86uwKtKmdMNwD0ednpoTGnxiijPiyu+8E
2VWfJMgv0I91Nw34yGTaYtOd0DYBIGg+f/5EX5i4CoUwwXDOC/NBIoxkgq3wMA4/5WkO9illTVbD
YjBf1oBHKLuLRKCvcVVRBQOwhqiDLIqywdkRP3up7zGZ6YfKGhHvlHN4Tcp+Cu9YaHYHAvgiX9N3
JZgkpRlXp5qp6ZeufW5uUJeQ2ZkHXOWP6NWqGWPyx+xlvkK8pAwLY336pBcXx7QuXVxSN5omB028
yqh9SLbqSA3kZXn3ktMvFRQC3Ax6XpgYcnjxBuY8xAqYOHXadTRPbg7NaE3o3xCWXocGDx83paJH
zlpXTpi6V1tcJTGUWc2Oep3Hd6KunpZp7PEXcIFCa8u8EOGrwZWHFl/M0r9+KRXWywSk5dZxbx9y
xvMaOV8X44o6zyuiWImmEOQ/mQZg0sO9j/Ey9fnrs5z2kHFgpxuomecp7MV95Uqu/rOm6DTpZX/Q
qD90eFeqn98eKCF/Bh0iMSFOaBP2FsZERgVJRano20H++yyBN1fTzQbkgSJqKrVppxY3th86oXup
YC1dB3RRlduVniBEcaI1ofZ/mKMF0+ydO/p1MdJP9VFIErAHg9/8EDmrkgVeUooolkwjRiZPIQto
nhuk7l1zxFwzjsSdbVtEmyBBKgfaO15T1UoSKxS4qR0dMtITQ056Q+58eb35lefginVO1fPQUJHo
RMzqtJ0sdFa20dZywEkz/lmfAVhnNXlrnnsh5QwFEp1gaCFubg7tyNVq3vcoqjyrxiaE3ofWklmm
30gDaRSA+rnZsoWpF/3FgvSgzaT6mlfBx0pSlRuhZvXf2P7AbvdJbzECKWXPnZc72Itoc+4rzvkO
vaERvYvep0f11AFWHlztO6oZJAy6GUte8W8YpB2cH3yJ8y2ppVR+gtI2OwwaVlNJ5BFudPaAHQ3J
RFjsydbhyClKUJEgA4lO2ni9ZiEK3TFGkFF5SaRxFNMwt/HMk8Kc6UjW9Dh/YitpWinFZuwmwg3r
jiPsWfIdG9y+u2mwtFgPV93rXl7ndrHotseAemSC+X9Jj88ID2mGTYaa4XilD9P5j6KhR/PEFx+P
XmeZnUAIYcgG8/EdB5tHccZZ+VPAeS0NybftbDQ0sh+MI3uKDF5dQJV00JQOSCC3UU28emCiHOyX
jRSFKK23qN21VLDjQ4Fflv1pMSvSpHo4uk/oBPcosZaYZjBEcgC43bGlKgAOfDwHhby5w2/0+zEv
MpZGCcOZnGJY/sR9P+oJVYbZqp3xim+g70RXN/DAQrXC38ZQRLER9pZdZ4t1IHC2q4xdw3iKRwEP
qRk+IbCiQkGn8er7hNMlwftfH5gv5EPN9gd+MkSNhIEuxdBIlSfHUCX0opM7PmXce61FWouNDtCT
TZK5xxflc7uQpKY4Pt++t46OtVqZAUUJqYU62LvgCyZiGv/N04aF6cL0XZnbAoEqSzcPTGDCHlhc
iwJBzOTajg5j6K6Ykl0mtfy/++fcZSO36bXDZng45DYJGKTeY0OHTiiXxOHjTOE/kmmpPOq+8ih8
+wdA2baGBPoOX1YYCTUwtTo5j31jNhINAEq+1DjQLyCpQtJLeJymbYXGfwrLHwn43A24XZlVuhMu
DaLfGZ22jDLgKvVvE3wQHPKqBKVutN7q/4Y4ai+FTHloxk7jRw7xPJHJ5MGf5Zpg2M1DUO6VaG/X
yZZX8KQ8r0lJOqad9+sYff6T3nWK8PWZVElnIY+G7tHc9KzDkobHOaek05re8xTZtd+ziPCFQUYE
/uOlQ3ZiJt1YEE+/D8/saO+NYVnwi0h/hKeTBETNes7PcYOopWJ5p83gls0knXfGecbhrNs/S3EN
uXu5Z+QGJveJz3t4dbIzdW1AzmuyEXhUoceQnCRfsK5pFpMSKwsJjiLoMFfXDnvO3S5ZWimrb5aM
fVcWzszRBRSmFLEbAyKYWQX1405/MwCH11JO7GVnp52g0133V0fcJ8cwISnU3ImRNOIyyqcI7LCk
xB+FgmzI6WyWIhYPdpvRpS0L5QbsZamLMk7rNazgSf4sIHXcBMnwQXsa4GFT5hJA6TrpsQJX4s5n
R7pmuI3ISGHsxhK7x50hl3klycqqFsTgcpuub2gBK9Yt/qQi+VQyAs4TWXttBhwlw8eU87mgGBLb
09WR44/yR4zA/iqIVTaK7jz/TtBCxKAS32tgshkeOWcBVergyHGGFff7AiA9Hv8Gah1sMeUoG5wB
mt7vs4rTyoIYRlJy5hwYfByMLIkJLep9GL4jx+K+srp93XtbOjfQ/1eJspFFKb8Ve41fZs7Jxhho
Hl0y4OT/+aDsnercB3iThlp/g4Q4bBFUFO5wB8ribGyQliSFhgzFI82V4pPMiFZDSpzAtLXcFhIx
W6aGf4jLG//Q2bRa0e8tCtNBQ4dTQNQS3W7CYFRM6IFsV+379+OMTGCWQHOyjkiNhAaqhgsHMLFM
H0Lwq0UlZccEQNuqHkWg+dIT/R2P/HpzJ9fgHwt5iWYmdopUzAwt/2gonNVFOsNNUpiU+MWJx2VL
esJ7FeOPBKpKqGPmlzxnknBZdDx9dhM1AjkAsXD0a763oqE2lycoHaajRB4S6B9XChHyO4FRaah6
g/xpm9caWOEM3NPjDfZ19yUs+UyiMzuNaZCt5QA8e/Qy0o9SvQwwuFBT/KLKmZsj5C8du68oQDY1
Oioob2G97NuuBIFOGII9SkCyh/Vx9WERpd55WrvgtP3qwkPaAQe4hnWuUNdY3iXRyz1M9iR1o1Wh
PchXt3v8ZoJCYyXCB1V1EU7w1JY5G0qbuqKfH4M/DT6Arwrfu7UVpk2/k3Y8UT58CCCzzX0PtkE+
seziG0Tk4mRHqXrS+V406ZmuCT6OXQ9eHU712Qv38wy3c8MQJLbHVe6PNDB3wDRMrSj54tkpdpNS
pXLqOEwz7nLzRqvPc2vfqGXCPkJ2/Bnk7nsXb9FOoLvX9aFBIylcrSgAC/LWTdgNm6Te9O4QyEP+
n4YaWpFS6TNVYTvXddp0hPzMAKJCEzJM0oVTjSyuALnaJYk3MoQFUzzit/usNYSZ5molwFIFnmUj
E4o1RB3lLjpqbDnhdeBVt5qfkfHnNS576GXqoycY5L4MqQK/b5F2IdoGY8JffBLQmr0WJHy2RcWm
s0e99NcxB5mOfIH8oFfKED15Ge+LCdQGqNm78j9eWDGi2M+yXEkXvz6QoKVLK5a7B+0W3OBnOxGi
vyGIHsKFJcWb8kX42xOiICK5lHF/6gEiA8o58H2hZuBRrUmVmsx9Wj7z4V8218LxN76KQ7HOSfo9
YJCLxFUlylrHA9t2qnRjRrl8RPetaG//QlukdwS3jJVO9BWXEQexPH1hpoyrX+YWkLUSGUv5fxJs
My9kHAbupLbFtP0pWKCpDgTFTyqqdugfCeHmk/FECgtK2R0jLAX4+ERyrhS0Z3KzONmvfXGPsIUD
/iFW6CNPwm2SLl1PDct+Mmc4t2JA1oy9yqSkTEbUHNmCKodX+0KyvL7y27uEhHGeyZqE0iMf6NA7
KEaK0gUnz+izzG06IRq7ZkhlLguUviFYLlvcel+aUOAed1tp5Svb4VnocRyynl4an2Mr/dDo9Lj5
wJB3WUjA98mlMfvBNfLSxMX1KvB1QbeH1lka8U8GEUEIeHMhI0fnEeQYojtOG7ojJV7gkFzftK9t
IEyPijZw2vyCwOBVPTxyTmJXwwcjlwRsFqYxvKI7oHjYZD3GcVum1fsncyqDUWYdrfI2Qax8SPMf
yvo7vVn3aEv2MqeVcUYgBjgc4R02/id9cBpg7fs+0ncnhyTQ1wceovq/bgPkfD1d/OqnH6OHJLoY
YU8RBP2fF3ESvAKt2kEFGjWxHws8DsJyZekzJe007YBFxgt0SGH2fy7kF7wRacDuc1WGdhZfyOWZ
ZtVMdri6Cb+w8XLBooOzEeATwPGfU24YHI3bYmhtQQzXV+bSkpQmIXTl7K6RvzATTwiv+//XfRkV
aLVOmonrKFbTa/eI69ZGrVD8nAwPCsEyaX93CGVN3mDJWvz90/WhHiqPnGmXI+ViexTiUsZbGRQ7
JBpFCF+GHQIPnESs13icdA26Kn5O+JzMT4OY4IIilljkjx1zE/NLhx9HhcmKc4cv3DlBLv8s6Fnp
9wqxzJuVMb4zwn/fCgbobxTonLKPY/hR7n+wYPhh1yUUICSxZDffjwer8NlA7Vb9XL34ShMnm4aq
Wvz3oWAD1zoPxP2fWdDjaMRUFvdtr5SI/pwn6apZljlhh8N1PJfb2PJ30yE1c8so326PDb5kbXZd
OWsyYDJzF0kbfdOfhkjfREh/Yp+2QNKzVYz9K8sAw2qdqBenuuc7lMg6MfbOZILJMvV3B8yrhxeE
vbA3TWe0rklvU0xcskyOSjYRbKJSO6NiMdN4cfp0VGLh6iOsI9CZ5NxbCBlLd76Maxks9JqCtTNt
2M4yc2uzYGVyOLUtqKr5eDq0pnEDmtDiO78xCrbaHV97EodtFRpDPakdYBEz8W5PJfsb8XDMdHRJ
OSr8wJblDRiKA3NR6yxnSpkcuiyXTBCxVzm2MmiG3BUUbKGNua+Mf3C7XrpIE3r0tEJk7aRjkiga
q5S8E6Qv3MAPwLG2ujwne48VFtc1zDwxs8jz6qe3Jj/F2ei4lY/ziyDZWIHOUgIu5XwlvSKV18yt
LDTrr7BIVZlvWPGXYNvQ9Q1nSnByB6I+0ss+1oNJRPmc76CPCFYkI/psSBiD7I7wB5sImBrCTzVn
y/fW3ukw56tO23EHAXZfz+RAXUranGsFZaY3uRkFUOp74p6X40TBHZRziNeawnYgDT5vTNhIDDVE
vfbkyisX6Uvv3kS12bQtbfbTuQAVIxdFC8BweXo3fOP2GSsvPGyr7BEYHny3pry+9gV1d2d7xUSl
rUVXyhgkhc7pSud2KWEhrH90yro1kCcfcNhDM1ZMKjfdy2+vCF4RWbHglugl/eM4If8/heBStmUK
Bd2SbJU1LX3j8B8TzIFDkGky7HOWl/Q0Xim2RMPUswIoozIabwQir/8jtVRw+O2JlB6xGYh00BSk
SXNWKAfrlJPrRXM4KyD/4gVJHxaLskLvn+RwNtxPDZXwpSutD6xO0PvnV8Jgj2j+gIwB1p60/HLq
bDxEmYPn8zpQOJIRkLQYW6VpxeFhyreAd2bZITt36c+1g01CgZ6BQ1QB5r5nZqOhcTzBJUHCD1SW
24hR9idiePZV+1iPz8fkb9Eeyqie9uyYSmNROZWlwWpJC7upln/EN2yqcqMFCRFnq1HsvNP204eD
NunP1j3ZJfoDrhM8ZkkdWUhoZndc/VYML4U/ylxO9N7GUcKDFHbjcRPLpYZeoKcJezFC41b/NeR0
UHrpRTjIqEMaMp/IOkV7Eb8LbfHo6kZok6K5hrBEJsflU77w1Vgr3wR+zgjxOc2owFNcR5Jyap8z
/7PBHq1PAARgnWYopPtVgWVIZtSnhX1+qb0i3x2OtPnaQMu06gwAI5uTMFDPROt1eBF18MaP5OCk
T57aFZfGYszb2alOETGoaUD2zZ3F9aJFUVIu5/yzFUzmvBOBWtNzDwlzK9szlNlJ2Trwm0iRqXC9
5olMqw3UYppHk1s/19jjuEH3qjUHbYZNaHQlosJJnLoJpGU71MDnZ30K3DLMZtWs1Du2FBir22MT
aK/6Tum5rXhDLPPLWj6bPd9eF0f7NA+JsXodEgwwi3D5vAZflfmobYP4GIcc2kCsu/EhyYLBFHLu
iX5eVSS0CCid0ATazi/JRkpGJT9tyj+E6uFojqaJlaCJkMFf1q+TECW8TwxTMQoFqN4NnkkASNV7
XgKVcZB/DZndWFGCX+73RSUY1ek2PVfn8MWs9G6tuNR70DE4Ut4vnHsvp9cSFaKOVXR+hX2zpgQS
FuWv48QEYwJ/2vSRWLiL9qqLbSSKD5YCnaZ6yRlI0g6pGqmBPiDWwji6/M592ql94ZI21jn/tqgU
/4WEx4t7c6OS6q6iX3wpWJlqZYKYitQBm+29OpKNWy4JT1pyWPz5ceIv4ViD3yp3F2ioABdiOj5Y
qo3SVWP7LaWJt7ZBdpxXEkluT/HBndErL/vWyfksWVRbjFKdrfVwy4HygeOuUXvCRWSLZxiI27AW
6ggdlaw6h9zt6kXlgLbMXMGR4D3V3l7S+XY3l4YUEps0uuULyrWfGQt74/MjGnnkZK2O/gNZ9Tsd
QLC/QKY0NZ/7Y5WtRhp+4jEFPS6/B2lmBmtnB2zjkwESbxN1Kq8kuhMPt7KjeiIHEhn4eH3kjDxt
ji4xOaEpZI3wlgz7gdlQxM+6zQH8YqTeXq332QwAAiuQuojJiTc4V63hWds24XxkSsmlc09q9x0E
wVBDLmjIagdNLTdjO5UhLmSt2+tb6Vnm578VvNo26Vccu+hzBN9nGG44ULMvCm0JhSGfno05mS/o
SIDAxhJIdfz/jptwPMzSjVUOqO4f5n1m/T4f8DQ9n9YHiKxjMdEwoP/S+Am1I1rDR2zcNV5sJf4D
mlOsoJ4SIz2JO/Q/mJ9TM37OYnc4hnOSohOkw876v0uO53XeUBX+83v0fZOvEd+8eLw+mxjBnUdD
g/sjy3HSJEm5YSxLgOurwXiX+w+vbHqJASNyTEgvX1ML+0LerxUkPCvfa7vaZjHZ1iS3Hbx/4fJ3
25CxFakynLfHycvj4rd6G4Q+/cVOhLMhp+HDIHGWaIjfe3A7Kfp3VuTr+cnWcsAS+VJBmTL1jN7+
K8bxYkLb5ZAhcpoUEiyrcK3U/CehDD306Kjdk9sl52rVvyEtVp/Lq8J+gfkgkoRS+MJD0wn9Ogrg
E6zqM5LKa0+/+Xf1vNufmrZHrD+eW+/hxzFQ7T8FKTcledyjMaUJg4glIOIYeh56XAMIsY9Hc/2j
V5q5PPeLqDB2ZI0bVzN7tp/1X1eCiTMsV22C4wa1zA8yFbO1NUSexMVkDrTEpi8K3n/zQhfwYFuW
dujkzvMQibqgNAbx7lvKDKYZhe3xTJMTbk1bzNbdUoHujnIWObaHxapq/z865gxZ9DNg0WMEpcuo
ladonbTrUUuAdO77/cQzlPIExXwMgB3h3ne1csouAH+uK+lyGrzg5gnJ1FFHjDA197JGBkC5JpxQ
KZ9A8oRDTFis/CejGh5bkCyiTHFsbaqzAT8VjgGk8gFkrCRmdQTWNkrFdKbLEi5GW/DYCx0eeuiQ
e34kNB+5iBdbNlUs1yeDz35uQkXRphqnbQ7Y0lMgWFnPNP0rMQTEXvxiOpsD20jXlS7QZuhmXcPc
OTpexMMN1/xI/6Jnkr4sKDrOIwx02QwS24JCGqiZKPXfdqay+gnW4bu1AjIQCw8FACyy6fl6GEfz
7cihokd+fif4UV1iDNq3ETXzHT7JbxGRDipFCH99GJswiCohdnhBsz+jmAXE0Z8OM3V5B7/2Thhg
/UCQiuuwRwsw+xUqOlUyhAAwoBLRf0ZQc1+c+tFT9JLZpQ7x6AwpHLrvYh0Njx6yyyGmPSz+EHEU
uv6f03KVPUTVEd+sH14rflDjBRRpUctkcSy+FDKYYz0d0DHGsix4QpRef+bzfat1V+fdm3R/xsZl
7p7izvZAGHjiM/f63ZKIYA+YJUvq/aCbOXtBo8WhR4XQYNA+i4F0ZsUk5vBK1vwjQQpGXBb1JfFp
qKWePSNykFC6TfAPl0HA9zGvAZ/jNDhONp0/fdR4RtMd8YjuoaaMMSYAAGzO2SG0vmw6HKG+idmo
sel0slIvsehirYKB53+QQWhUzRAWngFeqW8a41Z6rCi9d3oUJdUa1qmGE0khGChO4RY6W74Md2Sv
1P6l0wIV927FgUvmqtYqdLPtbJI5S8h4nvYwjFjYNG7QKzsvemvZ9r66cHJmEDDZTnzxbfHyzryh
OIka8fM3479zd5sFbNQyLcUDv7tm3p7o/RcR53nnjadV7mhjN4jfwXuJ7BadUwGZhFaWZyu1H1ge
rgX++i86rrfukFlMhFZBOUgiJn3Fb0YbUYfeJEF9XaAbP68uDHtABrlLwNFCzo/x+vtrXY6GDmki
z/MDaKvcOPRf6E515sqeXS27CpOafXkRCOIDsNC6MMB3d+YMG8ZAI5JZU5jbyP02LuYbzTy1Je1J
ty4jrymHKSfMqVMYX4R+/QjZYZyPV2nPl5y9eCuzx4zTw+J1hVy0Wl2hhe4tSN4f/d5WNnOk6FoI
tkhSY/YxN+WOQ1cP6yT2P/AoGcWYf/ZTnc6Ek8DHGrFWlxwXZqDH2GjTJQqjIO1MgnWSw37v07Tt
S3wHGrPV7GjheAPoTZ3plO6krlIehc7uJtWacuVkuj1/bmU+hpzkJm2KcLxcfV2rkTWoFQ0Ce1CK
TODauhStSUK7iPrYI1wut7zEXb7wsnXa6G12tLsIJ3rFNwGpaIeyUWQMyfRNwSOGAdr8gwew5ecE
k+0C1JPhqNPTPa7gJ1xMmGBygrdKLkSxLlZW2l0zWJK7hET6TvNCZlNqcw+FzeNTrZJ3QZVP5zcj
orkFsyiCkdTX7oVxIyvV/ya+ffhvA890/AUvgQbyCE4+dPCHpbFE4mMVH9H57jaGu8ZCZwB59eWY
vCm8yYK4WcJSEe/CRmorkC7IZax7DUNKcHic8EPVWKMY5tFQURkE8tnHPmnyrbl55ZFkcEPLnyJy
WP+KRVYIfdDEVrFevf+1DZgUSOzLtRriSvkQWqolIuseRcHZV97Euif/wKGLBPF0+eZCrvCtBJCu
jbWuRxZQ7/WyvUupIPSxBoygJ+nodE0WOnPlk08dXLxfIfZlAb+wVsa/hGKVE1gjRck1vFk8wdGb
Y3XzQghYst5OqyRZ75TUnOp0VaFZFRxlhNXyc8GoKlfNSImnLSgoc2Kd3G8Uhgi8Khib33rpJ5JD
pTDdTj3zLi9LH9wZXRpBpH411TZh9VEe5xkMfa9VBf71zQSzMV9ju/bByEwfvPjGLokVF6u2rA9Z
78CsiQ3KVadpKF6gzc8G9h8XdNvm39cy30yoQBRwG8PijsmhhpyLbfPGbsrVtsZZ1kbDgCaxttWX
pI0WXPSOzQAcJJtoQ5x+CT2dnKRnJHtAIMZOdnwCQLPVIOYe7usIA3DOLWETjdwEAVt3rBJ7wdgE
UsoUpDX/df/x1kEGAvZoLi+r2myo4YlQlcbdpOfXM4n5NQ9DXqiGJqys2I1SIbh3+HxDQy37f16S
EVPWrzsiz24AqiwT50lzgePlG09qyzWbjdxV2HJZgaobyfx7P6Ax1wXH+lV/iJ61wrxrZ785iGuA
dLJuAIkwRt6cWDFZEppu8J1H0leflJEN6we+NP9uzArW/XI0Zt+JxiCF3+C2Om9shjH1V/Frftj2
OPos82Xt9nzhoqXq5AKaChdr1Zm5oZPbmpDKJuwOAvSsoajKp4iwby/rROltATaUwDkUGB6z7SIw
8GJfUsciqRINux61Jus+JQzMtiPoGD+EfpB1vt6+oQuLyk/ePOzYuNHrvsdj5rUqxDxm8FXzbOvd
ZDq25vAgX2VPPLCJet6+TvRKIcOwZKHw8KO0sPhFBkcwpoiayjN0ICc8vwQ+44pH/pBIvC48U9WH
y47mWsv8fHpzszhJFy8BzCY959nDp7eW+i8OWUayCTIBokmvK3c2zqzO4nM+m91QfzOuu+TXmhnV
GvaSSmueU1UGYmiRCqn+D4Oabr9V6puxa32TCUQ1C65v5qFTHdc5ofZXkg8k6iJZXOhDTlOTkOgg
oML8VhdR/n9xUi/p3W9J2/SZPUoVRlkobqOr4PRu1H3WZiF4SgXP/j7SJxYM2gnD25YbJ33FbmX9
6JDjTTr2Eoe4qRB64O7vlZKcw5Cyz6zp/f24w5hXhpyGxFV7fpiFUKKrZagaX6cZL+VLp11z7oCw
WFfQLpJNfELHErb9+/2esU409p/XsV7Nzmma5F8Jj5jfZakrWLNCCQgIbbRJg/vmlt0YhXl5zFj2
XqyCIr5hpR4hRJSQhiwVhgXVCmJY63snHhu0jwcy11rw3yWW7ADV1xrbdJdlgg0m/2X65CNDd1DL
1JRsoW1nIdy4eKaHeDhs9mOUywqX//30t7nh0YG2ieULglXiqiW2wj2q7y88aE8Mo2Nqr2sEALGh
IjLeeMauIicGqlvY09JOxu52knRUpv19ja8ilh1g+OjuppsmtDWy40v5bCTYegfYPBG7KW1o8QsW
+Op4hqcmsnOzvJ7OF+8Ce9lzxH7bqW8eQYQZ5dwXmGu/74hrCZyD7/H1S7Q9GObHUkU0Fybfwa1J
U15+Zu0n6JDqfkalvI31s0OfLcZ1L1R7ObobjHf3ICIqxAbypScjIliyBoGtt/KQJMpcLb7APoSo
F05coMjQWzxGSmRfciZP78dJOzrqWrcsB4ZDQxAzlzgWZ1J2ftFB5hqBQl9F8SaS9TzNbO+Uj/MJ
a08y+S3GMRI4FSJg6+fkvfEjIpNYPqmwpsZggcEzKPNW4wBr9t2ZSm9wjzLHXPO636xjQ5OEZumo
1t8GCuUplRXpQFy8P2tLmFfkmil1KLbhtUyLYgTubiZztyeKj8hWeocCcTe71Ic1K8jkJIPcCeNd
XrgnQuH4guBSxn30XU5sOomOQtpZcZBe+s11FnYZSVdlYlBDJvL/nuAEjYUyzJ6X0/s9SIeg0f73
O21e+cMEH7hLyWzyULDMCACPFkwxLVrNYaPIl/zj/Q0/MgfYM5c6IFWXwut6ScFyLip387V5/jKE
GM5Rt9hU0CTlUScF0ZlAcxUBoaio2tTMBzGnuWhME7YIesUja5FTzOKRAQXoEXAxmlD86hgLGw8a
nlFPzt63Vy0QLXdyriNevzEQ3Q2eXZsE9MzJsNsq/r7wNBwkMsE6io0NalYgeGlI3YfMby0u+Q7j
7k7Bgx9LA/4cVIE5CF0q0yFitjYn0/y8daL/lsZP4sSAeBbDiN2fKVKHKl8APqnTOvmfO/vOM7gn
LnwQmmAMdn8k8ty0TEDKLjcmu81u6CDkd7Thdh0Y5V56f16XDVBBh7LWlJk9rFyaBee50cMPOVyC
GpFOw61QKmSIYKYFPrBBIHom6wL/9DDc1ODCZR0eAv08vPbS92jiY1mq8GOHwGlRkZECRnpYlXy3
z6+HzSOpM/kRUBE3L3pjjuKvGEU7Oc2+h2oDk89+uLxr/uVSm02egtDM1vhnQtzH1MOvfqvEjeCf
T2r8V+fReUGzP6Md5PPEmJA9ebQPo2UD8ewUJrBsb31A0yHTPKjo0d9ilztX9oo2gBeRKcE4KWGM
Z5fbX2QW8A98pT81SalhKv38KPu1yVCmhqFVeN2tUgCn58ssd2k/c/Ac6F/OjXv37Wfmc9fyFT+L
fF2R6BWk7hpcYX5SS/N2VOnD1Kb83pYGwkJNZRWVwSbLrnbcNfTxbdH/COWpiPkJ+uCHiPIETlJT
yADb6Ngbu6tKVGKPzMW4+OvSQqepbFKECeDK2hXOIFHdxMjW6D7w0ZgRtuCvoIq4eXVhkQpNRBeE
+1GJNBzFY6JVJiTOg5sT9BLVfPFlLgsvWQ3+kVzaOUtDMqKP8i5CE/6TLJtATIsN8tEDXN+FxJRc
pXI6FFRfnRx2I52aSdKY0wbTyCIgIjJk5UECj+7FplElrkqapdNclFKpia1PeWWlKnmzuCVDLIB/
IjrCwFrhuaijvMsQAcIYUQ0sevoPYCYLsHicNG0kpsDknbWu/KYRfj4aKbMvhPRNSZ44YpafMdm9
VBjw2uLSMjiPlBCJc4ZbFHV+6YJmLhAs1A3lZTnzSLcbHIwf/oJCNpdFCY3qorBj7K4agHFH6osy
TL6/713/5/Yff7F+bIxqYrJFRcnWFEkL/1dShUgWIK86cpYRZlN3adhNAGFpJ7XATkD8c+RhMLJx
2hAmTPfcN1/bfPCaJ3LBn7TZI9pD5z4ZDf4drQ9exZpHMCkjOrCfGHfyORan4hsb0D7xc72hXnWC
DYIOQeKNUT/JcrQJbOpdD412pf7NZGMoLtJ81pgiMD9hZ4euLzd6nd36DsaF44CT3b3qINi1HiTW
HYF409NOH42BZIelpngLSCIXT4u6WYTKfqzj80OEcth+UGhMd0PxF396GHzN15Ce2ec6q9iZUOHB
NBarqJ7wv6wuDYDvooSbRIzIWRwD+XrDFI1qJumouhCrbLmD2rJ4kxyx67GID/jH0QgnDhgC8bb4
xpk4va6jKcDsnaITmNAneiH3mNr/lI27vC8A53iI+3DOyd9MlFtZYxkT4B9zGMbUQZ7iHYmrxG/c
SJx2+i6WFd4slZrPS+R1nvgjozVqGBY/V95NeL3XT/dqii4t//3o1/dEcBaO0qlor6MSZ+IFNXz3
tBG9PxVAnvw6qI/Q4hUCH0PlsIY6TyWi6WhvHG0r0ncCsmYgNRXLOFdDTUDqYYjWrTnqXdL/VUeY
pMia9xfLGPSSdXReTBRmkmkx8VnHrJuKdrlcqnLAPEKo3GEtkLyHfiUE7h/0R5hxhMq9NcWpAkqT
890dXd5D5C5FprqK1uuEtdpXdpNecybRT4as/EcLTdUxzSJFU6DrV53IYnnftFf5iz3v2dhdb/jI
XRzmzkszr5THjT1B8da+F9biE0xcyyYnt4FeyCoz4CceBQ9I8k4KsiCSZ624BmFDf1xWvTGOZx4o
YembYuOkD98FeAMu7GQnVGUPgfsNmR8YbHbrAhXOaBWecFae/oY9YJWzsBYEc7VttA308UTz8uCW
OmhkA/v5mpW4c17gcBlhWEs3XCBVqbzFpPrLvZeykHCdA6wMJRY9ldlMj0SrzVjbqSfyxV/HvizH
C1vXMBwxB/8VlebMUH6tgOPCyDorCgmIhpZ9k8Q0nT9xyltOobFlKAV8k4k7DqMtdXfNH8qyDbS8
27g7j5HzUPU49X5KVUw7IjfAWAYSYndUyAvG+G4A75OLGQevuqmpac5MeeKyV+tMY0wGh8AVpW7s
TcvHaPr9XsSqbQAbIYm9SybB/q/4S94CzyJuPugE3B7l4udBtv6nmnhnuJOODM0hSQVh+ZiptyzL
f3U7VVxilu9VSAS+QzXq9l6+KyxxuqXl1+6RgPMFTFFknNTVfLZ6MRGMfl3qwnXyIYPPInLxkoqL
M7fpcZG0XWWftSm16cfv0Sf/pWkZGfCvxmcmGYHPKCEorwMjgxjBRb4C8X/+UIOaMmtNvRPZg1KM
LLxhYGRAWWW6RbDfe9+0Bxsnn3PimvUUYHqYqKd5ThzML29fT/WSZSoHenDaAnIOa5dB1RzPijvX
MZT7fwdkJANPL9RJT8hl2z2v3RQgHEk/R1Kvp6l/XCUXyM8G6ksU1MXGOqik69o2A0UbHZquvt16
kv233MIBMR767OMfGDMituQ5+q6xsDwOVHiYa/HhXlF4SnKzFqYlEBYJasNgokpZ63qI3aOUqrpI
55lIUJ1+h+aerGH7C8ouFPJIpz29hmgAwC89ZcPwsZ/VMUaA18SUAlCb/tZTTNORBzKE2zaUQh7r
nSWILJXOc19/vnyE+/ok1MxNJY81GJc9rS/uU5ffLEIICWXj2rqhDJtSGwNyb2f6fTQ3lqGv6ydJ
AhqlcQ+74jdqV9S6os5JKqcKfRC6XwNnLOJKy+1ZvqbznTD0qXoroDFKZTB/5s8/1JmYz/RL8fbY
YiGogiHAYr4ok8CFwEjzpEpEhrbE73RJCNzBPrEfinaSkwg62xceIqpLw2WQDAJxyDN1CBn88+Tn
Cn8VaAExopBmnvOlp4/IcgHpawHG9ulmfej3wr4+By7EcBjNWzyy+4Te+uGX8LKyFQs43anGprqS
SGQF9XXizjrJvD6L46WUT7CuiINuZUCpJ0FWe7eoN0Xth7LAQLgmeRATXstxdUiDkC0mvkvdqtAa
1CXiVPfBZ8GAoqSIPUo2TKXkLjkmUkibRqiCcxH/RXkuoRuz7yaTm2Nwv4A/MBsG6Zl+f5FL7Fg6
DYncjiADjLEwPmgrUzl0W0b8OEQJH94chXp/W3XaX4UHLmda3+QVWw2+aw0fBdYQbnLhvf8bF69H
XKrLejBWX7h1U1qGeqJhwh2lvdW0fGhPq4hOBwNtjGIPeCF7h3L1ycZaFyMEXFNqBVjc04biFzTW
YZaSBY2oGvtcqPgmlgUjPOGgBx/w3ecNcil9gRUVf1PZgLVYm0LZu4nsITRKOiEMKgiR+j85tqq8
bzUMU0pDPKvwYZhSckeYS1Tfbmj66LFRSEQX/R3zkxX+UJ0sa9/5kOL0mUhhmwSRUgzdxMDm6NBY
0b9Rj5WjRcclQVFxuoYlZDHrxj3KQvWGRUc4cofXtYgQrIrqWFJYpP6kaICtZBeAsjQrFOi8HB06
px79EfD6wpDGqQvS/o+aLlS5XylmEYmvN6EiSXEpIlN7uSkxEG9w0YPyzdI+Z0s9g3MdTp7YDGjj
C1wD+joYw2zwyHLgppPlo1UC+fHEnB4KrIbouLsXgJRqK8Hvq1co6q2hleT7ujjcuHO7wMimznfd
cSTmoH1q9ny/bPi8pwdU6p9SszY58wM45kQpebplwizYI9J0/MzN7LPS4a/koYtBNA5JDoyiniBC
Gn6i9hJ6TxcUDiZSodIyypNI/NVSlGdRTAKKoY3hPw24j6Jah3URnsGlH4lXhQf9f1t9j6NEX4Qv
w2HS5GsKH8iv1QRarnqsrpLhupa4dgRnV2WnDCUSO0NxCxBTSaFOBghwY2sACO8yNv7vzLqKZZci
tFKsZCnyph5F+xJhb8opYoyXR1f/4NFOe9ZWTgyRw8zqMGHeSIJIQLQf7XV463xc/V2pVful52mW
WhdJ5VZeiKsK1JeBoiLtW5aTlQZkPEvyRCSL/hEmBzHgsN0pktT0oj5wIsaQ5csHNkCIW5SqxQ1N
9ufG4dTSEC6Xse4e2NqwK5yzj4cqvFI1BpI2EUzQ02ln6CSbUDCN1qnj1Jbe2xGjegs38F9/9vw+
ZR8Kwn+sqCJpCtStMaXy3gHxnsPdmIbfq24pVecF9qltESLZugeqjjWWftZWDFYM9jYNFAI43rwo
4fym92oCgSMxZU0JsjTFRsym7clIz1Z/zVTe1NITerCtzlOlQmxa9iRrGIDhF9TnTFPJP/zYvIze
VfmQNwsvNrm6oVzIVoX6fNoi2eWWJv+iyyqrMG7nl2uv8pldb/zBQFrAYlo0aze1kT0SukGoqI8J
JmhoQgi9vJIx94p0oyElFGz92b+YvQL2Ojn1Cy6np+jzRcxk4cDAixzNrWMT6ssI0tGoA0ZIyFdx
lmHDoocXJNcmotY3CmEJH+n5mn6mgBYp6SZJ8mbm37GlyTrMgMQzv7xbYsPLkn1WNYRxceFQf7aK
ffxMu18WmFwUjjj5OPSGaCasSxJ+57pp/n3vFceztT++P5OhU0BRE/QT0jB5CTYfiUGcevnR0I/H
sxLSnh2y41Dq3Mk6HH210oRT7MBunzedhMkIhS3Jw9KhXnKsUzV4aLkFf7ZVqQkv8c5Gmyxb6fB5
FWKAMDR7Yyysx7LETY0Vm6LHdE/p7R7i4GScBno5yAWbiBFowYCcaYkMtjX0h4Dlkycc1edvOUsc
dcCoDCmpkkimricI4rd8/7qsBa7gzKKkrgMSb8VFCsflpse+r5vOEChIu4yQTVs+zMu28UTQIAzL
i2ETuCi0O50lh91xSoUW1t+6u62NnA8fyVtR58X4RJqoT56NsTvmiJC1sZTAyjDa+0IokZnW6+14
AXesYBIDyEOsahUQMlmfABM2gMqG3Rel9SupTCdOu7QBeYlnOGoM1n8S/BocVpOJIAOv1aY3IjTw
dSBEiDQKT/LKxw01KjVHxvNswPe9lQbCrkLJiOc9oz2Hjn+Cy6nrriH5wWl2I0/QW2Nh87DDeM5C
yLVsbAvn7f1s8z00+vZlPsiWy4U9vcjCnToF1z1I5EpJnjDA0CY47wTPFBFXM0LvXNAjU3YMxYBA
AJVXGOhyYqrxNZ/vjt8z5DeSrQzd0Le7uQjqYRmOL9GHPSzTjgijvQigcmgQupjl6O3feo7AYqRg
rTqvrNwY+XGD+Ji3SG7CJE8kcPp28CBZnfbcWAjw5241UVwhBuZVztneMN0/j19xSM1sjMsN8/qY
LnvuovDIt+77BuQ7jI/UX1c0i/exkQItkEG4nG6Vw+7rddFjU0MX5Uw6RZ/AYdu7XfEjEsV+FiH4
HWg+ztuiwu/A4GyDwEV8W1a6LoCJU5DWUIYB5J0oeRT/i6RA09wnH46V07HQB0sDH4krlLTu0wM/
fdYjcJ8SzJH8xIqO+tEOUXboJutpNntKluqGmkRPYw8IPwhobWTNvBcDHP1HhLkLMHxUBlqLBmbo
ZIgZXexJH7QS8M0oW1ou7JblYdD4LiGVXX8yjyUyOZZTVvsA/m+My3LWg3fSjPPGDHV+pA4sNgra
0n8nZMldLlnED30jVFY4wcH/28MmMWDRYSY0u0UkJ3iwoNtyVfJcZjqfCLZVCkECnAkTmKxKfn3t
IhkBzy1dOjbyE9vmOQ/R4Yf38KzCLu2Z9r/EPWMcQFrwZMSQM5NeHKflz8kAvTUfB5Kbs8oD4DT+
BXL0hu7l4pDIvPBzzU7dftiKLvN9GgYuPaQhaMcNOGZg/UkAeTXE+gVR7aO08zLPlV0st8e19IUG
ZIJ9raFL3egpkkSfrpHJvdR8EnjsSHtSb1rnmk/79sbSnn2QUYmVXk/ne/lPA7qWgp+UVDL0tqkk
a3UXm6jXTyHslFduJIMdmCD/olIgw+8jurb8y2wCBpJd9kfHR14VdHTyqD+ZskE7MwcOdZp+rNdl
/4CgHsvqmFs3OYeFl+gbij8nUBg9cofQEIGPm4vg1oazR05zUkkR9kqBRJ1WuOcm7dgOiFbpfhhz
ZCyEJ4VBykSE7lUMy6E/pm3zfGdh2DKtS5ikl6ntSn7WpILhSJG26H10wAAlPC+eD5wjUjH/7N+u
/1gLzskEmNSHp5fXFi1H90xs2GJF1uFNO+2W1sX6SD6aIq0XDDP+8R/hYQCUmx9IWNi02EpXqfqn
dJeI2F/nN9WnujYTaw7eA2FmpBh2f2MMok7FAumwY38Gkcd8yUkw19PzvMpg7kokIUOGptgVv1+D
23z8ePAemqnyh6mktGh36RuClVhDNUYOqIRTFjjKMmzunLc2Nx9vHm12D9GrNWdtc7x6hQqtuj38
/qLy6sUwU2Qr9N+vswK9t6nxNfuBTH7RGS2s7i/PLzZgr2Q39vp92NWWwr6zJX1VSXLVorkpsqSp
9qCFvYJiXwLT8V4018PGI5T4kAVA7i9eGjESB6do5mkISWnc21fjkKTGFUnwhZq94OYPh9Fo8ggK
1Dz8ANVNUDrpFROVvvikDWRmanpvuYloiNgiHDPu3LQvU4ouGvaIddLKbDNvnkosXj35CcVnMI1O
xK/hCNmzyKVcoyQtllfzMnZxZCfTWmAyiCUSMP7L7tyXHJ8p6rtZJ+hxli/puS55ocPBWc36UT/m
Yg0mh2VW/3ZubM+ruO7LQkhfpZx66D+IXs55H5vgHCFdXzRBJLpT8zWqWUYgfwtvJBhuAs8WDQfE
bvIcGtVWg1SltJk5W8c9eIVPoQ7KiGYtWsGDv1CTYR8TiZkYgOW5VTFHXAv/vOwPTYlwQBrdWNHi
+OlGZ4jsr1IP9Mcl9Qvw4Tj4TUBjOoTV89o+6w0G4Q4qOaB5r4Ew7lbVXDJjDCf80ChSCJUJqZTz
f9bQNT+ZC7+VzbbVRmg0bZUIResCXWKjMeNIk2Sq0jXkyoQSO3k7cAJL4x4ja12YgMqlgAKO4tgd
ejTicrzigNYGI83T+upCe3+3QzUbU48O19GgKv69+d3ofzlGA+5VCS/DD1GYictOnWZasZelBDJh
Jm6bedRmPgh/XR5Ng2pnIag3Isa/co2hml5j4hEUgl/OeiAQmqyvEQrGX5FUNPi9J0x36asEgZMC
oTskVvG15FosUBpCFtI9Ja9YfAxua9dXsk9XcKIH2dR3GQ0bEKO9FXl3abThlhrtCgv3sAtNukDZ
109waOMTFbweOh3FiXLUV8PZhAsdudSy5q04cto32yB85IDvzFn6oGAOPkzbFmGDM+/rZxoVJukp
IvTaM9kDpdPJCgifDVEzPXfA50TgFTynfCDPT95s0QoiKIhiELGEltH15R/qHNqNaRTa0BpxW3bt
qRujA3TIz75uQWbS8IQBXVBc1AXEBVN9DYT5mZYHhoDLBEM98hd4VkswJbkEOu2fS9QXoUq5JZRl
0Mag3Bd4WDNkyXJPtLrPSzfMzEynmdKIDVPfJ2t5TatkZtivYPAIY5E2ZpXC3QyGuINy7MITJqLu
mu8LwDAmfP0SFk9HaqaUpENmV6TTKJAJ5q13djeebiIkwecdujJ38UJv/jMr05oxjsZ2jBNZuqo+
ntfiY+zm6/19ncpdKMpk762pNgzl153Vu7jWhuAn38bq59+yaot+r7YCtd+fDv4KlpjXnKC529/5
kcDeYDUnSPhmp1oDN6DevZsXA4YWbunPJTSb0/qm5/qcsl40HD+nuiVz8yOU8EGxfqs1drgLCk+5
Go66zwuIciNDDHzarwfR3Thvwmvg6EgmQIifTmo6FfudNWJMyR7mjcYUzBhTEiHVqTpHDhf3e2mA
/zq+AIF1funlYVSCc4ijFzuFEzk7UW3vaLqNg6qvqbnUAos1ZwjhvW+ziX4LM5FX9VDM8c2Jz0wf
WG4Ns9Fc1K3j9BDblrLzLtc/Npue54/CeKWL5eEcdH4bD41lZy5+Ij6fi90qlw1t03lQ8WYADkgu
OqyhSdWpPNMNN1iPoUMnptdrLQoW+Kz1mWiUVmg62W7Ma3YJhma5ri55Z0vJcHL9+ZglGAteyyPI
Defw2veKVmc2MQfNKUq+1kjq4TA8xswla5JAT16g3qFvIFAdjoQHRi1v8aN+SVCqQ611qzSZ3OxP
MOLuYs7cDQ4FGrlwlAT2ygQoyc0lcEsekXouzgZRnZg9rEExigAZp/vYO9oT4Q26j/+X8sJg/EYA
WaSBXB1LpDuTLBjbQoAvZdH1YJJnNpy3jI/PL9qJBTk5WY5vMqfQ9knJsoQU4PIFa0fyP9Q1CjGq
FxH5if9EnED0X9kZ1W27nEdgoN10aeT+17a8WnLvLOKv2SwvC88j3EOI3I0O6AG8oUCFad2C2LEd
is/rnfGCWjz9TKUs8JhCBv9zjNumAi7RqD5iCcx4eUi5D98nCwcs8iSPgUmL/CiF4TS8OrSkOqIR
E/UXAlkyfQ4Y6xuqqi6JWAGJTFy23XifC9bHM+uJPR0vgF+vvUpezAW/2VV3gL5EFlrWDnK2cxA7
ud96gUu18n/5B2pBbe1iUcYrz7GooeQCyUPuKl/bpkOTkyrp+0g/ULGNDRHTAyzbpY8TEtf2cJ0Q
1YAJZ9t4Ut0nlDJVZQcEHcXmY/1ULnoPURB77SCf6Lfu1/jmTprErnzZD3+nTjuxRw8Ly5ucGLv3
sZvVH+sKNjoVv4gGKvDNgqGZKkIC26fgyNBPKr6XC/V6eEOvqE5In57rYQaWJe7hcWUcy1ng2NYN
uLzLwpynEBjCSXojVMlt/uq6efS3KLD5W02UDKOp2sIDYEVVqvy96z+sEJTysYtMSuBXiAE9aeoe
HLMcatiChUYM8LjnQWJN8l/reABEoLerXYdxhkcI+bb6DoKlH/oUyTj60HiL13hrSX+G6gJKZzds
ry040/JxMRG9EUAmoCiB7bWGIZQPF6j1RXuxgBMLmcIR/2UhEiGAvBFFPUbuE0bJHpY7ZWORPmX8
0fkBy1B5GzpcR8PsxOaF9vWi2JPXYf5Y7KrZo9dycRzaXHdNPCtaOaGZAne7lUsFK3knAtfnQYh8
CZWumHy8L7m/eN1p2f4uY2LVhTpWtF9y+QQNYcbkKaH3CainSvGE5AifqUi7QZH8JE0oy+zygh0P
FoMSxc0SjJ3PINSVTBHFvsFaALXGwtNYj49Atk5peIdl+uN8/o3Bvt6wFzSLEpfz072gBnGhVe9d
5yIGLDN6V1XYqT/nTtEVATDBZTymkGOU6+Qid1zTficzlOEZLg5CSFbD+WjaAfqmv9Dn3J2SkZPY
hCa3JTJMOQ31J8rj79/UMShX22hhydE++IjWpAa61x8MYic+vaLSrCv3WNiEqCzS8e7R6CFhCulp
Ho49hvB8ubfgjeB3S/RYVLA6wN+T6jt9diUXVYf9kDRbQYByLVOGaXAj7a8B9CSBr2PLipbInimU
bbKUj5NW47cnslIbXqrQtHI+omFhh/3DTNQOefcIJ6CFvXdQSILFRKxJbtzp8Yil61Zi9AEjnC9S
2/MNIpDPCENWTICRQnUXJJKeWlZVuPqC2yNOMO8P4XnpXzegtv8x2VW8wP+peCxdpVlypvym54Zs
CA0jbU6Jad97qZzruK2u3qqtH66Nn+spKcQki+h518LFXa+J0VqLgllzy3fUxl2s/xdH9EQxsoZh
jEtoGuR7H5i+X9qHWWNW/3ddkyQmldMAMz497Dph89zP+0KDJud+DguH7nrj8E/RyiqF5WMCvD1C
CkejxqWRTUeYyE+7ENVcjOggDNwrLpOvaAihymaHqRG+TbbSUooETGOU5ruVlosZc+Ojc4ZAEPZk
IrfGyrJgxKOjeCM8gHwAWkTT95lMsIEsQIMwMSZ1b56eA2YfEvVoh79ubql0hcu+HURlgxejbFfw
N+q2+3sNr5/OUtq9vbXzpX12gNKx/swMJsFCyhP9YAnL7xMrvT3mh8EycfijZHYz1BTAkwojVfa+
zw18NX7sUOBMTe/qGGOoaQXBzwRGBpSk+MwgSYgfh6RRKGqrA8r8NYyQAaJTfr4fZE71mn+rDF51
PFGvPnawWeHlcc0zBeeZ1FGCMCPySbdcPb770k/zGo+cJsC3GZc3YpCTTL+6wgio56d9/US6oYXJ
EYE2HtuF3gRVSdy7m53sU7pnpor0bKC5bLUZtcA3lxK8Q+PbFLoyens7mnYDXCMh092mz48YENa9
YwAWwpEEsdLNmR9WrT/sXvvslKWt/EaYCWnGikDExmVro8fyYwiV6GYOYms0ETWmTcFIDeEyqZMX
7CPPmCgtQVYY1r+JcqJ40M6W2cCAReuDmqYTTVjV/XRVI8LUfbxHMTO1sNGpVIF7Qfwku6hYW5zz
ZODzZJBiGk/Bkx3QW0rOK9PpDeH8IGX7tVQ+btImvMDvZNw88yrV+t+bN2urBAOmSQVO18ppiHvF
/8PC59SQ2Ebw4Xy3Srtr7nhb4J+kmWowSW2NU67FV7Yv18i9rl56fT+lVCwJ1fVX7HDPdcCsrTzx
7nZPdON1hXXfqJOFGmdwuny8QOcuptGApExlwmSs22w1I5E98GjZBSBiTp1QN1hg0jC2X2rn8o1b
5USl97szYnzQYCcaE4gstlVkA5NncvbQ4oNmALKFK9oD6K7eLI0Ws7oALASGCudg7tymFbgBXncY
5RplgXL4wBLighixUMRpilvwJNGh9+bkaDj5EsPiTNe9awdzjUSP6Mgy/9SPV5je5ZTqSjAJsjZt
y1tfA0Rix/rXCdoeRU8Vhlw38wiQS/ETIrRsuaSpE7b0+wJ0lHu7f40Aow9G/C06537BlPWiamXM
Qx1BKM0hcC86cfo6h5FacpwzLp9Y8ZZX2jpY91fKbJrelscVCV5b2t+VnWfFX/s6E7/X7SILZwwt
Cle4BPH1NfubuQV0yt9Y75EPds/brs+Mnxk/ic6TCKd6PaN4qYliFVsZ+LvAbMF97BbvMaw02cd5
Rv1J1z0FU7Xtht9HMNe/rr+Ep58aarYCZHzx+ePVBnAbOQPtroauwvI/vKVqIdcDsiuP1DEtwGRk
EhZZyB/3lDHiroEm2ny1of2pXW5zv6CK/Ldvj75bHZWlVJ4gYMQlO/Hw2kC08ji7fTKiCMD9fOw5
5fZNyLKvPNxxHZwefG2QtrBm8heat7QoOwHzdXvVCp8oQXty8iAC9vSeN3MofTZnegkI816FimLX
HwUP5yPhzVyKgID63N/sQaG5uam8Bnn1eHJHU8PNd4R3SQ8SCrQdNiymuo33msvnZd0NMuwpZFVq
y0QEq3pTeSJDyZBbwdfaaeUE74wrG7QY07qXNQL5qO6WsnpRWzGpXbnZalHcZmVSAh4MOFkCi0ZW
JqMBcWnIU9ItIo1IWcNXVUMO+pSKz5fRLf+PB/Q59sUyHAUMMvmDwWazZkM2kv8PLKxPamQDGIkI
EIbJvY4Eh5MhBH4Vgx6HTc24tLZwYp6wYMpwtMiRNmhhWb5YDc0xIuGXuvb/gh763QUEvjyTJ4Nj
SHG3qUS1EtxKVefVcmbEqoaKjDgRy5iGOJ+X2F5xKyv4mhxF6EQ0ceta+ghOJXwhuAu4koygMghy
TFJxAziLbqpVgTNgYkNCzN7xaVfyEnw/XwHfFOjz06kX//ZD1FLaU5vpYazmGimEc5IXdH5iEiYg
3V/+cTBPoAP6koCalO57PVv4+pE0SXolK3kjjUaKsPQ4rL62ijhYHF0RZtnhDp477pdMgytWmFIq
jmHeUgjI803E++M8Pbw+BBXId9z9+ONTP9iWOqRzHTEKK+6fB1rbomCLv24CBxHo+bikeav5g2PT
ob+9xH7PyerSbYL7SG1cs5ou9DwJ41OCFiOomsWAdmg3//iFIUOYffysydmyQ8aWmXfHNoepr346
+MgGXolvxs+gsuPEMD/68wJwS5gS1FCIRfAltPbCsS1j9Mlgq7QM0ENhgIPltZpGMufHKa8V+0/v
44FjWTkUxt9t6FtGq9Uc6DDcj9QypB2c9vKcp+U/QqpzghmU+NvcwuLm4eTDn/nJrZrCVbtB0mxP
8gFGG6IrBxSodf1RR0FCbUV8cNNO5sPbAJRotSl4pE1rAGyAaGU44EfzhBq5jVKdosvaQeIdmNoD
Wk9mDU19OuZxgxNhB+1zUWflzERYKkaI9cSNuRvmWIeklKzuNPJRfgcKV92JlAiO7GFyJAMyQoed
yv+l85EAc8K7azmHMoDM4A4dzf9gHdtCTM6Id6XGOFu8w859fLCH2qBgMhb+AKR6kgoCS0AwoGD8
9ZUycjyBtcCFK8uLumKG/OghCI+3zT4vxtAltvfsPzDDfNWGjDfgDcSq8DkMTYfr37pmlYEHUanj
RqB/5sjnav7Lh8U21NG7mew20m659dbEC4LVPQR3j8l56mvDwjJABz03AEgzbfVE24GRKMVZ1N6q
A2ER93LhY35eT1Uv1+LXK5ARQoa4RHq/cnHHjh2zi1YEvRzhEiA0ABfz9zJa3BnWOCQuFTcfiU85
GBwom01sglRMI1A/26PbIXDi+RzFkwWYqPQ6hwmP3gpkfq0eRUn7kRb4BJ267b7RX4u+9oThadzj
IqydyXJp7V+nObMCbFQ2+FSMTjUKD4PRya5NnjyN5cSqtkYBL+7ny8ad+FVwdLx+UcOAJrWcc2M5
dItkpsVWJAGjBA0vG9rbZNRsdn8YJ3Bahi2RBasWIqzjCGLrKeuwTkuRi7mPYv32CAXr3Bf74QKn
l9Loh3N8152QuzNYWOc5Zh7Ud5vybWu8JgGRbxQc0MpuGdAV2e67t9Z+5uu1FgyVGAfInbCvJyyG
I1eQo4rgK8piIsuR3AAC3B5RcQ+jvWTFN+L/NrEkPHdGv0MrP/eO73Y2jIa5I0agGSO3K+kBtDcN
DGUKs5VDMu0PD8tcOVwGSRnifSk7n985Y+X9cFnUsx9/9Zc8K2KVFgVnoHqxkGGHyJTjcujolGPo
KJVF12B9DuabUKjzCGf0psfnMVuy0umtwylLETTK/2W6N3xHhNrjpfpC3dLhAMDHCQHjtZOZr3ml
xDYM8Xc1D6uVnJ4RJ4ivUi3NF6Qrh41ITzNBy6gQI4k/wG3Q4JN1NoZsOeWRijpKqfxs3Jm3YPGt
FlWCZc938ACxjJRAdDTf3RnTPlcmT/hhdkXLRYkaTS3bYFPcAbtspwpq0oE+IT5bo0RDUf8KSD99
7iUbcmYz9VJjA8lUT8YUoxzTo/jvKhv8DzvaTQMHIqAZxJIKTwKKyYlD4qpn+PLCZgDK3oDqgSX4
r6s0Iv3P/DAJmO87IoJlwyJg6B+4rL3K/25/f9nxMwqctf9MhkAt0HtdXMCMedIWdHALU4uNSYIu
Emf6th1SBMN8hqt4wSTLP2c7XZF+L1cazZz9TiDgk08qp0R95YB8M7DIqIGzqtkNWb6SB22dRUzv
6KR2tHbt4Xyg/19GWubFsJ4eTM0EL/RX6Pqo0ll0naLRltYtTX0AHFF2L+/r8lR2m9vwzuLFReCE
CjdG/Fnp3v2wYBLw58qBrEub0qiH+nm1opRFDknTEO6hZdxUFBZKqgNViUxy47LSBeapvHWHwHBd
rJ/+KKoGB3wBPEcIEbrVNMQKBmDSEGrjnQcnYoJVXu5axZdWYPAD8IV7ap3FXRyFXI3cop0E7f+3
382tAqGTCaQG5/5HGgw9w/koOb+3OU+vPbgg2l0tRnyDw8IQcDWsxIu/j/0Z4jyyQ+vtdbUYgh3f
reuVUf1DnYJ6T/qwhDrRDZvKU1SPXwqaCJeiwRaYhA3/3XBE5Awf9xSMiVecUCZrWUtnzJrw2dvT
PUj40kk8BF1W9lon1itlZMroYPq0lQpxS2m6+ORA1pOWAPSpSU+9yeprY1s3ICRNAdyAi4Sk3cf3
QXY0wV3H0zaQo229Rpb8gEPsF8yeALOM+j+RnTA7QR2pMaGx9wUbi1Whq0VcVniSrpV+ll7kYJ/9
BATE7qKk555UWloZwzWsMLU5ADisvjlXl+ukp9tacrCsh+hOvakUQCVlgPYlzZVPXmWU4yzVm7gn
xq3Gz1CSKWaB86MunrxstWkBXkUKwv0De9AF5kbYQTFxI3OgkOBv8+UOoRHR8Dt8qBSqMrnAH8rg
Cj9vruPTExuvGLesQC1y+VkU2yHQaokPnWZOHVdwOhIz8UJMHGq2Hu1pKiLoWELqUItwq9LYs+mY
jJzuYfEuetuCePAf1XE78mgxtRqgJOwymb3qCrh4Rftfs1cdjKVv9WhOArKX17dz73oSjnaNu0S/
namaOIf6P/NzXKwCMqIJwWk7Dk2mgmBpWpYT6E7rnv2UNGJ99mbQ3mv1Zl68INiaoC3hgm8pfnCR
BbFIB3qsCTpywoZI9LRot4I0p8Jip9RgJo54AHf8Ol9pjrvyc5RB6HlIdPHhQrpL/IUCMrLDJoij
6eHJKt7e7YkZdy4lKezalegtfpmlKO/oUeGmqgt9WrC/ry8oKwWMMp5ytR6vgp0Nk/wXxuTKgAbc
nkiLd5nOo1Y7Xi9C5n9gAEkHrG4dRm0/Tk6zsX/cscjhH4zSyzBzyPgqt9y9OlE3XUJb8oXgbfFa
VSO7CPEV8oQ5gC6xHVg/XOnt8Vy4tTM9ZfE8euB/Ga0AusCE+Y4tEVMruDnFm70osscTJeZzrPZ7
UZrcD10wO/BVg+ZQGx/umufwpLhQVzjCqTiUrxwM39UXbETnmKc0Hji+u9obOq/7h5L360iXJpGg
pudKhA2Z2DZHcS/jrtywF+Mit1dzPv113Z8/1zz+G/OW/oRU7z/9A4qssV1+Fo5HLz8EgrYL1gqF
TLZqstovLUCO5rNvok8gHSnRyzbdCFfHqtu8M6C/cAv4pho9zhQqFNwJ/go1/1DqMv65UIpp6qZN
Qd2PeKwy05kCkGC9krVvNN+KeeIsAGBtEKTbcw7SX3XrHxND+FH8zcq6lfkFwqaQSCXd5pbu1KrQ
3nS8XfHAsJoFCrYDA9DOHHstDrifu2Je8ESps8lCaLadl8X24SszHbUesodeJ3rl3rljUlroIKvb
ldJY6sDPRMNhf5oPfq3UE4F/BKH/bAnJuwWVMRNR/l6G1Ka2BjEo5bPJ27qwzqJfJ6wplBDz9eaB
U8TtiE7DfnEwX3iYlTEVvjh3YoB2oyWQKW8rrKhOpkPMoYVOC0uyiOmM+wO8exv1ucELPPcEJAXP
LlIYatYsbBogOm45r09BGAoyCoK8KNfu8EhZniIm9mF8ND8CqW9Y3btLcvL1sdEesHRpGx1mKM6S
YQ+sFOol+GaxQ9ADQ2JtEcFV3EVb/5/Sf0mMYVU0nFU/rEc19rmfHcEAdsweXooBm+fClbhFTfC5
dQZmOVXT7nlQCfzIUIotcriGRw9URCD13Ryxcy/g+6H8dAouwx4XGVzwihWFIC6BJDkRTcHJX9+8
72WqiCF8E19DxnGSsryp0devOk3t4WQ6SwKjBHssrUQpCkHyeRt3dK29DCpEgsRkl8u4s/IdhgJz
Hbrpik6xRSJCb+GfS0+5lrxCCAkuweiAaqdzgA26fkually099v9S/lJhra63d01N0bH36B2HYHD
LDOalfUb3d69tLq81mgQciAwNo8iIwc7NFKPhBAMNew2flNkk5KdfjgzVumbW/rimCF3LhyZYCwr
FNlwg9i1rIctRC2pBwt5bKo0sXtHbQASn6hl/4Pit8BfCJOwAS62VcNDywSonUYey28etekA/y8K
zi9sR0Fx+JPX9zJGs5tvMfi8mGNPPczdZWlV2XsCEi7odl5EtF0fr9CvNULlqJbmZ25SGE1Gegbz
86BCzID2TZmGEX5g05Il6dbvrG8C/0w6KsXpNiyTP4MbqoQ57ctXAOJUM69FyecM/wPgrbbyWWZW
M8mMSdAHj3Ya4XiRibH93A1Q08UMfyPzSgB2CFEcjardkNvz847dwFkVulA7PwmeKML1oqtpIjvR
g/ewOFtpiWCNk3x6rFKUzvAxRI+91pcxsPxKKLcyf9hdtN3CcIFgxLpgvsVzgXWOraF4TiqUwaUs
Q29BLtVuDpP2d/+Ndwoq7jxDkKhufAIJmKrz/TDspKuoLI87+WbXSAJnelHXTl80neduKU1o/cAp
xPgRP1T8iVxeeHF+QV0x6gt+MMCuAKWQCdJfJabz3ZDTGkELzv7CTyNZwaCCozaPQ0cl71FRe7Nm
z2y5Lq4lFZvb81tcuJAQoixF5259bYaWyRYQNKuQPomohsx9Fr0NnjFxnLguSNPk7dTMKV/sd/3U
GJL5KaAyFUvvHiBHoFvvUvhb2jfnc2ojA6deMJBC3KWt8FURi+Z5cfyPGeEzQ519hMLXVMlWsW9W
UbSu/T5C0n5sx0hIa8VsnReAU8sYKaj/d3gLcFjXa0OFarByXjbfKb9PvvDBcyXm2amWNvG9XEFE
GGogHZK7Z2fGm4hUjJ7Jasf7jDVHCoqrJtgzAbuBG/YbpBfUPjl20htJinQ2V5m6z+PkIiVz3cZs
3iKpJlKl4m4n5xEblcjJ51fEOvFORVZxLDZ8WM8eh5HOOHko0uevEVmKtUVcTyj/LYgE1wx27ScT
qAX0qjUHmcFfkAkHAHV238y2mk5dWKFjBgI2EzvAlu+UcJeLc57wz3q0muDXRA9e5eDEpD/vWc4a
tV9ik/wTjpv7GHP8cIon+xKF4zf0DkFoN3DZY7HSXQlnT2+v6RfMsNzapZMz2Ff616K/xyU7kSNx
xdd6+XVxILFp+N5j4B8Bk1LKxjZFMbh2IDLznWu0D9qW2vKbXVPWVhPw/Urw6D2wPZAps8OM5T3k
LSb8kWzA7SdLctQHPNi8i7aKfnH6e7qBbXr1kLAEuvMkenj1WMF9sHIJaWHZBExRUQYIKRiLdSaV
SbvqXY2LkohxMol++qWQWD6CNhf1tGwCZXQndGu+1n4Ol+CHJq3UbnTkPckzkft1JnfgL5+Ngzds
fpqytIQD5xA1yenwpjJuCvBuxDbf/uumrOuyXkOZib7s9Z8JiBekvf94J2quiMi5B58pWjwtqFDw
qIymL5OFO6sypY0HUXjVja39vufu6aIkmp997YeGWO8pXJoJu3GaC5gRcnFVKAAX170DKxbu2U0A
oixSPiVFqnF87jdvytoCW8PpoK9YFbjyunG/NxbK9oqZrt5+EbjiUQyEIhGBwaKynjjrIEuGCJ+9
dKwLDpHrzT61ZScRZti/UEIp2wVmMUWZnbTgTdv50zxX4qZbY0l1uNPlAgML2BneFMtg42Qa3K4U
uCYpZhW8DC7GOElU2YKgpyvQLkiFozHjD+DRg98kPiOjM7vUPk701aoU4l7E8ryUYFZlMtE7VIa+
Uq5pFm431PNGPwYa8KBHZu16GpAL3GBkAmZCmBdbSknHQsmvyub8E8P0jBzFuzMFmmTvxvZF1pse
xGrTb5lZC4As9HtTrMYOvq6UCMS5fb4Rvc7Altip4MVTrCCac5AVdJAcc4N462V9WankVw8jr1Ug
UWD7VSYbyCGHjV0UELDWxfJUMTI/EPPqOEPo2qxx9LtzewfTkcr5mI0PYXHz/YQ5HUFdd/yYt1tp
1GINi65gWVdsZ5RB3IsFv7Bh21mbf4R2edWWbz+IOeMlbJauyXpFN+1gZI5wQTQS5Que4JOhrKUG
XiXmekG1Ch7K+gk3HKAhwdC5OsA86gyo6Ibgk4KmXvewCoMKy480f0KNc7lcZ9gRzxjXlLo6aXnT
ADU9DyFmZNoWP8QmxuVhAppt/5WFUYjk2Y0qY5jQfhkky+9lIX1+aV1qfkhepvVhhYV8dkJKDqmS
wYh9fTBOZgwSFq2hg+3g2aLGlSVdFdgZnPkKCxP8zTl66V0eElYcWG0gDauRjOypCgfKdpmpc/bg
LIg2ylGGVwKUSKEX2tPnEOBipAChIEGLG2yYgyVV2Ox39yX/tmhVfm9SiJwcMmRRVQyVskMT1Dh6
sjduwRYBV6xT4JmdxtHpVNM00w3HzFZO0DNeBgEV/hQVib8OjUYWp9aRaQTzqfEyqjydiTQnPZoz
rygh1dtKMqx7jVWIq2OSauAHTYElLhPzCqFikDXTSxkKdo8Si6P8Jr/VPFDwZ9up9w8mHupXiV8W
bITiT8WDoTphNhJsFs2ZEfNI2kqUr7XLck2VvPqrxDutU4mM0RRccaD1BvPqgxh7qkAC7pZ9BMdt
qmFLEhBygv/kyiIhc/CJkazhQzYXmQdyW5zsZK8F07rGWxucXdH6nwbjTUXUpJv8YXjML8wq/usK
7APfod5qNLd5iEtezDVYYAfuJVZMKEeTjL8Pn7WzU/lTw4NUmFXeu5unPaCXDP5p2on8pwQr35pW
4sDIGguR5kqEYTJdrCDxkSjBPMBO6DDFcZ8VTdhikwab1q2vp8spNkI2HVcU0BAD3zAas22IuG9R
4S7banbNgcPLkMHknRVyYVEoOEdicl0lzMz53l33Ys44d1HWvN+wlJGntgSdyMc5C8SaA/w0WIWD
RXVMv1cpP/BTGoIKOCT/dOCEHPUsXWM/zgbQE8Yon0QC2ZsAFf06dPWHOfwJhDJJzkjXmwWcVHLW
sCKnBozh/BfwMeU5n0FeIuKXCo1dqshbnN1uCFqT6YDGqaSqrv0HeC2gZmYpByqP8VHSpVxCDHjL
E1egkrRJTPEaw86PY/ZaXB3MHexWVytw1yiteaokiI21kxGKiC/M/AVTMo2Ucb6SJ7C9ybOPioB9
V53e1XYVBwHBfEd+ailcNvIuy5RC7btB+cqn9Bk6K6xao1BPQwHZcfXuGxudCF2yC1sNygs1rOWp
MYOLxLV4wyDS3npfTbU3eub0Qy06LGcWCepMrWhR9/4djR7N5g3DDj6vTMItOZgE6Lj9HWzZ1QpD
jmVF7Dep1u8OqrL5dV2mBu/FCpydrEsiEKlr3KUqx1QI3EGXOUXuDdi1Tt5F36VJWXk997R6ph2O
eQxmMmGX4dZMHw9+Ii8WN2o+0k7WHc87ftbYNNPkfedaX4xAhJbBEwlWEDHHxGbfvLGszrda0KkD
2lk1W6imU94LWdD68tL++JG1G9eDkZw83JjSko5Hpsbv6ntxsgJgUTaZTN+IYS8U5wbNfSYCfG54
SO3ikBiqjvBzMHmSITuPNiV/wWq+sp7M0bNZJ8FuE0EbZUqxp0BY3BHIMv58FpmWkMWAHfWAu4f4
aMndLMJP5Elp4uPSlNPW7+nfCqMHXmKliTeouxKqIV3eoMPZtb6q4yiJUaeZvjzb5haJDWcSDqsx
wMVbvn8zSQinMnBOealeYjbgnll5czOzQkghOEAIds0rjLsknyIaHk83Oz314DG49lD2/0UlnpMZ
zIoZzvHmVQyR35nS1oEUaeFUBNDDxN2EQtG9usSrQPucIj+waQeCGH2arOB1DnvPwssJKKigdQnj
D15BhenumQ0ZRL/VVzVano4km37rWuUB1VTwt7xIDrp1nSszbkJn2mhv5Kwbws17LgylaVS2ta57
dnPqI6KbvDdek+QvDdbc/G85PN7WrtF6jaRdWHV8AlLzEngAAurfeyHAj2ArwMybXMO277EXldQE
EIxLdxJXP/N3i6245Z/ZLSHfoYdNzEl4zu39VxOWl3j4CMG/w7RhIiD1zJBox9ME3vFvkUjYwDAN
Ea6Ied14xxPq0gClwXt5GTnHrv/34p5ryvW3H9mfm6VKNnvKO5EWKz9+3bts3m2QBH3on1Uec5S6
k7akG2mz8unNUIv/OVePCX2RWw8K7cz9Ef0gPUzEgszsMkvsiNno38t5194AuNChlYgvzmJzlkvr
s/y6G4sWQGkBLRTf8bOCyO72ArlD1RqB5d6tXN4Q63r4BV0/AZcJFIziq+VJdMSmodQ0Iahapi1q
AYeSF459i8vHrWvaOMNUXrxpFKYCPtZp3Ln9MqJyy5DxOOKMw16aHba2wyPTlGfG4+8aIfoz70G6
7dy1nh8gPWj3Za/+zNfi//KN5Aza1XbPNwXPyHCLsih7Rze3LwbSwsEEoY3bv4YN78N/8cZPRcnI
iheB3nC6fu4ci3KCj3Ux8f8WVWz7/XPt86Nij8lZ7RxQow8ElLsS9J9zWCi07ERWKNp5x+EXIRnx
QFz5vfGziv/bUqlgfL8AvdBWob9NgEIlHOqQQgvdLOdDt6+MDqJru5SzMzM343zckDih/lahQI0J
vpqt0jL4EISgo6Xut4avVCUS0A8JCEZgHtSHb6N4yhd4sF+qDouLfxNFtpNkG5+PNICcmp3K77LU
z0V4a5GD3BENdevH0SeU1uSlRaCCx+5XG4AFGAlalIWuKSmjMDBvtCjOSQxr95MZOLAp9kPxnYQv
CETKafLj12OrV4mRHHfOhN8lLxotWMZqw5/jHETVnSN/l2tZ4wQmMpzixHdGdXeReE5Yc5jGUzDt
mK+h579LiGkgyUMsPs2k7rpsKxiMlHAsQgR08FDHh/4gUyHnK5NCEvONAERlDOaCepBNqp261d9s
hSG0ikpXNaGZ6P2XxeCLLzDqLV605pE27ShuKiE4xQEFanHJCrrxBIthBLhtrOgvL7civNBB9tXs
7xW4An3MV7k7AhAcC9ZPil6AtejyAP6BOBjGYDRhKwLtcoRv7JvnshKAlxpLpI74+RPzd5/uUytz
mPiiIjAIwXpG3PnJr0Eyi1nt+w56PgLCiMqYt9kqPvyPMTCnGj19cBLxZkURdddhwYDISldWXaAr
5euGIeUW4dKSgzEWcjnbwM1efPUSXZV79qEAzDhsndrm+kDLK1sfGf7gDfP2bbrWAOC7NVY6Q4Of
LOSiNk5ZdFNb73iW11bRXLz2Nl3eT+oLUMGd7T/veHjmCpCaLvkr2GEAsPzeWzK+V1S4uARu1jH8
RvkUejpSZaAyiBZ+ZiY01nk7TR1MJnqz1Fh4U0iDNINUSKSkDltahFemqS1kE0NA/OureR/mOoDM
GlMhB6Pvvs1B/wGZc/EwgExPwjxopU8u3qj1TMSkSvK76LF3/zi8d9Wn9uQyMcj6M/Vdv3UjQeUF
5vvAhjHVjY+73EVdVaPJ+mFQWeoRQ0CrTEildyf1QZRjdAi0JFBiKT8AKIpW+CZJtdUPWWcQrxD+
D4SDox9pF4/sI7NUfsJ9uBj/uyjX5YXqwJAlemwC4+HflkhkEeqpH4rlnIOAqsTkkHUJYS06YtA8
axiU6eAAh2Qu/ryAzxMvk9jrn1Fq/+2LPXxGOBs4NfitXit5xBqh3xj9wwoVBMZZQQ2LtV1CcAbR
DtdGIMfXSXZAlbr1BVGUGeMlHXvZ5+rnY9mB1zJBhDp9y22r9I5ZXJVm1DXHgoTEYyDXTmLabOBy
TDAiIltQdkhXVdmu3sOS+CP1SYsRJtMyYYygxJ36KS8khzpJ1FMJZ0XkwaNWmfrflhhT/y79DVVK
VU8evQsCxxV+GJAOzWAxra/2vlutCNXpClSNUM7AICGIOBPc6JHswuyh3Ums7ItDYcOn1UAtNOkr
/4OQy6wMDQ/YLL4/Yo9rB9wxf1KNfRGWL7vKWS4UHedoXzE7qtDbW56Sx3V08O1vhU5XsLvTVF7M
vbYJuKOYoBZsm2Cda1Cry/69SZUhcvVCNbbNgXQUrSBqKcTlnhLv6D2ffiUsYbR7BH6QJhhPFVTn
6jKdcPuiMy/E2C8EoyP2ES7KajX2j3+IgplTE9ZkVh6oWhX3HgMMn94BwdJsXLwiVkZ+J+2Cs/6/
6a3WZLngowqELW5SdiaLd8BHPVV/2frw8ZzUYmBuOeiW9dxwjqKpLYlbu6k3XUBNn0dXJDSEDalH
3Cp3C4u/kU2hBmFAFnpaNxmmfA0s9L6UG9CEuZafkfyxR+JIaLemVAHQMFdeFhBcETKCiHDOmHXR
Dj86BTVKaULopm39spN3+RW/75ybk2J8RFyQAdzPDzZUmGAl8sk0Qm4tIDPufd9TmyAP5KrjsR1q
aH34VhSnSYThmw9ffB/CtWy+DvkCE55X+07V2am7EMODIqe3fwbpik0JPRc=
`pragma protect end_protected
