// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:42 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QxMQ6DJZacULuxKF+YDgpqeou1omd/lXsY8HHXhwBgxbqSpvRoGtNkDpqq0d662o
X6haNAIp+AiLSLUvqKvHgPryGa4Q0q2LhwrGTeQLHwx69dAl6Fa71sJCiMOBTeGu
ke75fqTRCOtVwsWXGLwbZmVsMMAe9U0UYBFna0cYvRc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 58832)
hVO9Q38tJqn6PloNSvRQMAmD0Y382uWMlGu5iQrGDg+saLZmDwbNPGl36eYZFq3M
BbQeuYwbSimcUYLtSfyRKqdMQRqOzY7WPHQmoBJnOX6QgWTHoCR7b1EIIgNMTqsc
JOtWcKo0wNixRS/SGBEXluzftyBQgSYkAnmcgWcCpD+VRefLVfqVl6+4GXz/ZOlh
WOCHNw9QtjLHZ9GMiTYsAyAC7GyUytpOrKx/WhStX2D3FxQ0Ld/IJbRG2rsTlBdr
Shh/TD8cg4hlFippmtGIz8kWQJWtl56kb5g1Z6LBaH8DUnKDK9WiGZbRrPyASmXF
YgP0znDO425V8uPDVqnjU5u4aF15bnsKAIfKb9QUE8agkobS7kIHyvF/NB1pPMjG
1GUs4LukT51YRB4Jeun8pH8E71rgHekk6LVwz8X/3TRQY0/HFK3Ggidik5KXo/EX
7psA7wnCAH/SjKhgV+mornjE1sg2nC+NxN0XmaSex2Wm3bJsFnlgLDfBXjJ3mOr2
drwnks6/g4EfxUa7CPdHj6rBYx2p+zZdkJyp8et9M99C7gA6e9Pay1yyr0CAWDBy
3aK4WL+PY/gl7vRMA2eq2Q+oSiQtIkU8D9Da4/cWIGo4iS0xoiubIHOO9CF5vJoh
oRcTAv/jmbiZJxfeHtjm4eoXjCW3Qf84qDPrEMCnaTCqLgZm9mPJGa8nIJt/x0n5
XCEgTrxUFhO2KAD/l36uorGyM3h451s/hlpZlRKa+AyARmKSnQWCSnF45UPu0LFG
/RxJOcTbDJZNWzmRGeyQ+Sg7hVWt0pktLu9jtgeELvWbMg3C0XMaToc8YR7jwd1d
BW/K+IutnKftUnUvvOxMmGEaaOa1DSUe5fE8pqcVj7R4sS6uyhQSI4fcbzbujQuO
hlTXBRozj6MOGFWhjVB4S27OHyFnE5SnoL2jC9Tcj5ZPQ7P1/GJj4aBPq26MNROZ
J5iNGnQEMCxAw4oBlea/eQh9AnNqJlC9hiE5nJkbV7wFAvCY8f27DTfBdjyHM3ZP
GmzBoJtmvL0ipFjdu4YgQRrvReKCs2ongMwoyrUCmYzMfNF4dq9+qIr9CnV8k72x
kQslCyEpmVKeT83zPj2f2JztG+tlC59ZyXNEjSRPPIiHxAcz13YnLq4NtUcKsFwm
HTC+W9oWwEfVI5KsxoGiJtLBSKitRnjsxbEx2O0ZqX/ZIj3I3CsINUY9yak5i81y
ndClwWCwFpujA37dpzPP7EqMnj+6oKZPN60saibcrGkw3D5wdu1udHZQkCEOw4HA
GnIS/9i+zm05Ty1gzb0u62+WI6yB47+kt1YXl3wKzfPArDYKfKg/MLjPZcE/kieY
A2+ViSqv78vYnp/7TYl9BtcOOWy4egsi/tozJPxgZQ1zVQfktvJgyBiD16FGgYjv
Qare5LnWEZ1ByQGFrQ949HQ1SG01Yx7mTRKW+1axVSLIEnUBp7UrMQTark54qF5e
47H1JDHqF3p/3jc6FRIuOfJTuUz3gJ1Qu0py9fOMVK6/9XgUT16kuRWPeWyj6f9E
pIZjta3iDVBa7EeTpwVvq0mAnAqKtpXaLo3kcm9oC9zAOyaTFNA4m52IqXjQucnx
kb7Nz2q/7hYnNJUn/vBv8geJH6VJQDtO2Tv0zA1kbC5OV//NsXSbBVXeMlE1WoEi
vdEzAlfu+9O6vLH5Td+LENPCzoTvZE+ORDX4jX+k0IMxnIeTD+LZgFZ9q5i4+8SS
McuOS0Us/oOR5BIrZ2rRSUe4DOGfMkNPEl2quVMvt/ZuUJZxCWE01qOZeYs5Kdjy
XpFdl7WjZpZqUnyUk2dhqlhkVT7nb7DlrDPNIxlX6pgSGOBpBsYo62J/CLqd+NIN
FgAWChSj7IYMkyp3Sy06chnoslkOoOmbPbO5JRRZ5McOW2YBLAOiaYMOT2LArB4I
bTB5XvmEVAOa1KJ3YcYMVuGahuAc6F+amMnUHZJ9b7NR1UJwBE1srNknFUxyRYyg
eObSlPRWEipTcKD48pglFpnB8AJcK9Elr7l7vV1a58CouA9rMFCXTXlfWoyrNZ5w
B6FTmJAegvwjsfKjXfVx9hiccD1fuODWzwbX2TL+loiKK8cf8hpad3kXORy+jIOr
OJ/ZrBKxCqXGWFBKqqkvdVJ3TbMW2aogVLTMH0e4uhQ5Fp/VX9dFbl79hfplXfjy
4kyStkmal0d1Wwj140iFoZILDsm4w/hRGQ66I4OvCjcM5coR4xSzNj6sPFZ/kS5i
ofnUhnXJUBaRH3dawAzaeurtamqT5Vmmss4S1jmc9bixGPJfIszDOpL01ORnssv0
u8VQRF3NlBu15LSEVUVFTmbTAQxyE9/RV31wOfIto+ZvtKqkEygMV+D1aDNwwHwE
40AreID/TFPThUUPsfYOufPKKMPKbrO2R8FX2/hXkgszycbX4dx7uyvxGcL+IKsY
Id4LsprF7hXUmxxCqz6Ir00bfkRS7YXaYeAVjMxuV1APzk2CBO6PXYlLXFleEuO7
S3Vm8B6poeNmBkFpZLZDBhbkoSQ7Z5wtpwsVxwr4fxijm1TSfldrujiQZWdoxH3U
p9iJ7Xf81LxHx3p5+VuuM2ucPf/VcMKVTNNChZjLhqxRLaNU3y6PeYICbS5umFFI
L+L1awdD92BRkAg/cpWUN8xTd0DryMHOAXZUIrbRpJwQ43UngPALA/JRRGm9/iXC
TWU1q4jc8OALho8/aLk837jDNPQfqAAEw6x5tnjXX5ktTyckAUF9eJLPseAcyyXU
px+AwD5sO24zz1hWU7Ef7N9l4YBTMCSEqaYIwVDo514FoGvHLRPz4UsoiMUkaShW
e4ePoq8ok0LpR137fmlq2XiCRdgrN++b5VZB/vluFWlD1VZ1m/6v/qV8LFL5XF3j
PfS0rqhxbwjEwc2t05BA8OY+860fvr9Y1d3O4K+BLJqTZizFL8bdDRcsrL4m1+Y0
a6fymAcnswzdp5PYV7rSaN1PKk9Dpna7hkXI5i1nDcZ+y5HG7qzoW2Y2XjKIGNfJ
mQD+7T8RD2DA7I5ZBKQ8Fbx2KIgxnVkd7sYNoW3hqaR3uUuR9P4T7pDtQM/+hDpY
cDLZTG+rSXayI/5KoZfK96PKthiI/YA6tzo/HcWOp6xWX4wKU7U12IpQdNxMOIXl
fTiDEYJM4/BeHYPQe6oyytqZ9CdaC726Pk7bkDiT+/v+68OWEGyp3T/FUaPyY0WK
DWIPhXggzaAH0GpK4+aH7SnV4Tc9b6p11mEDA1SMWBTb3pzukyxVeZFs10UMIEhd
9q1MY6LMoTmt46H0yZ4/dJft0bIBpoM3d9s7J5XWxisVvwGlwwXvbrdNNSLkI2ez
z5wc2B2f8MPomQsTFB2cQBJ46gsmIAFKk7wP04UvOGGpmE6B/p+5Wyc+CUPor+65
LE/L4HCsWldfArAIfdGZ5wY49IPRnm0WuD/uuOo8cpVOe1iJJZKMn+7xRxZc0Nhy
f4ThjfVd//YfDr59ucRZeG3T3uvP3x+T/xh7fBv5tQzWYPAxbOCm+Etd+yvbOiO3
jbKM1ov2Racv+sM16SGREkQbDHEeqW49AIySqD91pXhNNpY0H+D9Nn2OH3oN6Vjk
JNfUlhMF8JgCO2iyDthc2ckOrDLfgypF52u2T7h1tyi6AnlDd9rNk8PIiLGzESDw
LbSLFGcYsO2EKBTRo4L5oeI2/qNFOi229URNcGSuGsWjW6ZAxUbXu3OnHogg1X1f
D98UY/uH3g14nGgHGZL65EzYfI2sdBX+ZaFIWkmPvMnPgLOFUoD6GTUolmzvQHlY
ax3ICrandU8ZvXGPjzCjSdMx7La5J5nr9L7Q6ls7e7ir/xS+c2p/RqoK7FAznlZ4
UcHAC4qWk42MPZ81VUQJb0eL68HK8NWF/MzmW2owX95YXWZpUu6ejnS7TgYZ9Twm
8FQLMD6Lxf/AWXdT45wuMBBTgUcKg5y/gunDk88GeiMpf6pHMLSieDVg7yt9kB2l
drYhrC3b4VAjf9htq6uv1kVHSghFXs7Aj1rsF/M+UBSx7IFDwDn9kHhBZOcdcOii
MUDj3RWpLq/9JtyfrvVyjfNIuq7XiJ7uDqV9s/mg0AMarV1KWjp7G1EJOVHv0jw2
/vp+sBIooqNNe+NHzTlXpJX7Y5PGeS6jNpt9EW6JEKt83wL0SXQf52/Qpwdkda8/
hn7azMsNzOj9OMkJ1rGukTYSnhOYIrORRH6VeejCva9lJNiMsxZfII3yfUH/5fg3
QPcAi3vr1TrAjPnlB6BAA20CUub9d/wqccQ09OTcNRLBP7CLAKSuFt1L+H+/YU3U
gq3dzqixiCQhWCqfJ2YsWUgO2n3r1Wb15AUYtUMrgfCVAv+8oJnWo3mHoB3WVH4e
TMcqtSzR0eWIsaKYPJANfr2zwyI0ipXqIamx6oiO0yBthocCZG64+TuMzRqxt2u8
4KhfnFgEHwcxlFZlWk0UFxtgYefuzORv419EoFUkGCxH/sby8WSbwumMJS+G2LcL
NxACsA29YNs5siwG+kUmaiTwf0nhn+9/olHtAkwy3EzAVyhiaIKV5fHUxk4vQpKh
YKYMqmctGf6eM+6opc15SeB7xNq7uSaeSis4XT12IOk7y3UN2tCh0CtnQVDG6WmO
Ih8cpsvz1TYiIxellw2TSH0Y2HEdv1Gzhfq5roLogjKwz8s6BI7zZyXgoaqyCUZX
Sdkdmp62l8H8K1FozFAJJoEG1hRYhTsxt/MMRbwPZabGWIiSW9xDS4ori/ing3AJ
qoV0eof+PjwP2yCHYW51DwR0HtL5/L6Fws43h4AmD0xCZBSabykQtYs4JfBjRf81
FpYeLo5qa2pzNPnB6qdjgF7kTWXFGKgeTRcrxkLktzaXZ5blOR0hcxkuP6M7dv4F
JNxLUkPMl6c3N1boANCxxrcmYLmm1Bh4GXuC5823tVKEuSjBrethLnyxm4tP9+Mc
5MU/YkAxUpIEJipuy6VZ+FTjZgy3cl988BDP+1evHIhEmrFeDgnSK43j4EYete+O
loMH//YSVeaLgb3uUo2dC3hIFsUhEsQSKicmZW2eD6F2E/VfdohowMQtHcYsWN+j
112tNvF3qdWOs8vDNdqw33zge/G0yzc/j8/mttZAioyhCE/BRCMjtWeIoPSjLZ/Y
bLQwInrSkTSyzY+i/xY+rLvJI2dIpOHBFKN5qkFnlAZkdKLoXGBO12WJG3ZrUvNr
ywpQGmRWnj5DPMuIvuZy5S04y4pKgtZ2Jm4OUH05z4s5NU4M44ioa2ZAHBgGsC3n
BxjnRacdM4onRSqWyhjsJLmO+vI860yUVx+/6h4vbvhcfgvaJHpCti1tlhpjyy0I
CedYZmyE0kGB9bpTXQkuKZSwQFC/QBPJbx0h4V+t+vEV/ehQM4uyuKxAgdQ360rV
21vbGpEGUQcYP/hLrBJl6iHrYkcBI3OGx1M0vdTHGezLs18VL5UwGKwadlsdBpaW
uuRYWbG48grC/vOs+dc1alq8XAU7VRkXfCXdwfdfyWFbc+ctvWc2DDyaD9Yk0Yzu
i2t884uXG8fJWFC8Mwc00703xkSToNSqb1tfHcKrHKuZ2hUEflv+U9zTIMwbp9aw
fJ5RNyGqc7QVrdZzeLHSUXoZF80bEKwASwaaL5ZaS5Bs4dK5362etVrzvcn4f3uL
GKFKcjYVG8NNBoxSlVGGX2OJ9uf918mYQGqYvHx5xEULosh8n8mDog8THsZdsde7
R9ED+LqXJvHwzK05YBcdfUit2K0Pd4r/vbNNaTNSYXQ69eYJKq4l5UxT3yj8M+v2
t1t/WxNp8k/xL7i0UUlFOL/XBsGX7BjQuVg78mMEWpFyAZ/PT36ZdP2iitVE5XCb
Sl3okgcTTmNowuoRJ9Te5dGwJIUYF9dMwI6SSbo2kA4uFCKFnBgwiJEmlz0EMWcM
JCiObEFesatex0tOx91PuwPlHL19ZGO8aNf17wkiIlq37/jt+gBpWpOBRR7tUuRr
gGJfOhFb+Ru8+i0yjWcrUdOW+/p40zvaNm7P2Qb2lZ7scGAX/nhrqpyNL5l+arIa
DdLtiYqplNM3QfFZ6lNG+gnvCpvv0fI5K98gGhvlo3UJ7KgrNjoKt8AkdDQMD8yR
dBT4VfGw892AvtV/ufy8fAy60SUpabVh+in8uP2NG27jVTniXK9v7wvjwvhoDNTB
dsothZUq/jt0eYZoGrdpJ7hefZHz5i6I+4Tfl4skXyZhvYvD+21ZUcSBHmiGzztN
DNO76fEfvK2WwN+Q2pF+HafPQI4R9xByBL1m9RuQQ9X/YQrs6yQiPbsWqhQJoJfg
4/GPbOKe5L5Xkltef/3CFtOQbNXW96UwfHHMrET10J5pr4EwzjmkgNN2XVO38XwZ
zSIAGcPqARPTEc2AcUyVqEcTq5bYiWkSiyhYBEwlfWgdHUg14+1UuZQVWbNWNEZ4
cNUewIK+6+1jgMTFoD+u2lHzzolearZ6UQA8pnmwbniqbtSeKHVbpii8qX89q9/Q
5ShQFm3CRFYbocW5XY6MM4EQ3HI+KoE3JiEWVuzAYdnjVDz0syRTmfYNLPcHhhim
H3cG/2T6LfO9jlDEUBiHJ1Qu5vvfuif7Pp/TxCNDvWo8G6ZdnRzRuVCwcOZW3mAP
ollc+SgMHpAO9/P+TnTDK63sQzrr/Eh5b+cjMQOIe64AD8Igkncx56tHdsUGZLX6
lIRdPokwRcOTJR1HseBlqZVRkblitlBFqf3AdW5WISbK4G1bp/0pHtgWM1a4PJQ8
qoorjNTP/rpPYYrLVHZk/onJjVFKOk2GQch4bETXuPK8WyjZOO4zXypdWL+wkVt/
8vbt/Sy5MKHxZhxZswLVBLvz5o/qjbLNkhK/p6mU7UlCW/tjOstZq5fRAag5Pqoo
XdY8WNzjUSd3BJHCUO2QeLRwEFglm9KqITeIVu96owFOVSehfBs8iQtRIUqv6vhy
vuMTZ+DwLuYBQ8V0bd25k/3A6oveZQhlr/i3GeGzQPnWU2FLsqZvh8A5tqG09nv2
//01UPsiTbR2wpSvMErluaFnK1U0bIcmGC2NdbFeLi6EVSy+s1GDCFNDeaXXqRf9
NsjmiYm9sV5hkpwQCwe+DRVmXAwonyEyT086Mr3zde8Lg50+5f4lWRn7PU7I1o3G
qPB61cAr0N6GZK82WZ0X9Ei5OXfdTpPAwbr+nQTqsWggT6Rn2T4sB05cAOd9wFlp
BRwOSI7XAarDVbZLaHeW35RaPMSOsHUH3k38mHS0tV/6+Z0FKQiztD1MxAHBQJkN
jPCtdfwk+DwbzTlU8rSVSv6tVFpmHGdaaU5l31pFCW9kD+oa+qmftKTckZ6OcnI0
8N16y2fG3TQUhC7ZdPWb+akT/DJo/Zo5ACNu1dvATUCS7fTz3fEikPt/7N2sBdIl
5i4gQO1BYSljLcEAsoO3G4mQlpfLJdQltBICfcXyH2lecvE+NeGtR7jA2Oj33w29
kJp2GlsN65KyU7aHOJShtpsBJND/FnWyvD6LEU2oldhVNDJZVON4oR4WzAFhXdsM
B/6iMvAOI6uAZz1BbXVX3if8nWL58OSNRt086FuVDTp0vaxuS37oKSxBmxNuCZ//
tFHv5u6ZZtVndtuDbN2Jhjv7lHTllCWWbW+LRuNMZ9ywNVBf3401VXUN++ifTffw
a6BBJh8WiVAATXtVYd1ZvX7xkqUw6foZRyJLCrIVzUvui0WhCWB1Bu4nUAo3na/l
VOiAKqNUv/RptWPyMVQlkXGXZih/nteH14j92j3pUsIK8fQlJhF/13wp29yqKg0T
UhiktxdTbvp3LY49rwbnyK/kETSet4H+Sz8VU3p0+D/RwvC6KWWIuWiUUL4rX0dO
eX1mUEQYziUPg5sUcQ9wI8GFtUhbCgPpoBDCaoU4pgaFmy0Q4mGU+3+u0r6RYq1X
u8xzpz7R6qWLmqZ7AtFox4GB3OCsd1gZtDmR7ScKwt5n8bDtIKQHF9V0B/pImDpX
AorFnzaXcJOo4TEL5t1qVIlpGXwdLG5N4xQLE8/Pz5Eclf4oHlzgIfUaCnMc8HwU
xFIx9Jw8sO+gRJzQNKDFUI0ZDpggWMBnBLxcnsLahZ55c0dFp3+cm+UUW3PVKhAa
x/+PdoIxuaA31NN7PRVuZIlC5KnZhklBA/H2A32+wbghXmtiwQm5IrT6KDauxWxE
mzvnzcVUbXNe+HR81kiFeafHQ6Cjz8MUbpsBjQmxBMVDeuIKx0siGDw4a5nPm0CS
EZoenPvxujkFhYZKAv/T3nTEkEoUns/Rvn7hzcozI7FRlba7rNy9hKsejteB8PSa
6DkwQgtFQzKnpHsMpqLvo9lU00bBmFCoIr7KiaoAlN4RnJVmL1UdDObi8dpmru/o
I51OX/vZq9fR6U2Br/sA74JxgaXuRnPxaJsQFvHwHG/HpHkjeLIW88BXEGTyXiF3
D8cpYDOORYxAzg5dZAt7AEn0I0i7m48eG+l/AHr8VED6AZy1GDrNvrmlOzi8IGJi
7pQXvoFOWulSdUF7GIhlLQ0jTSJhWIgM0gZP8rm4H83PQjjaSmJ7zw3H+BO9RqED
8OQvhTk5P9f89rxLSpwAoTPvNVoEtUvmo9EV2GBaEsaWpcQ7wtNqnMoswFxJ14Qa
JrhQyn/8dklSehooZYsBelMyJBaC+5Cc/ZOnBmKOQqiWabR/8AqToZbkxC9H4cOe
eSfGIGgsnlSAafS239uP24ZOCnYfNBYGOQisNwK0Koc9UHuAsBbmS7BDte6rYf0k
c4c1n26SqXo/eFQjjI31oiWBvuwN/7K8TY72IHo+FopXOcKHzY6BKv8nHy47PlcN
j9Zp4zHaAcEnnFFZEGHRh4zkvO3zvo2yXC7uJso4XYQIgzEXX97KvwwZDwE2cvwH
KOAy+EIP/CJTHC7JlU70sHvikd+VXFEYXawL//mExy+W2InrwITsHBUu0HXBj9p6
Do1AMY5RLHSGoePGOtpUfAqm5X+WQ0zoeiM00d3n9FiXRxmi3Hoa3XB/9BKblHAQ
9scNUpmUSZ+O0xok7B/f94xgNRWu4H+dKdarRMC39XJzzodwluz7xPIvCWL4b9Yc
YVMK+pMH35fKpULLNeJOtbi+6zS51SsocC35kQLL5is5nfIIds3eoo36icxY7A7a
a1tA0FalJt3qUAMmmJEg4omD0HVwz4wVaS3p8vz18dxQshbqBk5VI9uaEyQozyFd
Q5qjGahcuQ1O5LFXvYUtwXHuzML8hrT/xwSwl1s8X1+UYZzzKsRtXD/uOqtfALM8
sbdb7XKgAB/uGhIUMoE1RB8/pyoJObmDXD264TkcaZrQyeWNONV4/1Y7XBeHSmx/
r+nm9ZsKxLdGvSsTJPSMcRCZfbt48zhIJl/UJFw2KEIbeYzQNRiwTIPS9S+FZR+k
nwDwt5f4lzLGl9FjGk9wPdXAiub5Z91LqmVePz2aXL8//FbhHlZ4CNILu78l12bm
z1DeH9mByVIMwiW9yq1HLwFFRviAPtiUmbN7OaHZ9l7smOB607mgRTHrcBEdaPab
8MEfi+fzo8Ab9OjkQM1Bno9SgZ/3IR+XuanpVtCoisbv1EququJmwWdwZGHX1gqq
CS+ZEM1fdXnPLbAqQ/WljNE57pVIQHA0yu5pTpS0jg60mY4jLeacL9gZrU2CjGJ5
22lF1N3kuN50sWgfKFqv0H/jxr7SU0T+Z5iS0v6jAU+5Ua7zzN7k7WMDs72UZLhY
Lg3q1zCu2zykOaKQWUaVrx8oBSGBzJDg+aa2D4K3xTpzd36nLdm9ftp/iRBaKOuM
2CFOz/g/i4434KDSSnr28W2UFR8S7ChbGtdhlM7LoT9ywLl55HburOjsMyAVm3Xm
82emUrgm/LIidfs5XaXtOsk3k65WQaT+JPBF+nSkFBuV5s8bWnw5gD9HYg1OEfl/
BQ9Pyk+Yjam/me4TV/7kb8RppdCuskg2AzqhFk2Bcn/ieiSYMkhvmCZsW/Cm3TV3
N5E9zKwnOLBU5tgUW8FskSRBSb9hIs8lxSuqZtaKUaz9+1SfSih7IXR8xgzBK8BT
TPY6rcEZe21aSGouA3owtcfT9c5tOpR0GpIP9ubVUdHoAQYLFjjAvEy/GRERbiHM
wunKjtDdmMqJ00LYGcVOaObJT7svejXuTKOB0xGDoFlniKjlO9qRpsGFqSFg5+Q7
9ard1RQfrw3e/FZUfW42KJpHMOR9DhWM0u08DiKpF4POAVaonMEknEt44K15BDq+
RRveE4uLo+kYj8jHpmZ9MnazjcSe9xpsAiib5yxjOotCnEjTi3Ptoo4g4ZVoJA9M
c09kPQ+M+c73EhwFArv9T4hdVehYfu6pj53spuLFGUpMSBxYe0HYIJ+/KIFTSwiY
PwzpAiuHmrenevAh9Rrx0S2YuN5tlr+bdxLS6ZgCpTj1uWIBUtid/zKkUvH5tMAl
Ztt7R5tXbMkdjX7xEP2iePSyA2Wnl5RTOjYClbRID4BLhhkS5SCKoT9kK5vVJPci
pvp95jy4yvzpsZvdWR+TeEB5PFWBgFy0HRDXntQsPPcXP/vrgg5Uap7pmmRDACds
YxpDl/Q+nY8/x7DhyAvz9iaRNaeipRoaaEKp+u0B3VSCAqTyGLIaJLfazayuXxUu
Yd8K13TWkvXGB1UTZRXZFY+T/3W9PqKVjhxOyW2Y6qht0kDA7SBBTPgOMRQ1s14U
63sXhN7KTdUapG/mYlGr+9vmERW56sEt5cCQJ6MuBNceSs71Ci/CFHkpuT8Bd+uk
bqyqd3wXMFH8EPMmZmvtMp8j3eQ8L4aR9KNdm5i8HevIAnux9qObEgoozL/5k11t
kZA+fW8BhRTIZjvAa+gBs2Dtdb2Nf9AvK9sy5YZydgCi941bvq7/q+0zT9b0+AHE
4Xw+KGRsC07PzLcOCUEsIAgu/6C2WAahayE27AKSzHUpp3xKCw6eziYemeeISdN7
gNcKkZg+XiE3kidofOkulnv2EanjV3/fg44G/I0Pj3Q6rc0jUQku+Vm7YQhdiXUi
n5dOqcx0bEjYffAFSjxIJwc7GB1jjF4Lp4S0RxFRnUmIzBW7ojXwjpoNrInx7i4N
QVUT8zL0kCeV09DMb5lMBj+FTl2ybBPw1p6A7W7EbtiloCPMguep9qVCum3jIQsb
cQ7MFgdqHllfflmxgtugLJujIlBcSBWofrcFWq+oL2NJz07XuoivtkMrUIDVMsFD
tNbNrttO9Soi2KpZfuDwmhBilDnEryWI9CFmNHDyoIM3IXe1+RSV4kwlQRjPvCOK
LURWN6jS+hkd6gPViVcVeYSD0gdZ84yEX8IcQfCrg98FVW7Aou1PLP7d1ubYeZat
yP98AjdKYPUNBqEzwXlAnNRUdoc+E/ijGFszfSRHLp9I5ItvB0zm9TbPBUSxH6zN
9fU22q6XY+03wbzz6QN6wxnpd/hKOplnu6e3giLF7qfshjoUCHQ+kbay0LyA9LX1
hpC6mNE43crLTyk0Sc86BBx3LxqCS9Vsc0EJ0rahPAuHtTx0zp4J1n9AfgOQKany
GGvAUDxwobhkJyzXNDYsrLRN1DdyZw25YKkwXdAn4vSCx1QTz40/CGxqt7HvRrNT
D1JsQ0veeXTbCyNHmxdzNsU8SpMH0kgNNllv54q7yDqQCVf8FP77oJXaMqdVrtDC
iUQVrsMLcQigzZyQLcAZYJKoITtJdsw7pV9QP/QXUwhn90YgVIL/KStkFw/fAunk
YRTMCup1KpmC6WTfvaFB+jycW1wZySre4OqB13pglWiOBLfjZHy/n5lJQArxgNfj
lRRtQshcc6YhE/QvmbrIv/RlDgDKOosm/he8+o1SfMqFWMt4aIM52yZigx4gP73A
IX2rCOWmaWtu4evhJg8VhLajckgAFDNl41MUL2y+eCpaN1JEhPPjHHC7QaTZeWaT
JhLWHfBRxVgdCMQw+kq91avY9F7lYOTB1ugpg2IDJDiEtvpcvJF064roBUd3fTpC
7GMgWU0rDCUCOPsnYPuDJjb/RyvaOwZQ/2ycv0rQW+60GuNi5kn9N9I1eWLImYsT
+St8/RjvYOJH7SMfmX4CJbeb2RJGYGHqa19Zc+3THbv4+bIUlwzVYTdf/5BAMnOS
LsTb2vkQEaq42ag/s3RQmTAHtIApw0ibNe9FwmcCclgVIjhiGZJmw1uw75L8+UMA
UxGDBmcriT7j8q8jRH7AVzAHWkYSDcxL3WEtqF0mTkkJirEHfwBFVxvQnFRyOK2d
onHBzbA+2ReQAB84e9twd2C/RIkt0tF53b/oCobSj2GROh+5t0s9JLl8e9Ko6dv6
H1W2+5TKiIvULKMX8U+1hzwa55vdmIc2ihc7arXjngdhYYuMpjuS1RCIsVmXaM5Z
U0BawxuljaocDMdK6pUmS0vk6hvPJsOvJkSGvb244MpKSE4+5b+Kw4Waq0h694bG
G0n4O06l3VReXCQpBsr/BILtEf5wz+y5Qy8D8uSQUeqJLqikLarxzqKYYkMw4F/Y
pFVueaPqfWRJdy2Lxi1xIo+vEXvRkDsgJeGd+uoKjdxDtOSEd/TD4J9VlsW/c93n
BHU6p4Z4L4mXZ7VpLzaVvAtZ/AKe3gIt3QKBL1lQOqqbc0EPQpqHCbxTuWitUaTv
mHphvk+eq3A2H7xhnl1YJNLLslug2DzFMx5K8eJr60rVEpCLmxQoXK9tfl4AF5Qy
NVxbRmBkyzikqV5VSqd/dQYfySMcoSO/349JelNZv60c/clioB2WnbQqqIvmYjkN
YV/wG6GJ7t7s3nC4KT7OTljWsDwUHwz5ZnYJcilnbQJ5hqRynJeJDdo1ddHKj95u
tR4LZVtE8qE2e8gYAtJuIZsqDYOS64qnb5JFJObVlAA+b0j15Z1XT6gYor2cAqpu
thZMpZCQLZRhn9RdX/I6Mt1YOMAjc0ETaithVBwm0yMxGdcpXWNtbLSFSwy2hGKM
S1cxuYwEhm0QjjL/blUmzYEKvN8tzLqtzXsUDsO306l96DbZxjDyPAe5QpoMe1/D
eESs7i3/ycL+VAto/tZNJ9WK83fUvSsW41lvEo4/RS6edDR7t4nF8wrM4gFJeBuq
O58x7hkTeubZb5lUCA72JKrovns1fKHssQrTc0fnH4WlzCHwFK0f9Q/+DwS1Hj2e
WjitbJTJ33Xqc4F+oz1gpyVdgVfgo1ZifN9ZQ3U9+S2QcT+u+XVMNOUiNv7FPq13
DfVmvE3Yu2eb7IObYv8Wx/GsFMrwnzVwc/d2jin3HjnXi8bAbrT2VXCxZU4jBXKt
TpcMl4slPeP+lqS4Nz+ajaAxv6M0qeWNigZiI1HBOO0YTwDl+wpLUu7ukIIQG7uK
0kxzqFOXaCly5KJAuSxWmUPNPmVG/GylKhmYyrECCL5jYphIE+/1vqlHkd/MaaTl
HZo19+FVCKfHlIyQnuUT1M80lwtxz3ViFM6rzgO4vnCUtMiBvRhEIaxLCApxzRXr
bPc97LxtI0uxV5d75kDEL2+HSfie/DLV40SkEQ4I37+ziCAuq2PAV9TEUGykGjlt
3Q3OBeRwkHR88FqZkJBrABXL7gSMo1h/23lHBAvRCdtEWxXEifQPW9UkaJzNNCcm
MZW5IasBBaX8HBDGLT0BvTA9HUzup0HXe/g1YE0s4QdrxzZs64NzBjLmZfLkbaJi
RS9WghBoTBAmcY7Geolgf35/wTs43es9fTmy4NovqokotzfLP432BZ1IUm6BvePn
+HaCZM5/zi4tv9pMJro/KHQBrASY+NbWW+El8MODyo1LEdqrYYhmgiK/P1jT6d8e
K1soKkV2g5K0GtT34UerXWQWHUoOUyh0oFkKHELgml9z0P8qTNnWVX1x5q+6dJ6F
ywD7leUC+HUyw1aPRbq8lDOnkVsRfxm7WVGglLfTmYBJe/gvYtJIq+xYtpb+dGDc
78Zr2aAmGpBEcGUP1ozCPe62T0HwbwbraaE+VS5n0pZD8fheOuC5T8QsH1U2W7FA
KgjhY7MmWpTbXd4ltTFBFa0Mo591KqQowXA6DPeBvVYLKkkgn6fiyKajVPPWJZ7e
YwTtNAx/JgXvcdHtWaQc2n7cAofKHOJnlygnfDKxSFX/82XFF9tpWD4liGRmFlYg
31NmJ+dPCxLbr7qFarN7KLH+mNfNqPzb3Tcob7P8NkoZ80UscHQW4BO0QrQ3NAfa
1TlRKDGXtbnZETJ5n0IIZrp9kNXAZsXvJqzUSM8fQ6EwLaSW3yNndZNbQ46pUnqi
r6WfNJqsXzn2I8bxAbYMdl8RGDBZSvq60m5Vbd1TEIEUtBhCa6DMvDqzDkl/d/eV
pWl59UZpafJzpsaaZPpLeKorxG6GWvPGIuSl8Vz9kFu9S9/Os2lZpvXHebpwwTgb
eVfBorpGkhdp3j9a3y8et46Yl+/3hsc9/JQ9drmpBy+9ETi6GDxPaDeTZlKB3w/2
qAF6aX+2YXAapjZ9mfPIo8iTQ7dSf+LM+/SEejFC7T7hQLh5CLnXoUb1bbnc9hTe
y/gcDhBmcGg7ydC0kTIEoO0IWkGC4sSwVfUz+Wpa69LHiAxz69XVlb5VKRXwOoj1
z0axTbYXzfL9q32er8xqKlX/eHLVVqaJ74nTdWzr+sKqXvpdDu2HVR5D/In11K/I
eBG1TxVxXknboEBVeWTmd0kW1vntmNaAbxBCBt95a/zctCGB/yc6/rc2o6gkbyad
EdkUpBvv71GeifS6qvvf57wHbFOwa8XTuJfweMtCYEmbCd4N1maRoFekbmleIPi8
KlzMGolZY3yYr0DVvHdyeCCMA0/sEWBJNvdaXt/e690A1yS+6N17LhLDV0btBloT
b6kebdlwxGJaz44RILf820AScw2eWWXda5MZizccKJ+fcci7JVuQCrIMpRkx9ucq
+X016k0P3E1SSY7nDXklivA1SwEWdtzY9Rqbwjtlz9o9W5ypy99VQITWrD4C+hsq
3V+byd3RMbl48JW2t8f/iBK2Waj9efCHRIQ9wuoqDe7KYJhVVhAJ3eMlEMXZ4Rg3
4au70ZPSAN4LG/m/odJa56ZDsSok5IwsugWmYJ6t22fNpuWUoDaBOiwqMGGxS5Yi
wt5n7RWx8sDmJduvbApdF2TSHd1Ybp9Q8/iF0ZQ1OFbRaR9LnufrJVh5FNoCmH6Y
ojDEmdHgB7bo9HCFuXtHxQnvBOw2Mb7Led/mLxFsJbaVNsV+0CPfqOsx0qcinewn
GdD06XtbOGQP2esrzSeJaRipHpLSsDs1YxCNkJJsXPau0+5ftF1q5CCLV49WEwMu
AG3iQ6RrOlXdLki8Rwfmol923Rv4M9H2pTjnH6cmD81USXSM0KnhGBDvgLa57wsm
ejwQCOUMmV4OGMaafR4yO2IAFaPpYxkm0xu6PFMZBtNPVD1+i6fTB5jqX3YiYmCf
pHk5uyR/WvUFnkibCFValE8lL/h+EVjOdDEesPhlrcFFNaxVPyQlZfUt1TtOHxc+
AVf5gVUzFqGXy4HwzdJ1JxVBBHVx4A3Rg03AlWUmJssVSBzTb4Sx7mISv+l4p4iU
h4QZ8atUZE9Pk5PjdbZ9ve+DmxrA78enqZFubwPChxp1SBAbtNEbt0UO0Uv4Cu30
X/adgCJwtXM/MPESOzUfJVnpkrOvn5IfhEXOmdTmsHeZf2rgeifSIpSG0dD96Prw
yZRPzeg7vBJ9OnBmleJEzsGUERrhAsCQDtrfKY1XfBsZKN+D6yZq1DBtF8Q/lgOU
plX/C22Ar4ndeaaFn085OmHGtucNS4Di8FXt6syMHXWg6qYrPxasFcHuj8xGuMhv
PTceGPwbIp4QtFPaQNI8hEetdFiyoQfNOwGNL38wOyERwXGPTnYNTLTsiF0nX49y
rk3TE1oGjNvkytOl0wcR6SFk84IuvZNkVgbKzLS4jmHzLyrr75sqYxnGMgJqQvW1
Gx3USQo5LudvGnyUrwnJc8eahEHDhN3oQfInGOs+DR5qpznG3ZEZygWoV6F/V3Sb
dAGQ5lML+zoWsS+1sRYeS46Kewu8zivReJkwi6FUbW1diZ26LRXx90ohidPFdjwa
7b0yS39O8p0kGnJ1brbNSsxmIZhP3+Yc5SKK89O+Qe78ta5NdZoMBzx8YGw84+ar
9vwZ+GdCxWHDztm/wRwZOGptCjl4/Arva2M9hfVBupjsxxanO9DAqXxins6iFgcK
PXNrljESFcAO2i0IPoOlVRV2m0WaveQsXt74wPzb+j+vV7AuJU7tzxydwcpgJ5xY
1/U57eyPLCWugAzZR8Dqt/oHcDNESdO+j/tLKSUea4xAkPHbos5ZFZLWe9YK7bUB
CLbgP/G5+E76Wn5CmGgjcueTpwtJyI8nfIwYr9RFNPW2Lt9FffsRnXGXlzKA5YLA
bE0s1aO5xy6MBg98Rvcb7yAFmDH5nG4QTtoCVHVFGR3buJgf+AUNoA8wg3/4MlUR
tPr8YX2Jv9i5lUM/ECHxxYjHOIXAj1RJ3MTVTawp6HEg5lZBd11wGjLSE+L/irG3
NNL2nsGUPjXicAD9Up6VOqj02fbZ4K1ZeBhrA/DSwS9EbWqnkiIHcKSWKq02OYAr
L73hhxsCIG+VlesnscrWLXLMw2hAme6QzvaoD+6xi0D4u8djHI1jnRrsrGItmtzX
v9/eQFKtv1tvpd+8sB1P+AxMSNnf8yUqFvuAqFGeePath3L7+vbCgDgMN0wmTsH6
GN14Vrzerdv8DNeCc6rGrvYFBNS5Twtz9UbeQUDtM8iePHTJlr8hfYdFUcNoFqmR
YfK6iXlNbADrWWzsQegnOXgKykxj9rDSSVvYq04qeenuWJhslI3dbNA1kCJDzqhk
h7pDcElNFeK5xeNqzAwMjnJtYo73jGgpWcndI29oMXGRlbKikAwDrwkssEYzbPIc
csc+VDJD3vbJ57ijlD/nKT37WaJG0JTF0tW7Vh5W82SQscCMQ+0Xup8adUMYXRyb
2SkeYmwNBtDtpG0NUbbl2Qbm0SMeZUTJ2Pm46b+QLfuBq8TyoVyUXW1LmrVP4F/P
ffyONmL0y2wc1km4YE+ZFEKPhBbxHvk22b64rUHvX4HaNb8S1JWMpr1KTlyijxqw
sAa+p41y+fxErgy3z+8c7Uk0ZokZ1/Ovk5QgnaVErEmDrZn8waW0sw3ooaoSn798
9x9TDIoK3EIUyQPoGDe3T3O1Ke2lKIAsRxK0MfFALUr9HSJZEsYxjiNgO4HzmOyQ
fH1vQQaxtuPDal6OuYDWgdtQj6DP3PKMIvk4etVg2XzPamYsOz2eFZiujqylaRfO
SAsvAGn//qCTQ6d426GAcl5div6V7S8YjCevg+/NsdTajtWrc6tu17pg/6sp1haO
r5U+ty6UKfBWypRueYwX5lpzND+Xh4o+M4iFqePHsZTnPD0rrXZQLQuS0qelh3KZ
FeAnxwgoclYlcEoyNK/HOhM7Obk0DhHyqzs9uJAYkjxZNMpIX3ARbh3EWKB51XM5
hwWZacZ/nGqmo0mEvgP+nIzhnl37WODuR9rEheA0/GqG0YGWzki0g9NYO3kXkP5o
kn2mcwaEd1kBC2Mdh1lNRKJ8j8tG6zymKzIfb6i4jIXPvliuryfkf8p0K2bz8JBH
ua8xoj0sGUnFx7xUey48I1hDDfWavGmVeYG9jtbPu0XwOWU989Ai0BYI1iVuGxc2
umjISNivoJMlOQ9nVbx+AeNEjZAn29xtDO9OLSJy+SG1abfDsH50V3nmC1bgxLJu
20MtuYRUKQpqowG/TwB9+dj5Uj2eJz+8JEIHmACTM290oI/Vw1ZPgt5FAGg/eMWq
bVIhNB4W+Q2YRr4oy43ZhIRjpCYcTcxNQ62Koe2NwKv3ioJV4Fod9bD0TZOZUDSF
UQE6mlglY6ojhrcxN39e2828vEL3oDDAYSdAFVoeqeVs0OFrE3GAAqAm21bL1CTM
pxnWOwqP7Y87goI4blrObHbx/3iccctFieuWUYwlr0tNH4OAj969UV/WO4eCsBly
n3WtD3lWFEZotnYF1b8z0C6WGkxwLDQ0Lo7I4KMH2zx5mXmvWBCnIVRgRoAA7brZ
1Hc+zWncRlAT5pteo6724n0l3nYU89uUsQQ+rqLvw909JWYMHMLXHwQm5SSiXZdW
+2WDDiLBvu/f1e4YBAaS1ROQdRCqC6N580O0C04jAJygOfhA3xZ5WWTZccx5BiWB
/ynkkPg13b2W3QUzFU3LVVWH+qyf8KYDulf6zxw/60h5QTH1iBInyc7OAzp/54lL
X2ZD+IZQZOVWS5N8GJQ1wlCG43OS4HDpbck/UWZEPpuAmg5jDrEdabFMLdU7YdVU
f/bAwzvg0X+f2Nm6giEZ0vnohSfQbPZb9WKbJw0VllUmcJemDZNG6nAtFMkbHjlo
5lhhVkzvJSJ6b9znpv5VbocC+kpeiyxOpJiySJBcZlDHZuOCvfAxATE8yjWpCMVb
qanWm5MD8VPEgMpfUCbXq79G3RJVRyS61NBivKMthHCsf2oWw1ZxbNSodgtKitdi
FIMuwq+YHi8bSf0hyLs7rvWDn9PwbCdV0mmhIorrJVrtYDqXO7rTxdb4DyEr0E3m
Y8DOeIPzWy1bxqz5omexXos4CXPegv4lWclHBf5AFb1HC58qpqf2dkaGHN//+SrL
BuQH/YlqmkyBV5gY8R2TGagxMECaeKFh98YM9KDBX2np3f3HRxIKgjLllKpKb9v3
narpYWEGJueoFnwhPC/WLu4+W6DI8HILNXF5iqwiDgmG6eQkUgyeTRRfs+FeWzdV
NEsl+hiuDB2c7tvsSVhOVTsgDHLiTOuk9tFz5xf40zTTxN4rALW19fywg6utUlTp
CqHa/dzN2IuK3qSj8foHWbHz+IWKUJBE4Wqm6XG3MjTjbFVSvQCzCr0KroF++ItM
ztiTi+SWQkXsU1TRiffPEqWnlxp4LrJPQBdbkz0Tl4qf5jqIoBC30okaVFgmwA+s
hELIdRQhGs27Ola1qcv541YdVrx6uOqTlUvZgg1juPy98CSbHsZK0VW2h7p6HX+T
laUKYnWWEAJ1nBLoL3JaJ1pKSB0epNUNtmJtMMixw0ceIFCa0Du1fMNGOIYzwKed
L5bV812VedTaRABqrjolMo69USXePknjNjYJm3TTijwhfprhR/MD4X9CmmKftSkl
7rU3wulybvcTofOzH5hU5QfDDd0Kn87JHyubjckb4AC+PEqFDUGXrfluv+Z5HtfB
/zuHPR8RKyZKY2NOJ/ONu37/TiyGAJiSAKtZEkqdpfp0j2F8ArI8Yv3TZmG26mYx
E0OgDew6itQKJcdqqD8iIlCb0aZYL2c9Ptpq/khvarNg1FzEBpmbaShYE0wRF6BC
hKAKdFX78Laxsba3rxY99CLMYblwjca+Uv7FdRBL9gB3gPGgO21lXNFWrosVDnSP
VQ8jdi/FOzFvcez0qY8TU+d6exnFY3AghQUDgI5rVBrqYfvKyOiy/w/GVBm/tMCb
yEiniRj6oQd04yEtHjSL30iDi/4PmNwf/KxOD0xgStj+djAF0FkU4A7sP/RcIM/8
jnicjCuI5XtVk746LWE00El6M91jtlnq9uf7gzTKwv0H710H/mQgQVzn/E2rCrek
hs7eVVzpd/x33G/kekPXQ4HepT5ysJiv0vEdi8/JeaRg7ul2svE57PQVsIZAIjGE
DVyDBgctagJ68gJ9a9/d7VrdyGSHYduWm79vx11RmKf97FO6a7+vg3QDGQnpJ1L0
HBQYR5fPYUmD/W2NXvMEepbR2l4c3kQO393BkO4Bhho7rIk1bZv2ZaV6PviQKxuY
xTDj1OvuZrEne0GAq1+zOmgIrmU49eWzVK1aHuNIYouLy60yUJDXyH9+U9VPZ2F5
8ys9HHKJSHGbaGH9qXuh3zaFmJxoKPuem727hgbamiJjdNZxe0zX8JzP29Jx4+zN
xoy3QKBTcmD1Z2HIDBGa2ooKF8rHzF2EZoooHY+p0gtGa6+yyCOiWn1FZVZY457k
RnK539M6yF9IJltKzkuVkOjDEmu1OyqPJwIGOObuk8Relm9MNuaxm2GwHnmwEZRx
BS90LpDRRdezHKqyh+8NCNyXWvN5/ibgdC3KAt6lAKXGSuvDFXDgaF7zXPRv6/x4
D+HnwagYr5van8AuiDPQsNDRkPTGjwKdq+WusIe9wy0mrx9cmpMVLsmWaWbaQbdx
7+Lc3F+YtyrmxIEiphSzsLWJ8c8Z1OE1MQsfWwgbAM8xxg/gwqt3Ncu3sXsnC8Dp
vUaxC6IA509dGdJtDAn3YMQo3e71oOK+T8XeDUSf37Igq9Rs8NahKMimvhp+PzyP
Hp403xjMTPUGWsyjtCH0P9GIZZxyM5Of8eSuHjUol8MKmuMRlHOLsl8RMA89HACB
sxHEa4sMOFU2m8986QSv6D3GgqhuPXEmtz6T3fdIztv0ALz/Y6Gj0f/qdRkFyimX
QuR8H//DNGENnbLMI0MBKHI49L43XYp2Uze3pE+g92ddOCPlD9l8glex0HloSgnt
urpjYteyHurg+SjC/hEi3AU8ACY4iFeyEgg3atXhVdK8Huc79+RfqZAEWBy+Gt9m
PNgYltCYlCbzzayxzQ5J3sXOILq5JZsK4p+Ca6c46ig6uTZvOfgZhimQT79FAPOv
KXWY1aY1dHZdwgKzdqXyr/XWpFPbbpbU7G5sLq624VZnIjDLZVA9n0MD8q6v85M/
smGkjcNEiucdqhp7f1qGRIxwW9mP8oRJqQo0Q86lPKi+H2OWtrNPZA4R9m3RDssB
FCo/AENnKk807OXKEhbL5scD3l1U2Si8tyhIsxzOoJ86ZexurRmq2jemWx/IXIB5
SfiX7bzXyT7HSMKbkndWhjUUcea7lMBn8KCOFnVhwe1yJ5ypPpz/XWKLo8Gv6dsd
RR+oasJhJw/57GldddwuDl4EfcRGRdPW6L+XqEYsUOu3DP2zbMAvW6aykV+O/4Vh
jtMYFx1R19YOFHKsqVnMGOo3PGFWcCwgWZXZmEWSWEHpotzrHLobC1TIUG/cy7OR
57p5PSgxQKAXh8s17EKxKHZmlKvO+9DEBuqUdWc5CU/l5yqvy3lv2yNnxkTEs8Vl
jcAlXvRxRczsdwQ6BJugXWjLPY4cnsAueMCH5JxEc8fs2ZcvPaYXwDQRQhuAHPer
dlrxaiQsTiUGTNOZpeCZHfW5qjadwOmgdmJVuTOpvjfwyl0Z+v1VC2x3bQPZ89Km
iIm/LoJM82JDZFVZTr2i6eIZox2MMFpNwY5LGOML9zV+pSon34k/q5xQqZfiWae3
R1ohCq2eec06+fc4J60bVCx0kovwH13VHtDXBg6PN/1ixZiUWXYxeu/cCkKjmBXs
36rp1GLdh82tQgN51s35A8xNbWG//ulV89sHtrDq1Mw3sfzeZO0nyn/qKFBdHyOr
mcmv6+jSsYx1An+nNDQxq707ukuQHjQuvKA8vcPnEY2fIc4DxivyDoIvJ14THMXt
suNBfAy9DPc7F8ku162g5CWtf6QZ+/Dr/MXwi9WnZUmAImmos57CZV5kU6p+U1dy
GDoiD3k5IppoWYd+eOLPbZXnzAHdxszOREzBU8iMFq7K9cWkw4aDqMKmwYxsnLUs
0bWrUmrl6WD7Bddxu5hDWSkLTO0J8MGFYnLRWQ2hzPxqOTgunpLPyJSPL+ewyJ3S
ch8dL1UwdpVw5ZIoavG7PUU1wBY7swqvL5QDiT+P/wcGDjoGI/kX4TOetXzgMcCy
p2FoPntmc3sLV7Y/9sJRzc0InNG/AVQU0lESYGv8Kwr70BS+hmiQPxcaAu0sfIcL
zEQDPYeHhstMJfQ3BZwXLHFv4EhTMmCYuvRhm7WDAsb6m5HkmS/Z0/eHT7+S5M8Y
msnK9G0nZvPaRBBdvi+ZxKhyfmeJ+j51cKpSXGownM/Ce+apfYO0NlT9hHz90zXw
ykFi+xpaKa8Yf7c6/jnWCZ4BUt7a+bb+zvfVup9xYCrUJKgNc9YKCkWDnmmU7+mm
adptRkD8BEs10Y9fF0yYmx7g5k83Q1rLTvQhQemwgVzzCXtcp51ryWC/AuR5/pei
iXTlr3BN5M3INBAX9RinOxntTIXMMosa2JcZWrXQZCLF4FD/hpVsdvIL8chu/5xp
CLPMjBbw5U/iIKe/6YfWOQdqu8pHsob6k+7rVGDM0DOyuNIxPY+sqLfEacwF20jr
Gc4wh+zofkr/iR1lmZjStvPrWy5aUy/OuXc43VeqkE4IBiN3mmyReuJO0P0il1af
OMUVgPopx39/6rH+zw2Aam+F0C0p45m/Va5Ao7Wmjf119sBEv+vC77HE8Sv9MJJj
zOsKZnddvVIbCBux4taHN0KiFHDUn8IciegvEORJgDUOvXMYtc8IOoRsa4G8F7aI
nGSI+p1r3U67l95W3M9U+NWW/oi99FIStedARs1m4SxAd5/cI9TsfO7u3xIYDcSX
Y3ENpNJjsdSOsGRDupkznFQcw23wg9CgN8xm4m0ToREvrIZaSbm4awV9um/rGXhV
Ll6dgOqxKvW5nQlK+inPmki5oL+oEgczPkbGfkdAcJ7h+o7kbfVr3seJ14HDXHL0
TbA1XigByMr6xzPvlht7rGZ5Uiw/+PvUu41QBEAIM2RIcKXmSSKbu5jt1h2ZX2EG
ba8gWMJopMIxB/HeOXKYDF4pfNp+LlQx4xJz9kZ+ghM424LWThRSDJpKmZwEBDLZ
4Q69MFRwTglFUGYORFxJEFdGQ4RHmRqXMvqB+TIMAAxwA8gXjls56DNR0jVw1XHa
etLbdiiQrv829tXmT96YxQqRrbO5dDp8R+aDPQFeZ4CPbFRdiiOa/ZG8p23v/yfN
PJjBfBHroXjYVf9AIbfm3jT8n30CcBq1mhFy8gIZZYg10QqQO8sVvU9XY6++yufz
2Ii2JLqGvnVEo8Q2/sN5LlXDz6FJQeC+/+TXxl6kF1gtGjxOw1/J6DzgPIUM+I8E
p6RUcWtSgQETiQXCzi9mkIGMYP4tQvB6gNC8InbHIyiI19C9/o7pNbeksAyzs5/m
5B5n4AWiPfYAjGlsYrCTr0iqy/Xbt8rDwXOvaVtcLrS16jBr9YDFy1DV+zUxXK8i
cdfApc0YI6Bl6YdlhOpTT2jkBUE68EbYYeXYQHWxT4QI+CceJyjqGd3jEgt0Nool
9J0wQL6Z9EsxH5SbtHhXXTkruLDxfKYlOLMnL7Nm6vsh3QKKRBu72flNRUhzsX5K
mx+MrL7RLLPUuJrReNcMzut6xsDB5p5LtX6zanDiGyitTOP/Gd4g8bwDzAntU7ob
sVP7uwM4BsERd/s4eTIAUOMRz+hmOyzEkkhFTEdKQaKFXFw6NeUhBfJCUh+bBIg8
nZHQpyKieP3iJf8rIbKw2QIb95SfkDEDo8q9IKNun2HdMavuxVwlCKo2lS/ZqUKb
2cQbB9irVbZu9oKC2v+PsHdTdasCw8fzxu2lLJOG84sXwuH7WlTYCOHLoQ+kGXai
sD0mMmA78sDNqm8IK1XT8rt4zpn6kICraeADLBpO5NCJy7rdZMQgP3tG7/TNhCRK
kK3Sz3WXYWLC4Yw/KARSsMW9LHeCvSL+9gNyKS0Y7rCqlDZOw0+BUrtYBSjMJRor
L6HvXNJtHrGA4PvG6be2MAArVmv/LTr0wSRCrcIClWpzEWA0Ir+46/x5rAVLzyp2
G+8ZL4J9Rh+NsV9QDHTtO94J5E0K/84AoX90cHMrAs8gJzexbM6oWxsV3KD0wVgd
NZTc0xw29vRgpBnENGXnHrwsEg2e9c+k2tRgjid24DK64Gap+TOXXTtaRQWEyi+E
ODuxXVzvDDV6/bNB84/qr/s+DTfeUvE7qnGvvy+h0bn1OumWDg1vtb7gq/nxdTpC
CC4kEs3nhxF/tZ0S12jaSP9smvtlwbcwrVyHDrrvS0//wVK8sNZwUkLXPN1FBQY4
kdSU/GyYukthfCK4J4WpBLTG3K5PD/w81aJJj/3yKiztjUntF0ROKyClgJ1Bx9Ty
b3nCfe1kBHW0DfsyAdbBpt/bRrCDQEinDgYnDhJuUvrc6sSqk8w9NGjpsPu/AQ88
yyJ158OMVdIUqN9sxVESHIaJN3ETOm9EqUVGJ+LOQqUzfewsiNv6XCrbLkDvP18N
TiOKmcg0ca5bbaUdtGV14lGl0r761lY1CWG2DJdw6kQTs/2T1T5CPahyV0ILBa4D
iN60VI7S04LJivV2KjWiBmcQM6xKg3t/fgClP0jzdxYA96kf31RsCNpyKMwxf2ec
ixzXW1HFvOrBfP7l60042K8175Dq+b7MvHIE89ZRKMaCvipG8yK1iKvppJ4beh0Z
5vonvE+MlgL4HEPMmFbk+C8ifrbGe5ROGQcq1RJJOijWYA9fb/3fFG5rMtT7KcHR
EUj4vApQb46cZz9CscsKGBcRRCnyJQQqMQ5cPwEZXtjIngBfdYcL2rjWWebOvZKy
tUHSzI5DBQ1IYrcv3kaKtmfXkgrkO6JapJKR+j5NqjLt1mMd8chae/+hNZm3yCAH
A7CBjf07b04GuhCpTIeIJnIDS9TKTvuWFyXkUILtCceC4cfc5n1hrwaTYC+CyluH
qKSLPxSs2miG9a8UySz672p2LnKPIZN7rgGHkdTcvNf37ZCH8DqXiAk2sND6jvSm
F+IzyJHa4qk6/G/8NlJf+T/UOZmsg8/JXP/9x2lJnkWxa6mBunpQIwgn5Q58RrBK
zMHZAg2zn/Z0wLQ4H7y4Lta0ipUX3Jm63lG1VCmRGkcR7VO2VcbublwykYJl2Moc
Ydx3ZPxt9OwMm2ykapS+P9e0zfbXDCQmfvNqZJ3/x5oaw3xLJLwX1OOZ9sf4w02g
t5L8nGrRLjcoNhIqqIebl87cebPWmqT36Pl7i8TGjvouV4WKUnU0y3yaKF+WETaS
DgeeyhSoAnS7uj6WqaAo/9Wyc3uKwNnijH94AqYLIkCtMa9Ecp1UFSo6i3HoH21D
W1sqBWsXVM8KZrnCATwIOz+MEZa9Ngsf9Om1jyr6Dfqf/F3fa9uh2BC6lYwwt0tC
lGX6m7VxwewsYxaf4W/3i674hJv51x3epXjgym9UDVmeFijDPO+Xnkze5KTVzs0k
l7FyDC/YUypSaFZn25IZg2yzqQP0buPJrKYfN3XsCal/FPbrjHRzf0ZIn7kVvyR4
i+hLocrbaNiZr9jY7tfuVPThsuyTfgtBcx3PPK1Eac5I7INfK0OwuD6nevs0uaG4
Jv0y97YLTKFrtZkoyCmYZLcqJrNx9E2qkHY70UuAtAj7vUC+AYJGMxTgLEBwyNJq
sdb52s0DKCZ6MsCYPO4/oSD0ES3AOcShZpwz0+k3MBZi5egSnZz0EJNlvlZWG3ot
pgIWfR1RkQE+YzI+4JvkDXXYGecnmsReBfk9yzUb9dS4eEMaESPLaqirVUTBYeAf
h+gt8P/C2G7BAlI/cYb2Jo3y6yCx6FocCzPAH+uwm66VOgOpnm0M3yVBUrXF8fwm
rC2lUerH6GexaDTGkJxRthqPme0e7c7dXrOPJoopV4mXCQOYKiZZVCuetQDst3e3
U9agcm/6p4BJCE3qRMAHbAFTyesiE6U05GAswEW12HbR5ON7AAQWlRlZszyt0ZO7
vwRX9A/q5UgxnFWu0CrLcPbQQ013d61lZ4Hc+ro5k4hlpngkN4Amz8ZEFJs3dfrA
pEfT5TCqmJDSbCCLWpfAwiuqth6YouZpHh/x49o7VWfSMPGa2P84UOz36h6207zm
Ljg8WUbeKUPceUlGiqrXEuU/2L04oseIYOyFjHvolyW5zcghJKY1WoBwcdIZxUBI
oAiXCAfqizRXqi36uvDOeQXbAxtcYP6Kr5GB4+wHXivDfdTs2VUMGZo4z6ucgO7C
IK/9Yz/Z9O7gpb2eQgR33ifXvQV0qJRMd0R7R37XcZO/TzDVdsgfiNmDcwqW8I4O
dktyBfJUhKAVSMwLv9ipxI7h+VXtRxI9lrdMvRTInsSfSQkUgCDRWwSyVCLKh/yJ
WEZRIDMyZ9Hb7rCJ+Bo8/4LWAxleCD63x1e6JdI2MDbsAdNos34gnc7mmPlUkAQ8
v3Uxe4KcpNZTrtMxsDqa4oRyH3SBuMf7NGkOtDAlGNWpcTkIHcflqwJUzXL4qiir
KWTHJMz8eDNg7ohS5+MCnAvwgIGRom3spqP2hiKqj76zrvcqaPuMexobPLnfj8Xg
mgfITW+R/Mf6UpyTWHzwGluFCvX2FBBcNepmwsO8zeS0yekceAPgOfvhc1SJ9RpF
q40Fc0NDW9NjE3wacAzPdjG7j4a+I03thSiArvYTliFD3Bvdu+/GJxneoVqYCifL
KKV4eC0Yu3sVd9F6wrfHf2Be5W+/DUqnrwqPtdZ3B2uVVUSO8sQxIFc712oIf4UA
sCbzoS0VsD8Iu4AFh+c3dgkhuq6OY24QevNPtmrxoUMwAhLi9Fqn/FqwMFSGtD2T
FjkMac3vUg1+EyoSGLHUOaP3xy+CqKFjVvfJZ0mjJZdOlToZb/3FwdEeh7tKDTM1
0oryC3JnxQ/xaN98JRCr6cWGAZLBcyPXnAGEUdATiOZ/XmNrHOO+05YtFY7ZYxL6
Jk2oZqOzRWMp58xOxOLSzf22h1nqp91D1+ROHwJQ/udrpXrUX1Dw1ambM4ZHKPc4
mKEv1lM3IObKr56FnA+r5ZbRxClG7ccH8uuE7RGFzg9/Ad0DdCBOh+S+NNwulaAx
DswGj+n5e7bHAFhsp9mx1LvHG2xCEe0muKmXz+BqBs3HliKXrqPAObofUVXkb3T9
YWA36s59plKno8VdmwOKiGFS+d4tGs6Yz1pBC/Ww5m2yKw5bznexC+kd/kiT5qp2
ll1QIZmZY/wnIf3qR4cZHRML16mBAb0NOA9IUQTdoeYzS9ZIzZODfItVMHL0xD71
eCp5uvP8XUcmlM22RL0hh9tES3zOL6cOhpja/5mKctOVjQvddWsTMTRf7+OEKvmN
Z/BGRZl7wwoUG4CSO+teXUauQpJlWXfk2L+OAcTkSf30p9v67WJiz6wmoYhkL7AW
bZG8y0Ejoiib+hVUNkvuXZOBuY9IFmT08SJdavvr+HLto6N8eZGY2/cAx3rQmmIc
DwRmHfdQy28GIHQABPJLYbaovHd4yoeF3db5J2NzrefmUcHREZvjcUhBgYXeWpQ6
EyX5eQc9K1XWOOUKgjRPHDZUCPl2nLrly04L3Bh9dsL0hk2//RNKXXpMH8l8h1Ub
HKNIJoJk1ppR5HyGBZtiqt2eVs1kiVHqTRKccg3lKAnvLsDV9vQMOMbmPVb9t8aT
vXpboC6OJKSM+E1egwmTaY0olSW358yvMfbjZx4ijaVakcVt4isG1YFYHUmDcz/4
H+I7UOnH6cS1rV+6zgtRjI3qyYn7cnVMJH+bPy71aeV4Ez2NTbpx+cbLiAamL1/Z
LEXFE1kgepr9XshpagXUiv2jbPAaoHfjObx+i+3g7Vny4oYEIfo0wKpnlw1arcJY
Nw+sGXHWon/Lna0VS6Sq9GFeycfLVw1HXUyPz+JS67pmTQ73hGD8HqYOtQf30poS
bC9VhRyhS4F/KIyMA/03+hiH+pcIvmS2p1Zirs7xuXY57+ImIGAedbX7bIoRd8Iu
ukYIlELJyiyLUcrzg807ai+YpFaMuAOwxZLEJPEJ/x+RRfmD+yxRU6c/G1LFiOD5
x8tHT7pL1ipBz6tKscAsiYV2AIz4jqnPTofMJOJxotO5kioSAlVhZuAI5+DTHQMd
SwwTMIEuYiPGsGSr7vUuEo49UyjGjEfqMQ9UoCpIzEXD0E9Uyp/N5o3SR+scTvtz
P7fQ6s2U0T67wFcbTMiBnLgzbdWMZKD1oq59SBjWBeR2F4R777MobgR5mYIPqpZ/
8f8BsgtHfO8VkDCGmsaymRvAhv2XRSivUmgY+LFQJ7/ZeQSn/r7b85Wduvs6uS7W
YPpgbNrm3QJnk2P3rsEx37Me9FwXYfEkhg1lkTSB/IpW3bUcONz+1fJKMaiAZ9Ee
PovdSucahWRpmC6oWAW8BJNs52AVypjaNuXBDUP0CoXE43iHHCuODkuLIHEtM98o
13QellC1uJ4SNo4JOEij86EReR9793G6jLU03tLjLWsjXrFB0vJZITzWNRoJ4CAh
XsSrRkqWqCXz4pGK7qJ3j4OGnT7v/mSvmjr99eZVgo3+2SaG0STkY7cJhyfjPvPu
guJ6KY451Mta35Ua4Co6ku9zeSYwOrsSBItO0dK9apQaOYD8Uwrji8B1NOKYIjZm
Y3yzzEsnr40onEhJk+dbbRhBDikaKHFDKepEJBKVDb1LB6MloEOa4am4ptlTJnih
aF9WC2wB8sq3CGis4A8qbdgG9X7jIlxM6PTFa1CtbKooZWZJGpFn8BYhmJSE+oIc
h9Oz6/r2xNnIDiW8ZIG4vSOa80Dg9t79wkw3b7cPGq0uBE5KNT4DGFP+Cj5yxKDh
EKTi5qQ1KNXxV39r5t9GzSK0Den8YexkRt5yMNaJusGuVsO15e0C4FWiLcX6y7YS
pEbpamJOdDibtGhqfKR9x0OREdC2W52A219lkHyXZcDVqruzhCmfDg2mWJ0HwAXH
qns6HT3S5iInUVc96y9d3x3udcQtAtM6TrCOQQWKPtxfNPj69QhIIUxnjRyC8trM
0mJp2/DHlxKUBju/vQVNz9WUL1ZhQvoUfnLH2ese1hyhZyI0LiTYLdGka+CCplrj
i9ZiMXeZcJdF8RyX9UuXfJR6IcKoCoiEsbnqan9BT8IFYVWIyhJUcHJ2kAqFWhhs
1pg5MPk8iS+aYViLmchX0oOgrvsdOM75AvbBuQc4IRwAfY3qdBzo0V3bQTMK2vPt
tdT2+eTEAsGGvXpjz5jWgRIzsiKWus4aCgq/m48C4N3omF7lbiHv+phMlmi8Uyve
GxJWd3Bh5kKnWEZ9GynDeLqZWWLUPAe876FdO+LHQaJaBHCzJBrnE9txLlp6cQ+V
omcylIWADq+Z2AgDojFRQ2Cg9Okgr+X7doQwUQiIax/XLqas9/WQoJdOZdX9uBq7
UBXRJYs0+WlDiRMxiY9rtDa2t3tA7wsJTVJg2fRAX2hQ1TDXaOt2Kzv8nItMM1eT
slA3KyqGqEmg+/cxCBXHA/TOmv8XerlwwBU7S1JJi1Se0V3T9MKqpZbn7sp2zTNR
CvTOxudXLs2C95aVlzQk4BRCgifKaUrFOoKQFhdPw4GsNUGjb3a9SPNjCSo5m1Gh
ZuCVpcbH7H09JCQIsnDgPcuwg/JXXu5VwRm9lAY/7Q6NHMRXNmIGJm25+0Ye8x1C
VkMlnOchMEkBmAaEVVXWZMbVEKMtpHYzPiLcJTEoALnKZCeNofyXzCLhj3AratbJ
EWxzgP5fWsZyRu2muu4Yqlm9/IpX880wXd6A+6eayFuQkRxr1MFeRdVxzI0aA3WE
8zf6G8qvXPYNmW8CFYInPVeqDBqEqkVzrx6ZZQluneHaiO4BVU6i8AS59aun4WmJ
lEPStWTDBD5EiStsEYP58yK2jkQHjZ52zwJwQoDQ6GHdtbHBT9ZRj055ATIceQzZ
BmdFOmJF9JYnnzvW48+/KJe3XC7hgCsHmlm0GgUobkhOD/cKG2mCwSmfWOi5NOvK
WWMisQLS7dtjjkYa0/w8D9GrFKr7H7aOArHEnraTsILx+lzpgMyhMB9oRx6vknW1
bokEwB4npti3TQDhvoPWqn5CMlhSyOM+G0gMDUqTfWyZczIbKKgFyvQtNmxGx5aN
SApmO0ZgWBlwnQK/bvWJH+Ycdj/4rqxgF0NT+IjVMhRiW89XKwVAWEqAXXIRKfJd
l0laPS9gMYH5SF0hsqcTekmUpsVWrVfCGW7/Blp/ksAGEje3A1ZHzkCCM9Fa+rOp
zJBmX3g3XuXJGIWpXUObVcqBFDZkVhXEy/HpSvbF6vtWMeedhaWCqnONEQRDJjkN
AjGK0YmTEb+j1DQII1GRSOz3iwKhRHBubTxYB6YB9JHGdV3F89mrfluQ5yNeePs6
eb8KXE2R1cAmugxJCR5NyZPRvQMCtU/um07fQ8nz+ZZkf/1ONITMsZCTCF9fgyZg
i+hobWmNJ9k/zeXb1dRYht8XHhhIp78BvEBY7IBCcYYyYJIWKPLt3Bu9OCb7jPWA
JT5K5fzrgn58p1c429of6Wv5YFNuvdN2us5Z41zjdBCmA5Fz4/fQXWLFpHtxawQg
uKIrO0IkkTIfER/1D3tx6E16UubzvueKaTX+y3+OqyN0zHi/oY//mYc9EZy0OGkp
/GMji2zUkHxHaUCkNZvIDr16Oet4V2murCwM+caoCjhTlbdyGr6JeGZmrCBbpOH9
OJvZ5meGXu+pjc0QcxegCaAtvEG3PilpDSvWYOnmzezUfxkOdyZeUvSJ5V/uwaOz
W7uPydPKyhml3KK448r0iyqt2jaHQI+j/FKvcv0TNIZqTJryX+zXSOsWGo0EFgTF
xGEJBJdB8kInAss/87CYR4f4h2+20hvTK4WW2cmj+y46P3ELpFemnEcnd5nnK8Yq
M07lLSKQP+34+uWCjobjKJm0S5eaJPo/WEWcApy/4sMochoiPdwEzh8kEChL652+
/iCEl0JDybysq1gcm3QkzDlxD6juaQ/xaRdtsn2qeIRPXMKMCCFU5yDq43JA+K6z
k6GaCTOoqjEgH1cMdmFN5k+OpUXvYpsO92KNyxxKeR9LYHZk/pqx7dAESzON/XBC
7vX20xna0wnFz1XE876Pab8KlgvCpDafbchEHLnjTEns9yFmZcD+O1mycVjO/GcK
7PWTDZJGE6qmzifrv6JjJNzHmQh/+sveqaCG8j0oFo19hZtNXnGX+YVVlgx/ip5D
y+r5qVaVt6YMIXIuoM8QLL3J4caVIQ3srJ7I2wpG9sPAGiSkr8xk0U7TFElWFmJv
LaU3xRZK4F3NGMz2aA3Zio1lSOYT88rVnuQSfqtMkzC1J1M2Z5JviOwiYHypU8Zj
/vrSC51SmCtRlK/vJ2R30tTLxVooXILf4ooA9s5hN8Zxf77RrxchAjM6v3Zh/DMT
ECkOui6ZDTsyXLUZLMQtanzEb2JcvM+cNltNUGtw4vaAx65jEJcCeaFIUATcdV67
YPUOvYiXWE/3IVKHhhNtC5fmhVyXVx422iU/H97iEylrNnZd9PCOH5e14t8ZGU7J
umLfhhWPeTucCC386O370mrBj5jN5cGKOiBKMJINMT3s6RwwkzW+keUokXiZBOCa
wUjkRV2ck5mLkonMbOG3m70ovDc9T7kvZE2wgdzTDL/ulXBXeDN2JM5lyDXUCWio
1sYDngqaSjiFfaRu8/Ibfn3V5AqdzKWb77amHqLc1NZfqWxM1OgugUsjSBncCo9e
AnjtWF3ctOvo/muy/vh1pYiurn+l/4ZaKvaJ8jzFxosO6zwRfmFhU+az4YGfwgfv
gBea4TCmFig5sQpEYlO5BmsSJm2GUYwNMhKkHbCdbGrQWnQbVTEtE9e5/GkB0Esq
IdaPhuIvIHRG3oxDEM0qVMVkrI4slBLWQhqdOPY8XdslWHUx0oYZe08I7uQhc1pZ
ej0SXvTmcYS1U/uW8zTzleor7VUaJGQi5Z8SfF7zY/xWUtvjd8v5cOxofeyE2i42
DxyBdmnjG/VENxnaQRBA9zgWXCOY2Cai7GRRQARd5QF0hmeeCadm/w9RS7R9NzRH
oJb5hRtuA95XY/7gkUioZDZZlf1jh/ln80Ts78aaU6+LgZKHAkP2FeznYdpXtWlI
Xz/tecW79uejxGBMM8yHQAvp5S3vUiwu2LNK0MN8V8C0cfhyhV78N/PYqDsyiD4k
Jj8rcVseab8DTZB//uaTDksCPHnyeldzrXRJ2gmHHdSkSrEvk4jgP6hEdme1mPjK
fsWPmndIGUS3xeDSsKi5EcQim0CTReo7R2BDBDpMN+PaZR6/1w/hT0JLY9cL3Rol
UDUhaKD/2MwMkYUxkXHUOGweL/8T7aaWZ9/ZHeg7KZwJmkRByK2seEsYjjsXM5vW
BI9+zdAycDebDQ0Ay554khDMmtmxrmowWO8hUhn8HucUZNqTVbzC/nzkFYSN5GHV
P7kd2VPSxvw5qcFiX2D9S7CqHALGDU+Sc9nRJMHu8jw4J28LZNeUe5MyqZPRFR+l
bpGua/og6jaVMmwgBk6YAfMnU09crm+dsjq+KVGOXVBKpXFpAPGt8f8Av5mUT7rp
GYDAOGZinqMt0dRZ4QsmEyDRuTT4CL/xaVuMiz5Tzqf2TjdUD/4DxSksZ9XW5/5B
QioipbvN+qsPd+zYex8c818OjX7YGX7FqHEg5aWDkS8++GRbZKO8PVZbLQbzutZj
ovcfASz4Bu5DTP0WQBRNHTEwrNgb16BrYfyAfxBHHrdJbe2lRHowpTEBiNb81WLq
9iZQvJMzXjyE3z26WsDvZbLWt+vEBW7oMaFHo6JfAjtLQR16vAkVj8fFeVKrwnVY
ThDU0Hf0/mUowJDnQinGpzFCBlIR3/S0ZgQtHFuXCdcNM1Ovh9JL8URH4g30eWrn
U0vleGtEswbB0tch82TvCc1n8n74N0GT2WstznjyyJ8FB0k46PvXrkQ5qcXD4DFV
yv+V7a4Cl5z58xmnxX4P65qo13p253l9P37xgmAODeuLoY9xUKuQoFEEqJgMYtYg
cLW2frrlFe65R0jjv159lcGaIxsHZ1jjib3FzyoCOtXzEaPPgb9eDZHaERY65/mk
aHrdv6CFYzG/dCUfn9H/3DRS8iMWMN6FG7uNmMiy5ddLafsDKpJFRKkq2KXpiJkr
PM6pqnQRWFfg/7AvHRcL0vlD9lsIPTJoZ8jSe1ei6euJMTaw4vuxhJn7L7KdbpQg
L3ygDJoM7zr4jGcVjyRPmVY/Yxm6DD1uXPx1wQlLVUOn2Ey+lHBgVZmV3GQlMXYM
/3hX1KM38L/ozQrDcld8MEVrwt/v84YGjxwrO3pHSwv9jUjILxU9sU7aQ3jA/1go
1MNRist4kLbfdNUo+jf2hrCv+FZUMdcy09SJwz/cnEEo0F7wc0qKwoSakoZm9CRR
yS6Rleaq10ffSfIQdvXkT96WibkiMbLZ9MiKzRtU0eCoeVjcsJDHMPItCSi08V3X
mH2BARaAvvAjsuMeE4rQnYiGXZ1NxNTOlXJyUURiufJU1ed7/6EHkQGWGa/ZjuRe
iv2mOQZ0mtUWLO5KqFFtTkCL75vZmFxSBz18e7nVwtQ1f2aIH0sNbSi1heSc2RUf
lrFWFJYGQg3uJlhZYvF4QkCN5dTTILtqCvU12qwMZvvvWIMDK33ZadowMJ686bDP
PktubJrB5wv+vgpIcbejnUochUkuArO4tylwnJ3NoUrlxnJU5IvSInZZs5bzrX2i
VTBEDxE76fgGYfnqG2Q7ABeKxajQmtz5vlj0kgKf124wiriUbXE4tdFCEVhzLozc
/Byy4LVtUChVkyBMQ3GVpfyosLElJQsVLygAiYZEPNIxTkdO5cgUSPYqbPzmrGbY
HWyBLlVaZIpRKeWRvNgRbwZBD9fGRzu+cIXmXJ0Sbu5x0Vlf3B6gDCr8ctS3viUG
t823FlSybqXuicKfSnFxTvHdTzW3boa7hMoV6zqg4hhTWyl8/3LPIhNvKepqGdWz
gB/K+1bGStzJKhd0/UGGIckDsDbpGdGHGXRaBadtXJyKSikbPPnOhVn8K1Hbs8c+
mMFXHN5IrWQpaYYAWlbwBO/YXCP/NfbK/kLiPhp2sH+7nkbLVGFxnWVJywZPWf3k
aFyoy736fwqvPi+VkN1OD1q7MuKoL6nlrHp4YrsNFIGcUtIhvpqp8kFwNKh43beL
DeFrtatPUOuJj9rnlRkp590IEvSfeOWFc+I887HnjfTSoF+KhPa2GhVmoGCukqd0
thfKyv3DtrP/hJADUbLqv8+Y7l0oozeLn3BYQ469IdKYSsJmZ8182tz+3P1j9YHf
fUeV3YxPHg07Z478diS3e4yjjz3zMYU5V7tMe1f4eoJqTutp+izZ5dv0GbyFZKjS
PYAMFcJBTr1zEPA3WZnUDyZcpJxu2/p1kSqC9/TF06P2aXaao7fHPyK/XXNh2EIy
bUd/PAqSTXnqGJR+vyswElg7qPnTPdAKDKQVSsth8UPzzdzDg5wXl0S/gP0U4n+K
2bX53i8dCs8upiCiae5MuRyaOiap5FHnDQs2taIOt2tBwGSJLDt5VDP7+xb1Icxh
OEy/U6391LRLAgPYMBrKfztuLAw4rrTqSSnpfiL+TouUxsMYHx3RkueNK8YkkGsY
LSujILbn/0WZC9DXeSK17aNnpZARZX9iMI1CBphDVSMBVSmK7wfgW/aa2Yg77wmf
uNVTv8gMHYB2AN05jqAHDzSo1oyrySNKR8qot0mWwE+J2W/OdRWwsUaR5aCOIZau
DJRwkLKc9n86axP+zXZsts5kK1scgQHa4/EqvgeATTph2e3yIG/zQgGcVquHxJAD
fxgNpheHM+NjXxrumf3T4LGLa65VNj0M2SmfHEclIbnHjKvvH6vTDwAgz+ZqvoJS
qpZeX+ebwDnJLtZeqSsjiyQjjJ1Kkn/4qZiCeJsA50DpVa6f0B6vJOr7V+obqE4/
krb0LF92rBtQVt/2QiHS3+F8HnOs4Oy1du7NnN2Z/4mwk/J2UC8IYYu/Gk+9vXKU
/fkbo47ooNZOiFNudWCeEBcTd73I9JBWgR1uu0oFALm9MzOwZurwJOe6xp7WkzGO
CxHVY1yjbJoeZEEUtm0X7Gl4fy8mI9g7VXosk63ZYebFiPxo+yOOPmE8oCq078ar
wBqkp58lqhmgo5nwzas0jg/Q5RZYg/sYguuHCg3s7CFsq4nmki6WpWFWFz/6oY4Z
/Rrh7MEYJGmX9Ktsedbj5T3KBUz/7hC2Uz9rIZwDc6tabip1TZXWOqR1wR25wrjv
Y3V61StFuXEQ3+aDLVd8wTV7P0LsLWlRJbSvVtyPj1gz9ZajRaDr8gIKlFtxq8+a
Afh4346zkULTgH8bCMD7jefv5beq57w/ZcWmulz/Y+x1QQjpC5CAouF34nRyPVe1
NIGuxgpftAHhlANTPd7YyYkUU67aqQRXNzUmYdWiNGsSa78azj/9y0uKRaz+3wLc
EHPOlh0LB4V7WuI9Udl5rWvb6m9EUR+yvMCLzE2+7OaClM+8cMFEegztP1Pl+BQz
CiPfSyrbNfiN+IPA5BVr1AfarevhyrT7+oP8T06UUzPTNWGwInT7Pwb0eOoHFyAM
95VRZnNHXMSjsiBdcFE2WdvRu+7O+zc9Bxiin5lyzy1XuNACMWpjNsB+kzEVR+uI
3fyeLOSEUAVNgEz6bYtIrkzF04pA7Yj+JzcY0eN0vYyeTw/9NUulOR2i0kdZyz2D
bTnJ3G4Q6ksHYl1o/bDERiEjba+EP2drgYaQvhMGGhP23ZGTevRL7xG/USX9ztLi
zf3tvsXEe8yIlfdEN812C4Zok3k0UGJPqpFvbZqV0LTd4CSFfZlhCPh9qauq5mZM
Bb4/qkMg5HewCtAEz7kiBfI0smwOr2ROTq6YmwosLri34As0pGqAjntuQf4ui+bT
Ftbx1fv36yzFubnKwORMgHY3JQwXs9EE6Gmy/fRVqkM2lwDSeGrrQ1mjjpYOL8RW
YQIkHApcwLXOomf8tMnr/kwurYtWd0zECQvcFxkRDrmrHDoreCmGCerCti0vakg2
ldzXeAunWpOdwKy12w/tQ3P6RM2D62eD56Ww30eNshTW6Qd9h1Tp3aekQ8EKJXc8
60NNQEpT3ulpwxQZw6FhOfC67e5GYQ7Q48Yfw1Pf7BZSuwhzN5DrSgG4SaTIbwU5
+jWOklVHoYAWFLkOzXeDX2vm0xtTY20bTQ2wMItnquPTZX1PtaIJJR0qKFVHG1nR
Wpashq8bTn0UcxneNPnumn1JQJzDQpCZigTMXonMF6u1bvqSZEFLq4SyrYHRJ53l
BD1LLVPVl1MJautWLp/dPV5i0iLdtYjHHcRrYNMzdU1hua5m8X4y/SA9kGO2B2au
IJlcGW8jxBP8qTo80XW6wXHD7xIaxy0+/dCtYg900oqY7a7q7023xgvuhiB6NbrT
42s/l4x2lCF7LxbUwNIJBln+Z6dlODOTHlOUnrHvG5NHE0f0R0MksIRSyzX9TRLS
X/77rV7HQyW05i+ZHC9L4GKPHprjU9+7fdj1OSoeSLVVoyoglV3whiAk17A81jAM
j+IFe/kXlfRxvHbi0KZbLKusO1rnBzhOO5HhUn620dJDeSldFnokCxIKGIxTbugO
6J6/B43ybzDVOBLsKDXtYxHy3qn5pYWee7lIC0LiXJ+QYiXs9puBxHKxWeuiaFE1
naC8Ta3bveXM8nsNNGOnONzph9IwSKOF7PzN9iEt9DJVxLer3nQfEw2QhAjUemba
RFY10zzSr/jV58jOF4nCA299+6jvSZ8oH+LRmG0J7PgSO9rtfpLh6mVO8lKKk1kP
AE/4wa+tXgZNxZfilw5nxTjLRxpwgp6gRHqh8DJCbRsKzCzL3t4B4kgU3Tw1Yhcx
dJ+NhfG66o1bgYQZp0nJ9aQ+EVYFiAHHCk7p4JsOg88gQOQxtmwPjKMVr851PFMO
cRADwJBVfDB5KhI2C52E+8WBaIYVpw32xF3TgxnF4KneWZo6XEmo1F8R4Sta7qBk
9TjACmmMqwQ9I7LMvuAwAcB2qEO/f9NXF2Xg6FSjX6Bf/Fcnpq9PPPGzR0UnJu18
0OSpUT7waORiqg+0kTmep3LeYA2yW/jLBNGdnns9M+a/gl37OQnA2lp1u183lUnS
vaKQd9duBuHodGt0DgFsVcdtCXL1PuphzJYbR6srA8ehJNGEBhn5iAEkOerNNVJU
oxLp5FmJkdfWpipKC0VkvMsest9dfbLNp9XyrrDyTwxGpnvJ5tN7cPr3l34WuiA1
2J37ZcYRhfedkflCVVARiAXvP6YzEQbdKB7IFFKw2EHJsBAfM8y0xNgDbsN+0lZT
LRZjj/ZV/7/f23MIUiyhtn49opEsHNUymt6OXQw2/PCvm/b6PHaOTYHfMP/ZZC9O
xoFsPICWDHmb1pOuHmQZ8152MqCUW7qigrZx9u6/tDLb+GAau4WOiGtmw3v05dYf
AYWmHEciEJXRCJx4DjYf4/qexJtZ4gnmpB+qIqzMMKQVQk0XR3ikUv7is6DGItT6
2NHxsMcabuF1bO44tcZ/SbnXcz8LXtP3Vy7uF4o1BLUix63GPWAXzVgoh7TFmgjq
LiSit3bgTF2SbwHfTu38IMwBt86WAf3OnpHZ3mHvP9QVHtywON3beaYGMoW/gVjY
vyWB9hUoWslc4eIfg0kkMpmzused/8eU/MYj27WtGEvH4RMRhm79DBEF/EOcfZju
NCPyJl+khbgPKdo1jUr2ZMpBc+LszHEOuCX6HBU6F7g1M1AmI/KsGLiLnHrVCyc5
6KDla0dQ3Q2vv3P55PIl70WnLx+JvHCdcbv1IVhrriLwZhqIJcqNGkWQCFjVaJYd
WWqL5VmoAcJRt9GvwhYze3SZn642fhwPocQoOKiGnGpXhLU3Q3EmngJmr5zR8Ejo
ELHGVyFp72qsLU9/NLWjR1QPIlIiomIKLjQNnMkhdC32/4bDP2YzZR9flh0ogd3v
U97RKes+teNqTiN9NcNO2+xXKgq+PXU7onLbIg4iWVQaz1NpddIxGMgsM6+/Bkp4
hMzQ6Sc0Uh+uH3kThWpW4WltBlolKF27q2Hc23JnHPpMXqvxvYGinBUmAW3Evusp
KhEB3U4TfD7EyCFhBUvnNbYie38HfybD7AqP4ezKpUlF3fNPONdB3I0h5vN1gF2v
94mNZMJw5I9LWGomin5QpoDODU8u+tLDTEwmqHVNsdpO3vGWimAzGQygZHKbCDqs
o0bjMgyDB/Ioex7vCMyk+/hGxyj5Y1AAy94sis8mJFZIyxzNdDdqyja2q2kA1EH0
09KVaaIZVOxllhDBDen5h0VcGqFUjwtonhP4A9bAfMl16zxIgRprmv65Wy8fqo8N
JVyhTlbK1QdUOkT3gULOy4TNc1yxVzox9tcPLhDe/TklATDYS2VRmZXNwDb57o9j
JLL/N5nMvscwXdEVMPXCQkrNDSITXtoZTqT91fSGg/8UVfLztJ3vwJyLlzoA7y9t
m6vMAQn/63WQdRZi/F+RSawdjBY14vGXAMweAzn2pnvlVLxmkSn549cP3SNHgH7j
R9lOMqQ6VCnk9VIfgh80yv0E73ImBzkLYlmTDv2FBTBuehFBaYvF9BY9sZpgpBUq
EBjHoUyA7oE1pckbffAdzcE8+jRMhLJ5dzOpTALu10Vofx2OFsdOUCUmX8F3Mot0
8qYVNFb7VC/uR7w8vyKwIK4TtvS43vix8rTbQkrWSaX0jx5IG3dmPAneaM5A7oqv
qX1WHkDPdc44wY8P3Y+R1BSVT1OJwIgmqFKLRKj9Ubacn8CWIUy3ugf0uxgkYZif
KX8H+V2kgLOYxeTP3htl36K1uB+AdBZcsLZHzPwRO5+pljAU1mgF7h4g0MH5ESPg
2DnuPI1++UcziHGtVdZxW9nJTWQ1CcZohJlNE72rY4C2CHpy/8j8nIB/ySGn0IuB
cavGkmLiBEa2ZQICut6GsCEttq7J3DuTT38fwgk16s8HQvuwHAQXKc6GSHk2fGqC
+Bi9ABVUj9hjqFSMdqtptHTE+eFZZ0IIY3L5fiEhAnml3/6yP+cyuUgZWn3gE4rQ
Xj4PhJ3T0bEde2L/Ryv3udflvRNOWDWfAJnnOmT60iWKfpxa5chzYoi0rLcb91XQ
+A7EJf6f8n1Wvie2dD52casDzcR/iQR7PQhtK8d2xtYOdNTfnpZp9nXRuxIINxXB
whXVDMSv3o0Oi5+mVrVC2DRgB+G52NxfKlp4oXeDbvNZxxO1pJEw5bDGsr1TkOeg
cJcEeAMDXrwRuXQwMf6NoR8VdhOos0xaG+feuhRrsYMfzupGz3oXZhlJ+Cmip8mn
2wMimPrlPOD+PFXlgkSoc3R3+5UgH6qsiSDw6qaruJPgmnW9CMbK3lMonrHguqne
Fh5ayHOxXKyn3cEQTP8fO5rZ92GryArR+pqLQTtg85sDbQ2aL60HdBpjpttugxOr
0+yRqBqITFgHy8r9vxqebZ3gON5RX97GSPABMHmp0uE2WIlRXhv8wx/4WgcsZuxf
5t6Us6mZKXe5AaJSriTPb+DzPlIDvicP1DPc55z5ZgxKCz/0csx6lDu4kkcd/YN2
um+GiZE+sVwbMiLcYm3N29/iLB3Q+BpjUuFK1N4Y9HzCtEBEaIKYe36HW2NB1Urt
4IX1P+qMUDGBQBCbFkwHHl/UzyhNN75aaFjorBfwU8Knp8y9WkCFRi4n0wDWbUKf
KHbjUzdX7J05PKBDrV58Xbq44dEU/cI5ELCCD72CwI8e8eB4/wEQKfpJHhQsTOWQ
eQDFSWfTM7R1R+3z7Cuze2iFGUiwAV3kaVteWpSfBkM4lz3wLWxqqgQxo7IkLFi5
8j1z7PAtMlHbtQcrmWzYkYCaz68XfR5BhDcGclC7dknduW/SRZLOuc8Jp53Qvzgn
C112KZbpCOaXjHvOU7vYHiRQJgqnnmQHKw5rTOYqB81iA2oENvQK3SYmxqciBpsf
ZDwQqKwTL8F5CJ7tTHdmxzNmYSSRXWlLU6CZM5H1ogOb3WHkxh4JN54/PEZX3RVO
9y7I8Hfukp7qiHzmRctZxVKRAEiQh+i98+m9An20alLJkhpIRPXip9g0oEl5HsUe
IAwmZb2h0bmofqs9bK0efosfXXpCuF3uC6CEU4u+T66uviKHAZd7lJBQRblUnP+J
rek4lt8Wn9LSRtut7zQQVRu4ppfLVCxyfftj/EhmVym9X0Xy9jysn4TK3wFC8/65
QqkSTnrBfoVIRCudFouhao4qkuQ9sBj8O9pZT8erbCvNKZdcR8VDCpIPT1Sr1c37
4hoqZEPtP5dCtpvrQyFdbb8XSfpaEYCwr8SQM0OZcn6ORc+kiJ98YwqkkPDMfC8E
dT6qiRoBFmOYZWpZ3XFwZsZLDZjoA0tmYzvkkZO6t0ZsZ1Kuu6azGLghoIVy0GVq
96O1olYOwH7dcekVId4pndmc4yPyQfT5lRdTvTP+RtK9xUhtA8/y8ioE7i3oeaFM
et5SWq8fmtx7AcI/6QZrFhen7Pu3ecCD19R4fT1Pe8/vHuUInO0DOZw+7oP8BeTc
S1+MNIh9OSbntZU91TN9JpVD6ol+H8njey1/BgV0XS3DDAYHa5bGTaIMk0J20UXR
30hq5Yb77YkNmYpCo94JDy52FOu2cRYW0Hcz+ZKqdV4ZMRKlygu0iFgfMaTGeywg
NvMKVp//fCd+q9ZSW+NiExDHj5+SrJIR+lMxXYgdDUlPaC0qQa2HRnj8HCEA5CYE
WABrfwp3uI7zXLCLVzBHs6s+innPeXNSmf4vWNnGsOmKQJZDQiiElvol8ZvSz4ee
NyaQ+k1EHIOWV3DE4qDIxIwko5qY0e5EiPJZnv6jwUZQ/xZVeFKyCbRrfB4E/e1m
NuFL8hyYyhZyPuVUz+O8GVSxtx2edcaiO9b4lvbl6LPxZYXGfccKHlSHnjPkYZsX
Qnu2GUJJ9jV84I3F+X8NHPHi6bJoqaEi9m/qQvyTJDpbHEyf6EBnet0Tqp84opMc
/fNtn2rf6hLBd2uaz0KIu+TZ/JIqcyDrO5wVF797hDoSqUDnNvIFoDQYccLUExMt
vVjRa/L7N+IWs4FcvtGy+0I+cXpXtI5opOG4wSV/4SFU+wYyfIqatFymf0sj706K
EpL2tl+vleeKySGnpcTas8kr7Z88+wmM3R+gYVCJo+N632arSCKo9qWyu7oW4NjC
yO13dUEAwAF9YyMqhHc/ZkVUpC3XtJPvnYLZh4Ek0YLch1J7WZA0tgBVyX7mhcX9
bBDRu8SjkBE1/3WCRAbIFdWuo1jeVBxAOROTGig6ngm0Cbs+xGqzkFlxfov/eDvI
3so8zbkxUSrLUeENoPQh2Uo9bWlHS7KuHa9NFfweB+0P48TK70tTamPwooaPHjkZ
tynGZytlJxixYIEVqpxFR7uHPj0WkRl6W7atTMNlCB0kjxkr3K9HUbJqfK3JezX2
i+TISPwxXpAiFlOeWEwVgtwYC/SBeMHyoLzVSHO343ICc9NZyNcXzkeKuYqYt9Vl
O9H6dXSDRjlx9WwSmbfjnoYpEh6uuNXaMIlRq3B91oYuOZA3vPMZrayRKqrve/gP
xPupTXLqSQ+s9zLAsI5TkkNFNUweeYyLd2AAUEC0aEvpoMU86NtyjMnf82W+zpKh
hNjyyoojkJFSLiASIfuocKbEYIepk28TgdYU7zfice/+SbCNyHsFXpy+5hP+3nBX
oJPTLG0VCdW08VME84NSCucRQUoAgVfFUHS96+Jgz0ZPyQDSfcKqcBoGqi1tkv/q
CUqH5UZYRPfH8MDuXhBn4Sf2VMVr/HdZeSkrJQFlST2SxgovaruFzioOBCYkuhkJ
iHwZJpukXN0RN43aiDfAbQfQ++fHm33ZsvsbsQfxfBkBHNpNcVVppfklNG1Zx39B
34HhZbmk+LdcZbbzKgUiVeb7UlUQ892cKRloJdsP72JRPhUPHSr17oBw2Gqin+RQ
LdD3VXldchX53izxO6zErrNyl63yZgMewSvDzv18WNt/5ioj0KQkxmDqWtEVkru3
YRVtc9XgNcG5RLAf5tC9BpU33fyemgvImAJwGn9wry1KHYThuDSCN9NkbrM8ZKeR
8QN3+tJjYbZXZyoh+6OvQZ3UyauQWZukftWNxc5gIp415NBgkvgk8BepUvoFO4d+
G+agVvitjBhyWCQHbbsHL/Y1uWk4TW4Je+SyM19yupCIQqNLU8Exop1WTMmlpSGv
MFACEzgtgDZcqI41JUkwME6CPlCzEfKWmCE6JHv8VIKPXY3TVtWX/lpZCp1ZdLCm
mXUNQAfOj+BWzrRYx0UHmVjFj7NJwChgFS9/RU804RM5fYDkpGczJpH6UQnvKxTa
pRr/aqsSxLenjm4DH9eyrRxHsL/qhRvGLvIyRyve3BisrMWeUsNZtEpla+1tAyGN
HL/cWDYWwEfFA8cZglE50Jaw2TdeTm1MGcKDlhF7rwI4/9e9HgxgwWYad95MKdBn
xE9ztK9P92gbNXsgWrNS/aomxZp2g9IbTeNinrFua9MO4baqlLZyCxTqCle7+6rA
ydf2eunEzwZNGFLaFmJ1fU8n3ygkljg9M347DARzc4ZttttWeLQ3RtdhqQE8z96U
iui3QaAx8S5UbuEnIulsL9E2adwPD/abI5lXbbGDKEJQgg+lHcbRfWLOhbH4gdIF
1Fhqbx6KexSs5tozJP8EShSwnOwEDJ/stcrCjy4S0Uql0NYbJAY1zr312Zm51s2m
JUR+jdYt/NlkHN+yjVWHBD1vRmROeLm88/AuTzi9iThOPD5ZZYNmosBAGeV6jtZW
gHzGQHMnxwyiy2QdYVzfdYSRfJ3r7keezkw6sBa0GduzR4XAMypXhcSi/e/qwkeR
8GBs1X5t2lQ3tHFscxSkTY275DTyvFOoIzGU6Bq0lraw4DVv3QgoSGVWPfqnRQqb
65uP9iRCPWJDm3plwMgk2ExfMWng6J7bT+R7ztiFeSVDwq0OqTWdxfqlCAQEtpyl
UxQ9yRSDRxg214p/oy5VQtDqzgVQC3qNV2PWQbNJGrVySGN32QemGce4vvvEtQ8i
jG3dRWZjxu4glmoEetNd2TnHVWltp+1w/77aTHcTe55tKFkTPrLl5vsKUfHJuYs5
zwCo9G4paXRUQ4LFaU4Vu63tw7QReCjma9892UG3pFGrsgjBdKpq7aBIoXYouugu
a6jJ1PaaLUZrpThZcmIcgGDIWPtOaft/l5Q+RK3zNajWPANHcRYzmE44/Wydi2rt
GEjPkK+WLHLPftiB74r42BE0It3HqDlwfqeD2CSmYBiWtsL983eDRW+8zu2662Eu
LgofDWSzEILrHt8dTMnoKQaUwVjq85CRJ+FjXFvp2XX0B8Us3Wf0/Mp+WWD4M7Dw
VW4m6lduSm4GAzyNb1VHwwl0o6Td3pM9stmJF7YBAFRMVIt3paZ3B9Fz/NzVPnqK
CYX31O71RT+7vB9uS6or0RdvmUaltm4+Zrd6M6o9EsJ9+d1JZO8hKgo0vLxsE/s5
mW5+TT0Vbx0QVF3OVBXsa5EBjDlN/n1TcJd2+n9DkV0vVUBioCW8kbb3h1i3cmi2
tDhCJbuGUA6Vo6mp61d0gvzQ3sJ3cuuuptRINkOckd87i7KvxYi1tlM2c/mt4MK7
Ssi4uXNXQP8sI4FrZZ5zTjIx9JKhKrBfIWxysYd25tNdbk0IfOxuhR06kKZqLxu2
Zu11gjD27riG933pIeSxb5qNdXsjVqqfMLhDF82MBdzLrch5aXyHfVcR1qBb8ecH
jryRtTgZIqU3Q6X1P66s14n8TaYICin3Jvykdqk4NgeARrWFuRr99vqDneEfBLYK
sqiyxEMUPyE4mqpYo37sGPfAb9dPTmuouSXA39hlj62ZnHsU/SaOpNoxDzLoqr+8
xwofdRJxptJj2VJrwNY0mStu7BWNRuch2L9EP4Dau7/AhobTEBHglKvmkJxNqykg
z8TUX+ExQlHENh+K9x551Uy30VlcsjmSMOck006xb5gkcG9AGshfNjtb3dcg3uev
JcqynNKhcSJaLAh+yIYc5EPnAnSUzyUzj9W+yZPRN4cVzCqrbm6bWS+tPSO9MA8q
pfdNVZhIxoAISXBV/sv0Nsz78AxxGZ55Y8s9mBkFzw4sUppKhgH0vP5ZYcu8opNv
8k/iP8Gcpdy45yE7TnjZPOMKUKFinZVoO6ZtS6RqzB5NJW/sMrgEbMvmoPibJfnc
ZP44NXgO15apKJl46SY7miHYXFCChl5xVmGWccM9g2c88iHEDHcQKGjtf5qTxxwk
2OWuDc0Cp8/pAOYbj3VmrRvE9oieAWAgaZs2YW+4cqdpFz11Ows5xDw0bN7gOAkL
+reTpJBaisEBeS6pp/FndDl3Cd1FQkhS0TqOsVkwSbeKpCOKwPesCeSVGBUNLag4
0UtQmdmgCqLVjUB2pUDMX9wxHKpuIKRT1W589vKSDBoInEjuQ8n9eSY/EbwLusVd
jCv+COw9dde6frqrHZnG9IVblII4BKz4bwYLKrUQlvcxwtTvgb7vvGjB5DnaNJCO
fnev8OzjUbR7zmQiMcFA2yaO/FuF4p2vOrzBLGC3F/DlcnFwD+NmqGseMmORVrsz
GZuzUsGm9nulUuI77v0auxQ3XzRzXXNhowc8qTex8Mbc8fQ9elrjcUd3OgcU0cfr
toYZccWZiziMrypM91Tk0Yc6JVjpZgLT8A5m5jsC8oV3x58WqAIfHnoaqHBpp976
MLlCpX6eDso9vkLhL2a0iNaT+v2kDSxf8ubRxVk2mKAo8jmc9t84tzBCF0QEonzL
jfrOD393iJhQYACkcJiPzjab+zUBWe6+84bc0K0y9+DPi5ckmPrjpCb5yu4iZzXe
ykzGT98JZu0dyN/PB90liI55TQN5QFFpo2WTdIS4vgAt9kI08lGF/8opGjDexh+i
njSIt7YrnsMZRhMWe5CqWHsc8Tz9FyH7ntQF3Z/CPuAJSpKRJXJ0YJOlSdD580Wz
67+GlE4C2R87SqDX7UKnZpM74N3cW6aOH92yBzq002hHFmnEyqbpirDAJSL8qS5J
+KlKkKHUhGEcLL0TsibXGedJRzTWhSkBY0WneWiwrLeA9aqwwUz7wPCZk7Wq4jmZ
nf1YN9RWH83HGws1q8pDe3cVH2XKW7c4VDwC7QE6xrAWRZRGXLTasvxtw58D/UMl
JcwdcrhmB8EfoDCF8vLPZCsk0JWl3h2GcjNhAnAN6yLsWUhptZMqAmj8X6USVG86
pxjtOjedYoY67Crq8j192GdJWCZVvGhHd3GB26xfxL/XreqKTRDT+8rFXIyKUg+J
j7kxbtD6ZRt0LW/bmFmWKOiBKMl4s7jb/dTZUp4b12ferYuH/rQG7/OE4Kr62Dog
abH8ztbddLM8DO67H+pQ7hnpxAGZNMhCI6Is8LcwKF59pdJQWnZXUw1itez6Wlfm
1uWFfURqY/UboUH0MDB11rtmfiE+YxXxWr0QZXwHMcnyoAtFqUK4vqdJmJGeJREW
0fvt9Pl+S7Jy5Eho8ezzP/FkBFVPB8boY4iFU8h0dNu1F28vunJsKBnQaADFa1zO
jmG3sTndSkXgwgO4mSKf1pqB83ZihJIl7U/PCqSAAwVgXGGFTmB8jsIRXiACWBYs
BNJgOOaWHep0aVaVfIvK/TncqV38Ei2RcvVy4HKE0BKCGVy2giqga+R0TD+9wGNT
7sbHHq0O8hsj7VcowRCd4T+r3CRGt6HzZIZhHCUBbVNlRVtwfnouY9MvHLPfaTsi
PnRTtIYeIrk6RX5ZCQaueyRWDjxJ+2JQl7EJ7Cjzk1ZvKM+z4EwwpCrYLOsb4bLk
0zxqsBPsf8l9a6Heh0vfN1aEyaJFHra0mLaEPnM9YxKkB1R0iI8DxJmV44Ee0XfH
2xlaZMKpk+03boaIierCKuSB9hedblEOqGlpBCcTCxg/rh88xUncR/AAlpgrtx6o
qMFxrbzAPV5+Wy1CuYAUJL/+spS5nzfig3MCgBVHe9qZ+ksiTvu+D4Q4IG821o80
OJ1HGM6+PLaqVp1AW3ftzcPmJ+eWco1HBswdjCNHF2idR2eHvJOS9ZalVZPaAjwj
jSMXOZ9kgwoXZWmqXXT41w85ackvVWo4WImhAIhm4i14dCzbUnWUNTC1atCcEYy7
f5mREXyUcqx8KxNaJ5qg1edtukJ07TQM5xE/Ag8Vn9cKvQ63flVj9qqsqty1sKFE
2tFkm0AWMOseNkXdXPLQtGQSDVyF4ULW2WmcZRtxxCp4Md33elvV8N19uF4+7gC6
Y+eTSUgco5HlCK8ScQQd7JkTZf/aHU7qDSv0wFbqAPfYvNq5Zd7Ul3NNE6nOsGtO
+2KsgjEMuXb5pe2YFb6F+SHxjFMVBxF0+C0DKwYeHrU18aDV3XH8p4q/SiQsFvIh
o3u0V/T9AU/QWx/I7KS00GX2JK99KBfMrYtTEl17no8Aj7N9F51IfBSkxuhdtwwo
UQ6CmVo0XgfUil60w3rQlZFAknCjvqKz/MN+ebhbQpp3nXRDYI9hq7ymzT2jv6Hm
E+tV04ywq7vxjGowgwvPJeNFcFxClB7GGJNFAPdQsCM70Mop3bf3hd8t4rOp69fd
NNzet0uYJfu9LhYE1nVKsAfz9EK2GsPaxTUc2awUXGgplAnIDpPuwo2wTJPTCeVF
kJzfKpKVHg4RD2DhRhs2ejG0sueBbq0DBf05OYgZguXU8M2PZ8rtpdLNONWBvkCr
HK5jmiVydbFsNeTEO+LEma0MYiI/mXRj4+cnniptDb0Es8697BLMKxuMt8woIdxb
HE4peW9cL+cY6pLz+/Qx+Nrb5q+JI5q1IpP4Od/wguRV01aWzpNfT96IGqDRmT+e
qC5M1DAoJFt3o4OTrhrhB0C7EmSaTZdseE2E0SjYr4Zw68Jve+Wsjqx6jwmbDcts
qo+Jprd6McKMwi1+RTlDPEHbTJMsCfHsC+blOoX6+CCssUHSZ2P0I31LbUSRdZvq
+VuFMfVi7L5rZxPZyEHlFjjBtFlVNqJ7qwJNQSfkOtPRs+GRQr64CTR1KVgTkSbd
Jrf3Q604buszdEvwijr04VnibUwdjKU8e3CeztIv0+vN1+QwJv827kIc1vFgJAwm
IbuBgf0sQ/BdVJhxrXJZDGn2oqtRcbDqNBeTSK8d/7FlJJc5r8dMh4bp0BKCmHzg
CFQZyuetNSBejjpeKzehujjmLqVm/AHRm/A8B+0uyZaeww5ZP6HiYTWr0vTCAmJf
53P7BB7R+8HFU2aL4xpR/uk1gNu5J2Fc6/EqynjQ4pWHszY+F5jTDkgiR0Fli2/P
U5ELjryJ3SulVPWOxcqC2LySv0JrX76gA2rcf/zHa9r792sVE+zbXUH5nD/+pViR
/i7GnuLuvtT5nngvwBgm+U6OEmoyxspWjRMfITLyLxb+oR+ttIK/q6Y7r9pTQjkH
P8x5DAa1ny6KiLwXWNVt8ZiCXOA297JK9Z++BQtKDkjuvwq2dHMTOpzZrl206xmV
QKrxFKgT5nmlbKSX/THAmOjpFXGBNvUXXFUMYFoMNi5FuUQk0ngDdnN2beddUk0R
aDi3c0aMO0JV1qy31ybc4thURaAmrVVmcX/41ffMsRLUELRGCremDqHXPEYj1BL9
//mWTa2BXk/TYQBm+q+SoDG/f4DIFr8BPAyYm4aktn9RvfkpgNvAvRypx9GuiSsX
7gXWg82lByH0rcnYTJXC4JfektALUuWohYS1GgvCnKroUNBsk1yhA/AybpeXhRsW
yUqa8vH0lAZf002IVeaRbG6qY3lvMB4fRn/vPr3Ew9W/VNnQmLsYfIW82kXHcYpb
smakl3F93TT2kTrKaBzeZOesUoziuaN6qmPmHmJ1gDG3Pm5LV0Qt6HlBDcsnFj38
I3m+si0cnWdfYQxUejfgOEpJ/qHkdak9O9FBgep1Ra3xFNln74hhDiG1dnnBuwRy
eq9P9hDYnm7R04nUb53y/vi2JRhVtoAify0qiTv4EL1hUNGcqfuZlQdV/XXRuaZi
hK4KJdON/GD7JPj9KXF40kkj1xfBaJv/fFmFX4BWGLfYA01S/EnztmLKEg1o36GL
hMnmLw0z5w/9xYfaY5yN6WGA/LogWKBjZXzcbUE4Yvt5XeCRXYvkABfqC9a7LjFK
aDT4eKFm9z4yEFa8qu3JXgGyc7eBQ77vxEeZfOn7JQTPEJmLwUNnYc1ZmDKhjHLA
U4o3eLp8v1V/izXZn8KfvyXbvUmwFUuBpyvHLzZp4Jz/tNPiCLcVEK83mi2WYRzf
IF2DTL6qBYgdIVmLG75tFU2M2Oq6RPr9cYwxU0pgrP7gmJjAq6kp4Jx22ILphyXo
0ZayeiTaAegf3ZwDdTLiErItTxxUzaRdKun7sQOjFxxVC5vNdDftEHmXk/aWH0Aa
7uJWB7sEZypNY2YoRE+4oH/8fcaLFA93kWid2iPMtkto96kSBuXSQxrKyiaeXUTS
maoESqLOcOkWGKAJhriwNgQ7GEACCf/DQjLqs6uxf9iJYXgga0OGLbyt4GzeUWTK
YCx0ntCrrEr0f+0zcJgQ80Ptn+uBSecWcWDWl35WRf8VW2m0Vb85p/gt4xfgDO8t
7EBDly/iIPQtl2gGX3pZpBa+MHRmmRKuv8AlssdVfYuFlCR8geJHZJI/NFlMHPU+
Ju3hEXmPAwW0QoHV6F1NpUhHBOP1Ly3QIln49vfbbHeBzwnoO8ao6JYoyPlL+F7Y
8GNUSVvV1GcRllg/HAfgRiQRsXF9BQScT8fLKAvSgt7j/3P/t1KI+nGL5pIjyLdu
GxP3mtQJMhLW6HX40bim1LCu5uY80s5mixXyjORDWMnoZJgMZqbMK/hYkLJvEape
j9kfWDjGYXxw7KweEyHbUN20gXp7Ke5txfXc2CN2eySSx0PbTkEhhXc+zlfGXCDz
ZRxpRsENxZnGnhJqU4h7easkfNcE58Mfzwy1I5bIjKRQjuRABofXk0CapAY6wC0d
7hxOIRWIIzS8JGGRpy3FBNWgpec0Usf3jRD7C4YmdTKZ8UqSwvm7wNhdEWYnYp6q
4ukUmzv0INP7v07wWOVU7CSxjuZ2/inbpPPRYPf5CARvqmUqGId7GlJtLAxi0ies
Yb3Db1ZU6I28NadpCTK72+/Aomf3zzLHe9GSRSd1tshig/4MbNBXYZanr5E5JaRZ
Xz435FclpvM1qIzqO/3S9KCcMxV6JJu6WW4041ZvWxpz/PlA+wzaJBRhMRog1zJ+
ID6FraujJwcaI2/8SgjVKwVhcebdJErx7UtpOp9OXeRn8tcBUebVwod+TrIMNmkX
r2HdBa90ZZIAmcKibKZBC7MjNLFByqxyrVZ8wJ6jSpAgqwhGtzg0VubphIlal4kj
DF2C3c7PJ/o9KwZ0BTzGPTIKvgxecvWihcucTfbBAodGKS+SDNjeKfu+8FZheFOg
JJhNmiw74YwAbDxV6J+gnyXO8MVFW30Z4Qleep+bgM5npmIBkUMhKyO6VaohtIjr
trjkl/Q4KWcTd1wWjQo7yPfLZLEpuGN92zuRIqiGeIj0n97aRk/xiQZ/rBQrJ3+k
bXAS778/SO5KNcp0bUk1+ZuWssg0EoOLEjrsyH70KTioLopksJZaa+coGb1GBECS
vJJTGhhB2g2hW3JCopTAQDCKE0cjM0tUPawphIsgvTk+35I47Ke2IM/dEqxUGS9h
EIuewEj6QUDZXhaQL2n+PqkKW38CtQq8c9nmSHwDdD55zsVYbVOA8I3/DtEbx6Gk
6rAEntIIbRxTYoTYSUZXBRbJPPpsatUjejCfqk1qyANeANaxvDM+joafckj3hOWG
Z2hKsEghAIvqn2MmZ7NSnFyTYO7MBU4wt319oYmvoDrbF+qB9uBjmdNW6QFbH2iF
k33jdPnYqfFL6xJuioucG6JKzd8v2A7h3qxpONfvw/ie+PXY84ptJLssym3xvfoe
biGWpjNyhg12y/kuXVJm+dd9puRnGV3QmDkDUFWOwBG1+ehmBWXm21SDVIZv2Ghq
gUITMFpm6ANeASnc8gdjqTh5pf/uE40Wk2AsRSHQjg2Q/9NiSYZqqsF3WWXqD7oP
9yLcuLLHhHX5ZJSAOt6MnaQOuYZJsIHVW8sZKvs0UyZ5opVm1I/7vxgmRb0A7YWZ
m6WjAb+rB/iSym4Cn42GeVWdjpM0j+Rh3N0l8RMkrAKDLc/zb7wSA+kA9zUMxjxE
PAUQ6+pU5sVKo91quy1USnokj5bHUyMwSAN1MMyDLUtcaIdClFa5pBnW04/w26ur
KgZhFgHcU2kUK5e/7BDg6Ot0Y1xuB38EuF2D3NZ3/0jFPyHHidHaAvFHBC6nzN0t
huu8ObEiaN7cCFXXtW2RrkA8P1/tfhpVgwRVzO4jxkKO01TJkWLHYzvF0gD8iPPZ
Nn4RT8rRHUbxLcFcoI8bZoikj+GINVJzN5ddeLTub7sacrJ3ZmWxUszuGzOKnngZ
Hxe0yrK3Uv0yIb0tki55+QnvLjIuV7l9KE+Kt2L4KMEpwsRazHWrOq/43WZAfhIS
7Tqvk6bH3V4UqpktlzLwBBQIrbGc4UMCkfmM36HNpfcggrJen+Hs/51jBR90A9/9
ykWpV/aU580LzO/f5lgmQW7N4kBM5/NumfC6Vyfg7XrnY3hUTMPLyvQ9r/39/1Dn
lW9L5oPk/s4sKlgPzXnRhnndgoWjZzt1c2Mwh2AqY3YDKi5epHhrovNZwNnPvB6e
R3FrBUU+X8VKPGiSeay5y82iL3vpN/dcq2lcojfHjiaQyGbh9afGAazS2jf0mgup
l/8odJkDv/OU4mrZLQjqUai1DSwqJs0BIzEUWPT2320H7Q7Hv7qzbKzCCrLXOjI9
kClQclJl0CiBBXGU7A/XjxHQI0oFGK431p4PLbLVHXG2mOSuiixR/DDXSoGeJFdS
ojTtCxxkUggNdyS8OH+vPwz1uP3LRMvZO+bJTb9dUAx0MhK4vLWwgMBbhm62ExT0
2N1c7Y0lPDGbDqiGeOsCKRvn68GjaqfdwxaL2Q2+QtvjYnfey9AePKX6BmrTkSLm
1SwrdL0RVLgd9wSO/u376En94YSeNVz2MWKjcwauvt4FDlgfV1y87I1Fl8XnVl4E
x6hof7k2c78FH/lqeXipyOZQwSGFrM/p7LdUUjDuDJKdxUgvOwNJywrmBOZw0vPk
BPMtFyyWqvNc73kstp0RfA9dBMLmCqZRYc+0mLrUYSNF5pLhgvS//uOaP+k9k1lj
NeyFIamw/Zpltzjd0pmkDmiZheInuxNb8FlfYdb+mkn9nobnWSfO1rcTiixDFV9w
imokWXa7EhWxi/yDQZbwgTMIu5/N6C5FJfa46JKek+olTDyDzXFrVaq052X3NhF5
MZPAE8oRLPUjFXShTg+uNo/05bwIQQ6vJeWIGmBn7CV9uoJhwtvVIWrS/ZFUCNAz
XlUndQngcBA6e9f5Vz1897/T+D2nZXkxwGvZYjWGi246YuMCO/J4HnHeUx83iagk
BDVALAnuXbBbGktwJmrNr0SYyumySmr56PrTK51imaNvXk4zyJUdqlqbqZhRvReh
dKxR5UwOFtc6NL4gutDjY/TeLGn2SK3VsAiNd6Isr8BIkXqJ2C46WyqTxZaC5SYZ
QaOfgd9PWA9b+nt0cPF9yzQHzIpopwpbF9p4YFDKTDoNt76pusHWGbQiK2w6snw9
LLFnMCVdXlNiRsspaI0/52MPKuLFhqhgevV30aZFqKQK4K3Yn7T0l3AbN+lO+V/5
QOfZxn+FMuOcv2ABmvzW2QbCkFEXthaD55LBJYVhHJtRgZJohBzlnqvi8pBkH55p
DiFJuTLqN7CWNgVqMXE/VfPipIbTtvB7o6bjuaAXlztWIlv8Kr7zrT0knDtm4XYg
BhcXk7Ldcgf1DN7/cWdN0FT+fky4XUZD+d/FIaMby8KfAC72c2AugYMVdO9kKOPZ
L98ByA0Uoaw9whSl0kI4/3562gDX/LV0Orf/DBL58p1dV2VZx9kdrPGGImvhtNtM
LMwd8RkhliLH4sN3TmqWyTpXlH5BxGVlAdC4POIxUgP+vVuwmXNuhQXm0HxeaamA
7qIZMB6GXqgEk9MQVRxoVKb+vP+Oxd+eV4re69WNKsyrEdzeZrrBShFS2Jbesbrp
4I6H8h0b2uPQIp3RtGthkk+u3bLIo4H8N3t+m4sJgOPmIYDmoZRkKL3slhFjuZQO
5k9HiHYStbitE/wFUZiv1H4taUt6OSOm/0W6MeEqNqIuHoOPO2+EVpy+f0xCyEi1
D0XyM/U0kASw0twzU+f3M6D+TnPuEejtFX6wdea08Pro15TJXsZD13acSVQ76UzA
ucmPDVJEYhYH8B6Kygu9Q9F4I/WLkQxLbYujNGU3kgOxGb25t2mk/B0wNQ/Lsiao
lWeP+sMu7EcMFuFrcyIro6iA1ojxhAGJiq8jInWTbnTM8HpNOxoRsQTJdU6UZpix
kEfXFYmdK1a7n99wC0jM/rJlZ4XSSV+RWD2c65K4CO6Lr+Bl4LwdEPbkNWnmiM/7
XlShAzTkkmJ7iyNwI1GbZLw3bVrpw/HS9+bmlQWY4tRu7rCKReuHUzGXOBfYCviu
JoULHCmeEgNWdIfCHVpuB8gtRWAQqOP5a1b8VfoT6BovRf+Kji4F0W09QosFK0/q
CdaJ3pZv/gSvXNuetkns0KCXXZ4ceMq6PTR34wM33DPgJhD7CSFI3QMlMtSbgY/D
ElF2Qz4VaMm0tsBlRbUIkjYRxXNKQidnWPR69lplRFpH3zxlLZ2yLapJvje0/er6
temyAjRGhGos0FiYC3KLBoXtYginXmraw66QPw4W3a/oZWqxAd3poCQn4Dgf7eox
M5QBZl9bP5ZaurJWXSDXeDrK4MCPw6Z/xYlyfj2hTgjXreJzzHWytExanjq1yZkG
JexvJmnrVlbOhQjr8TCZxaXUOsmaMTgEuTLOKTk3KgE8OezUHZep18+QWmgfImji
K95TQYpattcUGIt2Dj4pQ360hsP6do8jk0IB7Jz92nMj0SPw2T1b5DOe5llHc26l
k/B2LzOlvFyT6U0jkQcCo4LMvFYsAnoNvWYulVlVkca9F3YDpufItZspv/Oh5+w4
rDc92Ghrjq4EdSOXltw1XnZR7aSCIaDU9j7zz1pfr0fX7wJWXkPqUphVwrZVNcbq
euWWmud8qnAEzszRlcHPk0Z2ekRTD3iuZV+3xQDsVio6EXfZ9F5a8BP3z0pKilBq
RJBKzs3aNwvd0A67MX6Lcj9O4KDYS2LT1I4u4J61G/Xowm/HGBAjFX4wOLWksxdm
tvR108Uej2Y27goPc47tJEJ6aTInW5V74TUYeSFxjLpgrzdm7+DuKNzn5JLCS1uS
wLzK3v2C4VEnez31s8JJ1f/dhcJmv3IqwydKOS4OgQcepaCqniiUXHtdjDdjalqa
l9OzKkLsxCQJVEHOJVtJSzNBnSrPLEhsaFc3yXuWXRwdKhUYtoXKIhaB6OEUq+Ba
W6nseapS+Ek+kah8r1sOLIJuU5XlOreVjeNyZ5TR1dExmzhwEdNvJgsPA0mk59v7
d+mUCKsc5a+i0Hwir2X40ETJcdJtHsClMkAya+kXHAPXG6+jHy8678QTu2GoLn71
bHcxf4vbAteHhW1XWrPotBQpPTFlmKvT0F3M0di2aCuAy3WSwVSSyz3X/RtEu9g1
IZDdHmtyIWmou5b7aBZVsAW+FirpPy+2XU569Exqx7V+2UxQNPd5RwrF4t8jKS6+
72ta9+VWWrMa3DJGb0/jc6J29RZZDi6eO3/TygcQ+1JCfI30djF69uUy9Bh6NEKS
eG0AGtO16Ydc2Jkx7JTnRmrrYeVe7F4ySJnykso5OWqsTgzPLeBrIWsHgiuLPwpx
NLhnURm9SzSd0rpxeke4IazDhtONNTeqC0bgByw7tFIuFY3kZ69nA94rnBldaDpa
aGtlllX5N9eWwILQoDH3NEHSKB6dKBZRe3jK9p4BQpfZHacMvtR7DP0QFj5EabBs
GZ8I8zsk4I6QfVz4gNcC0VyHO8g24FLWzhx2N51xKWPJ8I6oITlGKmKRRovnw6ac
eR6d/QBpSL+oJTIaTwzG/wLUAkv0t2DvAL0Su+yRHr/Xs3IdRLgvXIeEeqFqs13/
V4ZyEB3a5MRAVkPva04bBGk4d1HAtQHVKD95Tw723sHBeeUUmE6ChNtge50xZLEl
aDZHQW5atAnt6xd+0uHYk7g2UgJjMU8f7Riy86k/6kXp1YOirvezJrGLQhv+Enw9
aOLbJaGWYOfUWoYA+pkFQgvZ9/hRESVn+4dAcUGYCNqaFvdB/Lv9iSJLNtD8mRWX
DHiLZ1QCUPsWX0c/DsNH+5LOSvtsz01e0ljKeEVmiJu+s20/l/Jccb24a8nxiNXb
TAXIGHA42dNtyOsUrKXXTZjGecvaEPB0B002CHJUb11CBIsRYxgyJNnuLEOWMMTE
ep2jfcYRS7ZEl75ZjeGKSIjODlPFqjsD4y/EmEWfdzPiGWRLKZiMz7rcW8U14BqJ
R//NjuyM2dr0ex9r6AsTF+ehtdmQQ7v1KZBMmSa51p6hBZ+4ZwNAmymI8zuBhm9d
zqS0VygoS9Tkvaz1PCzXUHKFL78KNz/5ZFfZI1vh2TtfmsHWsugC1ge7K2hxPxkj
FSnSQioZnqF0JU5+03icAv0UgsIyU5/6UvlA4jtXEBP7KDfwBInT3FOvc9iQ+zT1
ZLLDoPTIZQOp7ovps6A8zKPB0U/C5FsmUosS5FlmIPatq8RoGPCQYr7bZe/oRpKD
sxHcsMieQZ6gnXNJBrB/ydaVlNkx+Le2ZaKxJ6TZA9SA1xZlRXu199847q7CFmSR
PqOWXf+AkiSlfAX+/UDt8TEaWPtX0ihPUqG1hbz7MSmBEmeifi4WcjaxFzdztWwO
Z80rPS4ys/otwBUZbwAanPjmqE0xfZJFxb74YEk3t9bCFEXd+iLdiq9uUaIAXpZs
TAvBsvBuyspGGTt2/u//cEC/B2y7NiMiKRJbHkr2imG3uV7qHJCSMITF2nTzE1zR
1HIfPVralmxToyuA1mffDTVWO4YCLmVmOcrWw3gk0myJYcf0q0+1uFoKnpznT5s4
tB1V/oBOesx29HdGLKHwDmM0VdC0d/8/6ebAhCOJwzobVAF1L6QuscIVPst1CjLu
VWirxleuHU/AY+zghFWQmKUgEDdLMg2qmi6HvSqJwEwkkqzxvWM8/y4KdUeNboZi
AwLXd1furWgs3fw0pNKLStA8lyDef+LrGwyYtZjao7TwxZ0UuLHB7Zbp9mpEqoba
Ab5WlY/SXKQeCOu/L9H5EkBGv7uDKOFhrYab4wM/jwMnTQsT4xX0oVdP2VrMxkWm
mVh9c4eLK4baEL996eFOWCy6C1aEc9mzYlD+QKarRR8BuXice/YXEp9YIUCDq2qg
jWszCQeOZRh8z+qOAQtPUPp1/aPPH/abIJakvfPn7/5Igmhjg/MoaTcK2yt6tbXt
h/t1E6PSTNxBWycwr7CGvXRnn4OUuxXm5xm3S4F1WJ5jMVZjDg6SM14tHz1gri5L
qqhgZu8A/+s9ra4WqCSHHvQ2XJAJRMRCGSAEboZxqW9utTxayEpfNa1O2hWHxQB4
pVaFa6GMVZkei8EU4GPPgspb3x5aJFN5nH62WM1kRMdO5yGRwLqWPmU4JRU0YF1/
WfJS2vdw+FVY+mqKa70ya4NK4EcIvxA3qAoj5hRQaQIf/3PWYazCz0S5ZE3SZL3N
gDZdwTV2ufSFSU9AOUtXGdXkDqPWjMhKP530xlBrp8FJqSBZOI6UcYiOVzK8oxDm
FjgT2T8u9UCXMvFh+bQvykWTynlMbSQNYX4hF1/1Iz/U9ymSexc72OMMc0jiqZ4B
cZ0bH1d0dP2sLfrdq0ExCXRWVOdkPJ2HDaKBP3m/xefWmfkLnfvTHRgMQ7BTl1xf
VWf3ZpfjyTyCfQIVSLhHS+6bIK0XtgOk+Bztp2td/4nFiEwxG5VtkShpevXa0UIP
/3dNHWnwuKlFEiotV0Pz2chtc9r/cDsWfMGre1mWeW/eTJ6WuotemEo5yRMnkT1I
KGj+iPvl/B6KfAnPG/7/0u9K0tBZSv82V851+vD6KTqXqPvPaAfvd18yiK2VEIZP
FKvoocLmBaSb02zjaHi7n+pOpHqfTsZSOl0Hi/a6ZJq4TCpg+GjrGJr2Ftboq8KF
uPa0y4+QJhjNII6UlbkbGIfEQKEdyBIMsb+srwvh5KpYBEqWn9SxOPm3it5qvqjo
wFgaeI1lpA7KQnc+faWeGOTdBeGJAKrSJnUNE1b4Cr52dDHkbWbBryoWMN8NXDI8
Mawo4ZIuPve2e4R8mZYnAQcNePU9DTO9qxkMXRfO0rG3a+N7AEnjew9Wo7aZR9nU
W8Lt5bFBLEa5qTTIkkdjJ8WC25PqPwmWLbM9MbXazM+FYW3GvA4NfmfSc1iBGDjm
asfkj6fCEgRJjslo2S2Pjw/De+/O5p+34dVNIet75E3Uq1KWjp00u2k1zE9NP9NF
qQU2x7J5CXx348aGxK3XT/2FXGxBl8h/LBoHHNgmDoc/nVC7vsFw6tZlmny/n1Fl
Avdeg0IyMimtvzVaCdSuOVlNpSTY5QbEGhon2yYCCozYKvPd4Gs5Z/a64/1L2Uqz
p2m+0DdeF70IUUY2zZy03SDn6M0jYUgTxMJFa03UQHh652ROupchCwyvcqfGSZDs
fYdw4GFKKS/Vzzw3+NXJb70ql2XSEz8SFLNU+GVTn328yga/dF9hi4MPMTaDTwjb
WY6pLWZjecYDm9p2f05lsh/gEq0H3ZXT0fnaDWE+FtYZislaPUjgLb9340TxmGkQ
v4fa+XlIgDHvUVrm4miHYOK9CVOMN09LcpvrwnDOkkIIyQyxrts4b+6WkJiID0KR
GaoEVi2Ztd8gx2PgXgGskqhPj46lkBdMeeOgMbjGG3rPy4+3ATveFJwJLU+f6Z73
vPng8bbNwU1Mq/cJFrkCBV8J6Y285uT8mMDtcotK3gRIq+NKJbSBgnsmppRP8BAk
aiaR/YoPHnfLYaWlVd9lxqXJXKgjpIDH0nAL7gjsISy5goKW6FtxkgK8HJvATX9I
pn9SVePho8kbCW5FVstju7cjvVrWLh/uwdC5LsfzZPmXMgsuiKMS1cD/AbzhOpe4
m4LlGSRhhgbNQ/nJsTpkMpxfMi6by2A+lOXyXOy2Z/DUR62iOpT2rjVmoTFDpeGy
aHhZmTLKzmD2Rs4J2RfKuxgNVynykP+3X3jxhw1qY/zma/M4yTPUmB2g16R7NjtL
mZvd0tD6tFf4EzBMHXUxLS+nh4iQelJ/vfhh0j5Vo3DDWrT0H06YMbnZocxI+iL0
b3XH1KffoZmiFGSEYrCYGn1gxamx2qJD6mlchSNYWm9+b6CmMa9vHv/gNr35vR3F
JKPXUcWb7huyUnXOpnbhHnp8lrvd3ihTcVRmOm4A16dHe6+aKjjzdTMvaYH+0Rj5
Rytn+ccQ8QWiiwltrkLeRgb6WFXiSk/1+4oVcsnDeoWFRKRD2DkAP1u4L1GXolZT
l70YiyAq/cY5EJTdUJ1ZVcXOxhy6LB627v0sa+Rc+mIUaC1zRRGFwLaWQqyx7EcE
bnEi8pIGltLgGYM0lpJr1Iiyk2l7VeEmATJLb8uICJgZI4XnH/FaOYgsZ2yP7N13
1/S66Jel3Qh4RqAATztlYhGdfsELmevDk3N+rIdgBICEfIhOgOR1PhWp7gRTabNG
YQH7NNP/UUQyqo2Du7KC39AaDHXPpijSbrHNOOAsve6PswNbQdz0BgaqyNf3ZPly
tG6ftxwi92aDuL0WGs/owikdj3xiiGpAoNLG5ny4JAAzQX0yxYJxlYaB7q0cQty9
Nhb+/Be2oWcdL9NSyNyt8QegJ1YI7HsHa4AgT0HDPrDhwgmqoHDEoY6UaQeYO5z2
00yHJWO2kBud5zOYgbsbUUWviTZ72UMMwR9you9sdkDuOAMVZOzIJOYgJ6HbHaxk
BSCUsTMfEQ56aBsk0oqbHXrtFZRh4qEe6/MBzFdVdM5zJbNRZfWKbEaCHSG1zav8
yOX+lS48P4l8r+HSJgzvRVumaikDYcTyhHWr7b2dGwDFImiNlxlVf49tLeANBEoZ
IHUSi+jRGglf6INIvjwJixSj2n8TSbH15g8kKRicy57XYFKf23Gi6EADNqddPRNl
JPsPQJo9YNse8VCekJfRtIeCD+SZXf4UCYVw1vaN7xntP1wZzELjIlH6oGg6UmAI
UcVk4d4fwFiKcaQ4XXD05niUV5thnlwONrMBNTttwbcA0BpGmau2NUYQcPsca3vj
ZyTjyNGbGZbhCrfMNyPQEBza9OS8DYmjiBd+Fk9DW7R+9KgWDAIKA2D3XrJfanb1
B3xtvlnIszBXk/1Bvueob8gjAttn3+p6Af4KLEw/Z5//Oqe2XaHIuUM+bN1UGdz8
LOwD+S7vwr9lsinoqu7NdDTsowJEJ4n1zjiVsPAfPTe0qoQqYgqSaxFYoZIEosxh
L6SRQfOqBkC4SAYjs4ZPq+YUQ2zoy6GXFA0ylvyoMBFf8CK7bPP6FSb9A2p2x2hv
W3PlZNUZeXqV0INa/pIRqVma4m9iUJ9wr3m/x0hk7edY8zhQITLi7+7YuNCQRg42
SP32zqvPu8F/IquN+jTqPNm+4Ckku3YA2+4ZXCAs2aseyVFgd3aDlZhqPBWbTOVC
Bylyk/n1nx58zQ11GbumLMlTTiW2FIYdlTN4xJDvyy01mPw5AhJZqXYAU+ltU2NW
PQEeaSIT1z+I0NOJS5COZCRUxqUR9eEtaNeaNyvY9t/x/+cop0eesXixWgZeS6/d
9tNTAwQDfVPDgWEMrusYcYFrUwFFkQcUZpan78DIFjIco1RLr4Gzj9ccaARQjhC8
gQKY1iiWYrrjjHPWch1FCEj7j7LjXN7RyppNQvnz0/yqGi0J+iWJsSwtxIxGLB+b
wv7bwn7OwPVDAFWac+mK/joSosNLJztYyZe33kRyeoplTeFXoWD5XUFXGHk8peCw
Wbvmg1g0fSxKR96te3AMryp85CYKA7X7Ul7qJycOEp+MJkKBi9KS9l6K+c2ZQOSi
u5fwJtINlS28L4EuLn4zC1OGi7boAKOlSbSu4J3+EA/W3wObftsn5p4UaH8M+rJQ
CRWX/Pa5M6NMakG2Ok3hKo9ty3RQ04GDZHz4BYqtxs1oLvYx/TWJbf4PoNYYTTo7
2XyulPBaoUMc1aowBb0nBbecPU71TSbdYBoE5/I9gOf5DUqjUjFk0HorGAodAJKp
dW1/1QKTPjs0/y9WAblX6GnAX5dKxBZK6dUZLVqhl4hdY7gcpDNuKc3aCiVLWFke
VJ5MY4q/RDNpxNcLVZSNOteQpYgi1SVq2vZlZbk1EUBoLZgdvxBXDzXkHE5XkffS
L941DuWnl0uUfBK3w0EXbPQUgIP8liCEjefBgJLeHJbBMPtfSX0nRE5sTF4db8vl
qQ0qfr/LMhpy9ENyvznsJhWAGyBsCBORv9pvBFXb6Mpoo2EmIziR4BBTbGfFGMJ9
W7K8Zt/2MWHWsRHOb48AnITEc1vZ5RJOt49796Bpc2voAlzUbPJNft3lnnJ6+hJ4
ahDwHaoyiQYgZSrg8QOKi48iYPOwf4esGOgupMQRe0lvRhCLa0H67W2WwtpdPqNT
PH/YQS+A7CKdQbCbo0gg0kg3SEOU4C9/0yhhefFr1uJ52kfS+v65whNDf3dhEmtC
g5GsYUHirkhVFgBQwsDGP3mCHhp1Ll7OJQ/FrO7tNVwbXAbHamwr8gX+jMZByOd7
6M5BrRVsiRbjgwIQUdEAQkAMuJ3TvMuypJe7F4RuQyXzA4PEloSqefRJirY1EFWs
rmu4k3EzND+qqIx4ryD5oJbuh3bDzrzM1WPkWBvKM1wDEz6vNKpCblU0elozX5kc
K3VltsAYvimKs7qfQKgtS7rJVU4Pf17ocyhNMDPLX283G6e9OQrlvXl9c0Yg9hp6
OPPDGvjLuw24hAi7b75lmEoRFaJ2Gm5nL7DgrD7RPpK2HdM3Q49iWH79cEQgzbgL
8q7v8Nk1n+h7pOnZb0cpL8uyTbwS6YQYyq5zXZ1yR+QuoXPzXFGLuICNV7HMYJxx
pUMQ6fDzRaUnSz4Umo6TmLGGzONT+oynoxjTaZoJv2b77b8/kVa7EYBcTHdyrHWf
qeuKyNai2LOQ71JvoVIfRRIR7q+acUckJX2LohZv+E/EM6fGDQpz7CogmArlLClS
GZDQB6rL6Q38gQJ8kYj5KaXWSop+TmGqR7rdxhhcrrZbe4A3AH49rYoX+75y9sQ9
pn5y6ifL/5sr+RBGtVaaUOR5y+b/TFfsxTcbQDw1l2th8L22Xs1xFvGEna+GM/b1
ITpblvlklBrXt+SauTsZDsWNdX3As2KWjfqVwTSM7ayCL+ZPGrIX7YyPMSAs2aw4
+F2NONi4xMFvt1sRqMLiIuMDw6kWzDbsYAqCFGuNQChb+M8l7lPZrZyOMTNbfzGU
dxv/goW9mag9vyad5D9rmuXQbUzGbP/oSd9dqcNLL/JXkzTaPqLa8DWLWL1EXXex
P8bUFusZmODw5uLPueWfzCHkq6D9XUHFz3LRqFCTwdgc9NLmeGVyqU/ilcIt3z9O
QEPPJ5gqzyZXqyrJKzCgeovX96oWJ7D7Wll9SXCVcKGcU+P36ACrSRLHdKLkPlqY
rzsIjwTkYNZWc0KNHUC0I6Wm3iDb7hppMsLRbYJBlHCfr/LRlXGPXxBww4uwh96p
yJXiBl+Yiaiqx1RlDEuF0Xn758Y7k6irARdceO7Fmwghsjt95sz6Iiz5e9731J5H
BcsDGYBwgPOS2Ew5Rr2lBhLHYpGohwaH5mBP4+2kB9idJNrov2EJSsnTgJEpVmi7
tkkLXKTeV3rgslO70WkfybEvEbPLPWm2hWq0SGA62UQmDsaDyuEvbIf041zLjv7y
XdM7E2kdV2j8e8wB1LyYaYoIo1AbSWut9budZbGe/mhQtDwTZfErxpXen/PBBoEj
wHJKRbAiKuWNoZR+MdPUL4novtMzNfz31wMobmcmhQX3USnYcf8QgtX03L4aHwwC
z18CHwwxRIHkrzxymRONhoOkPWjfUcyW/Y2Puhvncu9qycTJH35tRgM2tuqxmV9p
oUds/UvfD3unSxFHDkSBauF0FfrJhr57g+IOMriT0aCgH+Ht92z73gmdnuoSQ8jz
GiyEosVlJrMqGOH2ytjiVjfGtPaASfiiDskQcpy+nnHaDWuz3Zp1kW5nJNGv+F4o
8p2BPewG4OWhtvgiPgcqNGLHIn3O/9/5QnnhM2PDJsh/l9dY/DSrn8j7+x0CIWiI
Ec0u2MQoOREkqsHQhav7sYk45/aBwXj9yXTw3JSzm3Hbv24A7hWGis1LCKbiyEAl
Wdq2dTLh4pdxk61USisz9Mq5zZTpXXSx6Iq43fU24EH44CFZS2NZE0LBtXEZfZ0z
VljDzTu5yCPJCfbLZmmOL+6nCuUdD7goLRgkr8s7l9TWBcpdrUmyjv2C8AQKkVFF
QIOOhV6XKn575PfR9JsXhbXbK96ysjSDt8WXJoXFIRGnh0ZWO6Z+9ahZdWy8PRqL
Nb6bZJWYhefORc091uO4x8xP1cpst2GjK/3fH6TbEEe1+9H8Lef74Y99XpinZ9am
IsAslD/s5BORU4mVZoS/qdtIdj5DKnxfYNzHf/+Hvzp4ysxalN2y9kFQy34vcfnE
w6JdBIjKAGl8jn2I2Aahh7bjLwKf0xlTh0ulvfpYkvJqZwGOLUFJG417/ZG/yGT3
g/TxbSmiTA2ZoNqNDahKWb9ORLt2k4qUlnNY4knUvwGfpwR47Hq6UvD2S50B9/zw
bJwISvtzCQHJmPmchlaC+6rshcw1MY2SpQ1TlCIokJ8pmKWWM0wycyYw4tQAYXnm
LQrAVhT3z/1jUUUywUUh0hz7prS2jTToT1uNND4jQIcm8mYmPCH9T2EmW3DODV/4
IrfcE394ccgy+OP167aM/dk5VdyYniMkXh4TRRbTG5cq7U1c/eS8t69Y8L4+iYzB
faEUovzIY1AiT50YEIhOaUv8VQN33CTa5osyl2TO3vzrSq1BVpSrGIJNolepcTsW
4o4a04muHa9Qnf7JwuTNUflQgpNvskDEBBcArg64xhzXLxSKpsLX6euD68st5Rmv
R6wesrzaEe/Zv5XCyAHTBQCgyBpZfJNYfQQEZucuTnbISV7SiUis8G9MuKfUkzok
vBNbfuZS2sW7uV4B+xCU4VV/Xj595H+Q92/rK+/ghLl+f8Q026NWgeiaEY8CLQQL
Uq75+ckZpllg3u42wT7snbMZ4IVBZdzVArgsneKKcrUfMilkCWVX1zGuMVU35tn3
dYJu8RdVdNpNwkqkjBRrU+7B5yCrjmtkkM6gm255sHiLJwBz3BZ4DcXxiHfBnW5s
W+R2ZaNHZApF9gGMmZZxqjzEcCX1I1WNyaUqf0SlfoLFxK14FqezzWqyBb03bkV1
ocnX9gJxVytWf5vuFVctjCculFGk3GIIKTiZLRB4FMLUVFgBmMTDaN4to0efuxyI
ckcuGyPEAjnj9E+uSH/Ue2AeEZpWHTHzHWJxHEcbs5szvAXTCcHfNoGSrFwaTiTl
+d6Ti+NZ00K6pd0Kk7Gm7CW6BSP9RadmiK7yCEdg7KUmTQI/v6M1W8XYFUZkwrw3
OXfuSQSLubWKP7CSbPyUk6ACLua14/ZuYv6SMy+P5TzxGx4cpyWp5d1G7xaiq6c+
B10iMelOaQ6xsUaRohUafbGrnDoHgxHnBGKyl2VssYsylkIs6T9HBdp3m8zEp0wZ
L/z4fFfhoBYdPQk//Pn/wAEE478D8VmfETACVGQ8tJL03V4aZxPHj6vY07XWB19P
B3HBYijVqRAryvbvP28NVF5otvEauTTyT0acMW7B8iA0VN4jjT+XLyijrGNDBxgn
G/8sa4nbvnDs4A2VTcGRgHryGzUJ9s2AN/tzf+N6WDykcKCRVGr17EebdO6ZIpZr
FxENbM2uRyUz5c1f00a/NanH8oiFbVW5PEM+ku0fsDfKdWvKfjUoaw2qBn+Uu7W8
AldAgJbTva9NtL/cI9Y1mWsBhgdkpq3tjC14rJfFbvHK9XriGCd9uYtiQETDhevZ
MlIkTOza+ycGPc1dCSvlkGQuLhqysZhMwxnLIkT5dkunJ/C9fzmWEg+b4TcrpWw4
b4EZ0fyg7ZQNXaqtigo/joKq05JoDEZgKAqJCLHJtxvBpyP6bThuHtdXNtlNRj+p
mEu2WbMxD1CvnGJWLG3dPmi8BOsos8ece+XlZJb5dBWOE2WyJJsWxmd0pD2bB+Mt
+dnuVQOmWGs1+6HBP0XlUDwU1Fx+9drYy5at4q0+7Mb8vDhcRJefepalQIBqY1XY
+hiPLPuAVppmV8xb9ayMH3VgveQbAjDDnNP3Nu7gNRKwOcKHg/0mwRl/TGD+xS1U
BHDQ5xE93YLaraRWrO6xzLQhqARPFiXj1WKFDM7UVQNoj6Djt1PKSr4Qcjs0W3sR
KW8IEEtbDL3Gtg+z2J4zMQIWgIZxOxPTiUMXWO1URLAfD5FfjnJ02nEXdy+soZzb
PP+QDAhRxuHEEJM5Ux1aefdVAtIiP5AT//zOVWCW43zD4tUTNctS2fSS6Wrup3O9
IbkEDJ47XnXqHDf+w45GiskcLx7F3pyb4TQMsPKhz3inJyoBvA+GsWeCju9YYxzm
dd+an7F89n+EN7ecgEQyJXK/A+AsCuXkTSaAIEZKk7ZruLiTsn5IUen64VuKToCZ
wN7Ufj0EDm5KQXtwrh9jPKgdt33AZLKOLQyBQ5YYOWcLkWyp0S6l4H+1k6nuGP1u
qnLTHpjdD7MWcxdIcbyZ382VbPDZTe0cKTc16cGXF1PFBgAUHMs2scc/ppj6d8Zs
kXuETvk1mEQKUe2QVWjvuzh04jjo4uFYfjKR11fcyCv/LJ/Tc5DTpQJTckO4arho
1vm7OmAQ8IrhzFB8Y1wsS0YObNoob6quY9RtdatW5Y84/+1f/DI7dW6NzOCoKdhk
Q76VCjn+1T0S8eJxCY+pyviP0oeqEaJxjiTgTICBcDPfurF3SbtWZBbZFQ+UUEBO
FQFOwVry6Z/by7/t54MoEdt/MVFJtSuuSkSDRCj1yaSswGK6W9Dk8EmBiNxFbSiE
9dPtazDoIMTIT79/Jwg97ePftpJH8Vx8fC9/iBCQx1z7Q8gi5C6f49iWOOQLiWi5
ftonu5hQOJ829gJeq/l4fjpQlXSvdnWH7J8tqS/sffRqQMKLR7F+gIVMFcSrQa4G
WVmM0u3EML0wkUEQTIhDBDOo1FTPmq5MjabIo1btyUmTSC0TrJkrqKCnpcm+nj85
DpCL45lOQCtAK+OkvC9dMAwCLyl9zePikH1ax5iPIsKl57w3QUFjTdOPKic1gaLn
UMLnz/20ANEHjADjlelsl9XEL0FiZF8f85lUIOdXUbeJREH649qvFiOtftfN/BHo
YUq13Alqn7qKl1kuJqQvqSkXpNX9667CEQdFO7udV4a+mGUnF36NnubpC2lvxcGp
BMTMt8paHElzhFdgnoRU131+ok4KCQfxQBOoNr5YTIVQVZNBGSEBFucQ3Zv2v/eT
9NdE2QKFeBqyt0EbRUFslHFWE/pjHRGo6BTPYW+FBIXqblMzC2yXgI9v5Z3eiO3i
hAkzEHX2unBTF9C74CyL1euQLG3GRcpbeRalb/u0EKH2mGOWrViHJNaoR8/V6HyB
iT/8HQjNwRrSVoYIHtsieGM66E7v4P6dcdwaNTDRCBLFlcCzNWU3cNMrOSxCIveH
UDYTkp9cp+rkEVTegWsOoy0zPxZ7OWR+Kjg/1BqQUCpSxm1SY2HFIEhxiZrujgfc
MeA9l8yx4HeQ6iwcyD3Ypjagh3e8K22LvOuW8dKZEr2AY8IpPJjiHKD92Hqbt98+
ZJBLRmrKRzVuQbwbFOCoQcAIN2OqTfLDYvUke1VJzVWHJyMUk+HVMVqM9uYNPLtt
TrJHyJvQXY7QN5jCCNV4w275x/tNb0vwNwLZGUs2Rn0uYNwS6Dq6swsCr8PIN+A4
n7GdID3IgqnB1J2BkByVi1+SBI+Ep9QgoFvmstuoGKaQVx/TdQp8solbD29VjT8q
+IkIm6XGQghoGXgH05sv1Jl7VgxZyYhc7YONJga0McJLKySHQ7P6YJr9boQ9z7nf
XDNAnVfyPpZd7lP54qqTwZ/kkF/0C1Xk6Gf4nXrlU3USHOwlLEl7s9rBcfGfZ80r
+rHTEVrS/bK5DLnHPiU4WFZQxA/mrTy/RUd90MYhF895Y6DzlCXbeMeADgyY6Jum
5PkoXXJ0J/ZoZapbFxbaqlfKCWUs+8sBcoMK+WZIvMO0WuLXGFnnOicv7Xml+gNf
/BKqDW6qMdkx58yWUSTnKNZmNHwxdYMZ4bKv2xYr1Vb5xRqi69wiAYuudEpF9D4G
P1iTTGurksCh5AiUd4R7M2xG9YNNt7Hy77zcXFmcKufLM25wAfqwXI1V35wJ1cmT
RYv1yAFXJreaZTffHEIPWbfu+pBHq4lkjE/i2QkJIoSfylrqhJi5iApP6RmMIXky
v3xFwyEdn3iw2qyTW7cE71cjCzDUY2YwYShyUr89Yyz7LhMpgcfDZcBbvV1ur5as
63O1DADRUWVCMCv6mJbY3TFQCMPKLAaUkQYt0BDT0KC9FQs6yk0y8s2OXmG0GRDY
Yd6FktfG3jkjPvv+8hLx4kxG2LgS30mj3qRaC99/S0piM+EtWib7WIu76AbBQCpE
UoG1mLwUAfbp2eE1pMOenqeg8oPglRF4LBPkefLoI/KHmXNj+Z31TjWEM+5OU6dk
2pNFHpKGfJhD29EwbxtECv8NVW/UIVayLFuFeqHoRNfDeUn2SLGzq3qanssXH+nM
vCbqU032Pl2jttu31rb13HnQJESBhd0wkeFa1sjhrETeC8cwG1VA1itRHUz82ksY
C2sHeaRWMLlQvcU+qBWKDqACnlO5gRvZfkp47SB1Y0j+24WA9lMQkbFOPQ9TAz9G
n8nu/Ap92nnhKQ4kb6YWZnrNixeOCZI+yhMcI6FFDMg5rKUfTP4/pOtn1Ipfi/Cb
GhfqVAZim38ESdmTiyCpviGF5M8fgtKmMSidEJoA50QWdjBSdW1eSmpXAlgdOLV0
N37ZKQltF+6v3N2fJ85DJU72zXU6KnMfs/+6gdyV0FgRFXzqnicP2EZTbEaTi2T0
MnyEacC1+DkQc2WDkHGzGnwvC6ZwmfAtjX//FkSGW7tClXdcjI/1XMhaBxsjuRup
UednncCLe8Td4hwk74UuwBizxehEMY0rm0dq9R76E+PWbH9BmMwU+1+RGveUg6/U
sdBh+6r42XRAZrwWykkolGSt9EuBfpu539IEyapgxtESAg4hWaz0tsSjFkBJCJSy
zEo0lw4P+77RFdX9N+u3ID7hXcDSbX57MJqlT1I44evHiHZAE+54K0g8KDu2eenG
l+RNW6//OIf4Murx51GQx88SEJo1EyJIEDi5WcO67k+HXYn0DqjifPTsDmYCzhLm
7k+3PO1dxuHR8GQK+2cN0NSBdzQmkQ2NqlOyy67LBQ+Nw+EF3Q+iGV8qEja2EnIP
lvAAT+w8e2Gii1FwCtjf/dyFUZiu1ceXf08w1+tRcm6AZRGfmAbfQEc8dR3XCLIM
WSqtR+wlctdwgrJ+IMG4ZlS+KXJGywbW+Xw0aigaxgX4hby7LmMhmlDeNoT+A0qf
6EZdHF/ZBoYshUVCBAcB3BNL5gnMAYPFqKkTxY6ZxbtnJ0aborxixogJIGT9ZejE
JO+3yffyMCPqBPl2stYynXFw5AFRJiOyj18StLOBApO+65/S49cQJiPvfd2jY0QZ
flX4D5PJqFkMbzjcdtLH+FUw47496huAzWnHV9Ug6rM6/arpz0wyqiYFwnL9xwzc
vwhb5LU9CAZZyVFlM8o2kl4zhe0V9AWUBpy6KoFoVIM0HEj2QPqO5OMKPJozpzXw
7kolz1J2/IvhYWHYLEw6aziHp2JcRF6rIc0fOUCF/AThjI/RDLcqlfl6ArXp3xZC
mlQWc4Sk0/pnZljTGvSDPXWFRltucmgCz5pwiSpP6Kek8g53cdcz621HMSFfIxg+
tdijbFG4I5sBg72yo4cA6Yw5LAgmIAnMGQBUkSN2SLZxaKFm4QJruu2TmGhBe3fY
kaW0K5kOWtl3K/3WVl40PGEJim0lKQvayx2mEvbDdtrSsUJ+4mNKOi234h6SptVd
DFPXCKxQgh7gDk2rckY4fBj8tNZvFXbHApPlQx7VIb4ymenxY7zPKnOHxI7Bsfbw
eRUgDDlSVYHOjWyTuqtdQl7ah4/hPVfFwlz6/amQwyMM2Nr+4IJqc6afWoA7Zt9Q
X++pXNEziStn+uyGiklkQByuEVKmhCVM/OE0FUT2SgL6IXm0JjMP5HtWoLnJFkpq
K9u6vJQcHhiAu2TBIlNVcWZHLU5z4B+tuLJI6apUnfggsvehO4tu946fuaTvACOo
yLRd1zhhC9mlNvP5cpYkRoUVB/Kjtufk+aXAWcdTucPZ464wg6fBsRXmDP6aktI1
YhoQUWJnvyOEY2yvuTuNuJSKxyZUL9tjcGGwtl6oZYIsk4hnbVgXPBNxEyvINVRv
j99j+MF+ivFI4Y1ok/WDfYGT/bYZZTsU21UR47pPe/y9if2N91mP91Lftqkk5QPO
qCWTSJN5SCsFV1gKH4lICY46vYWrhNFjpiosE53IEg+MikByokuKLNTh94dxCIHz
Eh7X1qHONr210v1QjMar3Z1mt0iLqQCVzwXysE8b1oYfrvoSpHP8iHRG4qJHAyLB
EPQrIXfyfNfwLYGWaQZl/3G8NBtAVvQi53xktX+OhzznDoGTh850JUm2D6VgoKER
R5CcCNuGheNWSF+jinSRuZDzpdLnjWyjz5NcMl7Be+6Mm0bJBC6cohag9hpLABUQ
j/Cv1J/B/jEIrA7cw2Om2KIBS6RMUqrt+W9OklT7vUTuEvHNN73Qbu9Tk+ioDhEh
IuQto+ixfdfM86G58nSwnYrw6eAIGUrWCF+Ix65pjpJy9UOx6l5aWDDFVfbSMcGr
3EMSqM+bjT6PxhwkUMFQWlvnr/qq1QShBHIfnDvJEahBGG9/cSOi4DbMpbKLvnUF
V7PHcvskOBa0fxIMPGX/dI7gI1w+XhbIrESCNIIDXYAkhcaoOHBqkkchMjae8BjG
/SriqkLoitUGgt6r+ZCHI7L9pLrHFKDV9tJ9/kmkdVZuvVSJlcGDlyolTVQyHg1l
F/EIy+H0XdszY+P3445nZxvXgvWB7/wtOR1ieMuyvLe4/aAlQYuHUP50i6oJlqfK
8dW48n2TRVEb2fmD/V2FT/1IaTvTzQT2ifYY+jFn65xHF4dj9fFtNYeMB0lN4Yc+
w8hqAcBXxRQn+PXAAqaS96KIBTtBDhKFHM4eb0NOU9iY6JDddnC4GxWuyizY4/is
nMsdh2XoL71pu+XIvFjwwekDDZAToD+6CdTljNP5SPerS6liNemXxsg9cpCem+qJ
9uniF0y+U60xVPzO4XmbOxbl14Z58JboYalPnEkw37hFYQSYJ19Tr5AxtqXcTiNc
tlbmjs6nIUcVpNPsvjkWhbkb5SoQpMA++udDzDF59meaMBue5WY6/zgrsBgsT45+
yuWFgZ0Y9+sMYbDBrVtEz8LKjuYET5nFEdPvZHnB7mcNioL2Cg3sQNe/xpUidjFS
zE0V0P8D7ev6D83ZCPgblmXmRPbnDz9eCADC83/bSWjRqkdcrPPt9k64fTfvepYr
HoiRg0qqVrp6RX3tnxhrR/70IjhqWJGMqvDqrur+mnUqZjsQMMCgwkfpVmNeYTqZ
EjEpFU7GhWqCLh6MRsHzi0hOLstGhPQnV8DFO2lnvI+P7Yx4ffgkAfvHh8rLPD8J
Wvh2c//ekK8y2+Zd7iPuti5WJb9EUyM6ngSsl05gCkpvlPpOsItjtWN3FzHrXv+Z
w2dzXbbPVSUXvkmuer6zQOCc9AS/In60l3wgtXaWXD4LRQFUbWh7GFuSHlceqWYg
kQUc4uqz8xhesbaBuXsjUPQYRo7zkA+hgjZgdqwju1UZSsGsaLaF4DT4P6yCIBcV
ZN0e6RSgkXgnNOPev2Amxs+5EI+c6ZgYfemNiIaxc0ady3EkGN5VBuB3BGvVKh8p
yjiXZTI4hJh2ux+ae/TorjG3WHa25WrYMBqZ79Z3O4jSUb3mmMX0RFAB4YX6TCEB
IYlxRDozyNFe5nEnVw/d45nlerqQsvn3G2ziFZO7fR9I2LxAXPriqt7a/qQIyqZj
PsW/zGPFSIIRrGjG1pEWxxgy4yv9uXkQnADbunfUu56G18brI4nLJwWBCkIPHnAV
osiuO/pq5wvuv3gjVtS+c6gppv8aK3JIN4yZKO0PrNuQBn4GLU/dklkd2ynhskuO
ixassMChQPT5PA9K+EA6YQKoRyOAd/aC3MEYotZTYn6UuqP05iLNUnW6vAlYymG+
yQaKWNmM4KOifTEuSsM3aikUQsGyDrPqTd0W+cJjMOu1soK2+Al/X8Jt59/WK0yz
ANl1r+2cgF8FQAS6H3n4ZlkqLOnvAVRcxncHenTSGl3bmDl3TOBlZJNHBL8kpjq+
RFiwFujwIgGrWzYKo/43macEh1IC3cSSbsl984k2q1t9OwyqqcTbsJfRzRfrZdQn
HgRJ82pUCc1HzG6IA+38mIgkuOCi8djEOL5ZoK1mxKrjRcCeKX5NunflVpVwz7/j
TWc+BqbhsYvzU7LGDPma/kdJrHPGCbFG18+u6CMqVR97cMuNl8BKdXW6ZvI2tezt
wQwR6d7qR+0ikWwgJhrx1gMaxqbdTC+Uu8TLc4DHoxrPrIHVWxGR5fSGvzLiXK9I
J9FHEOq92Ktbyv9K9ofxZ/uHmLQtuWHUyK/0Y7uIg5F6gn8qU3SEq4Q8sakA0Sws
kgYkn12kEDL7KI4MPMNXqpXJM89p1+lzByn9Q8H/nQWr83lmi0kQi7kts97jTJD6
jE1p62qdcj5TD+X5RZvnLD5WqyhrknplBsnMQtxKSkZwwwtkFaUJsDRg1Ndj6XmE
VW64sfxg0P0UDsHEX74GkJYpP4LaCE/eCRcRWF2ojWCB2i31GHMyJyVUk22IF1EB
JJskvke3jv3kdR9Mlvrh/XdwhskbqWYnJ33yhM3qXAnVHeiNVxDoX+64xBL4Iug/
eLRuvxTzGvzFkP5hVYMZOhtZ27UgMyrlgLE04i1S2kBJ975Sx7sek1Bm6kbqpFBr
cOjkTjdBOhtjhI7eZXituH4oq6FysPksLtTSADp7KerXVoL9JCGoTchrVPvNNMTy
O6MkjwRY+vvFpI4quOf6V4fncY6zncSsG+EOOQbPvDG5J0CW+5YlnKBS1FpwrcCf
vfl7Xl9tJ40BNRNQcwR3ioXJa3RuaRrIEFNLRqSGefKW5QSMYA+VIo0ZDSxslj+O
pNdDV0n8hVqwnzFJPKRF0eTZ73eZLcFOVU4xJc/1u65xrfvyu5zucbDl7fxsobfy
kfo0tr7wuYGxyLBg7pcM3X0tfQjwBHJuRRgCJNwxRdMQr2E/SjtX6afQr9C7yY7F
S6rHEUPmFb0s8klNBRPmMD+bGNor4s/xPzS5eCTPJIcU5Sg9X1gJBcOD9AYq6+Cy
xZlykTd+V6tAsc1HLQi+R/nYArapRuVA0tfxvPRO+sW6F5pe6DxRTWJJ3Z5CIf+m
oSyX+WRYi5NpYJZxxawXK5KIM6o5tsgQIE/JYLjOdfXCIiYUkDbCr0ojzuWtfwKQ
GJ+p6Soiv37kY0bTdd0PLS/xfI+u+l48Y8TW/YwNOjMCnxni4RX1gE0x8GsN9QBA
9IBwHhnYqclp74400Nd/yilUKzRHV65YCRAfI9irHM7czpWCb8iIS7tjUOOR62AC
T1UjRF7jUU5fXlBdlAjPI+u5M6+uCxg4rMuGqMpULBE9yUOuiMv0PoO/nfqBMA8M
Y5X4SVtZeUg4sx1v1H9RG0X9RVuvOgw40oxD45Uy0h0H1tJBlbSyUCJQw48itkAZ
jOtQQDr2luKhgHAngcGEqgAtQQ8ZZ6glJAHKO9FuO5GjXhcHmkC4fiF+8qMNI3Fm
3+AYibakIYDmNt6OEsdjomt0UrWXXDDVq4tlhFSN0WPPyu8VP69hGACGm5K/boAV
eWwpUuM8fDaftV8XRBIZmSWygLU53oJqaOpnSZmNwe/GKrJwbjzB5PnUO4TkCNXI
aPVaGv0m5iFQEAIRDbZ3a9uH1j1qI73mJSulzV7PnA6YRHnr4PeZD4JrA0DMyhcH
x0AhSY8ch8x2mFWAF2H26TnEL+moZko+8qULBsH5C0zdGo3KhoeJ13CbgyAodLfL
oM3/MFC0RTbF2nqxM8EcVggWBrPmlcurR/nGdMOTqWA8YlTt4UYfdiBdFlgfFswd
zdnh64Dotd9uLpYbtQ7NDDwHWDCgonXRbYh+d3h1dVw3LDhEFPJt1IBoBQBIKOzf
mIVPFsVlzxwZQhRLpi2+R6YyA+6GkDLe1xVILUf1sx1Ye1Xvymc5J5fgwKUUaW6G
uRnwl6go+pwh4+ybALkgQ6GJ8uR8+YKsYanMVjEn2kPioKWovdDMDb9ezXmuEyLI
gIFSFtaEehV2TuRYfDdbW1zci/l/xPHllf74+cAIC6WWx4x8+G3Cm6a3y4JFkgEs
eh5b9a4+AU0X7mKX1IMxzfD8mJcCm52btkZEl5O5MPaAlCZJ2nN40nsJCIkOKXJF
6Go9FfsPzEm0+B0rAglG00JY4rmrJJ4WfQQR57icCzaQjdDQM+OhLL9P2BbWg8hB
9hQcb2ZIm2q6T3yuYpPpC0g6PglrP/MsZKte/E7rDYT4I6h6RRr2pTvHhZA78nAV
DhcwfRSRN/AAPOT6qh0gXxstS+FedUEUAOQTIo+omjUW7vrlkW+zuj74dlKKowfq
lS0jEfnIEazaDGGT+R835jD5fhQGP9F0PtdCQOJ0B6/iP9pgDS4EcZA6qFUGn+XY
iCtRjFAAjZAfoagV9chKLNQPeX0ZZPiAmZIpv3AtzWV+tBKiDx09SIeHOBgxz5B8
PuOeMLYbOmz03tfbGx93ZDi0yPQJqiR7rxhvJVTepmfH9XubbXeUSAr0sYiSeJLe
L/8MT4UNgAY8Tk2UYZf4Y316n2ap6ngaSVkX9kXxoTMvuTBDj+UVuGa9pEGE4dml
hM2y+znxggSWmv3pUq2MiKVLiamXzieaZC8r9ufuXOIhpQxOutj9kqUGrTlkXq76
x7NXVZ1s1Ky0qfZf7pzhTVKLOOofITvkxAqIOHkEy9MxVGHCuuJ4f3c3d+L7vNqu
QpP7G/JvPr7muvxbbXrjywtbR0r0VZnbNoU9BhkjYo78FDPa5LeIomAGooAeCVkT
/2peHfGeNxpX/qADMCo1exVdD5Mgo+hKbBu7/YhYjyXN7BFVyjhlVUkPoH+yF207
PxqRmRZ7uNlA2o6wgDBCViRcOySalC0IxiL+O7/O3/y9tt9w1Yfdgg63p/dUnmgp
vbZwPLozfipyV0Hrrh1RVTUQint0DjRqQbYLnB6kWVDLAzj9Nc3Fag9AEI8DZ+IJ
Nbyt8DDUYz1cDYIfzwtTVMwNo4PpB6LcbznbzcMb/KJ3/HAbimnQhI4Eh3eGkOAM
vvEZt7RTTCdsuzrhWICLWn53y+nE3bc5wqvKQO3XdSmT7WypPrN2a5DDPOO+gf5B
HyslGrBm4FHdKge4oPUAl0x8nDtk8B8J1LadqvZSyHWuy1UIO0j57ZUBh0x26Rty
6C8/gHpNIS3IFU+ybyf8cjmk7l73Z5ySG2VDzZ9mUT6Ea6R8xwPgKM5GqSNR/byn
Xr2kNJ1/3uEFnwAe/4clE56+wGsFNulAPmNz+pIBT7EiS8Uz7oxXXTCx7jm722Dv
pnKbqszQFusMkh8ogulZqyH004EHvNw5EenQ6Cq5ip2h8Q8t3pzCHsTnw0gylfVQ
WimzApfdn6yo0+ZqRy07AFrb5nTKM9wG291mTlN3HY8DX/HHd+dgNKDiOdu0/uoC
JwoelHPPGK1vMek1BPydeH2TjlIWlCWVvjqZGgzPnXMfqQB+NBIJ8X0fwyYtv5A6
YppPmptpcvp5cDBGWt7Xwb9yyUpT+5n8Xm7ZalRYUuJwUs/notzBewIIPi3ZpxEQ
02Vjczr8o4g7LNzrODFzLlk1U0O1id8JTYAodvZl3Ec//+CBAp2v8lhvNPf5Zlgm
SJS2d216v99PQ1DKoCDHV1w1ucqw+2pvnltMkskWAqW2iUdgb4DF08TXlcuKVv2O
7cMBsULCaSynUjnq2ARQDYNF8mzzWPgyFRiZ+5zCs2doeFYccnRUnwvhrgvYZYmM
FbQVLUq1q6nOZyWtCOKbIaloJ3fuYjCwsBVd8562Qw0RL8y6GPP3BCJ9XgMtwGXc
1Bf2LXtwpNEuZ3/ZHXB3IgB2Bx0BVBR0j4cnuOBZ6lxxBj3268NvZgEdtnQ/ZHuF
PeVlL7dKIi1qtCauQVt4eLf7U1jqsDZtOJvIQfN5bD03/RFIworYyMaTGMwnZUOn
8WjjSw1GeJh7DUjzhkzLlsM+nfZHowlGjNVghV2XzLpDloHNb38P+B+2svzNccGn
UAoAg4S3OEkQp2vV9pO0LHcAPMBtzMaSndxDrKQpcPyzsslKDaT+K2zzkbySVecZ
oXvwou04bHw11lxJ3gUQ2/2mSkhMyLJ+F7982ugYw6GE6cCc4NbpiAjrIhMJFA1n
pzONRj8EOKbxvtkb6+wN4/vKC9BiRyzc00B/5e31s+UUV94IygWS5eiu1VjPoasL
DivuqwI2xz8spFDrLOtpTLXEka00SMoebbgNNw/TcatGozI1N2MqPoYFtigjlSRu
Uo2+Nuf8jXXWZcr35stvu1fSsudTTy9E8Q3DIyb7Ar2cZUVfcy6Yvp5VUfDeiZRR
MrbvU/BxaWc7vRv6ZX10iprQoINH7+5BmRwah3DN2JW2zGM/xEqhrHn+GwMBdLLv
7vCP7Z4aDJPpgJKWAJSUk10mIiZyXXDD8iKkpCxurdTieR7s28IvW2+rHkdvi1nU
0L+5dTd7OgUieHZojaazxDhwOjbdWELDU2ArjiwHMn6BDc8nHgUoOYl3su5ovBx+
WyZs+smOX8NQ8s/EEN4a+qiZXqwOZzKPjzOc3qg1INaErgaiiasTEC0Orf9qgAKX
2mHB7FG5JfXzHG7Bhe0urii9AUyFEWc5dlnj8AU7T2YTUOqaFrXtj5BKUfViPA/D
iZcBosglIdukmBfVRhlcLlnfeElGlnfAfMUI7fGwOoxAWcO791eCIV0A9hdjDypH
Yqk7dlJrWmYvrS4IteNIExqncYJ9t65PDbrAMyFT2wGrgGJFM2uYgBnz2CvwW9OI
g5Rs726eey8y+p25yLfl7zWoIpmKqV+hTuOqf5zIBXLPCRCdGqxzoQjTsYWGMQEI
SpF7tENc1NHhS6Z0lWUVooCI+t2oEQNLreyk6+t2BhxZ9FqXW1JL13slhQBwqTN1
It57FBAT9D0I1eU8gKZrMTi95EZ4hsvPsMZN2BEvXX+Y4aTn+tufn1XUjtLSyU6y
C0F2zRVRyh8bajs8M3IanjsCwvNM85tCIHwOPBjBa+/11jTbHZ1alhecRHNZj/3X
Zp8gHxGfidiljzJmnxcAG2YosVVaHDlnK7jiLJkSwwOewMZSw0/pop/6hM/4GoTr
3hOPuFnorrfVwtIO3yQqU5KNgi8BG1b9XBCdrPlu0QkC3qOpPpQzmOumSfvzRPD/
KO2bDgsqdvEGgGCs0l3M0m0FTT9N2oq+D18MvqZevtKbkb27ZLuj+EnhiOcFMaZ5
9CK9qZjI/bErRHXzWYKsJ0aPBSh+bT9ofAjl7aDtG4rJubBW4dzAqQjYg9EnorKy
vnBKwA6KsmNmGtHgvFFvZ4UwCC3HJBC1C+XcmxzkSh+6u9Mu5iNosB/qJZXHvucO
Tj509qYpx6ht60ATFTSs4Oy/wE6mnx21zqvWdKg6QCX2u14tLlKljVODN5aCcqsX
ntIixtbIvn2TfTCMABQfiEYs/97eLq/tUi9mhsZKe1T0dysI7y/0S/bUVbmt0KQM
FxB9/fjjv7hrGe9vZhu/lFb33phRrt2+DkfiAaTPD0yxminUpU1C6JtNA+DS2qZG
++cnSI5N8td5KycA45K9i3qa/f939fYCBUyKtKbznICpvtHcHgePC3PR9BOXDnqD
0XHVgDbWeTDe44f8TqpQdSnnkNQtwElR0+DQFyLoNZJoI9PTaRmvv59FlQc3e2rQ
EpxxiXLkhFKBYnqvELj1cXtT0Mo4Jd73REuk1CqnvdpHVXRtyPc7S3U2/69iDmHA
hHMjlVW3J1Jqt+iSimYJIbhQpCesCT1XtsBcpeNZ47dF/wQY/zOIZrlzcspjg+hM
+IuNyjMK7Tk522/HrA0MOO5cVyRcWI4bYAfc7ggyoccG3Gs8BngQO5sI43RyAmON
V2lvJg58ElMyJsRBgjJA3h7sEszj+neSrxYygPsSIALwo6oagfIW89kP3q9XTXIi
XSu982fgEaWDHIyyNhrlAbfxOUyq1uhkdMpZZeqf0wmYj7dBa44bRhGPZBKATp4M
P/u0UAy2w+EVhzT3OefWGFinvxauHFeQbNewoVHTp0WlhkJ7OXVdO5w3h0C1FYSu
lSr48sNtpQXNmyR5KrJLk7yqygYnauGyeG7jdM43LbdIOEvF1nsldd8BR9Kb5oMk
5tEDTWe3gPgDXVoEsMBf5glFlbZ6geM5t5qYqVeTVycvBFMdlS5o2u3ZHa2clVuf
8auKgZ9T46vZb4hKKrw1F4/SZUCf37oHq/1nKxBqt28XX7r8ATbEbwBItIcRRDB+
Jg3AIkf4rFN9CchKWkhDXj05zKWVWahJsD8yDNnJPIpJhVAVKKVsbdvYgzIxQppM
hjFLE3DPpKn7yaBl8RqRPk+j6R5ushWC30hIK8WHGxMejtXdq7+e5gRDTD+EEy8N
jG+nk0416iE3A1DllUYgu2HEciZotjVCEB0FfQXlWC+w1rETn+dnRl3kYv7GEkmH
K5kyZCcyFik5vKWJann2bjEScmu4SwqxE6+IgLAR1nes9CSGP/ISiGVL1lVqmB7M
1hbMgObEI7EVeHMm5pQgNwl/exXMPW8O+NH+lRPBFK08IJtrCs64tp1FNhEeTv3B
fMMkyV9xTEmaO9bMEseKe7rICqFTMpoBi/H4ix22AK5FEB6QwyhoqjO/rig3NH1t
fIne1ztvN6IiumBIovQjwmtSnQjQujP6ze/MRR7IxArNNCHPPblam29waJ8z43IM
JU252aLLEJPm9hlAvO4+7uKS0TujoaKA1BUie/LMykcXD+oTv10sV/GWAs4Wff+F
P8wC5SEQAaWkZSrTCe7YZTJmMJuZC5Kbo8yzcyvYp4ASdNzv1s4i1zf6r+lC2nfK
fJlMNP+OM8OiD5jFdUvVHY1HAzaSbiYkqtN/Z1eGQigilOQKeW5h9qOPRV7Bbn6H
FNGzaGbyplK5OESU3L950QRe04QdM/uC4QYBZmK0pFqs3fmSkMvbCiOasAukffzm
KcGLRYCrLVAWSDMTgCwY5oUbJsyplbqq1SgjRLW04CCvesAUdtCZgGVGUtF8k+G+
fFn15vojHLZXqHS+uXIRRo8RDJk9rDvn8LRTn8szRv460dMH7TNiGBmivImCUOum
amh/y6bSKr1sKTKwhcicSdA/yung4M3H7yDt5OyGZTQXsmhx7PpeRRm+rrhxU/Yi
KhjT65bB99ataKCipSQkYVRQyR0mmC55u+5vpEwH3V3QCGZeqoBGBfVkkoNM1wMO
Af0kNLKBFFKk9mltvRxP/ji+hhmzfefGPpPM+ycDPMOQGD1qAgjNiDMdyud6nKQj
LkVhwApY/6vrzub8JnfxRnbHo1MB9eCx5e8fwe4BfdvlT9XTPzMGl5z06ev1hbOT
q+OwNbMMypguds69OJDDC6x6zOHJFPax5FXRwmQ7JgfkCDvLVRqDDzDl3jwkxeX/
tlHbA8jd67voUeEIMJN1zQxrsCtflZWc7t1vzm96qjaL1YauDWwDvVnWUKmE4fQT
HEQKcLDxgmJtuVDY0czVPjuU2pEUseJqi//fDkSEtin9nWqvsEJXr292Q6Xm0IiI
wtzkgdYL8AsGOuhB7E7VLvNBeRFg2aOqPcbEDiPPeQF+3/NNRiE6K9mJCgaKTEog
Vo8x6Gm7wuzMX3ChGpUPj3mYlino2Oo88knqfbdw+YmQZVJucy2o90sJfnB0zSsw
hT1uJjQLYv+5J7/OHA0MhbTCkUXh3hvy6UEf2OjjFPt1excoV4O2gOat8Old0Ss+
5EMljmYuZ9zmOG/o6TVisLpoj6JDWwrCK8wnMqiNpvBP1n1a2h/leWHDuHYArHz9
wGUaNKYlT0EgWaQjjaAve0xnQ84atMY3bk7u8M7+fg/f6NDZ5u3TCO4EY3ZOGQzh
ByT1OMg1kxlL2pGKRD3lE5ZCVk9GDplkyHnVVH1cwHq++ppGwfUG++CCOvdmqJfT
nmxtVJlNl2vA5PMF/8GaAvwceB00VIJLrRcf0a1X/EqSRFzwFbcXXisdDUACB1se
glGOCgfnwVJ8WVWCBtUj6pW3XhNkxqRY3N0FqEevsD132ImE5I6j+7i5YW4MCsLN
ClVZw3AtEuJ3HKvRgSO7mi+AZGEZUWfyiSnhwY7GWPcj+KosLBMsU/DPt4WAljYc
NOxPp1NgMl6C7PFBl7j7jvMJyHVASH4t0EAxeJ81BP7d9ZZtRhvkHpxEsCrY2rt6
gE6nsstL6Ll/FoMr4wuQt3d28bjSnJPWHMAWscBkY1Nj6oUESaznuxCehdGcSj1O
VrA1eRTdoPOuqZd1A/G7Tn4aIKMBxbSIVuQQzrauwdql9Gd260b/VV0KaEJIA7BP
Ti6bWYtoLb9rfyFIM0bpfBqgwMiUqxu2ECPgHWI5dzrzXA/pHiMGC7nShnFkoH/5
wD1QxXUnNq0cKLSr2pNvBvdKyA/AhHY89fS215lABgSbWZLoX0kbsJNBOJFYvzyn
tpOZ9FcRvjZZE6v8YDVV1LXnWDQk17ZPIAYab4/sgfs0uoXhNpKND14N3OJcwK/S
JKV1dexsb/Ow2+1DiRNJXo1Vd9blE121rNcfDQ4UXF263wPorDo/x/n42Rdiumta
+jJzvGmPEqrJFMWrXJgn7X2nThC1TMF9J4xpXNKq1J9/A3FkFroNye2jX8QtFftJ
+1mOH1GDcsFeQZkuzo9CLfZtDb8jmAKzI5JnFz4QXwTmqxB6VBr+Fqi5KHQ40kCo
pK6H7h5IHAKjCjT2/eMml50FKnS8+qU7HElHZBG6u0z1TJbVcRCFcNMnZg/zEYAw
puWQNxV6RmPD5hSh/6vhJIXqtgXaTRiRC8o6/7Np6/wnYjq2WyZumhnoEV32n3q2
VtAOoDp6r08awb5lnRk3BecgSNWs0IY/Ug19ZNlM50l2vlFMyZs8ZJMCsKhVStQA
dpOSUUS/rQ7Q5hLZbod2MA77FnoB/bKpsDv3KKXTaGfJQDF4KpK2PeZAUB/I6Op4
QzO+yqiE0xPX5/GRCN44hR0NF65GR3WO9si3fv3E3102MgDKz5T8l2FIsn4R5cU9
VgxbuUrVQfUkDeu3GSAp/U2JE/YPSKxq948VM6gbXLpf4P7e5k17UpCsDgbHhKgE
Opps7/N9zqQCVmprMKxJw/YkYWsp96U92xdFNVrFQhxqHNGA4OoYHzdoAg4ZhggE
+00zjy+thoNYK3nkCB+rdjOr/AC/uTfTfeLGDyDfpAAA+g9N7IrT/GUegwJVHhfB
Wi/PvsT/UPtoHlsYuF6KyXAhvO1b8DRmEYImoC/qmF+U2G56nwOrSFPNjoQFH6td
XoqUL2nWxlLNei4CBk7hhixXl+LF+EzWz+rgApiqWE2lddPnG9SOCZ0GdND/3OyM
TnuvApih1EVuRdW3xIuNI5i2NDa8sdq/OQ04NIwAPVKXDe3FV9hx36tzDkJsThur
FcBeOShAFLeBAFCJeeIYQfynSowDbuzzdXfyKxWYntT1HAYG9A1OpraOYVyrZih8
tWPMySECpEeiGaLaE8qmlgQ0UQjthgyhtc5quPgpwNPQ18MguachshntOZQz9JKy
H9aSv7DhQG0eZqebGnSmmsvV4Wyq5KLOG52HIWORVX+TGeREPuiXFBtXjx6bQPNV
/0YAGaPDYhRcN7xXby3O2IeKBNIzkIqaWd3sNWFzyFu/oeek9PIfwzSqNkIyQvGn
3pzLfrUB1SqSfD0nuzhcxWThW59+TpIIuaTLNah4Xio=
`pragma protect end_protected
