// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
lr7Tw6wGIjnat3MbGaWkK2rhroGILy+7AtWyEVY3gUDbuakjcl3wg3nafk2paNOhmqOH59Lg5iGh
Ge9ZBlPf0L+vKGe4aoZ8mG8bvZkHnJMBYTgum9hpFDAQtgjXSk/wj78jWHeCxQAaMHfbypVddhew
f37xf2UR0VxQZM8Cg/lhaEZG8gtdydIQYTOe98Kdfod5iypChghETBLBen83aZUm6FsOo7Hjn0i5
OyE0+xt4YoC52X9NrrSl1aEeRR3ZiH/RtrTjITKWuEXBGa4njytIbu5bIv3kpDHvXZ/iln/wbQ2n
2RfZ4Zs26B0JUUIxWxYGPpHdQ/bNpygyvMUYCw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
SyWsdc9HfYX1/CLCD3rvhxunX2DcpfWDj6wTsvxHxWeJQQIbHwM5po1R869fo7kilU8aUR1hnYZT
ztHUR5hLrczAKXgG8kJIS/zc4lg8iPBsn7Ou6KN8IdaByMYwZDmk8pznnm4+2yHDyxaUxfWwXh8M
yG82V74PuQNDZ8VbE8dYoQviKQdfxvdWBsQYuDixPeEWRtYHdxGnLwpp7dGeR1QZRB3ZQX5wdF1C
wKlmMovQsoJtQ0mwHzoldpCdx2hcGyLRKhirzRZ0ew3d7PoKqWK3Qq2TCOhs8+Uu4uMebSekhyQV
eAy2S+YnBUPaRbXv2chaBxihRpT7vUr3XPAjlI/8JMlIQ6nArJqIaKddipoH5y1O37UMwDJQkP8R
fjFYZXJ0ghaeXQtvVH6Cbrq6rDdg698p+rXKkCbkuDTrtgdBT/yfohBdXpfVOGoSdUZk3qpSECaK
S+H5kex8bjjlWyaoI4Fr4Id2DxfkeQwMjfYh/PHbYJ/82sF1e0FgX0khSHm2mSmWXx+KIcsp/fq1
SwKChJI23w6p7jKM+Va/P4bH20iSU1WdB7o0wZBYiS4dcEaHujWS/eXiGeMM7Nd/6fjdV3EtCfe9
cVaHC0ktvat9t6I8fM/m/fApqu5ScVyzvQ9xpg2GQtu1oyQSGgztJLSjkguz+VPDwxE1f55mBE2X
9KHCmGfNPXnMLeKLD2ypM/xDjySQfJyENvKss4UuI820Gyk5d5yFlC5OFHbcxniktnZCmXfi/AYJ
BGefVQsauK6Vdfi4Aab0crTrzOUEnMNvz3r2BBF5BMpUahmyLBhTOhdiz6ZznIJ2ytpueq2WsWV7
B5ix3H2iEqTo8iYwxgbWp0Ne3DntFUV4TpNBh3FKu+nSisanKRjB6Ux61Ta5ca3+sBK5DEec7Aar
bkcUuNqdNdftevLRdk15dK2XQ0zBGzeQlsdxLSu5DrDaCy9+VWTQOsqBphxMskUO8qE47KqhafzT
RXxjD86jvFqeEQDt38K3KrmfsVDFcMg0zJy2ckqrddfI1JL6IpLxjF6g4uX1VVO+qjQu2w4fCFtt
dj6cF4U0oumUxwl2FKLFui1xDOJV4mYv0R00J0vjhp1zLTROYna7eZqy3kvXD0B6JwdactypMc60
TQ70sxCjjurpdB5zekQKpE7J6udJ4YLPHIJWUnKA2Soh9C/aIs4zJvG4ysdg2bs0KoHOr6UTU4SB
RmN1tMvZ+D5BdbwUsYF14MeOPl+1823RrNlyumC4sddUPr7wQAsnmvlSmWiXpYUsH/5eGDtCSJ9y
TRQfPyxbAb9hep55AqMm2flq2YXUjkQDiu18KzMeNN+hMspNGVE+ZDf8q6yvnTmiwd5gxxUJdqyl
iCKGx+p6+OPZORHHbTsVa3l8bQbqxy0Whi5jBJoe7Z4Muvt5X9u9g4SYI1Pe3KVbcuZ9ytWjrdnQ
OzARivw6NXptK0JN63lu9LYBD2SdY54GXuJrZ2NE7lQHqWdSSyK+yXS86Y44LRsovUflp42YnIsB
fOFGDVtbG8IvhUUdSkALLgJjNdPRrw6SVQTlguO9PzYrMoZWWLklzEhHvA0pGXepyLiWeza2kw0z
GfDIKtpAaaHZKJ/jho8HotSyb+CXxIqXsY1l5VAJ8MegIh9MNK8nPS9+//tNup+zND/+amGfFQKk
leHOFCZxCCFIuC8cl75LSjShpo6LN0WD+NRXuw5o4RG6FbJQXjPBhZkJbZ//wG0wtbWixdmSuDfJ
HS8TrDyHt9zF+a1CWq8RaxBSocJ6rJ+k3oaFVTWX4oOajb7FWvB4n8UpwgahB2gdCjeXWyVlrljT
dgzgHBQ7wTfCoTEHmDub4IqZZTIVbBLIQtejisHfo0VJqkk0YzSPvhHMYv/uzG0mdTpMIj/03czw
RB/3Oze26wdrShbKG+fmXmcIEVnZwug8P5Ue6gIMNXpB4ub/PL8C9p51cM2695shPScUGH5QxU2U
agmdAEwAeuZcC0FmUTr7Usghp/pV4I91vKc7WNgSdf3Ex7kPHCSW6Y10MJU6b//1H92J25bcdBiL
HI+tjr+YukstXvub7uyKfBHzCOa3xxwyFk1g8N+1pRdJSEo/IMLnXhxRnVp0FNp4aRMTBem8zzhO
+SloNmUr7vP0drnfC1LL8KVH+dUC/KTWXSCxyKEK8Be9vRamU3g+mwYZPcu2T7JR1vUP+4SWLkj4
XHDF4dkcKIROyLeXTDQjMqfGyeED6vKFObGfAEpXJ5ft7x7r4cs8yhZTfX99gksM4U6BFx1CnVp0
qsD8OAZ60HCajv6ke+/AveEujclYSyWjyKSvL2C/vZlcPdcVr5AXrZ0veqe9X6c3q/v+aHfTSZ1D
oKxwaIuq9F0zQKfgfKGIarfDMYpTwzBD5oP7OzLu54vDCPlOnPNls80EdnxwWeSjVr6IymFQL2uj
UulD9YRs5gjVjFHu80SArQoQEF66OkR64C+YNQMvJTLUb3lvOwwbi1Zm/3HVSd9UJAwpxW82coFO
svzzw/tMU93SHsnABGEHuHtdZ14XD7s9v/lw8r6jstex9Y2OkVFt3uqNGgTpF2RxDgs+MzGXYM5T
8SgTCdBNeWaHYuFlmYPA245ODhm2G5QOeo/+7iW9hKpOAlGWt/EphRcyFF8qKw1XADtIccMRSjBJ
z2z9NqMFyuNz8UQovVIvfbYORfsIVOJ6M+xDZ/m2hNW7gdrxLisvPq9NN6GAxqW5CGQ4m0o47qER
vwCfO7JUxXAt4JIwB+/ITqDLCD6PxMcu8eRLg91ycPvq0nbbyDcX43r8FthG2I/OH+8ixlX1xbNq
9yOEP5JCr1r2LOnSyVfO0C/OfGwizhvSW/TlkXFk2aH3179EDu4O6BoTuxKRk8Dnt+RHmfTzd9jO
5j2Pr1guse1dv77a7oSjU5pcboih4KiVXneWVb0z1V174VP+lK4oszHNCvRpzXGbbbOy2arFoAbm
Rl9azMykOHCpIz0gPxREKX7Qr/y1VgQwyEU+UrIa8YSPwzds2+1qgQpebT2HaczV+ATnVwBsI5XC
uN5pmPj4QTO+5+YNHio+xqvFvcpH0RXRDy6tz1sILuEDKPv9jqlYOtV62y1Q0WuuZqUAn24NrXkF
2FNH90FXMbiXKTOD+X4lIuF8IFlsh6hn50oSXcnX+nP7e0HaGZjrmU6O8ENNzBXOaFF1xcR3ELK9
IMVHv7oTWLfi1orf3CF38Y9+H+aWIOkduuBnWbs7meOqSJy58TuE7ZQzIZ5fGZ0P6wgHhNl/W//K
mPRDqGSd+9p2fT+1Z3d+Cz5RsAvn3hhQiQ8t2VoT5/buqRz2qfnXodn7UMEeHQ2WNqRt9q8rwVKB
F7pbm3BkokFPenYfbjEy5r0PrAmFCivRdceXm3U/nFKbp4OfmKL0ErsQ7iwEfqv+v90B3Fv/xO4G
7HoXE6EoTLYcgsspe0m1JDeEjZy7f0usMnOFnNeiA2qc0ywDs9gSPGiYdKaaKz1hk//jCvVEW6ou
rH7vTMuj6330VrATOIOpqy4gIysGuvioWfjT+zwvgybakTPWFQL2+mhaXw9F1EvcqCmlxHOQwhRb
yTVcg9aUBXpqMNDfShX6dLufiVsf28RALewrD6Z7w85ElKJ8DfmT3dRzJiUlxe/ltRqQf5hWJ8tA
Z9emhXaxJg1H1/4Y/fPASsD/oy0Ma7PuA1jVlz74kdz9dFId8xrdFB0JpIQUCaec8X1AGwhVf2Nk
L3iA91/tNjjbBv4Mrw1mCn3LHpIOvDiZN+M7u5hOSD0sF92I3H0Kfu7APtk2GoMY381gnamx7Slg
GZHgyzWtgHXJLTM+69e82aEmnAf+0QaSMlKzPLu81RTJnq6zw2Zb4arKTEJZZ+VlXf39jQX37grl
PVDPWslSy9yAILIAmLCiPkgUgG7P28u/oMGdeAhjtni1k/gU9cwvO3OXhtF6Y4sWGj7DGAmHOeQ4
RN0ROpj6uprxkWTWabGUIP1uYOG/1DA8YgVMMYw2SV8JFRK3r3QvO9zImeJNEYooKWyRWKUNsP9W
P0BUMNIGfIxybD2D+A5FUl91so0U+qFaTQqd3o+4WOy2Uxu11N6l3OpJ/QWXADfBXfvDqbEJ+wyv
kxnqNsXaJSJNC4kbYrULiAFS/WZg3+DVPNHOB1ygLRp45e3JKphZT3pfAbhYfA7D0UW/pK3XejCv
9vWw3SZWJACEn1CYpwIGKfBzjNUERYVuFfb37NV7/JSyl18QWtnTJiFF/GcfcW5tEgxlgVbX3PZr
IycnxRAiQ9N8yV4huuzEoal/RSuMUonU/0B28YMhGdeKhASSngaQGkQX1+ksuEcLleP3ndVhBVtn
DPn+wR7ZI6tJEeby//Tq3PilokAXux84chIXS1X8mJ1Kwk79rOFXO40G/YdjEzr0JYukeP4yUEYe
v3bGgvjmxU6P41nJ6wzdH06ztzsY3izS0W5OploJ8O40aNHLmNIM9nCiQyNqwPrqMhgYYWiA4iSN
N6bCp6bfS7/nI0RUjAz7h3AYro9337kdgS+/0Ww/vInGdLLfixLYJc0dA1xKOLywBMgPsrHg1dOC
a8Y3GRuqWrGItAUMta+gB0VLwY/ocilR09SlR9p6HIJqmcId8CKfzi7UcemCPyeMksM3Ufch5i7d
xt8R3rdEYcy+8mVpne2KgR8VwXuGYZPi1butzWS55ImW+GaLhzuq0P6j4LpKmIm4f7ZLaPG4Sh5j
wzqQEkBClw4Q6qJBmw+d70OC6ain1Ma+sLK+eCG+oUm/BQo/tHBIOKLQo/7IsY9lwyjbaZHGQSV1
Q0+75PRrtk5gr+IVc7EydYvHrS+dEkJpdnvAcGKEOV1xRCviMrAsF2o7GLD6YEqQm6gelngOzEAv
bDtLxg1eH4PgAuCPXV/w6mc+kcx8APCuGSfNmaILMUfQdj+nCj7Z7NyUGBO11PkITenWRz/ko/wX
2ADSVYT1s7N96QQdXy9mrYLT06N4Yc75IrLNBbGBzG2Sx4FHxImTYP37AFD0ZBLaFbvrakdfFPcq
HKxu6xsOEeZqy3yuquUhAXpv4FNNmnzZ9gjVFxttFYEsmrbdnkdddUvOzzc5e+dgFILOtoIrnu0S
UgV46pIknKGbzqNtV3AaH8z29SbiiGG9Z889cqMDghm7dBpjcNEngccV7IBYszRJjyq3hya2xbwL
V9nu/Oxy49hOmvnezxK3BDTlvPb9jDHWbiCcb649fnQZTpQGtDvpiwVlQqB0QFA5nd0Xy/Jg0J+H
HbzhUzkWhi1gn2zHBxShYBUkI7huoCjKJKGu+LofOLufmZ/wvvr8cYwjySgPOPdcBVBi32ZfAu9k
n7aTSyY8vqB5rg7IkfOSCBtAztpNam0LNTRaF/SpBrC2xH7Xew/eou3V7sitF39eWw66GmHo+GI3
PAr5GwgfW4VHkB75/D0+ZLfS9X69WCnUF20vtn92LTS3H/gGEA1+wBD6+/x/eWC25SYahI/Bv8Eh
R5I2LHZWfsRA/Xkh6LIZxy75R7pAFLYcKWtousnspOdDaktZG3vD1T8rvCoDffhfsu1dXN65DaEw
QdpK9Oq3elyalYHNQzaad7T0WBhhAlaL8xti0cHWNlh6X53fzRacddqas53FBrS1jJyD42wIBFKE
+fckxnV9TUjhrTQsoGFqg2exA19LKk5zRuQhJ7vYWO9tK4sfTFwDt48eSIhB3Y5xoTwQNKMZADrR
OtnGmICRRdqe+PiqIrVUUckKjrcnnE0vx9XsnmzkjvB/oaNOuCMIFehrs+/ktKXqxQsSj4/1308n
NceKBFZRtLadvGCO9tIUlskPRQoRLj0PSd7dQ9pvfolpWfV+km0Q9DuDPuX/p+5wypNMiPdSdmD6
lXpgmA/2sjJB4XXmlQRijdcVfD4KRnbP0MbTaooZAfiNqRQY+MCUEYeNcrRj2FKC83XdabRt+rSy
QZF7FSlyQq5rEmNY/YGiNhmumdIYQSHc9Qf4ZTfcG8o3+BYo8hliVyyyXgpFplIduHqmqMLoEuvD
bNYUDjh1a0Fb2xmrO9hkotEOKZ0bnPXx3nzKr1ZCh0bV+AU/WNemxlwh69C1ruTbkFMDMqEH8A8+
IY5y+sbAVzh2qKaN7fKbkXI3UznhpbX/zd4gCD0ttWfTdSXkjTjoqaph0ugx+MtgA6mTpTyGG+OV
HnyYFUxmY8bd/Ul0/X1mirPGMg1KxN7AZP1wUXfOECgx9hhNCI2MeTNZgKvv6eNLSvxJYASbg47+
BWusWJiQz+KUTX9GrNb+eHlhvY7YqrW1SLgPCe/dno3DxycBiFl7F/xNEpTkx4Ep/nBX2EI5s71P
AD7hIPFwqLet2WfB7bGeALOC9+Lx23G3gcRktKwopirNdWuyhVZzO+jtkTpn7RF91bZmEUHcXEzj
9a7e6TR4F6oZ+gYBCwwy6mAYO8caM+K5/Dw+IsbyxBmD2JhNNrulQNTynsTA5MWE+B/IgBPTXLaq
Aq36ff9Pp9U2ZFoj8WIWHRN4q5Kd04hR9uFmWZ1xJY1SCwcf4iTf0YIKPW7Z/TK78CEEN2ET612O
3974VrNSi+yiJD+Bf45C3eigtCMl+dbb2jE9ZIqEt4yUYQxr+pmWqRXgUDRi7ajSsQkeXFryw5au
k8cm312niI1YNJyF+3T0tm3aeOiyUAK7WbcQEhzxpz0D5FWDtttJuQ9O20pmQJ8sWcbsrSuQjS1m
PODO/dwJiVr7vmp5vMJsB5Dcmy9+zWZslIDfgYC1zvQ3NZPnD/G7NzvCX8ggW8jBsZLsDcBzFpN9
WFi1UstdKBwsiYd/0Ch43iOl+ScVHpSxQuVyMIoup9XG3eMAU/LQB/Ai45GHnotDG2ijcursqY6J
DPmqxv1zwnIBCQOmI/tbwFihl7xZdJS8fSPx+8EtDhATgCFH3vdRw8UVfQ20SiT4Vwcime6LReky
rEeSOm30gORTUY8h6UTb4b6Sx4gosaK/6FSm2dZWKJSJlCJceKqRcmeLC6f0L6LyqjYMi463DYWh
heO+xPYRNhu6rQUqF+DhS0bVED1Qz0mBykAncypRZV7901qZedmFA0yLkNS9epLTWq1tCH5x8abP
CiRRUGLybumbUplGY+yY1msk/QShmoap77pXpD9D+tj4z+LNWLoeoHO0s/G1NtIokPqNLkGIzL8d
MJoGWGBpbw9ibp182MmAO8aoHvuMOZIEMnOEGKCcLMRD1db4MF6cqdKhpn27xIqrEEuWaDajqzI/
X8YgIOharntymjTP12EFMSEtuKRzeNxG3Q==
`pragma protect end_protected
