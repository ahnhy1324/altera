// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NCbWtWbWmANJIpMHzPoP5ORUd2lSFnWx+UlAJhhuenHS5dTaslF5mtk+xzfF63ue
f59RSrrlTzzS4XK25OBCnyRttcyC67pZRcr+9SOzWJ/djYiWi/oviaO4umwIVLgi
Ta/gLxduTaJLfS/fguzFC1Y235U3L0ldyo7bXaXByNA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 62144)
HHDvhJP+QgprDFLnHSW5ZzIZSxMKF5gEw2lF/ZOMF73EOGZt/SF8R4c6RHCaiP5t
CLC7zpXbGIDJfQeZDqbkmNpnIoX0vlumrwJA24x14xrLvFEvAFMG4vY3DXoEjul1
H56L8bQDL6nne81++qSnyrPp8VRKMPIJL8Ah5KMJarjJZarL4Uwfhq/VoE7f+cNK
Is+pkexxiA+fCmKxqlqZ5UDJitnysoQ1OwsbdmpOMK5+9GByotRca80jIOku/qNo
K+mucXyzWAmgs29dsfktTOuIHMNFbIyxN3qs2IBPMMD998qWKDqsx7fMfV94h7I1
e3dwLWL5ig12w7a6LPUSqGVRQVxzD7sZm3UTzO6eojT259X4e62MXEem/iA27pLa
/eavYd7MoDqCAYiPn88QTuPpOUHv8uDNS52DdZ0NtcCP/BlAaYT4Kuu93QKloPJl
irhMV40yJK9CKiV2aryn25YGOF6Oko2n1SsgZaaCwyQ9u+9VEng9pBTKow5P9mgU
Q9zYGOmelrNaPDhR8E1hk0E2WHjPcdyNYQx8ymVp8oPgSSxBGwsM/VmfNnxV7NdK
KSDm45y2o/VHqFV6Vfm/FCnAZzC9fj/1a8G5OnU6cIrQtzUumqCfe3lQJ/gmTGK9
aEms7Qw4AbfWBExdXlwCNcRjAS3Q+9Jb+J4Yhc27Mp83t77dsm7Hyz1pFhyHFCOs
R4pywchi4kW/G/f8nHFfwwK5V8vRuuh8SzLqBh9vfwRG02ew7d7deMOS8W8l1ADh
AU451c6q528USADjaHtmoh0WoPbey6lYibRgGqOfhHP4u5jcAkG2o+k5UgJNpvAP
auuoayZVQa0czfaYXZp9zjW9vrxYbYGz+XavS1LFiB8SQxmX6tNCYg+5Cy3xSPrz
9OelNS5fQC6l/CdxET49uZ+9GBOhMb1x97v0IYIVmEaTpFXJ0lmBtDKen8tlM4MH
AU3+9wgEM1NOzyJFaSOUReNG4csDaIrOfyiqjT9535yWp83uOERFJP+B7GvS0AbT
LVF3fZkouO1wu6p8iW7DEHcgOrjozbZ4z/WpDYP0aHfZTTl2BESkcmtu97azybPR
+piSEcF8trNz7olqC1gLrEJRf92qm/9Xj0g93SXnH8aPCauFW+BeHihYljIE3dFW
nzCYbrjmNGqJ+RIT2dkvJ0dn18p4qWazTZNmVNPCG3NucbxnkXmtPsfPX4QH0bPK
jSNdA8AiwRFs7N8DHogoyxZzwLisz/7I265QTqs+pSNetzkMbw/m792iKONmmeSQ
/3YTHn4g4Ss1YCwfGkRroBojytwd+BOHG2JDTZWHZWWlKHexAXQ5OrcXM768n98T
zmbc0prt1BbZZqrBXTeBrfYyzfK98Hd/wedzaFZuxpCDcYlhpNmHrPmJ/Dr+QCxH
AI9++avVqHWE9iMQyX3ZcC31vjeiPAwl1FIMct+8T93r15bDa1giQTNkaKtcUXcR
amwTpHG1TGgyTrtuo+psRapZOvETbXozClmETv6CT+IEW0b8A/LE2OlF0k58hy/d
orRWQx9NMJsqKiGs72+y/CyLuYA6tGiyiy+jG/w/9dOk1Etl34UsjwwbcezEG4zt
RKRQai98fJhS39ONnY9RBl03H0L3ackccwlVXINW8SrP33QFVBRIoHYV3yLVP+A1
MUuk2MjgnVS/Oj15McO74xZAhkfp0YIzxK0d0yOlg1vjCpqPSDSbcql8QJhY2w72
LZ1gTZS8Nr8/3aD0XmXHn9FZfhoiqT+iFZ6xP+DFUfMJnbP3O/q5V/yOzdoNJE+O
7ZIudoHQswBcgjN5rK0p7dSkOljt1nFkJBRWtIdmL/49EbFQHxtQqwhJ0s8A76QF
w9zgiNiCVu75FoQyKWqlAdF+gOWJpBm6SI/bhI6+JjWnFmKit3DuA02mbnonc806
qoaWAwjF2qV9GbI2vz0Qds3ajs7lldE9jnuqKPyc/PhGgQ9KHdbPwKj0byclR/bF
6H24RRa45mpYp5XU20tjJNhlNhTvgyKRgWrN9ibM/bVOxjnLU/2M06rfN2nA3SAk
QvuBtriOZF/I0ecek/JgQDly/ZvKICGZwKrvLo6Swq8kmoMa+VtaaMaiWZTeklLv
xjEpq46ra2nburPf0P01bMmMnUjgvV16qkRx+pI/lbkcvUO/ZrJ5JtOcHYlolola
Gl9TfIewS67OdEwxSZqUV2d8Nezfin1KcVnAyEUDMoWmcR+5Qfr4gVBXgyPJcKfg
Jdc9aFVYiYVY+lXFfrZIGgyPczl3JL7VHi9Q9gY2qpkC/yqh6JE2NJURnkWGrAYT
kjYuM1dW/vbrdkBZyC5/n06TPoAUj+JIk1A965JFOzKaNS110GRVFSFRS6eacZTN
bbhyy1bc5UA9q591a7/Qu2jT5OwIfSQ/aP8Ygx79WLY0df0kw3e3EJLhEl5KF7F9
TEt8GNso8wT29lmwQQytYbPT1R2JpAfXpcJBU9wDF5Lr2jmlABzbzjG7BE+GgrGL
imGrtJtyZyMPCzOZx3y+kkvRc/PME7pyS8fKQ7QWmfZlOeuPkuYpBINWpwsG4Had
tpsMsSU412tExFMgXSmV9E3dQhDOmpYFd3kVNUR4R9lmE8esLVSUjujsJB7ywbaQ
kQxA8VwrbdI3gSYf29CYlYZFKuBof66TUGR+JFOwU1Tks0xxfVxMUgg1g6BksJtn
Uh5TRC7FVgCmwON6PvzPySCf4ppg+XBHkgbdTm3K0t+R9jC/S+a0zjpuay5uIQaq
hcyh5Atlnj8MAHZqvTpvP51vzH8q8//zXc/0CeYuBoZpdFMVXxiYv+CiBpGQ4xlQ
NpMbKgwTtC8wQ9ExDHe7zEr7afB5KE8hxHeTDCtt7FDE1BbmEdv6SOiTHSrpHt4o
7Bu7KRWXhkse8aSqc/JgBPLy5zOAn+FhAJAiZjmJA2VxS+8vQzodMjqWsnFGIySU
ZQqvALFtFKRD/aqMySfXTxjYHyisOjOnfBEBwKQnxtGJOgOJq0e93jL2wYf9rVzb
q9Y7hScPfzlKr4dqiulW9x0UQ0P1Ny3juxscI/yvjdLcCmVLIISLq/5CiHqw5qdj
yZxbEF8piv9x8/hjjHLc4A0ce33CuSBFrBSs6pCIuijAWTa/p4hcPTES51v/cd84
Z2n11M3ogYV3EEw2a/I17JqusvOewCQYoEyvNspL+9e0i7GzhavxQrRtuRSi/q+P
whiYQfrl6bEWcQU23rkf/RWUr8GCmdDkhfycSbygrtourrzT77sYL54HMpAH2kiY
Iwzx9hMxU5oQiuvPaI0coCK5RXVHHoduP8XZdUFgIeqs4TOxU83obtBoLz/Nti8Z
FXQaeWWl4UQ7KYq5ABnZTlk4+3YNxbzq2H1SYiKnmjQg2CqRpSLdzbiXpuzBClAT
RdPYrXQ7HMGQdN2JPNGAvliNPDRPIlznH4jvUvXyiys9qFv437YPAQleqPZFgEt4
JyR54mvqeSzDyPa9kslrx6qtruhkXGgDquFERFSHqteyomIh8tMxKg1XRbU6/Y6r
afR1GI2D4je78j3rBFJQZnP+Ydkl+MY1OlwLEfCtCeNligStiZE39TTrklZXweWc
4fP9f5vJTlecljfzka11u3+Eh/HLNgvtm3Wc+VvgZhMeFRrrzntyACm960drtuPW
Nn1JjJsHt7v+Ga6Z/r0fJ0wGYT1eczAYSUmJLX2KyXaCdz/IRFqGSb8IuVVOi6U2
7nmn4FHIC92PGIK1BjHeQQruzTdbPur2K/ThRnQ0EJPbpYdHkQ4kLj+aUeNLKnRt
tuzb8dHcAbNpsdqdvL7Llxj/n+l08tyiS2BAIzIZIA8VTzw1tiqdY5nPE5pB51Ub
sDS2hPs6fYVXKBSXm5k3Mq2hWHD0Q+qFxh6IUYmx5oBUnPAzmSyzOSI5OiUO/nq1
RWxDFEp0lKVmpqcu2+uW61tyXvJGZqGEb2pOwpVkMJBMNU1BaQl5LUj1i6ozy94x
mTqS0qjRik4tZOmeqxMhXrCpNTvr+h/+deNfjqdT4Ptj3j0HsEkHLTVmNCAZtph4
Qc8vwvdTkRgCggfZs38rZsODkXRCwRGyQkHAktX5ntsYoHRRYJEiB1zTQ7vaYagY
KE5YBO7SLMXVolAiBV5n5NF3rfMbhiobCzEuX1Mh/wGSTC8N4UQWmd50FJXwCgwf
oinPTKkDVnRWsT972DZyx7gj+Z6twqqw2r+KQ/gGP+5ORUjjrtBoaYnRpoADAkNX
NK1bwOqWokE4lJ/EP0aQGgsM6Jjgm3ElOpvLyKb/hPZsgmiPqxlBYhkukopH+pzs
KrRKf3Kzi5uz6GN/LqCsq6C/L6YSNcOHJEXhPn3CtUlGvxs8q7ikXGMonvZ7OWD7
KC5/SjknDxol6j1BGMkpz+hlUK5lepK4Xf2NOraLt9UsMHjMaOkWNxFdtn1AP1fy
crcg7aboKKxzGWwoxDP8Jf77Afkm7kz+W4347UkUpbtJu/5PXyYxe5q0N32JPXXX
T7D/922x9dpBB06UsrPW4+JtWjU/CFNAvgE9tiJNCdBbWqr7BwCF3dBSgbxrzSfi
9x5Vn4mCXLaWNex7KMCwFJog3De3KuFy6H5WBr9dJSrc/Js48ROHkixJ5Tj6r5Ej
Y7g4vjfCGNuO4nbcVheVSf3fpfSFPnrTMwtOS2LSjOwFGoQljBVmcotT16jlwvja
On6N0I8jVbWSS5bP+K1fOBlEPZyhkr05HqE2pdjUl83eSGeBYI4NSRFzRdfh/TML
nGqn1pn84STNQILGhn22DrB6KplL5XHn3kK/Ya4wV3BCUoXAE5iWuUDKaTN60ihV
5aPk57MqnSDZV+rvOvCk6IK0xsXumIYb9G9cOKvi8o4pOeM/fi1M/hVdEOkjjl+g
nWQdZLiBFySoxFWRcSLaLb6KyoqcTH8FrwK3M8FwQ1g7D96IBRnVDOFpSzOkGWia
OcmYp1pvZrEvk9rLTSGiji6kxTC7e2LrDRJSMfTxF3+dWF6KEZhefWoNSrTP93Rd
DxRiRhmLMF0iV9l/smbMr1hHokyN/kApcODbxGrtEEtc0REMcMnUyVfVjym+chpH
vd4kJuntXXdgQy3WtJ+R/VRNzcrn8KIsX7HWwNg8AseGdVWnVVCPe6Ki1/sAzOn7
NSu83jsRt8b3RizsnfE8XIKtUvAsldphIVLcSncSVVMJgle0ko0PFeT3QyzrgtDL
Qr0N3SbXfCWzi4aB5SF3FBzXKZGkLtwNESFUhBciQP8mldn+pa697d8W1DRAWw+7
2mJsUcu581YpouUAwyAMFOfGN79dGPthsNtn4EEjYMLGpbwu9MIPJqO7Cs8ivZO+
bIR1/b7ODVlXqzo2M7/dJXg9RLmOrwlAEMcvK+mfaFgTpzxcYU3XD0SjggLY3+w9
U56drk90wXiH2REWnyzVgjF5TDkL3pU0mruSBJgU53eJUZQkwc08/Grjm3j+PK/g
xZsOXBPsP5yriqiW7fgU1NR+n5EAgLhSbOHSonOQ8fz3JF0F+iPon4zYtIJJd9jm
IjS5eIns9qaJDRAziWgzSg4BOmV7PMr8/JA3nm1BqTfF/Jj2UGe54kJHUedlph/S
9kquqNULssbdFiKxDoSeMqIiZPfaZnyn7jNFG6Dr1/p2opAoR+3643ipwPbl69gP
+32Z59AjrKuvTLESQcJKIIIkqmknRwM9pqSI2EXVFTQ0BOioriRJvNPLxShLzm0y
/kTB+Z91SCqrCtSsjh6aPdAZsFZtpTiS8LXu8SjWbA0onOIJLgTdA2eVLvsz0rE4
fjmBCOJjDz33eUirR+CAC4G/AY0vYOvBcKpzl79LUKCKKSr3uIRww3NbaQ+vJbbd
WXXZtc2skIX8sTjuo2pzvWIsbrqkybAWsxYIlsBbss4GbNaJz3VTrNaa24nm44IN
FykEDk4Y4hnxMdP9c3Qyz+0JAAVMlyNFB6+w6wOp4uSYdVeyYb1q5P5ZGIq0oBex
n9soMaxODPIZ78ILVtHekCpJOifLQw9n+uZXee4nqk+7V9lZ3fCbzc69+PW2lU8m
FGQY5z3CPXO8kK5lRAJCNgR4+nFUL3w+/vrMwN1e+G+s67zuNhQ5RO26mC3DojoT
k3XNDgrGOB5XFUkWG0MROuA3OUIv3Jx1NyzBh1lj0KMH9yRi1FQpz8pUQJ9Imvzh
gxmD9NzZdDdk4VdpPCqZsYgo1vmZFqPGlg275y3b0EuRedFjuPC9/y/tkgVIdxht
LoN0/ZBZO0kdsyDO4ufIuR07Xcoy6VqVS9nSCX6yvA2DEJLx/H2B3pBUNstcoK4k
bBuhkTUYOtBw72Wu2S3+Bci6hMHsNI5Av+bg6TF0Y2579YZv4qs6jqxohb1EaPwv
bMyO6OcQUJfvZVWaHsscjvXfaijwBjy9H3ZgrJSIgtfKLU8Ybte4U6LsyNA+qSEq
7ffEVtloGcNxyrVqaEipj2XV1bgGQs9DHgwCK/+GM8W52sz6nWjqBu1t7B7cKW9r
dpijqfKm5TktroneTXOLoEXpA8ARAhebaj2i6KuxX/z+VpqrqvLYW7iXFTuzFbti
DkAhvlyBW9z2XhLRt5b8SUiG4J1+UpIaswQnHDcnBw4QDNYXBHJQmdD1a+iQpS09
cQq+TS+azJGfczoFeu3lo3TMrq6kTCXgIOWr5AwKlZBc8wCQqZH0VmYqOqnvnVh7
WVvXb3NQlbtlm8lbPi3z278OO218Fci5wsfaNNY7olEsQkjpqPw0Jb7v52uxzcRB
0wxENyGxsmqMcmUMJAbP7jikI1hj0AGF6VfxwE04kPIbIGSbBxJH7qEL48gUNNjG
RrEWp+S6h0nN6QaVIF7Gx4VtLap7obKOLChbDqbmeOVLmVIN+CxRvITrbvqM/6H/
IxuxMysRzbdyn79v1v4nB25q7bSMCLLAyEJV6J3TCQ4UJd/id1LYJpcrep+LJO5V
bQfiWDiNNeEimLgUlnfCcEt51McMkg0OFXVN7XGvMfVCNDxiiTHn94fKqpvYYIUu
NQYPidyyX+1u8u1kj+7ERfUoncj3zwUXqec2OTIb1vfgVvKvxyhhSi1q3ukZR1rf
1ugdygZOhVnaeEzjGj4HneLkMa5TpZQH1rETz6nJj5d0ynWOAx+Y8dEVwOe02f4R
PeRjs1RqwHxCGCY6xr8KrjqRbrSOse9fj3a2pmzDsBepe9owqRNaMNZ5rRxq52uc
psyvH+w8YiTY3Lk/iwY/DGZPnhsAW2Z7trPA/bdQd3oq9ZGrSJj5rx1/gmY03fBy
tzGPpVJGsMDNSzc86VZob8dDkJWb1MTxWTueO3mhv+IfcHcpSMb7l4VGFy3Dsqbx
PyZUNpfWSo2FdIS0xKS0bgAKtIusq1pk57uTMjkzfCrbZ728rLhhN65PLMiL3Y3l
aYUGhXVZ0vNlhEJCdMeV9T5+Dd5zHzaCAzN19gydD0CFz8mqo34bcPPbA1IP5Auu
2nszHH/Np1e/EIrJf2wrJkZf9urRLESUH8vVfmCupJW/EY6Kkx8HYc32dSky/GIl
bFyfJSdlUGKVngkevTAIPaeEjNuuR4Ci0pCw0FRj82VMQJ1PcgCbTFipHlQHGXhm
nDnQ1fHrlPWe+d7kTQqVRXnzgQwJAIs9klImm6OA+jbHOLa2bHG1KQOXL6PepJiW
+ds25QO4iVC7Ye4T/MAhmHXW5v17/f1n6m9WFUe83wuL2lvanbSg/HCnpu7ZLJXB
fvzle/plwXj9OpFqFvd2cVpAFqaXBszYsKlxEZck1ezXgAicKAHqLjl55Rb+n4cs
zFlt0ZOkZVk3/Sw5G9GnCpx/zBMMVfkxrQ885bXNLBkdZ9PAk2cc5DjHMYjixUsW
8/WMmgqYqkbIZ8Lxx0knYVcGwbhOvQkCJP54GzhyVaoc/n7f9WC51iBmAkVm3BrC
V0VSWn8zp3IXCipFmP8MSJOq5r7yOsVPYDu9GQ//rFgg3gCVzA3mM4Rik0ZZYcoV
P+f6TB31p36ThWEVqPSGTQplF+Efsio2DpxmPEmKK4wLI69nRHT6UUm59qQjp7gU
6HRXBP+OzGhbPugipzBfx1xhetHmlQpf4Mk9/jNlvd7kyG7Xe56jaKMYbYcU2w7z
VUPTF29oQOVgj0sEF5y3/T/Rcs14cWpQmFj2u4cuTrRdxtMpWtxLKUI0ivO2iosn
gz8sJd+PFxNzt5fhM55pbtoioVYBA6RSW+gTkng6E9RCwKVHaRx4yeJcOgEn5kzd
ii3JoAUJWXnRcuUqD547IwfU7c43Xb5XVg0VnDh+gfc08w734gkG2onYknQ7Yu47
L0n+J8GfSjZQk0Pk/sJXg4JyXJRQAyug3YLUZ1qoEIRP3gbjHZHrD30DZi9W11TO
cjC9HvLUPIU6jgZ1ztF/ubnoOGsl9Mfy/hCKem9DaBRvckTPT/LbqIz8b23t/cWd
/fGR0olTxblHY+89DoiRdYxrp6NuJAXQ1TJL5YB+4qxb7ZoSNjFVAEIBJLt+BaUo
AGDzDcKdtaGPVW0JMlxb13xX343xYIzK8AymBJlEPisIzgDC4nPLpaDJV3cn7BC5
i/rlLWuHYMRtCLxHFY+h1fhn2mEtSYn94tolcqslxweX1mUBbDcpvyYrHcOlMieo
WGjMrbZpURwGUkZNR3tp81bXY/Ic+8u0ZOpbdT21X+GnrjhABt71cOtdY7js8OOR
PnlZDEv6zSk7nUHfXVL6/6JX8KWvyceONHOyHPxZu8+h+1B0+DGjDhr9OCKzApa0
w+6CIG4Eun/yCHEVUmcs+AJh3MMe1RUUEtTQfiAER56gI5nzQOYMuJO3n9Cop1zt
hx4VnR01ddBUpX36V/RdthtjEeX3XMAcUglJmQGokEyPYQ+uyR0KBB0V0ANEXS+M
I2Y3nXTlHF5cfj0c1w3AuhSx8bkx86mg7RvKLQ5W05DPYfqL1wkJYleALgw6STuj
uJ+QCSU1xNztH281lEmUdSvff37nJU6z0EldHcnPI27S0F4lkOQwKXgozzaWFz3B
Z8HWbCCY3w3sj+pl713DpkZQpWYtiMcW+cTV2p+3EbkGojNz8D12aWqhZP+/x6vM
psQC6bMIRRHyt7v4Q+zBCgeb1UaWvV2Oz8S4MK5SNXbFOj9YYE7CE1Uh/zLYkjv8
DgEAiPci2gMHz3m1YyC5/DAdFmi3vekoFE/ecuORkN20Xj8YGN5pIUKXVEOEFYoU
8dNJ4qTYq71+t9tg7G4H6ZUSvOVv1E6kAQjN9UWt0XoKwARqg64UrOokqIHsz14I
wLcidQ8d6jnqgol2nZsoUQAF3FphFDb9G15Qu9B4QiPSla+x/O1MCTgy/kWDRswP
ZXdvl3IQnh52ZTsyRVy9GWemmKLrJskUKO0Ln2qIqMmow8bLz4+2DYc7AeIqw9Gn
rPNmbjDw7ZlBNJQEB+oODHafOynVGCfNQh0/VtGaPPOqsR66DZgvbcKTeFZ4JWGW
rv1PQ142cDMFt49Fk7oLA8Zj/q6FtNs4L7aOlmfRZBhv8S8Fxg3wCM8QJWbt0X3f
UKS6QYfKLosOYFRW7WcGz/6upv36SzX1UKCm/19tnc7W7RTvfNHBFsj1+yjMj94v
Ah75KrZkikInNaIuITtBdIcno4xqnuwJmoAdLfWB+vNlOeTRi0WucD8eYiG19EVe
xCUUu/290EBFfARIOV6+0Tp/Zh8Onh6lV3YOlIo5DfdP1K4f/1VgfrGqxfvVYbF4
YzSJnOXL8WFfr7bhZYaahXN4W4reqNzveT+7HDwxWzC/pzayXw4E2va9DtKHP0GT
n/UshiCvqSo8+mpzA4E2XJdrTo19Zt/pbZf6AVieRL+OMhnx0CtxpsC6bF7GR1xm
gtVuUgDZ2/fPfzPbvLMO59B8PLVeBexXrgd9Jfsf/6Z0rYWwR5VP+6FK27IhJMzK
DCl8y+Lp3Aq6nmolZ+iAiL5ka8/XSz99dCfasxVxRuVYvYtv88407PHufI3RdAHb
2haXwuVKTi+tWHebN96tTT3a+L5f00MvcDJWitRJHcozoHxKnishW1Tqr7l53EgP
1UZZFKW+94d83byEq2T59x42GcwT+XHeg6R5/7bkVtBenKIlKModc+r0/xhXPo02
W7OBldrf4zcV1QZNnXOanAfQesK2lGjPOLQduefVqv34u0qkQ/USTGV+cN1rYdn5
LARwL1wKV08tolnFMtyDz1yyZsfFLYgo/j9m2gSIUABd08Vo/Gt3+fy++6LBG7iH
7CYIJMED6Do6NJILMMd/d4J81fmgDxWcEkyYumA1XB0etAqneUr6Kk6pU/asg3LY
5kxeUQkaKRLkixGJgJ6KmE/r6/om90dXcFAyPOt8bL3Hi3M8U78INQhvh1fio7MX
Lyewy2mzdq2WN49cBoH2HLl8CZoyekesU3wnjAzPRWFYNXzVsW/bKvgPMglGOUu8
SKszTo+Z2NLKtrgDpGKh26Hsxh9h6iWeh/H1Ku6ZT5EHIQ7mKt9vET/zFzM0BWn8
d2XdyYAc0fFtGRrhQzvOvIIOGGBX9MbuOfufGnoMKcHTAdMgrKUW7yp5Ax0/h5qf
3DYlHERB2rj/PX0zQJq/MBUsdbucYv+Tvhzt7IbJe/TnFm3xvvYGtp7NjP3EPlmK
fvvK0LPPViMBd9woRlDGnrAVhR3xnGMCeQHTHpFXPe7OuzjCm9Gg0CSSYhjKHeyU
ZA1rviEHmNQj8uWQeBWwOePNx8rptTQ8Ps9LScRghKQ39xnAnobhYOO4p5pfoPte
WNzu4yjtikmclp30DLDK7od7fhy++oLrkcRcq5agCuK++wxb9R8cAqAPVOfmbXLL
69hBaMUAs5AGfSK3IlB+oxPPKpi+s2k5LvbEG3N0gW7p2yw4ywn7yooUS7jm2thn
xiGH5sJBwZDa2wL6TsjlD4uHFliXPyt0yjlw7CbPDp2m/RWd5/X0NzjtAi/u3Spe
s6u+E/R/h4RIr1oOnv/d2FS1Qkvw8QMYPrhQxDw87XQuz98Y28Kz/FGSaSiwB7P1
ql5VoX8VKjri4k0DiQNQye9C7o0rxamYG2/6lxbpOogdwRcq/X95l5ts7oeSJJgb
EvO7zZOKK9xHsVGKaAzD79HVBXeCu8wxq5IuQlRtQN/SV5zh9ryBcfkzQfyKZze3
N8rAFyJ/tQPSdHeOcFZhkyac2SBIjHSY/djqgX1lq5x8nThDRwGMBBNVHOmLZchq
2kDGSQtftpsBTm3qSYbA1HlO2wr+XkgbuBe4fviJuuqz9dGZlC5gVMrm1216M0/e
82M0O4NpGzL7EQiJf9Btl1TNTgUG295JiTPP8VZDGdLhphFQ/Ovo5R0Y7O4bjoce
hu59JYpi5wr6vngIMYhsX3GN+ig2+wDehajmVQGwYJH1hV9083prOj2J4gt029lC
NPKtCH8VUBTPcY63XawiBjC6UdTn87WORUwOo6/NPNi/vOJTDVvzgRk8C7StV0NV
idkzUpQFMSAw7reJIxaGETXZsEFHWHRZhoyxpatlUkB2zPcqFOkP6Zd0+1C2xCh+
6KVPJbeahsQ+XofRT/WEFkHadbnDfnCy2oNEjPNDxIfBkdC0SNqD2x2AFTGDf23c
dTtlz1UFIAHA+jgyD2NPelAK8/hDs/VCsQLGbU+Pyqv/NwXb2TwBNksJlvUmHHkZ
W21rYJdwwG5Gdinb1SH6IgXd8ARDQft+u/txJ92dsQtMmeuGuY8G0bgeRIPecwzN
S2+rzHufQTaEoPL9d+bFdMpPE8LRNE7CXIsWy3cnnnNUKFSeHJL/UKEzzc4E/KcQ
+QEmMOp6WklNoZRluoygX4RgvsdhZn7ix4fs+865iNdGp1Pqz0s9mUYWyimICjzz
xm7UrCZ3GbKR2BWrvF4tvWycQBOvnX8l2xoX8VJFkMoeNFP/Ao5aGdOI+wpKovgB
m+bPuC3pMp5ovCO/6hn9dPaj5w24uHTEKbf2M2XJlMFhCYMm7MA1BnzPY9PZkITn
kBvzheR+3sDiKjbmWjJ4tsUO+V5m13jWTX8EKFg6Uf2sF7pHV+I3HgrikAt9LjAZ
4Rnxv9aM0odrIApQ19Z5EhA0QfC+qCrDjrRVloXDUWHLGz/ji56RseT5PsNnG/aV
yiRmG2cuFOZr//CiK+vnUTQxh4J6+99I8WNKkT2BuQ9+Rk50hJxzwQbRWim8B9Ra
R9OmVqFx6ciwQGFol9bbCBIatiJJN/zoVfkANtvUq5JIle7JeJU7vD2YtRBRYFx3
fOfJnz8Rg8iUebhqrJiI1dGn2A503BFJGvaFDSDsQ5fpP5brA4WEH07kAb4h0T3v
VAWyUW/LkxTLkZo6TP/r8pyncetF9QungOgrixPWzPxliEXnVkt5mtdAelosGXTm
kTtYD6TaVUhhjY7UiFXVNJhWIMhnI7O7UIxf2mxWzTjoiMH2bB9Gyj3ysoyez9DD
PxW8VE9i4GgBC6GqIReU6QCLoijBrdC0dKPqPq8PsrXbUPPi0JNOhgvZQBTrt/aW
UWmxppUrmuiy3jQ8CaiNs+DPo9LeNa8sKbB3CW8gqiM2IZjhhP2WZ5dusxvXovDI
cGgRwrEcIi6TEyqE6qC6jspqlGpKpbI8oNi9NNd0l9l+CKgdfOeucqXRJqYjB+8I
ivzeaZtjBk7ogGIuRN5bzA9sJ2OQQbikV9tJb05qtYDpTzTrta5Cd9x+xUnd2EmD
HDlI6+ep14VEk3Mzun6VjDiyfsoCeB70V/X/uj8CVHzCpLAVkkYnO87EKJXA0o/+
nD4CyJd9HtPZO9akIhDEKM1AeT7WQKiEmysZjMHeU2XGjroYWqxH9Zoy41m66NLY
X3J1VxF+t2PYf5Q420ynlGLi073Zta4QeTKx9KGsY1NHb3CcRcMfVwd8FAU6dTru
RR7QH9ORINmEhz6P3ZRFQ+/dXmZAqmtZwS8nYkF2Y8XzdlIMRdcVRa5tDNKeJejO
AFQDdYbTbwPxQazB93RRiPPL4Y1iInOgBI0iDHrEsjwcL6u51LCtVbIs5+17hFj0
RyWoS+ISDuPKzJuyZ/YWpGRaqaoWUP92ZAezCIAh5mjUUL0FKiehiD6Sclf+HqZE
EW+Lai3i5q8G6SQ4NlSn/OcokcPW1L5y5UV28gQmyH2dS2Ui7wXPqN0SW63vSC7U
6zBjKwxdapOCqokhhK7PIy9+RkDqlFMeO3tHq+5yt15w1Bb4XSGZJp/XlYFxe2BN
TVEDdkpjuIyZ8ox2TY7oC+hemooStfDvhkWFs7iGpUyXCI7Zzzl2iayZyCJlFkKM
Bh47FavKJj7afa2VU0TlGulITsmvzcNnHifBZVKo22suyDt576FcyEDGegjjY/qa
RTLc6Xr3LxviY6gYa1+MbFvEKKLePQFXUEt+Ej5+V9GJ2ukcs4V7Nb20pgjyp51t
EaaD/p7u4SKC026bbuRzX+z9jWUJVGPFP90T43zEP3Q8oeYRNdyv562RBfWd4+y8
3n2Mt00rCCA6QrIbqISYeHmx7gGoslUSugIIHDqiUz2Qz5k0Y/tC9RsqpiUmk4Cz
r+KOzH0sMchEwZVBPxZP7HF6Ypj/5wGW2Zn07VOEYTxkQCj+0HV2DEVa+TR0IU+Z
3DOAAQI2B8BcQDSnzQEEXgwSE3/AptkMbkze4H29y0GBHK5dGQOjJuH0JJMZ7wHI
i1UhegdxdZ/ceaMFQYlN4yqZhm7/DMGIE9NLLq1tt2KNQUMdzGipCBgU6lbjp6NK
g0Ksz//RF8St4l5yGun1+H18xrmUp8LwuR1dvFRaEkOsVozJEyf7s0o9Vu2yKOLi
Zs6RCmPjFjw8drGuQN2vyVT86lv9HuWKHBZl2LgKNXLFqhR94/shkZhxxYmYmsnh
wp97u0a6oYtMuOq5iEWl9+lnT6PeOb1+GpR9Q50qpALLh15Lmn9prip54tBeWCWa
zJo4/hSTzF9uNaMhd8f0hE9jlUq7HwWUNMMOBpfkNYECegd+v36+5f78U5YLqbz/
XTispbcwr3ClYJ/7KfOOLyuNetuVZZb9te6SPqlQsZdTjaMtfIdalU48dpMWBcCX
4yxKFm7PDBqqyxyZDqEp+MFtdPxlVehxN2jEqvzW5jOHhhHEDXUVq3nnmDmO2eG+
+4SugjsfkjdlE62lquBAUZH0iNiqDmXzvELgb5v1B9ahaRfFJenu3PiHvRMELi8T
oP2LLBJ1w43aThQdbc0XSqYJHCx8Ok6ZNzauQbvMqdMf6TWIZaXgzCPdzqc76CAL
wZGnoKalGgaTIXl62jzUvvcvexcov8wuc/5oWNTq3l55Ym3AoCmwFpf9pUcxDIEs
TVM1wiroF/voHUCLT7H14Nv+sPbRpZ7gbU0Jgf+GkCfmP3Nmt0qoWF81UpcX5Osy
MHGn7QTUSdKiSTXAKIADG2xo/hLOb0ne3H3UwQUHfT2aDKCguqyXUJPixHn9UWrC
faK2qT+MahwTyAiVf+rw3sn7aAtBuEZfarrRjsNCHpTlp00KT7H6UJXLBdazXbbA
78eOKYDAsl/JMnzSgwwqD7nUUD1LunufaifVlHrvpqRP8iEti8xaYtefe0L+vx2H
cpN59u0CVUtCzi7INd6MYIhWMiHKcURrO5LduSCZ5bD/Mt88Y9aRvid/8oDx9yS1
wOiKsNvOYG+v+6sOMnxoDgCLQBvHpeisC1MIRG5zfYXnABA/vDgFqvc9lIg9hggp
IVcmuJhNCD+I/bYs4XqUU0z7EGfP9NRw1FFrJo1if+eNLVZnbe0lbQgMXWXvVvN5
EZOmNbZ6qCA8Kw/13sg5gN1QOujBJyFer4ToyrcJ3Xtozz/zLN3PF2Vwon0xLiRm
nyPbb/m0DOHf/SSwX8ZywxWXoze6ZsUFO91K1DFKEci7wpPOFnLuFh5LgwEzi/ke
m+Mt8LIBmtYTTpf9ix48uJ/GLGG/5rTFiJGMEz2NOZfyiyMSInqA6Qd10nSbw8s1
ueiE884ZlMGUGrEo2xBtLutY8jW9sjyU6N/Juw4kToMjQmGSYL0JJydU1PXTSXvB
hmV9wgZLAfWK1G1RIOfJooc5zHL3JgH5HS9l50JN0avTs1BYDd3kY0maw0oGjmta
X2HCZiCntwaEVGnOKAcIaOsU0gFAdw//jecLP6k5LfBcwYivasBUNdS7Itdxd0uP
rqb35ZsF2DZzQFsKuIFAnoxXljm+PbSH+kqi61D2wqJcKqcsQPxpTTopRWGlx4Qg
QnW4lnAbaiv0V4w20eretmL8dgYkZsTreY6SY7zAAOxjw1hx3I4y23749cNVo22x
IYP22TgY/kcWMMmlrQHP7wBE7uh14zMPLM3PcQ9cffQc9/+CO9tyNEubsRQEyPAQ
8oEm+tvz1S6ehIUWO5j+yH7rBKvOO9l69N9mOGuxXV347Y7BEy8vMh0Z5niCA/CO
n9zRDPbPN7Y7JtHxCcKPLx+oNvJu3d7+Ix5a8zj3A6MzyS3XE/ckkXuPerUGgCVV
/Rg6yFfHgS6rhSwdLZYbVNcaq6Jy54pUzlsnbpofbt96hLqHK0OxjtfUD3uS45nu
dpUemqu6Y7Mmvo+wqiteodrPU5At+pQ/LOMJyi3Z2GeHwzQ1+K8C/d9vLPDqqzEa
nM7lEo9O8TXzueOzsQonW1UUB+NbjUGMsxGipa2E3f4SCYqgJgyrHtGahB1y4XH9
UxXe3uteFdV3FaDDRtBEw4jzbma+hWH0HeKKUG50jyDb5i6FL8ifevL2V9+4WjBa
ISSLYidS8bLsFeJQFk9VqMDTCV9o4Tome0cn4K8qlOsJWMVrcFkLS8ZM5TeBtRj9
CzoS9E6hr2O8tGILluuS1yZkyn+vvnwAoMS397rBibDig5gdHjW7yLAXE7vKorPq
kUnRtL7SIbUHRuWJBR5wAdJcWavHUfaqTOTWnAzsZa0H8DTy0l5z1EPs1FEIYSB1
xqInstqalWezZAiTv7070u+x2NuTy4EQ6x3vH58tXhvh3pRVIi0lSpgelyCyt15e
82HphbMS9H8nLdy3iAXe45NdoAyXfw01UDPmV7UEMuYNJ0WlMI1JHcUFGG1WpI3o
4CxV55609a/q/40QSR7/pMR+gnI3Wz3bkAGVZU7Rz8k1qX/I/TDI7fRdQfqzP9LF
xcuwO8c2S5M4owvHShl4wLiXYeSN7uiz/MCeTTr03xEEmKGYTGso+rPqrE/M3sMC
wxvfS8rLRpw7ktuCM7WPltE3/X3iX8WHfNYsX2jZuecYmwYN+KQp3HyQAPb+MouT
/Em/pZyDMwYuQET53eXO7t2/HpOGwE6xB5EPWkLunfn+ygE6poin3A69a13jqvb/
YUCtxH74Kxi8nPu4hiUhfEowg7ZNanRq1N/ThIr5h41Xy0KI+nYBfmcoa4elKf6E
7rFzGrtk+z/Dy8IxAhfe4pjt8/wRhHhX3mxrYwx6EZTVa1QCMTEV0tdou3eCUtaw
ikhNyBgPqtV7XHlY2Gc+GeSX7jDclRDjM92zUtNbU+5XWBKYNR7Oxj8Fe9ETO8GW
84PberAE/9nosuJLqHZd6NBkdjhjc25Wgz0h3zEHf6ApiAN5zB+IA8HaHjCaFO5J
tc+GtTWdZyUd0L4NRjUFUCefy91iGM5DqZfJkZ2XNeQMWrG4h0cIRzOP6U2zHWlp
z/Zn9FAgY6dI8ei3iW9amd4j7+jG7foAGlLcVh28iEeu10Bzkig8gPtI9dyTu5Hr
t8uPNjWQ79O2FDsRr39diuSW9JO79RbUoo8G+KLIbg1fYm1X/vnZhLHqK11HpGUL
Ps28bDvlwejUxIT/srlB7FUIF02kUaZy7Yp1L/OwPt5ALKCHSQ6w1kgeikSDFERO
usBC5WdA+YsLfccQND27sNSl3CcP+H/F7Ts1Yicn2Ntqj/eg+Jn6b3y70le8p9lk
SmSckVoVR2N2qp4kMUn+MpH4UKfS35I4O+DtoPgiLC+u0+L1RFD7szmV7SrqBZM9
wBihXZvKQZn9Q0c+Cc9+t10ho2/4wl8DntI7wgOdR38ItgdMn3NqeD4p/noPNjSH
c5nxwpcPOiffvp5c8dRMhOuXV8+UE6OS8sPFLkTpqOPcPrT7JKu1Asb74/2zp6k6
b6S8jIb1O2CvjvUlaEFVEjFxNuf7+v51ht+DsthyRtkNMRViS7NSzolxY0207Ybw
SSyHzj3Yovvyl9LUMzERxw8Ar/UCpUqH2T5Ut5DzOnNzOnrGq3ZK+px5/BXFQNVw
i3bVtakNBOfv2OS+FElmnRw0FBnKtedFlcKE9jd6DQtlyMDyAE1/SuObO90kp8RB
cTqra8+lLK6Cmol9kz2R9TWmxzacYBGqY+kOwk3JFbd1N0vYr/S4UEAGcvFa4yci
0R1Png9KLWM9lY1S7A68rITXNLuRrZhp81jy0Z/vPlqwk4Qgq1L7yVADCrG/K2iB
i3IHmlpTcM9ayR9q1G5lx0TQELsdVIQPXF4mWfkKd+g9UOxKLbiJ7RRUCrXI60Z5
i/olDNykzLO2FEQRusgak3WXlaYoFp2RSGQA3S0+TzbIuI1wZUZMvBDsV6G8tAFL
7IEKyrkgaXRn0EtxHlV91zmbxYCyUP3kCYSNGsx+TbFr0c2wEZb6QAz1lFmUz+fY
nsv+qMsCAmJFCNtWeO7/nomqQRYSbdbh/xTGPlcic4zGDMiSw2dLgIPCjgRJXoVP
nWYCqVvyt5boyyMnfTQ9jM8mgYbIcDkmkUNkXl+xFsd2/IFH0LFBehY6JfvwiG5a
4UWBIujtJyOMirlUconZpLi4qCcoQbAIR+hUxZg3exjPSP6w1hafr5ElHuq8tTxl
9TOAgj6dTCL1tUphFgcLXyGRdJFIBxQcIYJ4mEYUvliRHJUJfxPYNUVJ+8lhEtCj
9uAs9dwz1Z+9SNnqGmHIjt57r7v+NAC0FbPdj8n5hWBlgFKLOAtPnnLl5tQIvGGj
udoFTLsFJyLNwl9orw+NJyVHa8au0PtpUroFEOoaM2ZyNz6nXk2HFmwkS5NoZ+cL
6KM6gtiLU5fWy6+8/1k7dtwItdmrjmCAgsMw2p+ov5zGfx2fDzfP8PHsnN6V2dIp
sTbejtirWvcV6Ttfw3IfUQqmyfB+9q32Wz6OQF3fr5RgrHD+Ao7hBA+G/kIsW8f8
DWt6pz3FhkeEPm9rOyBgXmikl5GasOyNpZo2obUtWg7VfvDoSFmSvIEzWVO8yprz
NrewVFD8qzFjlggUH21XEwct+bsUe/k9ezQjmi+AGn46XxcfE6pjXM8t3dI5X5Yc
v451HcKSTLjENjgZGYJ09J9B8xV/UFx5UWgWs8UpfdeZH8RMuM6Bduq4bW/TeBAR
+oi3DdpAfwAi2v2QOAknDt6/VmeuVgIPNiG7pE88fhs5b1RBqlri6JHLl8nLDGhv
xXz61eFipFkSDVHvv/sFpUMR2fI74/sQ24tjrTO9H5QKFJ2uDCR2XtdQv4E5FrsI
dty0lD6p1BWMl44G8pXC7aGDn+EVg1DKowMViOYGAf6O/nOQ40UTPQ0skzWO9hUw
E5XydccAEPtgSaZIWfFZcN26t0H8YxgNBVsMqFulBlhGr7bz0AZ1WIgfX6kHrSau
5KXgyFoK0PVqEtj7eM5UljnafxKSBXVTy2NtOwHM3C9lLmsC53uutcJ6yx8rTVph
zxJkj80dabb1SccA5serOnp8D3ra6ob3t6PqLJZp0rivUS4my/Cct1QFYzTyYSt2
04SLgIa//bpkrAGe6sXnQUXU0qieckcHpoEKLvbKLGtR34xCnt1yvapE6rgULJX8
wBtbBuE3hcNanvjcxD7GbENmRzZG5rgdIyPNSTBOZeyeKuIVG7OZUW6LWP3HhUxX
gp+ku/gpjrUYHBrDLuwU2ur3+JfL2iYI38omsugAaDEAT8eYYBYaOGaaLJuTK3Hh
l4EaGbISj1KOQfrtx72daktNPBnzGjKjC5mxYzbb6nQCyd00QR0zx0nkCugcFZll
G84sLq9llGlO8EPEF79gq78cH+9lhNogtIoqK9DZtkDPlcL11OFjtIMdUdc01pO7
oN74qKYET7S9ZE01YBYKiJ+2kgY43SVMSXnM1DXgbhrwcROPdYkFzluEAupPQ4NG
qOPwm8mlILFJMulaYAbBqxq82cjKViFffjMvHnp5d+tH+oduwwxBN/4bgEjGgMU8
ZjaUMjxmKq6Awwv6wYi1wiTzO/RcLdNa+5Hmujmj1Jcn0yZIobAfOZgz3FkVZwVn
WujBs3ep4TiQYdNZ8Plmop+lj2vNbCWH0Q0A3A/hZf7GF6RLzp+u/mEF9pw547HT
WetYq4WP4/1bP32DeTM85Vi1LfNn5+siyLN53Je8P6uv8mn7HLWLhoBsJiXO9XQ1
/xiIZKW9n2w7bQI/qi8UaNafUJFXQ6UE+/bdB1tKnjOfPqUJGXQ6s5qSIbUYKV3P
xU9sFWAl1nPxeOH5mmwnLQ4sx1Am36WfPTv8QSimfGF2sFnm763+j0gXtxB5BgwH
ot1ycW7C3BPsWe+rRvM9NTXecj+tOVVlvGoJW0rbYu0UnWoieXhKPwN1Ao94twcL
PnNxTgFRFhXSZTtn9DsDHujoCcEwJEg3Ite/EN81FMGN9YYXhtbKcUj5gJOT18p7
DoFrVDsTciG0zPbMbBdyQrxLxzAiQjfF3SEmMcN3Ml1sIU7z843MFEJXfvv73MGE
zxz0IzmYdSK3BICvAJ1Jzj1SjoXI8km67QCzecN9FVXk9SpT/lxuWHOmKy5KZFj+
RJ2tRYMhc1Sg7cb2DzkQBOgSvpiTd/zCUAMgDgTUMfeEVVjEOu+xVBCEGnwDAr9A
rAZi6df5LnTh0d1dv/1b1vxGYflrZjtpkzesmOAhaM7iAzEqt1mY7OKJNWdJqkp/
oawkWRyCC5N/y5EuoYf4yZ4JSJ5xIaTnKsZMUV+IUdS5p/J3DXH/nxXiA3FM1uYr
s0pHfBQ7eWjD6Paa4MrKiBZroqjmBqRPSoQNu6ENoqbdp3CleaH3a/3dLqczVxkA
c8mKxzG0espojN+LxE+yEWocWkjcntIf2hfTxacrZ9X3/OD6jzpDkVAgjdjw3Y3k
eaTN1T34dTmlrzyFd9Ou0kKjcP5ZIl3YzWfYfp6I1ojKbv1gxY8jLS8Jvr3qOunN
uOZx2I0cRCmvb9fJivqgOpEE/d97RdA1SW84N3PXb87yyMywUeTDq50NUc6hLpLU
JJkbRmGgUzsO/cCqfyi+cOPtgQqtPuiDwNl5Q27okC5DdP/CF8px9y20SX+5BIem
od/bXjOl3u33x/UQ6z4DuYcGfeuXOLPNGPMt4CHG9jC0Rr2o9b/dgUl89TBU2mRv
CEm5h3+04xSRpg1b6G6hXKqrSbzhPCVXKy4z5uhCOcOSnofePraMxqiUoN1UKGwx
FJ6+HiCHwTNFj4R4SKWLBkgRmBR23DTGEMx9A2sNALlkIX6qGLtp3B4HRb/6RzcI
o1i575YqO7Hu58n0zn957KBaKwHC+HatDbojNFDdpTgd67nT4P0Cry9tNiCrgkHX
Xah1BTyfoYwnPP4+RcsCmI1r6vZmJ+rnbvAfLss2CBUsc4KSn8L/QK746t2EtaIS
d8VgxPybIqrWxlCMXlbtgwV3Ojw1gL0vF9z1UT+CQ8uYL7yO1E0h/ZMqFRAp1gHl
DUDFF+mhab0sbXNhV0FVjFhzRN+I3jlf2AfeE9rgkikl/dt2Y+W01X+WdggotO/7
rKxqR2opeJSZmJEEMHiTtqsPyjCpz070T7Gt/bvEi9/cSo2FSADCoJRQ03sqMNIP
l7JFQFK/RCLNl+WZY31JDLCnuQeH8veNlD2Sbu1ZmjkF04AggyXzgEC3LZiiDZBa
heGj3ozpon77PSJFkb5kj3SJ5Wc1wuZsa4Z6jofFWxw4ZVw4OyFzIDt7HqGhWzDd
tEPM3/EbByfxTFfCXpfI+4ZgP3yyOMJpSzaHZakBZrX9pAUPdQ553ugjnCiIcGJd
RXuDzBLu4sOBrhvEc7kLNaPEhorb3NT5MfbiO69D8l9WpHSTT/Fs6yBtposaXWd3
RWyNWRj4rN9Kk+BIY9B2CUWnI1gvtjNRNj0O6yQ7rgVqHAdtnUw8iTD8cohrM/jo
fe4Xc/4JOM+cpkR5G8zQoyA05S48dekVA4IrlFcQPZwlYUxH9ZHCQmVpWZAIJ3Rh
dRf2aVftXA3VmWN18jv5MuBrq15kuzQ7lEQa5/Pmkb7UmJBjOAeBnWzMesojCuQ5
2yLjfWsh3jFOT4/sPV3Rt1NM0UASNZ2o3WJeYoKEFhvrqJhM4kN/fp44URDzV16p
yP/rt9aiy+0xoIg6DNZgEjJ7c6FBXqa5Z2t/jlnjU3uZSu7PJU2ncBJYko9zwWQ/
NTslKvXqc8TF+6KxyStUYF5Soq/7iGdYRAvoodun/sUsqmS5fAkj+LTPQjG0i0jK
nnikU5tQ4XMJDcfK3pEyt6zS8t2hls0IeEeYbYZ2ptHl/ZfCkehfsWvaZ3UCexzc
xVkNI15yzqJN4V1vbqp0QWeV3m+QGU4aIkBoV6WVR3+lnf4eHdXr8Ki/uU+lxXnc
bkbi04I2EtbuIZPuK/RdDzx1Li+ovLiJGc4WypniU3X45qJygwmkh/z6jnfzl+4a
HhSvvQTnmvyCvSfYPR3t+9Pj0ao5l7rmmSqXlx6zWibndYostvTBBIZQ01urb26C
qg5GQ7qxBtRt/PzcSDmCtRrTKYD7jCYBu2yxwRrzDR1Lw7/DY17TDx0Im78OwvGe
zWUbSBk5vIPkB/OvOD1CxLIZmqu4MprnChrL/BRAjBxwMdmHZwF1W+qMXJ3S0PI/
cXAxknEJfdXgvw8/0baGUz45e+zQ8p3SySubIqdxwhHqy9oQFTYi1EOnrbCWl/6w
gpF+1s5ohP1eZ87P0Ow0VsfZRBo8QA+ey8iUy4uilLiJuThNzHzUJL9Ixtr9dr5G
3bYwhn+85ydOfkih1ESjmwxP6ZZadv7NYsXS0EIQ+cy08efy8osrCFE0vRN72/rC
YY4Jw7ewzMjeBpXy4zwWo7grPiSeO7dljVcxxjttyLz6dzUIwAI2GXcd0asKuq9m
TkVnmeQ8SThUBfK69Mjx8dfK0mpNSQaUBHiOqyfI0J15tDIp/Oips3FASZqxFRlN
yKojqF6INzLxcJbmkIKAPyn+vUyq+uQ2TIvzvIRUbVbt+n8UJS1emiK/IKYHQln/
p6IaN6ViqSLs4OyYfadB19kEDuHttUv77I/5R2pmjGmxTmtnOZu1Cq+A+9j3V/eC
/L0e1EDhXm4O8vwebDY+ciXc8fGLzpSc4P4VUknrmjOGrZi/zqD/T3Cj68w2M8go
cpBiqASyXWjKK75axGkcXg4gdKBT4+t5NTT/RaY2ZR4lO/tJ8ao4FosnF0xFYnCr
RVSBVJk6M3gTRD7OHO5fDiFqKec8LcVzGJYSfFvnOz/5TY7F0s+A0q61KHbHo7oF
A92Lvcz0GSAaOMrOeWtSnFPklOr9NtN46LCb/HF0C+KnWBStXrPunFwlEvDeWpPK
JhdvEKTCyiCFFlOL42x0kpF7XkDZ4cWa26H1L8tBZYTNY/m0GYRBCkifKqSP/xke
azl1RrTp3cypK5cd1tkh7Enaq1ZtFRS0sWk6GQ3NKJuAMZ/Y9hGds9XMj+e3r/YO
G5D0v5rNNNeBgXLDdhxpt9pDb9NTVKOoNSzgLHISyv8f4yAvugQnFAocsUZo1VfH
TKzM4KAUedsKP+CgS4KcGjtDAMXQzDIj7drsuEXRhbZLB4FZQT6yitnL+4DTqpq0
fc6qXMqgWGaPUGr1JSO7uVfEJAFyxQpuYHaaVg+ydUK1WaemMdjVX61PhZbTepFy
i5Y5GpPZwSQQwldzRE3wzXf155RC3hui0uOfwp19TBdDtB6Tv5HhZ/eka7SMjGNO
KTmTPeoXK1BBoOX9SG5vk0gs//XPwW99ko6tyDYo9sCquJbzyLFk3nQHH8+TZ4fZ
Amuh76F0A3CHUciWb3oGgBj/l2Cht2YlzMw0euANb/PGz/dDeU2KMpOMTXjLFuWY
j2MsRM4RpqeaBd+wRs3dOzlWEHlasjmx33OpWmhkJ7IeL9LwNU7ANXGwBmiLVmBO
Ucic33MEGau3JvcQWxp5yrwXs1EYYN4ydN1uT+5r3XrdFPtspiNlJUvZNBcwxiPW
zMpPVuSm7sEYgisXi9U/6azvjC+dRoiwgELXtGCZY2biS9m2ciMYCFSMvmJRXu0v
B5AGsPM2vNVQyn4RCGp1HUIUwFugTNqGHug77BqN8Xi0KYO4eitCQmsnbJA9uh35
+3iUs64kgqNZfvUG3jhkD9PqOfzFaxo9f0NiZgMLYoI7pV+2tQZJj6y0iWmNGVJH
VK8VnrH9WBiKnxVqR5oH7AWZZYi6cxPWZ9rvzUMPkQar83FvC53HoTgpLAyTfGuA
E/1Rqa6AiuLAdav4Vbz2AgS90xnFvKSaD4gIpZB4sVH83PdzXeqZR4ZGJZHNzhRJ
bMFNnUyI5WqUCT7JvMv0mSk+yJoQMVlmpmB0YitrF62ytHlQwjmuLgrAi3WqYZjv
eZUDwNIV8PphbwpSZxNfl647T5bpFF2Qns/lb3IjInrDE/fViF2qtZDZUbCt2PtT
fJXEIk3TufZMtVZQDlwxTwVVMDz+wOEMup80pmrhje5S760fsX5S464udWXRPhdX
Lm9c+XD8E0+sljMscvvo6Dyylbs3rLrBhHooamxJKwDsTy3YEc3NAEvnYwwXFSe3
lH+bitn6p9PRyTgSzZZiFzYo1uDFORzu6SmNHk6Lujb26H3RfRT3ODNFb1xAsO1R
+OLL91aIQ9TXGjMiS2iwOtste5t5fDgI+9Mxj+IKv79cmH15LBZmUGQ+W4UAe9+O
4d7ClJ2jKwrLfidzkWCPuKpWuRflC4S/BXw2lAzE/FtkhwkV73YLInPTIKq+BmLR
sAXWG0HboJFc1mjmrXIDXKBjLKkW9rXKv1QJsCtxA5i7GZcXZpdEvZ5pbFl2nkLB
IE+jbnNRV9W18WHSt8jf4qi8Q8bhEylQ1KvlFFq0ZeLgrGk+gvqjNNWE7TRG4d1x
8AkwwCBacFNclwmu0oNsLDMSrQI//l2JcyLs84hYzmcxh3y+Kd9hbBKd2fQ21F7w
oGVJ4TMZWfhGKUpWg98qQH2EQYvHzb3JkPXIqXzgX+WPuznHxd2Odw6Qp+cXEX9G
R4xRM8MepQ2kKTYAAi+FX4HTZLaUKC/ywgi4QkI7pXAMEdY6vo4iYMGyUvEHVfCV
UNaQqJe33SWl2LC0sew9kxPg+dhggM+QwQZK9RkClFlLRixp/vZjQwP6vg/6Ylqf
Kv92QeTCheWQJCzMMBQIiRurWAZxxAlEUx8/OEJOjhWlBBSQ+zvutwLl79ymm+2u
Z3oG6Py7RnPuZpWIRKH79kPAYHeT040KiOfQSnFBpOHxcIaLxWEgsF4v0GQVJwso
z36PmfSKXCURWyzPUv02ZfH+/0virjw+mvS+ySOoTQD46bzAO+RCVTHwpUPpyba+
CesnjfgquVQWgZTIR+Boy7E1d/SWhpQG5J8HVHaubvFb2JSbZbAjZ7gxfzW7qRX2
wB/Oc0k8EyO3DiuLAg9Fq9sLOML4VICs6JUxmNK53W6P7A6zbT4f6alMU5N3Wb7j
slZc6AlmIXXASm5nMEyyMbUor0HzXNuzNDeKYRa64yn2/42pBi1WUSgkl0ZFizTh
qa+sJg/WnwtjZWRhZWFaWrqyUjbRFwLbTVOq3pYYbQbLV4veIRWzWj6d/ubTIezm
hyoe82yj+SNbeo6A37hfgscRFbjANBuzs0yUsncfIoQIHCEh3AbF8Mzzveas/1lg
dRVwXDTSa1En7ilCLUhgP4obWlH1uJCi//SQYLjq+RXVu9HzaWRkvOqvxzymzuFD
KYFnW+E1dSFo1eRYr7DdhJTq36oH+Doxe4KI1HFK8RKrE8GMPJ9Pzyjx6uuTSF+n
BSzVme4OzwcwS8rrRBBTY71tekbdPPS5Gty6EkZzA1rCB8+SW+uEKu3sbT4+HLL4
+aYEUQZzcBD5w9afWFDhja2qlwqKCtzdC1Z4zIzGL6ZGrNnIImGW9mKCugJIA4y+
bMBbTn6YpPfJHmjVZrz0ljMrYNYgGgdwICHvfRskhl+8bgoMR5DAFG8lIwYfmk8G
vEfIUIjA/D4ARrZVQO2IsIUpjZDW7pKJCPOyfQjkAkhU8hSO/5k37hkk4p274V04
qShaSfuCg1w5VUMgVPcwzFM8Emj5ykRoRoitmqTu5cdsdpUxU3CKTu9Ufzf46t4S
x/1BCQdJzxtP2P4/E515bbE26AyslaWte0RzDwwnxVpPF0qj4PXofwSeAwQs/YXx
oDPaXSVSxSGWsXGVUh5EDXM7BEZ/MEoAYyFJ2MLHzkDc/rcSsyd3bBoSU52a7iSB
wBabkJzPFM/PK+u4HKyWGlQXlqxH12KsVuMh7b2Lp7Kl0V5spy4wQujP2poXNDZ3
jjT2BBiIRM9WJvxrRd9RqrxcBFHhJp5hX1b/6UEVqTHQpOxLz5h0hYgNZQIMxTDz
refYwzA7BxabBr9cfPEZaG3QQR4/o3U+yVwqmoBZDf+AUdrTha/UBWWtdLr5CqAO
y2Cdf8skco6UczQkoFVm2PeoCBt0eFcJsyF9vrtoTBgdU35u9qSM7DK9BCgklC/x
XWwtlPlln3MwrtriocIvGFOHI0p5AC2IfCU32KEbHLhFa+vM+QgoG5++t+5WBck4
snZR5kvezNjx+GA/H4Mf896aeYBtSPJJAfluymMbjy1yIEGkCh6i6AHmFN+lQw7D
/htwsAo0j4uNKO350MkKyl+lLnVMvaM0OrYQ9ZKphy/B3vZ7NC92rX3bH10gDzwS
XUxegxAyG0+zDE2gWNW2nozhj0FUvXnAb1JOBRhfEczkCaS1SiyzIgnO2C6AgbRr
OErdVaQYHYIU9WNW4brosnnkuq2m9Ag24Bf8OJPJQCujOdjBSjFJ+4b46XpEINEZ
UBExNqvW3t19AnmRwaeKX779mJkhGmOGWl04CNmHsYIvyDTBc/PpsUFWFrSA1yCY
v9WgDw8zpDrBAWpoJjyc00hOp5rKzbvZmrUIUvtSu3T3dWGIsbZ1uQlS8fIptDAZ
qMnGZPt6yzH++Hd9UHLeaHlozAN8YFhRJeflF1LWl5sD8QIlzQFN9t3LCm92qBeZ
sogFc3TrIevDAv7z4ZXEHqh5MUg2fwboja+MiBuFwcsiuGbDqG3GzZJ0uJtDLNDB
dC8BkZIfjkFUFuOelwnibP4asAwt0ntAEZAfkHdN2gGtZhrLvsFCyoYG6vt6c9gd
skj15VjZ6ub13BhTXQQr6BKG4FPGBurGAxxqcubtUa2K30pOP88WaN3IHxqILpAd
EsfSb5yW1jQ9kb58AsSXomBGd9roF6Ik8tknewqUYrZI4ZKog98qstgG0mszOoEr
X6t5pw9mzWV2t0ZhxQIlKCLz1Vat0qO/4euBqduZlUDt28g00Lq5tIcLDO/b8yHQ
spdSnHAAmUvufZXxAIbXeXyudINwngphTCjr8Jbry3tIyswx3OY/HsobFbmw51mQ
eKRiMvuStGF+oGg8NQlc1UAxIbAS/xel1inTZ0E9p272TjzJSRl9iKERjqBSe5rM
juZIgK5zkoqnspGA6P0F78rt7reen09YxjjYutOiwvpUgTb8zvmfwbSut7+zIx3D
FcJF89RXmexM3AUL/J+h3kTKyyQxr/7IaNwcuasUBtyF3sYCNqK7ueQBNTos9Llm
XzIh7jw1ZQTJaybP5q+B+sRgHe8fnwAxcqQA1Y025gaoS3vglWEHTc8fPhu4qycf
m8ReN0YD6fiBDIiwKeBF5kgJ/gwMJOZ/BveEHr5K4yq22TNM29ci/+FUWlkiytsp
OwQfmnbu5ojdgMzSsTsoz8NrhSnFsz75k9y7JVeTFnbHKb6OBhYn96jtcidvmtue
Brx2Mgpak8AX5VFvVQ7nKtm4cNfbqXuLkNiN7qzlofQzMcvuUeaeHreHeVhc9oY0
uWjOTr+5mfrF/90p+RnnXDwi7Et/ALhe/eVUcnCjH3HZpp0e2K55LYx+tI0rmVFK
qW6rd8/L0v3xbosPYP1MwY6CCEgak+Dm5S0J/yBl8EjM6+kLo6kpxwM6P/N5xrPI
DDjU7yQNs34PIIlqtL4+APssU3mK+S2UUwbQ4CEpe01DKiXBOMXXniHtI1SXDnUD
YvnxzHscYyF8ydr++tGhLAC7vXyluH5ZwyEF7Z7KT+Mfrt4MvRxs8+SOnNw1B8vz
1d8RXC+Os5iyPkoxsr/MGVJxfyphA5S8YjnrtWlDbOa4Ju5ISdMXdEDF/fKv1W+E
zl5Kh4lz32h2Btn/sVN4RRIKFIgFnGdWCrWH+eGIiiYyQ/jlozYp/n5qgWDbESJx
XycivTOLvSIIF/n32FISd3o1tXtWCeb2VVXNjg0FZ0yMnhCMoO4SzsTXewMJfCj3
lOPk1+ugL68hAxeaBCOb8LVVFjpcf85MaS5LV8z9etmWMYaThmRFrtlET0DqJR+b
0Je7dS9SYQtgruMHjbOq3QDDayQV8/pJRiixCqyU8RzeF4c2iPOswC4AsTjwkZOn
o+8t5nTosfT006j7eTCQda+RlSgdLqgAtY3KisVgamE9UeVC+su6yhsQCKG5AZFM
IsajKyf7yd9oDfN138NM1o0BYEZxDkwKGh78AwMS0/cjWYL+JSmrl2PocwyRW0lr
xcDMY0hNz1gT2gLoUH0CoXuu6nTBvSgTcGrPoTZNSPJf2FC1u/ZkODzz/ePDjF1Q
RuNjLIplhpgdzPa6AIDIL/3nip65WYAjo0SqnT6hoISbjqdY1miXEhbMVJqHvtSu
FwPUIRwWPnGM4vD1rpC+CLBHJZ/fK4YROVlrk5vPUAj1pREpY+gwMPvO99g+OA6U
mbI6kcDWsYTWD4LBMY+wtAPWwxzLotHnsz8BicK1qdW2FIzFVH0wFDT3X4Rq/gaW
Vb6Poo/FWPabdt/LcJnWWrQZrM4o11QcVSO8J+UHDv55+wUcqxQFDpsKu84Ym5Mu
UYNGieTo3t1bLMjhdFxnfO7Iw3gAXv7OZihdHaDw4oMBTxaixzyJb8OgCr33YQnA
PIr/equYAqjvyzLuwdd9J26S5D4G9KtbSMHwFFW3AABsHMPB0izzD+neVpuaISlc
hXt+x2l2Zg07+z6CkrEQnkkmRiolzdF1H8pIarEsBdiONQkTuSOsorGkbG8/3tsn
Hy8Fo5rPrB2GQ8vyKyZswiWPB3t7wF+XyuTx20jD/4mz2kCaODymLfZyzZDTTcJD
HrpGR49geI2jrKwMkZhJRZ+Ik+fmJ7MauLusU5VjWTZCuP0eJ51ySYHNrBPIVx5O
Q1jQertWNqA4ArVmREhufjs9UcjlQfAutzdLtQh5qSoOsBf1fFutma9aVB01QG5O
ji1lsY/z63dqLHscZ72L6iyWCeiEp/WrfsmSgQIFHfcsYBIsQsTwPVMKzszLJyac
SiTnym685p2FNOX7d+OTCeKeSBTw5zRM3cW2OUkAJwN+7YSei2yHfvdDjsj1HAKw
pInUXWFd+cf+uxwClRNNnVw0ttwaPJdyDJTTYokodFKRMW7Cl5qg7qE6ALzqUHEd
5xM/9E0yhkx26ml75FzcyGT73c3xM7UjuliJvbZiRsalEuwQpH9BEqHjfmA9j6Jo
KdTkwJmvIumih4gLE1VbQtuQE6K2ayJiCz75gbWwVenYUtj3avEAWy9DtYGzuP19
GBIjZO2dX6j9ahSITZM319v6qF0Qy9DTm7KcHDU1ApwzQBd9Uw4y/TQJJUQ8u1b+
xSBScIEmDYohwwwydVXP4nxLzNxvYzQkgA27Wucuk+/XT8RnGdMyr2zuZ79dJ9mJ
IFXjvAqkcyOWk8h6WIwhhs/NLvoZtwiXCLftf1DJ6zjxZAr1kOFcMqFpwhzthyJj
4NqWdon+d5arPEBzV8SXQPzeLr+mzAUwBlKDONE4Kkm/4j21eistN/6PJ1l5+LzN
cIsVP04rzoUuwSe4tq50/2xYvWGY+zd9u0p72DejcAamEMyawT2hxCb1RhHUybwA
OREjRMaDRh+OxGDwPzV4iXiZl9pLCqFhlxnYb2DHTPZsZhDJ9YC9wWheanGYm+gi
rKFZn9PYhmH35cgYFTT1VTTehc/+p89uIT0lFYN2LOGZsXyOiG4LYXbwEzADh3T4
8+hOuk52gY+VaGGssKB5SLlbLpATVJ4Tv4w1UNsk5yMnoeIMxiivxCpaVM2Z5OGg
AISnltzdBtUFKdiqoWJVdTzrJkJkPHUBEyx4Bdhn2bUJZXNUYxcR+T6dF4sP84xI
ZJxu0lMi8gxMmVApVR/DblQhnRl7kY+LkDM1VrmGAKGzwaU8ZsDVW7ktCOxdXLaD
zXJltVmNCISoaHgJWnC3Wi5ySS0fF9zvVAgIl2qw88eBuEb8MfmLCYTqnALBbgKv
rOEU2mfOkGYpHzif9vg6Yrnv9IMmgjkoOUcgY7ie6nleQryVxZ4uIrN5iAA9L+Ri
ju0d9GmBrp/s2+NswvDI0QamYAPXO6/A6odPT9f68LFJdJ2HQK6zUOWxQRakv4kq
MxD2niV1KzAF16RMWlxTFj7XKJOfP3vA5VDiJ0YpjVnmkN6xnRq1yTaeZMraaY7n
TzgqYCXvzKCbJIFpBWLp4s8OAM8Brv4BujTCc9HVFtsqnXv6d5OXSPED8pHP8Wz8
i2/WdmujcZfibazRb3UtvhY9qXMO+RWEyL01FxCti2t6tpcT8RgYxpbiRY9J2AO6
tU3qZuNOFyP0Z6VJKjDAF/WNNUOHNJq6kfBmEzjSFwqiLa5CubDZJ799f4F8UBrF
uSX6Hmzegh7Ik6XtSUhNE8lpFNr1HUIE6/aZGzLNPvr2Sj0NTM7Qlpj/4+wqZk8/
Ok0REw/KBM9DNCKUaQLZL38ttooacdJqIbnR09sQyxKMOMgOoGdRI9uMHS8kI+S8
v4Yqda9ATurG5Rtk4mLVH5z8c6B2ku6PR1T/bIQKeTicotYlsgETyGPDC4tIUAx6
tgEn9kmJhB4GMhe7t9RnDpERvwde3XI2LKKkKgoXJzmM2op/lnRxipEi0fZgsOfb
5k5Cq6MudRtbmnRpL7Zf8eTlb80Bq+Jdo8yp4NgEADOiHsXa/CBOxnC9k5wfjz9L
JAcsXZBTdgua5STbrlm+AlP3ShWaJjPCv3b4CA85rfbjxvqZ0M1xKMw0ko2+pEjK
L0qgz5x3nuCMnB6Xxde5FqAB3q7+tFeuejKWWmQXn7y2+/bDh0Baw2N9n1cl+hen
y7rpv92nO3f6k9kc428sxeM078ENGeZDXctKNTQIWHPgIfiGhxY9ReLqlVzNz0pt
N3J/xMAsQpxsDA/gtLmvV6owTMje/f4UOzP36QS4EhThSYDtsjVX/2str6x6GluO
CLsEtdha0IfyZos7s1pndt6rzf6IOEkbsUe1MdPHnuY6XGv+X+mGc9n6DNXQDhYz
eVGk+Az0XDKL82oH2PJiD4epKY79SmFrasHatM+L0vHc5wRgSPiYmxHJ5gG427vp
TZnQDH6AQb1+UQNUkqh0UUCsJxODVn/mW5rdQlW0esZufaDfmZfzenwcqgRJVof+
MThqOGD7BOTWHJgF198nGCjgyyUbD3G6Bq14SO1S+y8Q+DtiDQgeIbLM16oy6Q2d
uh3g78qQMWB3N5tfM3T8XPnPh6gU61UVNI79inBHY+whVyZeJk/zSwgIaxc342r6
p5OPvQoKOYnIe1KgTC7Hh50tbSQbvMz2UpmHyXmxTyHVjCEdgB/GlXzNGiWzOh49
iunhUNsQ9cu+P6X76YQEx49dhKRcZmUsW6Ht9thz/oj/s6dyevcfrRZMrkRjTQ+q
Y464tK+HSdIEnBqKp2Vfi1vff0YUvZK5oqkmi8nq8cxVHirWT50ooDUoL45a7D7z
4rgYVnRMS2qccaw2STTwn1/nUIhhAtLWXx1oeXVV/e/AfBDev3+UEBf7HdU6fYMp
L4YrpsxWpMLhdpRdk9Hn2wbHbAQonrtdXuRNOmVLo0Z8tZaUHmvUZjVxFY0g592e
UnJnbH5Maa0Hhz7YWHj4NAffLZyjr2P2De0ab8EF1y5mT+GNNoPgkgzLejwjfKut
sszktB+k7d4EDfred85NpI7LHDVF3/avG/siAyDEIFvYv+8eZV4QWyq1sHk+mbhj
rpGMCsgwGKmsmxmaN0WLdB01IFIbA41JmPoqIIZMMZGVmwd3fnbe1mGeTIWNoDqY
u0M8JKtBaI5OS6skY8zEvKILUKaYL76mjDAKY1X9UriswQccarGfKl6w1+Mg3VQp
TJWkqLhnv2bgUhIAufqok6v3WzXvIh1z2soev8cjVrgfUhp1EPua5vmaR8GchHRg
OfJfkrzqUhKb3wy8tkbcjCtlUtpsaA6aena1oCycxy/NXlvIDkUeS/auYzGf5ttz
N7Qg/cS9TZjwqhdaNBP7hbo0ekrEelGkdik9OnnijP1c74xIZ+/zXclDZo2ZAQh0
o3LsSvL1b954KI2uaUqzLTjSr3Y4UG2UZILZOYA7Mt6WOJzMbOQwgmx8kI/Hi5e0
QpjwTINqTVhkllrYST95UxxpdykI6rrtnzQF2FhkiobC7orAwk0o+OUmE8A8I/Ug
IcGOLlfwL13hSIt+CdDnIaoi+Lncw1OlqybxEOU73blXQhkf0N7/4E/40/V7Txp4
ltK2B+y/HoVjCQL4kBCj+mvSFnEfPYms9+xaD8RAqMc3bIKPonjrhWUelwAf9Raz
mzC1WfvU6YpKHxIOiFcZnQR2mXFy8PSmJqX8tuzNtUMtwIHgR1sVBmkjeDeYoq3r
imZpK+NknDPsIiu3SavstWvZFG/QvkcKVzExYsFLb4S66JALIgL0H/lFjK231hoE
cGxwETvmB20Sa4kB63p08PEzxBqyP3EBYOiBIjhhNwr9y9ux0SVh6DsruW655dQA
hdAzd6J9TCW10W+hEwxks2g9bGffITNcu0SYmlVr89Br7vc5o6CLongqqfaFIE8i
6liiPUp6LXdhM9RmyvTd5PVgNi6oKCJXgLZLR2+UosF0vepG6FXomiBzPLHEuPL1
Q4F6PclnIYlcbyU5nna99ibNElBbSGwXUdwkemUp2K0CvXjfJmfsQd3/cKZRTkUi
sjJUVGPuzNDCzTEBRZt0YrNZmWtmjAbJs6KBmVuncyuet3jmUUnpLWif3sTpE9tS
FAFcvikHoWfKRlThA6kf8Ae7O1qD7xvRG/J1oUhKZzatLYe+p9hEZsd4BaWSGjf6
kei8qB03RINTpSuH5WHVt0SoUXMvk9o+6CFtgFAi7td5Nyf6OXZooQDEk719tKdM
raEwXajKDpTdOE2HrPfIRUTkFMM9ltOKBwA7VmBn12Uhk0jCdx4HdYZPGh5uIVbG
sP4dzgOlr9qlhheqCUpIDRSm5yjy8P+E6mqOVm7Z+eIV9dYBoWGoGsDR79CVd/G+
7qnyjocCHUfTN4SUYAhVweHwWBiC5OiTAyTWmNJmMTgj7ZLIREOpxcwG/ckgc0ek
D7vBGTR79ZVLM5wQ55oYrCBSbmW1Jx3L/L+1V/UyM796XsvmIlGWYBl6voIniBm/
ifm68Sp4pVbvcvKAkc+UtisFplIQob7SDh9WQIhLJoU1K0KbYKFdOKHYTnCHU+Rx
+KBrG13rg1sfK7B1wzFN4VScxQaHN3S07dKKyxEWgirgyhptjuUbm+MlDqNxJrxf
SOneNlgguRbJLSk72UiFv61hhbeHa3kqKyaVgBNR525xIW0yIqrK1O3mTxzVwQ8W
1MWrUhi3LXLXusW9/LXOrTYhXvt6QxazskAI3cYhL/zO9KQwn8krcat/Dt9vKH0W
kNhsq2nhtUiELtUNrJK6jvS9e7PvQNRfG6Wv4X5ZhUJQK1cb8p1qFcMIzge0rrfi
fb2RwBTwZmUdTilyhpJftUsYkcOfS8OUaYWkJJW99fHVFlhAvLPBP/FLzwfej9/1
rY96J7j+yjAbFUjDVK/aaEYcUqbrCSAm96aXMM+1OgXfOMOi+pXUO0vSF818Pw3R
Rm5g/WrhvvW5x2Es50PCgAVSiegVYSW8uWxPLBYtGOekG9cHe9UOfLPWgeHDub7R
3wimNKvBI2Ph2OOLFZN+T47U0VzNmW1tIbGkQRbu7gMiUjqPByMwWoJ3DRBnBR4p
cTDzs13K73xPfHLzY7NxaybwHK20wQLwxUzERwYpOYy0DBOsp6ejKRrmF1weh6jW
8YlAqc70A5PdCrIstZamfJ/WcO/+Xz93T+YInAc0wSx+5nFGyOmxwD5KfI72WDj0
Oj5iFDupC1VzFBVtrZgfW60EhStr05MutzBfLIOZ5pzvlVSgwFQAhdsURm9O8WBu
6b8RZGxtXmXWRUz4Xlyly5WL8BmGmkP16+pe+TWjFWe6OtLlB4JOkzKeVKCvsP5l
QGAjpE4xZvCWT9inQG9iLgSxyVQ+pX/XhZBe9M+URyDL8pnLg/L8a0/Yg++IKXAp
VVigsYcf0uDbCG44v9Io1a6c10CvsMW3lWKsxKyUPiK0/ojcszKRdyrcfHV9DNEJ
oPmDkOlgI/vDUlsD4FzUtKOXtkKPQRZNglj7jv7daLIMHj9dooIn63AnGL3aHbAH
31jYrusjcj6WWbOGVtlecysrU7WR51k1yU62SWXeGezY75RzJ4hunmAHZTVIJ69i
jH3xSFIj9HKb7jqawE7McoOitMEx5JBwgqTAJ+9tsej1F68uOiq+syeHVAj66H/k
fW1C6iHPmU1K+rb/ZHx3oFvmtP+iSBsZvre5FtolYOsSp5zC3BRUsEFhBt7Jvgql
qm6MiELrixrlx4bgrBNi3HOUVoNaF8+ntvm06t70M9PPtiTWlxWZzJaDJ4ebanRy
X4NL9fjsv9i2aV/FNHn0Na2zp3NLDWGOTNUwaU+sxh0vuU9PX07wSDLYTLcTgRpl
ODHloqy7B/stl4aaDKYkzR9TZuySY+pdXIgku00YfSHUaojO9NloNFEooizCDD9B
GhbXhkb5f5e012kbXb0oDkjC43eZnp2uxt6G6aP7Dxj+HoEvQkpj938t3owV+dVe
JBM78oe50yGfmwiKy+beQo+yqkmAghRYSQ2MP6JZeaznBoMS72USQM8TbrdClfiB
mTUjkDAIn9xYFf//DLPEyjr+jQHKIJKg79f8XkwpUqDZgDF7elWRVzVO83dZAm++
IrGGXfjHa7JRx2y8uwoadsq8xLGl2IUIGItga268xxzt4OoskAnS0UCUCm1cTbM2
W9sdWg6pKfiY4KsTRoI8S7UkExPcsuyacK67Whg3EtNHveeOXiBUQ0Ng3/rtJFvF
F44eqcS+agCySs9EVPyIMnYw5QV3JhAnt8XvqwBUucn4HOShV3SaDvLWYaSsnUPh
YsJnaqTEEVsRNvtDceQml9/qkzUULZAbt9gIHx1OOgdeS//8n8U+QXiza6inVdLG
wlPNKR5QFGJgIXdO+kg2C3smeT1oaPhhzjejEmc+d+dtAyfXDXH2t29UDzPN2ETx
2ARI7a+ZyyCwBTTV2XdVJdme1zpKAWAOhTEA9+yBRwD4cnZ7bhFgGnEDFHJyE9mH
BNqB1TrtObYNYrHjuiasOIwW63+Julqr4t4P9cOMRgirM9MXgz2cQ+2G2xqG0MIN
oZ8spcCeP8ESjAZ1x5MswNe8hC+QM/vLM3xtVVqD1cTUBt5CEIq3PKacBbDtZAiB
ckz9jcSwrU+FT0ZsjuDl2StfitHXqOGegd1ED1MW90AKxjubG+udpMYLeJNqVryZ
A3jzl+N92GmKHUE4uZHDpT8qYAbxLVGFV2m2leU2AlSU6Qm4Qi7sxzDn7BWAbtZb
uYsDXdG1oDRmK2zsRWPQ0t5IqCEPAFkxlym0+JWMK5WXv6N4kO0GNBzFkQQZAjTl
UbriHQWn/VhsbuadgKD0idWlUpoMP2DqjdKGNmZo2ctXqLOQ3zGLNXz7FKGdWSEh
WdDf4ChkpIcVlvzFcUDkN9ykTFKWQb2hQUMe82SJOGZ7Moj8tosnj9vajQXmpl9V
4VJa+Orq/jKZZAA+q2ZU22xOYYbiz9GIzgKhX0W0m2mhw1kE65QShhdZvF4Sb/ia
G3aqX5kv/A/vuq06wuFdg/nKM46C/SNqc+u42gFffjLu2X0VaSrHod0mh9kOvc+D
5JDF2g20ILb33ZUEVsSylmzbFPCbmoPvWMkZVESAVuiPbumEu8NywdCO9vwcOnPc
m1viy9i+UMgh3RhrCiQnpv91ykpHvM/GaSSySiUzNSKqJcL08Mmyi8KP48rnJyNP
lJ8Ns+JR9rv6agNw3t9T6A17a3dibkFBWDJhmuZA5tg+D7vNc5/HdH5/iziCUXb/
3FjzNipWwu64OjaGtN2rbNKVlU4f23QqVnigJYf9fevzOzjIODAOrkqGcwiZGq2T
1PZQY/ZDroxdsLlcxW0v21uaBNf1yAkCmJPGQuGWZgBTfskmL7zXXPWp0uuyOtRa
IYkoFhDvM/gl/4n/qqzVnmTwopWlYd+iEtlX1Oy7bwp19Upwv44KR5z0QAfRglKY
BaQnBVhqVG/sIk8cUFi22snc3cttKVYB3lgFH2vtJjtIpLwc37UBN6Bxu1ExZtO7
mVUCNRCp9wg9/D56JimAv/zp61IbaBqk5/KOd42m2xpvW78BOEs67sNjv2+bTY7P
uHM/5geHwQjVWw97jiNqCpfXggbBMhHPMW1UL2Le/xR/eDR0Sc4aUPyxHqZHJ/Fu
GyqOZfrFK0h97houKu5prQPyQkGrkPxH0g/SFlSw2aoYrvdJUaos7QMLny13aQuZ
40ilBNz1jYxZP5mxuGRhwUixnmGmNxDK5CpT5SjapEr3YcXGh78B0uF2L/Be2rWY
ilM6yGp9suhiFygzIlcjsvf3Ecy52tFM1YB3R7d1jF9oRUnSLNxoGjULnakcvyKP
ElPKU1OVIoRx7ibFt2cN9JgLGAu1sSlGwVYL/Todv6ZYYFcQIOEC+/B0429ttLNk
8fWJeDcEGG00xd3f+nCKQ70cmi/ZcoKl4X/9t73kOQsQw8/gNBM+XBzjXHDp93i9
eOGe7fVSNPW4lBjW2gg27WSKd8N2Doq5qvXZ2+BLNXYOe38DEO9MVvqCbSc4gsVg
dPnVJgutZnN5hotVN98/5fKyXaBH9q2pbLiyUTrMk4SsYVKEJxrPgIvkTw8OX6Sk
4EEa+W2ahn8QYDnHWKMuaqWHd5TQw5ape0nuNkfC72SgOaFgBOmne28b20DZQLim
m1KeIxJHqo9YQ830M9ZMbsBGUvbIxyhjg9WKPOmqZUnL21b+g3TePe3AC+hufTVc
a4P1INTmuwaVYGYC+hab4JzUu4KTWoozMJLCIUwwATnW6vjD8wD5jvAPCrRPz8QB
E5Tu7pkglgUKzPLk0XIRF5X5th8jHUf6xAkVzHC0va9BCiWBnOiIZGP29NsQ133a
vsrTgMhPFDAIZ32uO1zqtPEFVcVS58B+Zr8S04GIUKsxsHo8v3UtHq6bOMCJ55ik
9AGdJmncFGC/fkvyZcswJ/7HntXF3XwNNj6d4zvtDO9dw75GyzaHiUH/dLlTzC0f
soJHXngA5Dv3RjLxLcs3MawFGMH2j5CLAv8JJP4u0r8i5afa6vp89aGOa41QlPpi
TtmSEUlRCv1B8/ymYYaTFTKv9X5LHtANcLchev8lDEavOFAsFXqQRKM3TGvoZisT
LyHx73EaOoXQM0Kew63SSMqygCWDSmGYOwDnGimmiV1+8RlNzr0a402I5t+wz1nJ
OxUGUwq2ZkRdqIVFC7K/YmNoy0GC8Roh4j+hnNo8O4bkZsWsYbG8kcR2Jl4/smZg
x323PQGI0ngDdohKMp0d5sz9WjdZ1nKd94hpnnrSeUFHy259X2u3sQ0flCfQuVS0
Z0FNcfLwri4yDgNJGmh/TsaBDvdVAJIi5f464w091g0p8jeq1SvaH8XM6s5tSipl
sAzaG5khzl/doDcLBapIrX52aQ9+RYD9F6eCpkbIvussdIEKS4ELw2B61EwBXuTU
nKRmi8fHQTs0svlB42VOekeRye98gIVSJAnrbREs047t+GpthAVtfG9t7mJGdzQB
sOOaKzz0GbkBKIi/jNm5VYX1jQEydD18REUnESAwgVWBBtfqonzEuylySvwCyrIs
J7SP9SEGnbaTiyAGTf2oCRmZgYvBkeFR0wSopQxn2lii9W92IVewN4T/HLBKCsco
6H3bW1ZVLGJG5IJ4hBpBh4a4UpCHmEmGwhmszjBqEC4abz5FHVZ20Uew6NuBTPci
77SGU1yvzA1tPjsq/llvoCXXdCVL4vuSsWlKrA7Aw96dr7VML/OF6ZAxKZRZyr3a
nszpXlTX4jELDiqxfjmysKCz08H3fKvOQh+4Tunu2AAEgm9iLMILKZoMY1UoAw0m
tBlXtjnNOeZA8uwyUKp54li7k4tqEIJUBm+uDNaUtvUvoBiZeMicxmdAABTb+RXL
KIyJy39167w7eIuyidPpT9hJ07k9vOu/bHNe4jDIFYsokfnVc7uFJRh0dzxzrXw/
IqM26C/c6ENeC2m4tUnhZjHeaEpxpiuymu6gO7jyIGUu6j91vKmRYTOJV2yJUVNy
g7Bnh75tbDnIpHzhyudgqQFjVxQSmdKbdUo4RbFTJQiwMslfZMm9TNiBtu9t62DI
hSFRau7hF9JiVAaTdxfH4WGcN8fnJNs9geAY5cWFO+T6Jd/KnPpTucg0XAIJPtkU
HvZ5muNpvxo6nGNJCff68SDHwl1UkfYU7LNckSi73uhkin+j0MYO9sRo4etJiIw/
njF5oyTE5LLp4PVD4l+HnncmlYPf/MmoOXufVzjUHosewakJHcPjd2x/JexUL7WU
yZYcY7jqdSArrSDGRJlljY8KQshSpXgYWT6uen+SyYXcxZCZJNpMm1rUa/PgB02f
yNFaIUsOf24kvhctnQfFNmhe2vELVY8tlbCOF09Fn6o3dTLVvAGrV/ZjHooAfRJi
dPPoD0eB7Tm87dNaBpjfKaD83rDLilpFwOlumqAilZsnUv3gjhukS7rk8sNOj0v+
IofdHBRSaUlV3QRxzpQTNyKUk7jmcg3l0a+sEPMQhXO0fRN6JotZEb6jQWvDvMRJ
9Na1ObBRrYjhSI0FLs0k7eVsHwHOs7R+iSEHhhJFmB02s22BztCCBc3Svt6uD/8r
mT4wo/EozMvg9sbyPmNcjs8/KOL2UpjUtzj/N+RUMbyyuVMQXlZXvahPbdwtNud/
i+3m5dngkHP1sqpBQ0aZcdy/9FVN/6+AjVIyu9+MYPjbKEwaNSj859lsBk3hMygt
JQA6TZkh9iveRUpi5yectAiRld4dE9gq6bYADmoZs2Bb3M4r6vMACcgKhwZgKdmw
0DX6KSf/LPvO+nFpD2rap2cUgxGLy5KSgO7lvn8w6XwKPO3cfyhyXtx604D7knlK
6k6zgAh+AvxVClz4Fe5cZm72FCkhi9FaQ8wt2gttN2+RKbAbREnynFTbaRtGvmRS
F6DFlRtucr4tPlGiWQGKUDYHXZWKyTDUZccVg+J5cdTXjUn37D3PIbq6y3h4jVD7
wO4PaBlG4ytzGUhNohHDZvctQvA4MMFBDM16o0qgLAN7aeZX//j1KbC5iEzg1YAI
/kTxSlTpg3jWPjMWvpVFpf9eSFWhPssLznIC95OoHQ70l9o05UaCRwOLAJtnF2lv
J9DBqQPvuJIcejQQ/AepDCStQEu8RoTXSUeLfRX0MBTq3aKYQX2UhJM2cbmGN8w2
VRsxhS+20OGSr9jj51iHapHA0Vok4WKoxDfyE+pDcDfS1qZdefxu/BIRG+bG7ERd
Ln+ynRrIfaVykzZLwHQZZVwcgScMOusoC6wOU/aN3rUznavpwKW1IpPMXTzd7jRl
f9zjvj+Q2V1mKDAuS4CeM+ycdxBx2in5jt5nHIOl6k83lad4SMsM3wazV0WmxpAS
MhXv5hjrn7PIuitQFa7yXEG1tzGJPi2gOPwvlJ0+fnJlOWEiN62YqC/5bIemYvyo
VCTYIta7tygD/BuoSj3X1O89ZY/mdXkEsVrnYfBeaRU11f8OCrFr423oH5TBqBxl
UR+W+/VLjai4cG1m+GRBRwGqHbYhsTSzWNtCRE52Bgz4SzMaUAazbdRKW+1nsBTS
kYVDq56YoPQWC9an4+fQ6iPGvt9ssrbuIqiEGHhDUeJw7SaqA/xm3ZSzkmRiPQYQ
SnI5vbQ2NIHWHNlMhz8MMeG3V8WzGU/lifb/yPFO8hCPmmsr/DaGqXFdkeyTpa8M
jMJDKmp1EJzrPwWZjXxEW7SMMkMFFOw8zTVxEEwLwZrBmbZ/K5tzkmYSvENQJHf6
6Cy5CJDRb8wp3x41FjCxlqUgwNX/jZmmsA8tC46hBcXkLdvAue5o/wZIVUEPQ3ww
WvpHu6teCEAaT5ZOj77QOwyxnRsh03dcQD7gMJ4qSuVzDzuCAmH98YhakOHVe5N0
CjIjTW/G9xS1kFfV2dgYCTXu/+KAa4/rGR2rqP4F0nEqTuRzEHM7ZUFVYHVIHUi+
qdKxCBIknQBogKtM7GGV39hrkV09NREm2xFgVOi6vzMBknKlFP393tEnGbjOt1LB
EZ/GqA0F4Vyl+N7POwahcN7GoWw23KxfBV0p6x1dnOj05McCA69mQIYpwNEAZVUU
X5ZqbSb5CFe/0OXFlB3iSBYLT+OcLde8vQFm+gu5QGSrTcxKMEK+OL1n4PBqx8Vw
HaXWjwKO2Nv9AgVN5lJfQrkPptHZJix1/PxzPt9PamWywM67yIi8xXBshpumbyV7
O+rFu3EBqfzoG0nbkz1D02WL4CXSVzXtH2NBwzSFsyQwjoyArWMW1CB9cnZ/FLIC
659ETY3GOewX/eMz1i8sIHUAucxvDJjLhdMJNlVUzaympWBWFvxchoJTyyKKSnJX
WRX7FNDP1J0kbz91N+CEwOOPqDwtGEsXsgEdCNbFQ5gDJTCXdTmdUr4zzS6lwcAZ
mMOshqSLEz3pooA5Tfl1JozGfI9iz53BKhWEPPaviDm2lJgmFgw188UjFe80GoIu
PRJynC+EvxZHMm5U1a3cyt+HxBNzzQWisMt9hbvshJgkAZSUNfzsKe1wdQ938UUi
Y84ugiOvw4ZtDINDlocVKIjkWKxnDN67bbvgeLIeL3ZpSyJ0gR0Rkc0D/UH0RDzE
843M1oAUXxQlhfuBmG1wsVHW9JvLf+l0Su3t9UZ86f9nAQ3NzhqyGsgONPgs1h/g
OhCEBn0Mo5W1B7HXMgBLr+RhV1F6JZtsAkFuhUGPhz0MV/NCdKYJQY705jPdlD7k
f4nBikEEEn66jKaSldFOA/VDeT1MIooeBOlworPMDVzbWm2YCKM2QT7+foQ5us+C
LY/4HjmTC/AlVGk9JXL8pxdpSk75fFGIS9IR1WXSXyLxAioUdZG/S51i+8Kcb3Lr
dIxE+I3KiQ/9bPvKjTua2mmChyZ+E8SxBC1c+OXJoqUyIaziI3TbsGtWwgutt1EX
mjJi213dpSbdq4YGe+fZfG6U7+htmAfxeqEvTA2wJtih2ECtLsgR+rj2bq5O0eOh
K/oEMT+gUgGccW0owdOCmGvbPPj6vlsehmjPDomy8NoXOxqLdZTwDNvl74a/yScA
QLRU8D4pshfIw3dzBK/7qGsHTfl4/4HMHzyLlMEfDEtDIzTfDo8upGomOKNfMISe
lpRLkapAvxxBFQ96B3xoO/pd/+0nfFDAsrjcf7mNPH7VxwGYoS5WFGgFE3u1GIUa
z3feUScwJWPfNoRa7CJFgzl0CMsGlD+879PQLFNLgsWcs63VXMjtSSGlDYumcjXW
0j8c+MlnBxAcFub2gblTNnEyeQ/WeZb1TenBxUdlWzGV9mSajTrJvtcB3YqRbgas
3fefx+vMBbwOLWYaDEpAWimtRcNTMshqAL+Ccgfa4189mOJbhxdWD0famUvNXUzp
Y/xXKzG3K5AwrsQ2a3hGglTVj26CVX8j35KlUH4/mlawZVbO6KIC8DuFI/p6Af/A
PzZlNXi7y70oe8RKNykgrhk+hJhcnC23xavnkfVK8Ah4OI1gb8WrEIvvXXpXq9J1
6ffwIHPd/llfMlea0Rge1mZDcDc3eUeUajz0IiXUlunsCmc6fVJsyQnswxn0WJz2
UPvWs6DFhzQmbKtHgap25WmtMiz9cbo70Nii6juFPOH8t57GOZLimpe6XCmLGM1R
JKsjC1repjUgsbH5Bo98tMOI/Xu/xCurdK7AH85IgQ2uDXt0cchnxtxS7m5vhYKV
9BLrzU/ebsINWxNATYKAgSOMlR3jV20zMpKEpEtRXsZzYFWj+LOtF6mEr25ugdf+
yJbF8HuN2vkoG8w8WlzWiZK1tc5m6v89K66jZX9qKPiDodBaHdb4xOjXa6c89dl+
AoAPYkdHq3UcVCOjvBvhDtVK26gU/LBC5BfPEig2kGoIKAsHrQTMK6E1nZRAqKG0
vcLV8VckWAhXgXQCbyGWSqtCTtkUq7i8psopmjvP/7RDu5qPXw5B11JhjT3kJxuO
DYU7B5KOcX6aDByJlKyqhWGMt78XXrCBIp5vZ/eBjTzwaHGsDTeLlTh68GLJKJQG
OOanQOVzibaaZhUvBrNRAwKDyWcpPW4+LZMTEiIP9pz6xRJtr6awA30CtCf16PFO
qRyGb+8f52Q5M+mNvYzYUps5/aUJCQqk9cmlhIIUdi2kd+Nr7+Ati9oi0JMJ4U9C
HdvrvHvwfKnbap26OFR9oOZuniWFIBYJCekA+JsnAOIpjVsoIVEOXVqYHr3gH50j
E7vAx7hnMgtIZpubCHM58DDn5bZS3aD378Zn+nskrEPBbA6fZtdcDJeZZH9yO/q1
1KqcwLUO30NlXuk4dOJHdDRMIR9Cx+WB4c/S3LC8iGKwAqy3fEovLZfuVBU6I5JZ
ZYdR1VbT6DI47K4aOoV1IV/MNWtMgXbN/td4PGzenU8J2IEdppdFJSQJ6svBwSQv
MKDmY0Rxd8y4Y821V8lOqb+JxUxgpySBCa84jCXI0rb2poLp8Ae8LX+QfD0Xxq64
zV0HLNRZbyqpLO4PxznfHYYotxyjGw5WQDqEGXq0p3TkMcldKACtD+Wgr3q0Dm/S
W86HtGJqmFEcLIOd9246O8mD1hyWI3G/SFY0bgPDsSL2eOSBJq/mTfaQ0uU3saNk
4DalRqSOgeRjoDtrPtP4gXREag7/42RL9bK9PYqI47bVY+DEklvRfa/z8rYwmfwO
3Iju8xTBw+JmOoU6aX2f9E67UfFr87R/M4Yx2qSXprd17mZPw0CLnFXocgrfAt+i
Ajy6pO7si3+i9lRQ7nQt3XVv/5lRoKyj/4pqDQQwav5CWGiXZR36ahznqsg9fAqu
YFryy4c4D5AcX6FHLYChpqLtoK4ld56+hEYSFCYW8w++A5wcOKd8oTaJvgDX1b/0
dzrab6aRrL/rPZ9fgQeX5eJp5f16GH4So39tVAtanv82rXFXkF9YnLeEhl0uJt71
nIVu6rNRoVNQnsQZm3hCwdv2kJLyiVMGqly2CT8gAvOTdEngc9HJ8obB+dmLEsD8
fl4liM1y9eK1H1mWBEjlq5QWJriMstgz0gsnGaOwC7yzE78PMYIy14Kne0PEWQn/
Fu0mkRwsvFpo9zfSlhYKaAe+LoWcaUQHv9kAZ66JJy5Dr/a8KvQtdqgqpKN2IP+C
iGqGkIPVugx4MDQg5OGB5eSRE4ywDBUUygJ0ww0cTzzrgdfUO5bVF4gqSc5cBodX
v5M4MQAE+MfqJD6pBt1BcQxyZhUMTRJ09byXyO/nFPl2JonIjOcs6CNzrsRjC1/g
gNKk1RELLGW9rCQ6FKAZyE6DHf/8x92Ml+RsiDQCsa/WBom10RmT8rBChcYZcF4V
2Rzvm52EzAS1r/1DbdEMGgRCt3lJyrdLGyTu5bgGy3P/pRWYzEK4oxgUCTz5v7Db
5VD0clIll/QyWu4OWhg7HBeWI2CXRMpF2susG3c7dEAYHtSB8J8EiNON9NHmyivF
YFcKkHiQ853gL9jlkErHQAeDaqqZy3yLUT79pX5wTq+quZbfDpNmskb0Ae47HyFi
A7fwj/f5D1wkBRjrZ1UKjzVO+uRwJtGqk2XRdVaqMinMp+vgOSlpBzOagRGDXcdk
yH5w28CwA9B3gg2urQvs0yKNeLxA4NZcUebwL1DFtGW+S24taI792QAhBhrHwZ+T
yKxQJDfC1yKYJhTd1n5Tv3vktwrALeqFkRgIO4b3D1o6x4Z8epfrO87+QBFXSKMp
PPDPwIaxNcMl1cLsMjt3L20nGXge6CL6ERZnCmjTsOfWLu261FtcMvxmza5vIELB
mX1vQ+bMFB/LdYKdTLRJQnfrYgjgieJloRsYXqDzo8wIZjm7SodtUVfBxeZGIlVd
749yI9pyCaBCbrsP3mA78zmMCwlyzGmkl6U6H8vHsx5e3vNd7Zka2DOBxMoKfhpD
iiASMFAfuULbmVjyBcPsa2BMSivS7jbk8UUETZZ0XixFfcAXZqNSgi+6j15QM/WN
e2Nbn+yEdARqv/qp4i+fO9dxOQoQtxmZBMV/5Yu4E0DlSja9TbOn26HlKrO/WYHO
Pe9FS7tOSDuKVBHTggAvRlwkDW7Vd2FWXkL0CGYWPBk7thrvR5P9NWEvIWzSw8RT
l3OKjxBQ/Tcb38KcLISmOBCyqYjRukLzQPUFd3gVf593EOlopNMTj/0RcG+8FKZY
ZpLjBpP+VlxU6i4biygFL4yx15bQfm6C+QdSjll4dLd54pnTL0RKdIEpLVdcV4vu
3vro86HbI8XCl4oSbi7WfF/x6NzvnBTsF0aqWJQEvSCftB5UnIjg9a/A1lGyznvQ
KdKIo1Z5jnkhJ2k1NECQVMzeUB1oIPprSqAq/W+/Dv9q8lBW8YNiZhrmdxbHFtir
MdGqKkMQIlERmN+Gk8Q/pSYkwvrTz0xijSslYpqMrHm6XRBvwCvPQWhS3EB+T3NQ
ZQHOTtu1LFgT7EbnFs7uC//edDRrQWqUIc3gHbBHkQBAVxQ2CFkiVT9hi7lu9UJI
hOZA2gGwl7h1lp+vsX8lWRoCEBW/Kaf3lw5yn5+uLBfrQYRtKixb6UZsAXbiJWoS
QM0zlRKKTHj79nFRawkYKhoPV1OAbUmu4DFTRhlPWMmJED4xJVRCrElQTosvT+zk
lSlOgXIVJsIqEg71Bm9HB5PTJEW+x7nq12e4eL19VZcEzcxrcwPljz3cQzs6HVd8
5yT7ZMbxWIN+A/Dz2//qgREKSq3Sx5RydILjckZcScXJzKzM087DpxbEM3oguhFZ
1YAiAKDL97hAAdHbp+nqfNEPRjGIUCn1QAtkzrebd8B3eSvq0wsWqK0M+VjFMHag
Z2pplE3nSfBC7rQ0ivWqHbSjUDQ52VJQ4TsymIYLUtFWHO8pELEv5+Qp6n3TfHzi
fSZVK+wIMtnl+sovkFhsrLPejq0QENCKVknat69Lsrn19ieoPJ+pEvStaHyLuGoE
7j1eNzJwEYnIDXh0pGuovGaHDPcdLuPo4vxGLAb7AQjXKxyOBiY3zfpaC1FkSVSA
OK4ENYVtTAbGVaY/yU5yqke7xOCkita7K+4UPzsEYxapoa3jThhWwdic3MnOtD9j
jmjqwHgkZpo61Ht5682lwr2jqEVldCN7UXUGA/CmQPOfn7vqGGUQ9L4q7Y5d1Osg
ELlNJumtmF5QN1spy24v87LZ7yskgLXQQYudhi/r+wxTWsGETf4eJ5Ke6AjwkDXi
hvZJCMz1I3hv9a0wlsuL2bD5229byGGg9cy0BMg+4MEoPVWOBKFY2x9bK6em01Bu
9+f2+Y/qUIEB1Qebci8e/3WEriiFhBS+2Z0UsXLO8sT7r4CcB2gG2m1GQvdLP9cO
69iKGEQZaMJFPfeB0I1x/xbkKnb0sCqZh83kRgqy/E1PjEVCxL4W940AMk5RaOae
U//ysslzi6daX3gSrQ0pLY6rLFp+A5127ndo/yE6/mlSHctrooLiXwN71gfdcnRZ
bsG+nSbAbZyDvnb73wAWUUVOvde7zSIV05Dk7R7erIPbHw3t79htOt/eCWPIwSit
Ki0KlKQON38CSvzz6ZWFfaCDBqMmPUJ3mWJVfX3Awas3VElXMcbD4weDJKs0dn1V
Tu3JPimaYznOzumUndXeaiHE2zjpWHDE/1HKTpRaUqCc83AlYPyWnRkbw4B65Uin
aBYuhHGpNGOycDyTg3Jz1uCsvmXBp191P9CCW8u4+H3/S5yGMJlzVKd6rfYX/Nba
GAN8EgCOPx4FcYKJdc8gMB5VTv1/AgbSddZny/Pp3eQ/VK3sjSfVP2Tv0gQf4sPN
9DO7My8tafhuQsO0hyzkg8lYNaGs5KkgUt3TC4Iw1L2pLxvXYl2llRrFOks1QcHZ
k0B7O1bus7e7+MIg6lQw6sn71fYns8pZ8GLOiPC43OJ4pBMGLJIMjrkQ6AFc+t4g
7jbDwP17FDIz8z19nW1SdNt5aJrJocY2NoEAY2iEWq8FeMacFdLftWGbachQn1jY
RjicVxcUo2sxQ4jiXKXQE/VmNoqpGtswyPI+Wfkf5anARHKnMkemsJPejyV0mFle
5LTNQ9XELKoyBxrYhd8C9c/LODL1mmLGhGbu1NfRYOiyjKNpBtnJLsi9mNjQL9yE
NA/5jh+3NIHjqgggpO4wSZyH2te0CQq/2hfqsRve84SBOxkNg82pKzjxCAsVkfy0
JOr2JTsJ5PI1ggW9Gv9P1idx6ZVmUXn8DD0fzaefLPMcR2XuZ1UMJNMm7BSgJs1D
ZwO65SiWvEGNEUevs88bp8fWWuc6DQ0xx3muoYKDi6WeUT9D8g14tg+6DY5yi95a
1VYj8l5ontAuINZlJQblhlR9lcCn+YsZng83zZPrb9XLWbPtqnhsbrQaOUuytqz1
LL3/q1cU6hoB/21qgg8e4lAALq9QlNztlOrLU851OrSVgE6jdzJaNhbS4EnPvsvo
qfIu3Q3tiBTFqNmkBZn68qeqNZDzCKy9bjArbUyQxo1uVcmsfkUuZL9ihioNGe4o
iPiYOsodUsh0wUZqNM7wN2eUiJTYTzmM5WoJYVphhN+GA2g9mOHHJalePFff8t31
qxhoVzdYIgMVPLv9OCbwJa8+EkFF3tqoGhWxMsiLyvy8Oii9U+JbSO/0vNOCoWMm
1A0cdkqJW5uDaFDVX7Ve/svUoTQlh8kBRj9u8v7Ky8mcbleK8jhRMi83rCpMdPyO
IbgRLWsDRNHDW2iLAY4vpLy9ip1r0DB7utx0YJKcAaKoYlaCQB7Df8mBi7P0J0EM
G7M1qnfBNWCDoX4FovfUvyysyMlg7WJCzaFrh2u6fIuMdLAGVVE3r3Z9N534hcH/
+iMWzgI5Or9NFlMrviDzGxTTxm+GUkw5lzyK6Gk672W8+SSFYVntCwXr1WArHoH/
kYMlzTtMr8QvEKt87aHgLbxaRyDIJGiGJzQqJ5oM3JzuhyuxpZRnBcf+woZzscLC
ermMaCWEclf8NqpH6SX8fB7Se4QoaRVLwX8h10CyvkvvQ/y8Yd6j6uNJUBQg91C/
ZL4GbbI3rmLJfxJ/trqNCWRPpP0j6leWNrFgDyXc+qDc4o5/svR/oby4Ij8djgw8
trkFxYmikE8KYhHYTcNx5of+ZX9jEBCs1o+1LhG7I0nWRg91gGU/lRrI27X6YbeS
78Ke5WJVkI6xJuu/7iFfwSVSLrUfdfnf19c1eO6uAn27Yeuiv8bET5NtOv3uhZTb
ZgD3wpxr1pPccXdEFHtP7QpsTNSlD/mXT2/Dd3jBiSAt/Q5+g5s9J9Lwf1ZVhpBb
KQl8Yo8Kwxm+Vu4+RMbbnHqEgExsA5BkMTHC/iPvLnLIoCzSzByFOkZqaD4De9x9
YGMLJCzGDj1BUcNXomMLM7x0ddFbcZ0YJxwpVrsLUtg9wCSVEoxGhoxOCiLNMJdE
R1zCDITndm1JYnm1XhH2Wqpur2ClEeKigda8IBnusKI1bCNnWHfVG1r7uwdS6hc1
SgRfJOeHj6uAPXfeU6iDWTmnY93vi2nyMKhATaBY9lqcMkldgze6qVfHfM56beT7
+MmK9GO0+oGumXZYLn0iaXohDMu7eISybufSaIpr3y+i435f/r4fb4lR/gkzzX7C
6I+RQ/ocVIn0jEx/FMiHCsJhN3CrqYFfvGRtPuv1y6wNvihPshUy33bLjQMx6gtW
6swr9yPFiY8yBETxtmKmbuIewacE9TnRFTs0MOGiHNaLg8MoMp+V3XPOCTGBBY1x
vHGCcaOhuehrq12vtjho9b7OUxJl4dErL93YnM0PD51opnyZZKKFCC6FY/uQaRCb
WQZ+smNAaMxxX8V2ZDg8nVzWA4jZ4llC+Y2d7MY+RiBhMRLgK1JXIHeOvv2dExfk
QpPdnaMXqTMjfR6ruCN4aRekG0kPG7Y2Ho6QhmXcVmXWTKdZSIMENMtuAp5TQuAT
WXbl39IepBsjT2W4LG34Obn5n0PG8AZDayWOzBbAn6My86OBZP0HrUh9G+wd3MV4
wMOW92/d7eYT/GLttt7jKzo7sbSXPqFGNPND6tbuexzlGabu7gU95ua4/cLx7Scd
Jvta8xam60HyrM3/gRI51E7znypM4Y+LcRg21YJPIs/hVtk965PCA8YyRBnILi5k
1rEiiBdAZLIKUGCx5cS10RcKewFuOvWzClM6vhfje6nfzOWhVJl4hxCkdMZRhvu4
OduqPD/RinQvaAVabjwrxiP6Wl3oCoDZoUtGLnbQLkqfoHc2BkwoAZkcZW6amjd2
vedOVngyXLbz1KkgPXq9uyj8e9TldKM4a+tLEG3Cy3ZE5Y0L+Ag1P1YwmkiRPAfY
vg6IR/yNB6PYwZ/qSvmVajloPHaaKKAim6oGI0zJvWkZnazjnmmIjwly8nI31FAP
YrXDvyFSJw/O7yMwQqXkG+F4iY2ZHGJJ19QK12rr6SznjSm/5iWDLUJwndG5JNV9
8USPrd8Ey3/OHiPQgK63p/rV7hmL+eXOVgy8tpFlE85b87o40env8w8tQheIWy58
ELa25TM+MfBDLvTSDqbh1+oouCx2lWuzy3U6fZJ5Z/YrQw7WMwlamfD2NyHT5yQx
zpT5CvttXGp7GTZAVnR45vEysnUhNvHdN+//cqGLoTSuCsnXZQck+oqbqFT8qFZw
FGarBW8R7MOjUqMCYqgTWFoyKsOvIB32Qn2vB8ELjf1aRaSALnnGAbg+r8lZxT6P
GSdB98w+Fyz5bh5hbwY1ABrAodvoQMWoisPJ4P33B+fuSx967XZ1c8HWFwB5l20V
0ww8l+D11Qmel4qVDQRabVMwvEX1yKf83pib1xcRBVXqnmcNRcKs7yWw+yECv0LV
QekhwlZ7M+WkGh2AJ0AauQkd7uq1pZ330O4P1F9+/oAdF4ZGJUveV1LO38Zfg3Z0
i+jI52Oerg5itc2DVYvHv2F/eXs35GSG+/sNCZtXsQQjM8HbDASBTGkpwNPSn7VS
DXpvev5QG0Da4VJ7h/DWBZ/pujFnIt6tEQL8uqcrcAvkhe3sMEOEAyubSEfItiyH
Io5B+teTXKc7iMSqVtBzJUa84pHZjogR8HuXbidkTcay5vtmlzm4/JGm8ejPLANp
a9pUnV1us1ej0X2uPLTs0iugmknCsWmaSp413A4JgsnXmRvIPpjDceYndpI7gSGj
hCu3ABeBIaVTDVY2JCUqQqmBsl0V1653RswBmEmLcBKiM0UpP4OoguZnWt42ixiU
op0YbX2m7EEIn31jXq2YKa72Xj4mN4JaSuB4sJfnCIWZ++STb3E4GKeabGQQxFxI
oeTC3QIMc4kvin0+hhHoGauFLUPS/+hFyANWvVDh+SH5YgxRFyVeFdgvauSQw3oU
2hrD3s/5Ts3+geGpKW3vfvGScmFKpsGlK/I2zpEWJ/Yj51buLII+D6x1IOr0OpU1
iL2PIRWsjS3Hd20HELYdTvN6hR6g0DklhH/mPyNA3r0v4pOSKCsEcsHEKIfcjLB5
sTAraCvvfMSgxCfbLGtPeE8rqAVuo/43pdH9QV3kq56ih3q/enhMb9t25StxHT/u
43o2lCDWjxSr75UFoUvHZ6UYmz9sksGGABEJ/rxxr6k2DKf9rhxAIkZXuOWGsWW9
jtAff3L2KWgAUk5b89i35fv/BTx0kYq7CVyozzY2QdoWUN8E9HOsvAr+pHsenC4t
4TtCvAwXTHduxqxwpMVzSFl5kvVp79EJyscrKrGEms+bil0L2DHIpu+Yse5av/zI
GxieyvaDYgJgt838j9/NeCToPmR5gABdjjEDdPI3GyDkK9DW2/U9I5MW2bHJ7/D0
xkC2ZW9sO1GdDyNj2PD9Hsr37qS/8XfIhw/O35VR3nlSimlToW2aH4D++ULWqZzp
9r5tmSMZ0/MBcqt4DQMKC8Oz+AhKh7Lx30QOhzJO1qB7xMC0ud2xLlLO1ClPloWv
fjFhLzBNseo3iofZs8mf/L6O0rKu6fyGeFnlYqP3398WVVyX3J/axvBe7Q+ZDq8F
pwND5zWAnfOtxaeUx1d4fnRmpOVtfrL1vqGpui+zySqF53Fk+uNcLmwMwh84wlkO
v+ZyjI92EVxc+w0K6p3U0EL1F+omXDrKw4q8ci9W939PNLK1SFsu8k8332yV9cf4
9dBJcFauVbitpr5HPlWUaM61c/fJzoo3FCBJBNXjEk8YF/h6/iCGeMgi9kqlF4YW
mR/FMNQrRmYUwynacNUOO9fiWzrze3bIsjbZuGIjrThXF8iZ6G1zdL8hdylcK1AJ
unK5kIXAenApIyOIR8pbcwqZxFGJKcQEpjXcsyrzidL4xpkzxyj0QU8WlhupYHsN
0kk5r98T5F2XX4V5ZUL+aMno9ttyEDpqoCvHL77z8WyzhoE9Ko4TqiqKtBeg/pNh
oTbAc0Jj4aUUgPgcdSAycPLRcwb0rJr41UYMIPH22jJqFZfAbibR1WR26nw3uDi/
L0epJiplldGuUxwB2QXO6odWuh+TtxbqlRNdB5t/EPQxT03ceH2ZDr5C26l6jgL0
jbCLQ0lfFlbMmQwtTw6OLRDRSRnWbODIUmLgL6KpEvubCa3ix5mN0RTR/Jjwk5O6
HE2GWKOanlJVgbHs8ixcbC1nzuBdr2hQOwGELsyBc5B6LnkwZ14+7NUDpN0E1PsQ
htoOs6V0XMcTMIdcHF/UqEIc5nLt/59Dl0wt+zzgNx0Pxbb470L1gI3eosp3zmD9
SOB5kVc1FVa5J/ywEnAssWaM15yHIfN1HvJFGcTyxY3cTrbRF2oTZNQ8fA+wQfka
cVWOJN2MfuxKPdXqDj7lhUNKl4uprKQv3hAErP+jgfuVPQIPup0QoGgh2L6ARlTx
Q/WyDDrDBO2EDSPg2V2kWHO1NamnmrJM9VJWiOV5k7rKrvanxzCFcw+2ODNyY7aI
2HlrQxrH+3F0x7uyuRYRiVjb/s8YNYbkR2UQgTp5cqpLOH1cOhrK/QFN0iyGlBZb
tNr+qZriRKrypR8B6PaeLU0Smk2ZWsEBrmHPJASG5xxPlgUS+tc9vXrGbwmafB7z
f1AC7srnf4ApMHWWgLUr9D2tLLOJhxgCizSiAVNOdef07lbF9aaR6IgoS9LzqrGZ
cKS7aFctH1Pupu0Ac2fBko5RWdrfDjvVMygfzlTQIGBn3xWg3KtHHtrrJKTHZ0Qy
EKwekEzvrBWduaebaT4Nr3106MLvdmHfFmU49SnmTKiYM6ewhouojJ1mdk0oagdN
eKpOwtUovaH+22rMh4Wl8QepP81ACCGKUyxP5gEDgRPRuvIPUmQIxaayK6+rxqxu
afK5Uau6dbrByLtbtsjIBsdplCjCT0nfcH089Dstz2IcKySAniX8DHxpAAVe37C1
Gex0uFibk6v2gnAkQ445cbSwl2sbCgVt7nWKX/JJKSO3nmH9OxRbNA2Jc6TmknIg
/BFuhQIbm11YjefXWV80alBScjDVXa2BrFR2Z1azbW2KOWxhIIzcl7qGr4grGLD1
qqht3WnJKig+j/mts+uDndqui/RH4v4FzBOKXqu3Y1pD7KzOLMD8akM/MaRfH7IY
Apzw4VApEI7Xkb0AE3BrSX4gbeC3QtWcBh/OM0cxP9UZsxdlXTSMzxTW0HpFKTxn
mUNZTDRE+6frmMBDX8Brx/fhmTKyD1YkenyspBT8jgTFKDFOaprByUJIZMdWIivc
QzHcHJVQ3ZW5FvE+kOCUerRTzic9GNzRF2YQvZSk3mN2fK9ack3KtFdh1gAI+yXh
EfeqoaU9BCkj1hn4LTAs7cywuIcv45vtXAooBToMBPMz87d8oHMnqtI8hoPB96lH
0wIfSr006kX/2qgF2iAx4zxT8PXWuocdJKRiJmH1p0/nt6+2PSQOPAFLS9uBZXS4
CIpbvgsyL5NpG1dws6EFfUc9vTENMm41MXNhUnld8We7yJVDjuayl0kHtptFM9WK
oYX61h/UZkbAR+xwGv/3tTw+hM+SiUG2kWiWe6Y3Ffx4pz60xUReNhbH3N7KIv63
ht5cZDeyFPcFIOMslzxpmXz6qPIHLlvJk5QQlJQmIHOXwC2WbxhO1qNldwM9K72i
fqPgww2w+OxpTbDMj67ihSqns2q7tsQ/DKrAghkRotOXQMGk4zI8jvn+fU0R45+b
yYaKsYGFE82qbSXUVotU0GMiUQnDChlk+MmgPb34s46hntWQeNLMeE0bHpI2sYCo
uPPdGWm2Ap/BERHfa1sIGM9zXgFvAzoMs6l812rqPnbpUtU8xfiov+Azep1lTbAA
U1epYMl1h0nFA1JGr4q0p2lt2fL+w0TNBZnFoKqaKvc6p6Kkt5l1/Us+eK8Byxd+
AqzCwThXm/9IRQiq5PZ9H3+L4oaumd6HqixoOwQMws5G5rxBUeYHfeSNnaZhZ3WJ
jvUedgynQq3jgxBzvKqYEYBjd53NnUcw4tYE0va5xQ1wVGu+HnNXFgqTqM1Qlbw/
MRXZYQ02WxIruO18HRCs0dnvLR7riuA/8Ye1Q4iD+OWUs3KotbzFe0MWi3r5taZs
h1pleurxyGgtHBPjtPbVJwoxjFNzTTpUOx67EpSiuK6r4obFOhqMyvhi/fIab0kf
o0UQZubKKvNOrTs0ZIVjSJ6DS7srXjxgyMUjy1jBxcln/GPigeArfQhZPGceoMdL
RrXxax2LuJGymNqbvxlRCWttmvNcLL14l1ylZNDKKFAzWyJBqouct2UwS5u1sMMI
9H8eRMT/5RjBF8KzC310o/LC5BtELGQpCEAyB4M27v45UYVgudb1m6LxGGANQT1U
+OQgQYvOKuJKS85APSFT2EtMJnXSDQLTEWo0QXH32JP8RCfPw29LajZJyfs5KPOO
5KsIxvxo93sSTMlp2HRSRwCFHfU63G7GDrIquNSbiVxdJEbGPSz9VtgQF1PiRf0j
iLLrDarkeu1BzNqKN0g232xDQRFr9+IPcmb7dkf9CVssGunB7a32m0oil5DYPGjy
oWNMhyf0RPu4tKd5bmJg4Z6yb3UikUJH7E0cSOs5VCDk8wNlj1aYKClBFQp0wTXr
uOh80CwAbhg932Hpk7f8OqwsaMQoCeVmZ4gB3/mFcbcvHgtIu0fhwyk8YxsyZTx/
6IlInMkybXnkfEi5V3ZdAvBSJY2FPmL2ogJKjx2TmApZR6/fpiR4SWqErgTvYOrf
0oDyrXCPCDZRt11vbqBt5o9ep7fabkOSR5a6Jha5lNIQw8sdA76XlsKppOpIxkeQ
mn26AlKQ6mRTvxsaKpcfxrJb28oJmN8YHauviZ1ngYYKSaqxvYNwEDoQF0gSymrA
jMoai2GPexLwFZKQ5dEBlNsVUORvSFy7HVnFtRtc/4hTFSPHz8ACM4rIVB0arJc2
KLMidXSigMpkfUK6fporPDf0RRx3sW5Bx823X49758zr8K6/zSlW+L0QBQCyKK8H
Rd/fz9si24XlfuYbcJByHl1HmUyO6BAJVaoAybnJzAzECnlTahUozGDQGmKomCGb
IInbVpfw8A4Y3Gsiujy8adum83EuuMzWcLzrgon3JAU62BHxhDQoc1V7wlKMNAMZ
Wh/ObEAZJTyiMvwp5WzHk2Fn0vWIkouqhn5b/PRmWoiUhCTf/0P1K57ucFoXlEJa
Y7qNs0p96BUN5j3ZnG59utOlzvPoM9pJgeSgkD7K5WDgoiRH5sVPEXxczZXFPn2u
AWKgyNAd1iuKwXXjKp+wmar4xyFj9I/aaVoQkMczsQDwJVmDWbIRwnmx0aYdMUqf
VVoOBzKdh/tc9nBNFQFlTKxvmIskqL6dpU5hioBErCL7NaI0H3gfTabNfKMmxX0D
1iposv3r65W7TsQIVsrsA2q0jutDVgL9Yk26mTeescVE+m7Kk5/XSu+nQCLGhxgj
or0scWYb2b9D09lCNrjUpIwu4nkNdpMY6Gpnu7ZhOjvaKrUf745gnobJU9F9bMI1
6+vusEYbHOYAANjTyPHnl3vTvEejaR3wuPofeo762OYwIBxONpDAvOxvVuVoIyqV
l4d1+bhyeggRaeLS3tenv9LZD00GgTGdWhLCsZdp/s6+yn+w+82uH+cuP/RU3Hyf
ppiINr1J+O6pixxxdoIe1t2P9VDeICIPFgJgetclCV2KBXOUcw+TH1TRZ7na1PLQ
QozRib97ZYwnV6x7AsvgoS34O81+DFoMUtOD2+NIM5tnZaMK1MiNHd/6fl2VJszN
ugQWstcPXHVA1DSe/K7lDOir46MAf/RTq4IudcswXqZfTS9dEzcHA5e2KBf5oTFB
MI4VRXc0iw2nYvFwsd/Vm8lvlfWkK4YCQp5vfgh7EU+nO6Xb44EOhr9v1cNZKQuq
oPz0xTL5SKebs+ZQH9tuzT6OGX+49WSnMkLr3FxcgE0LY/8Ew9fW+IBL3kf5SG05
kRTSQuRVM9obfz7mR7Fdb59XMe6YSQC436Dvkq6cw8tsw9Mq0YoQfqKIb/1U9z4Z
XeR9p6WZSWs7z1JGlqtov8bdqq0j8TzFaItMw8TppT/KDmPhFuDpvfkBz3NnVMYm
jY4kuPY2C8haZzFU6GDvT8ynE7C+v+lXmmE5lM61UMRA6k0a9BuZlM1Ws+XtcGJd
WGhcqfbA5D2k5D6A0aV91xrv/t5KKa32BDkdry7p0DaIRUoo4lrQ3OCeU1NQh6MD
wgbkBpWwzTFphVPWjOZBMC8h64wGd1mCRXQpWhVYpgvxd86PRFLDti8owbXL7PAO
R+eLS3cEcztlisNHP48J8cY+hhLxe4E6acgOHDgDLaqEkpL9YX5IqvRZmcaKrSZ9
CF8LWLV3t+mDMpY8sKfrJv8VZrgWJt/5p5M/hdQdUMvtD+NeoMEVXDLUsoGw+wZ/
Tg2HA+DbjUu8/hfBCxxq1fEMmyUK42W4qYlCgt4tCUEFKs9vDLg/LsbM9mYTqNls
UmQK8btpodZ/To+ikvjOIHFXwuiIcFhJM0H3cc5gz5IyqvfIbSKJV08a2EGwtxaO
LsYEEQwDy+IHyMe++0gUH8Z06BGRaWQN+2dGYQ0BgxgUNp4JxexqG4RGVtUGQISK
RjMKW5hrmXq1XOOHbm7OseQ97Iu2R0TLTt+U+Jbxw+N8IHMcKSvbXxpdTFpY4ifh
Ct/l9AaeLoRGp1LKPxwDhTOo04iZoWrZpcW7A3dVdktdQXIwGVKWJ2x+n99HVXaM
ajZFbLyXUsP10qEt33Whqt/OX3NIRrMcP4Cr7+rCHb6g7Y7m7VFDK5/OhRp3hbYU
XpiKB0l2IWI5x7wN4mip0fJELW+4qMsufWOzQRsZeGv+xKuH/UzzQMqHxrOE8iFn
Ry25/r7ED7dftSo15gNXLYWtYXBN/aueD43fHbPuetDLpiZ4JWzD+A44Nj8GTgIJ
jPFNWGIBx1lc3Pfnd1OA0dSU6NlnmFi70A18+G5M9WdOvbV4AlPeheNbYfiSVPQ0
1RTA9I6QTfkWppv9D3AtflfOCvOu/kZ1fAdwKiuGmVpSZPaSm9WoQdTfXkyqGZzt
bNOE/vL+rmIlU5FtjmtYPfjm54e7+SJmdf9RqLVXO7i2JJGg32jxm512vAg4R3W1
cwSpfbzpa2lG5AvsIHQbVZr9i+UpNuZ+ndagd+Y3UYZKlwy0cVI6Vh/jY9RAHixF
WgxBKcj8TsVODP3oDzD2RbGBt7xaZgL5nUlWSYWlgz90rNfcYcSLGYN+WTppci5c
IdOe+Lvz9FDpdUyd3at5ujvWGIbCBvdAroO1pFMIFJXfXa5njIUEGfVe4hfev5LX
6gWrMNpwx+J9pwvb2/dwhatv7OK0mWboMYrcI0/0cX+nTR17SKDVxKW6yhldonTO
8gjsX5adH7YIEZPsDnmudW3pahXrhICMFq/E/WkxinTRWtmLeAj6/LMtDovBDpla
ninsVoJXZmnSVJiADgk7zw19v2oHEzFI6mQ7eNCRgZC4ISWS3nLo8HqNfawCkJhT
/XSkeASsmUV05EJg62+u8XSPTzfzsOloq2wyFnf70nPwWmA/opH0tQc41ogie6jS
Z95Xfl8zZeyhCtrYpLq58Ac5VnlumQ/aXmTMmdA9gsaYCbseQC0p6PE/40qv6rq7
GlFS7iy7zpriQBGqD/c2zD93fBQ7j4xDgN6DvxH/TnZ/p3bf91toEVeQvtSSk0As
M51rRscIyI3Goy1VA49v1MOAeUhMLz7olNC+6CGzr3z4aAQ2ls+X7TefVTSlNpZH
mLn+8VEL65Wh0eYxWdtVeDVEABtjQ0gcz+jC+kJDnRt4Q26bNpyCKQhh7TwXuhXC
acYvk4UG2z61mLDcPJ3ciaK5fGWsOhPL76t1UJOblBpOYC1OHdn8kjewgnIGdttg
CIBCp9a75q6ZNMmq7Fc4b1feUlpf3AYgv8GNmwsVnSDw7BRD6UxtZJDoelgghXpy
CSvkYkAduQ2F8ch2PwuMX72bKiqVLN7WG4p/NjYwJUKgEqHa1YX/epd9kgzTGH6P
M0zOvS+ee9BtN3i5pPz3QlTGb7jJ3gQxq5N3xFx/Yq+EyMoY6ZqlNL40YdmINdUs
GhbiF3ouHAm8GfeDUc4Sq8fQmZx+1jEVE/pJMK3zznqbCMDCE9lKU8LAxKz4zP+a
n66OQAOyyPdtluVYt5NnrclBLl16BW1NM5uu8Rb6fZwwYDdJUdKyV9fcf9Bq+wqU
U4tM4ZwbYE0ZmLhc13X6SL+8ns2qHaTJprRBCNPkJ41bldAljjPnsqUDEyB/Ofd5
U/T6LX6aNWfhq/I9IUAe3WHXC0YoBNlrDXFIKMTS5vZz8OHVrH44Jec20tIb/DPI
lS31TrF07DilaDjju1IF/AJepzTYAHSU/gyJzYEBBKMsIaRT0jAwZJzph8qSyup8
cswClQbAGenPsbq4tqEAo4zJRtZo8WAYw1mZoS9g1XxCdx00tt3IyLeGCDLZNxtg
BW46vjhQi+P9ZgMfYE65zDG3CMFh1p/K7RGhPEJw5ES32ciQ2jsKnXyK0e/UHY8d
yrqMp7QDo7LyzvWOjF18bz4sEsJxsi9g+NWeDp27NI0WEEz9c52DwskHje+4YQ00
syQF49Hdy2FxeYZDzSWwGJ/YVx7i0iP8c7cZ14pbkZKNsnb55D0EQYZcmg4l7jw3
Gf00xro8giO+HOYZmGjbQjoaAU/+zn7oFG3tL++h3soLEKt+almPh9IzhnDzER7l
MB9bG5rY2FL3qN91DbcuB7prC/FTOtIBYdxvj1jRVuXBN+eBZiwuL1XK8bWscurF
+CSErKD8kqTh5ygeSmdsyo66i6h95PX5GylCDTP2i3DE/K3dlhzQWo5qnAqnqbPs
RBc5YTmy3aTNuFEfzeqHvchw6r/V0gNSv3uxBigS3XoaQ2zsOjXTXYMh5Hz0dF3W
u5dinN+l6GNFfqADd47Bpdbo17ErnhLwLZC4mN1ioOxHdWppmVYdpzoVOQ9MzQn+
yHdeQ7UEVswosU38/XZzOCaKetjPjumu97HBm2Ccm/wIeTIH+22MZl2ro24X9wdE
VCebEzybDd0sJ5C61kd1rTeQ9sK9VXUFzUOdup9a9rvOo7CfkD6spUsq2xsrh5Aq
u3lRuKQrFAkNMkmfnrR2XTfjeadszTeUxxLXf10D3OKbG1KENqrB0wdGZhqidxcx
HJ/BWvyytGXzMpkVxSXTVttQn//1aWtbOQTY1Zi5dLc2/K0WXEKCbsEEHFSencLH
mPaNbTe0h2q46CZAzpEW9L4uSBkoTjs3Eki0Q8Axl4WRvR1kGDGGTAv9PK/BvaNg
MgDzcLX8Zzopz3ebJdZ7uUCKpVijyPVcgT1SQuoUvjpAfBn49dNOWy/N8/KUX3HW
utNGAVh+Ltz1+Qb7RFhsumcr+bOSXX/U0HJyt2eVUAr/GecYxFscPZhA+AomIrHK
GeA5AXBOnCDEFsQXvlk5gOe1O/ngRKd90XDojZ8ll96fJVR5IX2Tl94TIYAaZdfT
CUwxJ2Alt5XWT2ddusc6GdR6Nrxz+bkWNdFOEW3RjiLgBr+c+XnePtUJfE1/6Cwf
UJOex3WOHSStDw1avuqQz/TPhSYQUNgWiziIQ1vaab9rbUzI9JAtv/wSTGh6JuAd
9rkGWrWTZwOT5xhBsCfFfAaxAgUu/jrbdZe1opzrQpiLyz2GRaXtxIlu34BK5Aop
2ml0TY6Wl3/pwoi+dnvjIAnRpeMBL/VCGQ1QsyRiBhr9AuNStvK8zbfJ6UHoYa0Q
flUbxjlDq4ZtL2xTvWbqb048OMsCQ1byLMtxiqzOxbRE0nWnBcJU1e6Qyg7Ep5PW
Tm1q6oIYAnTlyKcAZMTINnGpv8BXW8QUiZ+qjpy8Atse40TnS1Mqkax0YvreM4Im
Xy7bpck268N0t4Sr3bg7V1X0h0hPRDqwa9aevA24KwUbADn5G0A/Od6urin2ZHCC
C5IpmOZ+IDnL+mV4GLTQieqziqTbOz++NVNeTCLRfbBQcw7T4IGxPUmcG8lDHDtK
G39xceYdOpixSFBwMLoD2y+d0HtQD/yb3zaqZ9K/roIddIBoOckIkO2ikpsvilCC
7fODq0xjnD/rZikc2MIoRLo1c/utuQkby+3GYyRjSoHVNYdJEaK4KVvrhDQrYDrR
RhQ9SfPFz3swXl85ltMAU38Bejdfh5Fc62zx36vLkLXEtlw902jDx2u9jXm1mzAa
Fx3P4EkYNn+JIlHbodIHHCqoJC+zEMT7+SJKdZnQE3MldBzJwH2jUoU6PJIzrIgb
nyyhnpGwgxtrsKGwdQIDzUkJJW3Vp0PJ+HmEQK605zoAViMiUvgqpB1YcCecntlL
IBPTxfKp2w0DOOIZ4oPNako3UP0xaZeOtgnGkXCgthzg3A9bJ23kUnuLzxU9oMEG
/2ZEfF/JMBMsAO6BtbVe0HYOrMPpK6GoQuPjo1/78uckkGu7dfu4XTuJs5/kpATA
O8ItbMQFpUFHzukEZJgsQ5/owENKqAaB/1siPDf7qJFR7vo2PIg44IozjURWlJkI
tTfM4fTud/AZ0spz0ThgMXlTEEHA027o2ZmEG6sFhdgfxTyDEYqrawbiXXKm4Fa8
wNnwvdFAHFFiMmV+ZzasRRp4w3DWFK/X1/UW8UL2MJmMVkIccS8HaeTIrAmBsnGT
qr+6u749yGpLMPvrAokPFvXVOiCEzEqNDgwFudE0nw/jxb+kMdcN+9PBK3vzTvTG
0Pn2wQOWhSY4tlXgjBl1zuoOjg8xKx9eCjUa+DWa2cgE0Oq1lrVSzs7IqF1SpBVc
1jSwGnoQ2NIBjvJLVcbv5w3goUTijgIrmWc3IqPBaF3Y8vumHzYjdycWS8zpL9o4
PY4Xzymm4RdCN24xFDV5Vw8KtWhqoeSjbxSPMSWUcEQorpfm5HY4PsMazbxP7KR/
NTdHXhZ761AsVWi+lNdwl6lq83OYPB3/iI1sqw3pXXZBYKwMt9GRd3TgtCZSvb8x
RMsgW8GAAcf/TGbyK/toX0/EqPkA93CUPuxFzEkbKWnS7o0hLCd2BwsrU28+96hQ
xnhTgPiaa3xaWNcljSwGdacQP0SmmeUwFZ4oPEe7pQw/iJMmJSrgeeeFiw43fUpq
AYpALfHD5sN07YwcBSwc4wzZXZ8/NJNKH9bqrqXaw1pZhbVSkCEy42Eb8s9cXkKq
0zomIrVaa+i4w1S6aVyiudwVjzsoChLskDuEjH9tCTlRSTTGoPRFIj1zY8BO+EZZ
vFBVvOEDnkka7KdGPEf9PhgkRZUZkQOmJruvaMKt6dX92OLGyJnXQ3C67dscrWuJ
wapOm+DaBDfGON9TNIuRqYnvc/uFXZKbP8sljKeUHiAhXM+ZXjIjrZvrNZqReBQ8
cilBM75RU2iHrG5TW6/5O/za1i1zRnJvTXE1xct64XJn3yWOoqh2x77DF74jSIfm
lDmki/7DU+SXUmB8NZPgZBpMoEmxEcm2Tlf7f43vmoagiOoI/MHzhIbPfiBYvAsO
In0Ir4jyu+VmrKJ/5k8Xmyu7BvTaocz7yA+OPHNkX6+F4F5tK2huDMEppkCwA7m2
Qx4XAClLuWMtbL2cE3sCNUl/Q6tn88d/YMZA+Naf/9XBIsguFz1WaUxt2H6pFRr3
GNsK0iC9toL0qJx4fMaliAnc/NegW4SEKYkFgnmp0f6l9AUmcvWiVeKjcOeGIYcC
agt/oeOFzONy0XCazIFDOT99McerQtT15PBIqgeceU+9usnuMKwzJRVgZtYAsSC6
Z21nYFPGCDlBWBcKYvEgb6Jj/G8J3GFMjm5z7CYtig+8C183us6qJStNUqT7giUB
S1XfXaT+0xkTXIKG7hOA0IzVAigJ8AZGS0BX2Gn7q0/NmLBTgtI9WiLp9YlyxwN+
dLjXWGfjMaF6HX1fg6dpj89O2sE6sK/zS/QmHnXNVOtvgav9selrqwUNUPmKswqV
IMCbSmCu0vbECYRBLTbEa30vIJD0xVdNwMhZfz3jyqVmQsjqsgUiTmtRxGnEWjv9
JlBVSgPlxEuD9J2lKVh0dhsAHIVi9OTQzRZtVNoT5AbPOgFtQLKnDAXIkGkLGcf/
D/uGEM1dADHDaWyKYUlfQnVuMpHv4I/FAWY+5CoqOF4oUSa/M7ZoZxriokrMEGP5
5yOeCvu9TvlhiduBw7ugKNjDAqfwjxS4GNY0/g+jC9hYHZbmS1/AyW4VIxyafuXR
aR3Ioj3VTD6wxAU8DrGmaf6LjKebXqCSsdy08Er6sLYWLeY+QPT26yaro/qhvPL8
Yreeux+m1ckwI9zxUeoSt5fSxJga69hL6xDGtP+y4UlH43nZeEw4h3gRNjpK/9Ln
TAXHznyVWqWPxeFUInF9B+cpUTIm71yhrrpqUQsMUDUjUITScYzDTIzWfW+GOSBv
LAcsS/opfUQ/wbcMRf69pCBmk3UmR0Q21+9U8f1idWD91goL92ulp79Pp2GXwPPl
7fG4B4KUJZSwBp09WuVRWRDi3WV+wn3cmzRe1py7GLsiYwBKAUg8Bx0iZGnrtLGK
lLWufcrxysrA7yNTIHkIvlY3pgpickzwOOE0C3lPjDewnUegxkSTWRiDhBAmG3LY
mC61LuT3/vQrXyP7hwqHsW3ArPnviUvoyuqPtt6TOaaoYJnJ1FSj7ocNIWwG8zhj
b0SbWecfJGUhHP4f07LbfXEbdam6e1ttKYNywG8zVsnJ7K+K5Z1XG6pa3lfNVvx4
sv5dKBHNiUWNumCGSD0OwZ3vMW3uenBPgkUnMnCXTmRf936hvKXUDaF438Q1DKKj
pBuHJf1RnrNZyVHRc281gOXauLSi9IDVB5QMA2Ki6u/E9xasAKnpYAYmbyuQdp65
hYsi06DGqvHL8Pwc1mYEk5O928ZJnMAo3QobGetY2O+QZzEAAQEuGRQYRoWqOLht
RCV2ZNemDIjbW/I1i24QSyXiJKZM5WF3FFU/FKUHkb4to69gI0okn/bNlWFvRyn3
1P1ncplQZgeLTZ9/b8uuqZt2BGIQtt6uwejy0+fbw4yNkcB0saLM+0OdBHWJ80+j
MbcB8DKOqGafr700SB8v6qID3BiOHLCgG0PLVfCtiuPeKD7DSTrkMYKC1huBRMDM
4aofe2h9NCnrvrXgZxguSbk/wth1zL3nK8THiJWVtBMlvVfLl3zZk8MDW8OF77NI
rZbXEJiJ8EXUA+6ppRLJjxx0slXfALYer1ftjH5YRQAspetE/twVhVrfBIxm+yRy
mIUwezd2swnKrkooJ8E/pY669XER/J9igxKFE+2tgEXsong4s09tNrstxUOFgKjf
nKYNeccB4jBKYVango6L04SYsgV22NSxvhVY+ArZykoYnl0G+idLIcIL/YJvMR8Z
PIHXuznfcoENSuV9gQGOWwHOxCtrrkfvTusnVCLCxmVOY1kY/q/zb/YnVZPUN5Ip
0I0mePLOneZvjTwtKSGCzjrxW1AaY75A+cHRNSdZTowgPbog2NCyITyJOxhCXN3I
aDei2APcxFIp9KeyVSJG87weB8jNeTpZCd9VU1Ys4+Id/iAYyIxUJk8PfhNFMZNf
0hjzKSnYOE3rhxA7WlWEnftVicG14sUbY7JVFK2FT4fQFwyBZeEsnHBAOmIEqNMU
r0Sovukd0LME7q9EzaHIAj3mt7Egpd8N0iXGvhtKJc2/DT25VYN2emPVft/COoXG
CosIlPikMFZ12CHTIAWXHuB67qAdmBw7CK+L/6yjFS9zJpEKF0xQdaAHB8ETbmKh
2dDnLNG+kyxudhHWq8TGiTk+bHpeZ80yaMMxS2q+F70+qcXVwtCp4lDOTD4Lj91D
iV7p5gZt43YSZJ7ppMSlMqlDmJJV4yfqHSfNyuJ0jM7K8lMI+PHmFbrHUdgPv4ro
2S9kRSv10y45H6I9LhD4finG8MQjPpnx5M/JeL0LqIWgLnW8X1MOJxENGuG3NTEy
2J5HTyMiUjDISjjJ7c5zRpMWKQaQFHir4OJ65ROZySQpfi+4xO9i9VuT9NOJH/5c
Iunk7dRtO7elGLu58R8B0QzWnPC/gjzrpb/iUqtVY6Eq1ERE4sI2JIntur04SXkG
RB1u1C4DRU0SCl7944C/efSCPt6Zbg4t5ShDdYNQt1GnL/urxVoeItCIJoVycCsN
8G/z10i0bzPH/uQyNJ96eLF6w2DW7dDqkUKGX7ICUFoeNxRSQ49RDgqYPUcrWAFt
YjZJVZkgnpbOcPeaAl6uU6wWxKP+6UGm0eArYZHQlZj8TgEUAQ2t9rABgtSvYqrL
+iKQjaLFrl8xezvP+4FZgLP+SPet+f9b/uzjpGht/O3XpVJbjw79uibZCJVFGXP6
iOompTNXDgHwQBBseyYPKUO6thE4Zh+UrlAqnXEiP3+toWiVsktMQTtUk+GmcRCa
2yZg/1wtI41/pkvQdxxHerUVjzS5w3zN6BYklipNclzrrRRn5Si14EKAx3lvGup1
Id1RSMMDfne5GzmPuR0cR0sGJrld5wh8c3A9vdjxTaPIbqbfj4nXzWjIXr2YGP8b
2dM3x6FNIwCuRNpis1/jBmWHzB7WnNqhHpm5fikBd31Ti8iWhGYoq+JEPHA4aPmG
jWgkinEW7Oey0+eKQmGetmC5pPZljXv/1WKo6AF8KsfvFgc3iCXE1Cr8wJ9wKQIr
5I9CbyOJa0jDILf3FLqscgW09M2Acg01c36jv2Gv6/PvU52orHmn2bIIGaAGjtQL
IV4+yCLx/KbNIneVyH6w1AinUAz1x7QhhRSuseyK3xZmd9/fdeYDVYLOrGT3V1Oj
p0TGfdfweqWP5aBEQTl8BbbYAhCTFR0j0rT57tfHSZSLFSOqiASamQwe+e+IUce0
PPDw8616/SDb16IQkF4K11tMa+rqrNbm8WgpTeP/OgNe3CJgNHcx+Mh36EJbG8RJ
oXAsumIQUUfiIDKCe4lsYzc3R9fkNmgQnuMmSBpwncw2KMEPUK7t1v5CMz6YD+EI
gzy7wic4jvMmqNxAd1Oqlxqz7c8QNflQbQL+IhEV/s5TPoy0lpMmxuY2fckCGEnU
Df4P27wS//hbQyYxOq00OYvkI1u1///DFpsf7r+LID9/Cy8juW1spO0qxWsKV3fC
krFVya/bVfWfaPoezLPeBBpEx4M//ZE3QEwmvYt9QeDBlLa1CUUL5p4l8pCzhJvB
lft9bdLL2e9ilP1RHsR4nbwHi3NH0CzA9zAePOj1u4jTmaQCyK9Z6vCcqdFkN/QU
YrQOItA5hpVTuIgGm61aAWFZeyeUio0Y6DpYde+XCSDCYOYLvW4L/hfknIdeOouL
BPFpzjn2e4Ddjgi3nI/7OCdh4dVgj0Fu+liPYjks15SkJuUUQPGnrQzRilM2zvIb
hOJ78HqwRvS48U4uD9Aa+WQwVF1HxJSh3yxyEOyMULSJmW/7mK53pIPDRF6x55ea
hjL0CGkNDKqgsq+6+I9vVhXClwlshwB200/TuHyNkgAFyUln2mweqxKeTFNEuKl/
YDNpG5B6zRtvDVN6sQI56b9K1oyiLpvZnniBT3p3w8k30ijvxEr95eZW0XN7mSyi
7J1FGrqlfVey0mtPEo4u4j0dto8soIaB+CI4wd27kyJK+ps3ZvShYcPbwiRpKl3S
LniPqkA1Q6mbn85Si4WHYLJsWSaVCnYizPj15Gmb0xwfEtieiQ5dv/nZ57WpMVzZ
JPsl8D0qaCNTX85/yiEmfViZsMulBoZIvMeuuXGhu6LH2ib8yFx5Cy4vdBO1xaY5
xdOcmns1fvnsyCxN82cVBlyPsqHqnoTP8F6wQlsHOOSxcfSsnTIVD13bPgkEz0Ly
YnnWzivOLNUSl3l6fzzwQIURhjak/n6p/Z/vRTFtp6lXH8/QE8nttnSoJHrZDeQK
NByx0B5sEsLxBGFFXmzdznw9oXn7/kqosiHY4LdcL6cBeIjPDN5ZiD5x51Z6wnI/
rp4/LMeEJhdN5T/fpyHaVjoJ4e91B2+C8Z0cy0Jy6r1Aj7euy5U/WdD9CrABLDVe
gsZy58a/EPxq9Iyw/w0/oNhnK9eInR9GVLSsf7W5geZi/Tv5aPkab4HG6VB1KuFI
wJotcjIVv6NyIjjkqouCx07UlQ3r0RO7D3iYdjsTX2TL3YOsAljpY1aAmub9rOj6
lwyBrDuPh/Lf0fmOrPtI38Vpi5+MxdmBpIUhrHUt8xYOUlo8Ib2WoWb83uq62ElF
dp/AyF2uBPkTWyfBEGj7K86M89sy/ejIFiUPE53EwCDr38O7+JldJHSaVLNAYzDT
FjU6FdauPVKQaxzFtFfOJU5iusE2mLv5WsENLTiIB9O9X00L38dj0oJ4cSm7RM6r
qd65ytdtaaXdKx3fP9nAYYIz73sdxYNTXmCEPL+S6d3XE4Q7F3voVfJRrwpHkecn
UTW8bB0G60HHBaeFvawuW8bigx/qqp83L8JINXtfryN4alwB8FUFXffBXhUiLaaW
8aAxzhbNS5p58nMKkUBtgKbRPXWttlvgVqGbkdz4Oy8NQnBH5Rq9DziVBb+BaqnJ
yzaIm+oK66TaqlRD2g3cNJbzjuNBQMhAwA6cydUZ1kq3q+P094fvxr8JURmjhOZp
KwyQFI9PDWTwg9IyPVKm99E5fjgeKaU7FGWAMG9+bq8ueYuGQtJK3Uwro3Aec/fz
GtMlLP4ANBWzRiJTwLQrIB4Db83/gWrZttj3HtqSOBLG3nib+vBwczjkiIlBQWii
qGj6Wj0o1DyNcKGTbgTVTeG/gkkFVRefKGXRo4PBd/ZVdjOiABhY75EaqoXZGmNL
2lMCxw+ZiFJsrqPeKyQBVtQBKjMOsk2BiAyUKMPUo3LKX6r/CTTryt9GHRW6IycF
FOYjErDaUy68lwLgVtfH9OoT4L02W7tr30WDXYGiYSDiM+CicFJDxc+aNytFCs7i
HwAsuEtxAN1cxkyEGhuefCfYaY7SCHrcU1Z9kIzSHjAot3JzqXerq3D5+T3RoInL
DR1nQ6Y8My5oyHbLrfQwtPxWGrL+fqjZm0GXRn1LKSmCX2cm2Ajqmc/MFnE6W8yP
gDRjYrpzOe7hm3yw+aIqFKCWT7fjIjsJcuDUluhHfgl0H+zn2xC4KXLvCxhmNQoQ
n4h1vczG3dm94cpsPrGS0LxnEqXatAQlLYxpnam4BPeE9KpUBiv5/FiZaXdukIV/
nzuotsKIrEMYClg4S/pVO84JoihjmoFp3vPfmLZ9DlZGbJaRPi0fKCVpBwVlLSD5
uWMSHk8fPBFGmnq1R0UjKZaok4TbXd7fPuH+aKy2bWeky8AaBvagWAHYZJxqu0Iv
D7V/MEMijai0+JDuhhOVjTeiavxH0tAEmdzJZnow6ttob+I3yXbuCRUnkrB27FCg
BWa9oN2IUSLqs4IES2on1jhWcuIPp8pkeSCYBphYEW3FpgGtqOukdhq93K0DgoeL
kd1j2Pr2bepaCJYzc57IK5TnKD6nyGvGK9aNukoM79gByXTuDfoVaFJGZF9hNpVE
856a/aRS5B0eZTDf8/M/ezXWSiiwe8dhpYuDYavYndpfv36TjeBu6fci7c7k6c97
QJ0/UZV+AXUH5/hcrsE+KdDy5h8N7oZxRHlBIZBP+U6f+Np2HgMcIZMJB3vNWsLV
vbacOdJvMJmHJXCgVWWZXyuuiDfTjZdb4yv/Clnt7t26tV36K4W6HjOIpkFwBqcR
BRQqVWTiVz9I72CsghJol3sU/KSz0/Pjtpp493WYrTPsg5S/29CSlK9jbRpNeS6U
YWSooLP/VAeQ3T2nIoAcE25gb7iFw8/o3r8a41wNKdjmEifiArMPgHaAdPSeGtM/
CyCPzloFlj2B8qdSZ6HF6hOlRVL2uMfGgLrZ9Hn8vgSl619rpVgcvF5A73paMHFq
Y+zw8dPhwOt2QV9D5Z/0JT1PxFGQ9qCiHeJLu99QbYKJqPKhMgykOI3myuWBcoHa
Ewoq8Gu98i+IVO/KUfOn9wFZ9HrRlj4+8XYAEskRgy0FzF2kDoWI+3IQjmQX2Rkv
olzgxNigb26qnV1vl5nrDxHI6PY2Q5zZEOZpqv2P4cIvtE3kjO492RgjjU9GsUS4
4gKQo12ZA++dIeBstbZjAYpWyn4Kdwh8UoAaM5mNSarWx+b9fJvk2qdmuSPoK+wH
LJ0+Bej9W5PZL/rQfHb0wu//yvuQjlCg2W1xxjW+CceWkfRbSiHkE2tCoctOv3g1
wEN62Rrld/GfdwvjDVcVVVjj3GWWzdmlhsU+NCj8/A5d2HSIowmaAaZbd5xnz2S0
rUDG9O1ZCJrPakpLztpRX2FJbv0y9cPc54+0hhE4mykBhjxtsWHopBLC2CV1WNgC
eNxItR1JLMB8c7tQ+AWst7+aBIFJT1z5bVBMaieTegAUaYDT9Z+ux8R9xReNSkBU
KbcMIIz+iFP8PB0g0tHi250auCq3Oj9AIg6C4ixlYTuxrJ2csBxqWYCTXrchPctN
riI4fMG8WYGoHxTifm6ecQvOzV3t9Da1B9J2RswBm6HdHrI74zMEPbXEfLOhC46o
hciDwUKQNO2Q9xoiA7oggP4FcGGis7bTFjKomV4Dx/FLOkTddXx8tffwzQlaDGBu
O4gY7C1AW6+Gj/UamP6HaV7QRPWcimfRjoklDAgOKrro9Yj4IeO1dtTS4ZyweLuq
YD1SbMUYCSpnTd2Hxnk1PiwH1tpLW1Fzb6Pef6BmrlyyMi769LGxXOePEo/hvXgt
4UZcUXs6PC0E9PqdYjxwm2sSntl/nNcuhmbM2qHkpxULwIQjZ0T6d9SaiRYn8W6m
RebfA1DbaZ7RaTEH32/dxCOBpl130CZqdkKpTD2n8qPE9LxjfunehM25OAARSq6t
RAglFfuO9IzElxgRYVwoCHAAwAfYKzHA7lS04zwIH64OyfekX956fHbOvBjGiWSB
ujpXiQh2ZbzIDAkj7fICvXkDSeUm4iX91P6O+rv+zsxkvxJm2xYBvqb1pSqF5Ta6
sRhVOalBD540LzL9fQCvLtupMAHSureCMjTtWJYjzhSSxPR2sRmohpRHrD7dtbur
NloX7/8znzHDbGRzkwAooxWR0ujIqjIPX+guTpIZk04uSjNJ6PPvRWzHwk2ZoJ3S
L2zpR3DvXUi+N+5fJP2QRhREAgv125jw0OzFO1dY8nVFSEPdIahykXh5nc3+hDw6
hsGu4hNkPs9zuOpIku0n3e1HedxZ1mrjj2AeZg35rlSXSPlJXB8bBXVD1i7iXk4O
xh4V1Ld4p8oeRQNbU0P8Gfr4T7HZg/OhLzCA4Is16QDOF7CCRPVLTpST/AkpN5U9
YV/8FOAjb0JX/oJ5YU11K9G8SyHpBU2iL/qFJ0RLvvILP3lKegSBcUdybyqQPuIY
ZU21UQeDEDGCOv81FRhcdzoNnlUsytcSbkUvn9HNxSHvwS8LSGZj50Nka5zlcvxt
8V8OGsIwFlVvUe5wfyWP1bOC8t75otXgrw3xN0FtEX/vvz9XTgLumsI12xOt0In9
EPzdDzerbIndDGJ3to5pTQiValTDEn39MznrDDlvYfv5fH1Yv6TOGU9tkaQH/SoD
/d+Wv0N/bf1RLBV0a4Rimd/kyLr6h4eETs2jS+K6vGU65dpuhyPiJFknwRcxEM1y
0Sq221XROvWgKnjKKMKQxgL2ypLXWItohsVpJlrz1onPpVpbCYE7elzxj53YNnZF
ZAtM2tB2AnQcQPjMI66od7C6URJ2rccG+0Z//S/bJJU/6sEYpbtNDrf2zYmAXznL
fjnThypGCAMC8qUvvCIM/JP3KU5v2BnUoOzSGBDNl8h9YBtUpxjrUsk3+Bo2IMdt
fcl6UPRgt6+ATtbv7ZtXvJbgsOnRGf4sftixap7JMOhl0W8YGI/XIUH2fL/oBwhK
rWdMQ9Ied7NsULSDUGi7ODxHWqCmgdKN5DlzBn1fdAPsnUDNj99PdOOtfuWAkVNm
xvjLpPAMtF3IKjVmCyL6/G2SzhQJDiwIPzmUwi9+Ovj/VkLHO537tRRmkYlQ3ND6
m93zuAA8AIgJHhGpvHONbv60iazJEx4CVQ+HrZa8ynUO8PShrFtisuibHP74F28W
sO8yIIZ8NORpu0yrrqs71x+8+2xNeUxC1RACtIeUSLP6MEC3BmOGTS2/rEl2hsqG
s+IipMMW4rsImLtjaHbSaulCcWZknmP4NvjDOHnJ6OtxIDd1yq7cBedjjiwjjJyu
qSSvk6kwp0/T6c5QjeasgCXrxKwfIKGqFPA6gN5iq60bHF92vyvlt/bIrfnWmkvf
OxjSyHY2MZ3e5NFRSpa1q4I/lHd8vyjFz54FcadCu+i2RPvGTmVFwFsdS1G2vHlr
WcSUIRk8cIu8nmxvVB+xcjk3pvoxEt4OGVry+J09f0m6rl81Z+ImRS3N0ZqSYjgB
dREs6qMPbV8S5JifFzG4aWGBs27cdziULc+VzyMRqm7LZlWoV6t85djjL1AJtfqy
kJs6aJ26JCVpJ9021T/RspInUZt8PS/e0x94XERDZ9Z6jegVRfpkTFSn+lYugCkB
eLDcBUiMyxGJhLdhNsQ11BpsIejz6Ay3qv0frnSuxvLrfn0Tb6OwJhXjbFMsQh02
M7KK0js4tRd4wCLrvsr0tVBTxXTvV5yUWO1dkn2cvJ0bjRFd2jl/OCrnwnspx94z
uQSgmi7EKuNXqKpRmYd2YbroHdTCSPjWVZigtP2NfaPmLBSfbwSk49cR4Ap19BW5
1okVfQ+q/zM8Y1nNUrACbrLw4PtJTyTsc7eYB2H6qbNtz2cepkolg6L3QKHA194D
L0FP3pDQMnETn8+6rtXYZk8ARsebY5fL/Advkvq9S9rAqMTXphIriTDsrVpaA+FX
l2NuYXmzh0pMpGjVxZmVvAZgND5nRhO/HbWopi6XbJrY+lAksKD6L5SyeIdYuzxz
HKin+x4o0CR9pIqDzW+7F4tWR+7+xEUlaaVnPCiQ7WIBwvsRi2HHSw1I2+P4vVVQ
Fhpv0I5bf0PM51SxxlpA1g98ACAmjt5aTJdsQg0uNw3TYGFejZR4rQ+1nGaJveY1
Vj4GWhJ5iCwj3xjLAZKUYhgurGSvdW1EUjp5lPE7gkEAaUBSZoLpE9i5xzhm1jcW
K4xyRONZYmU5OA6eNictDDfrnUxIvfeh4cZFVwaSXiGc+WR3zvDxbqOps3LA7vpk
ax6lSvM3ooGR5uhONqS6cAZevKhAL0+E9dT9mj/sfEx6WZ+nuYnTOTBNS5WDZkLO
QDWgdtYolZ80bRtnpxf99EvpzVby1E/ETNbh88dU7Hi5MXwJzdWotpGQQNKIhfMd
Fyvcj7I1duWD7tTEwti7lkiGT+6SoZW1CsXnDHHyTpWuWLOuaVOZ1CXB74gpyWww
Y92b6GHsgTHSMBnv5n/j9Ni/VhjHWDzD+cCRx1JpJEh5/t3Qu4DzEXspARzwufJW
JzgnvEk84PUeK5EEpxSgqvWGTGZKkfxfgx26ZVIhUTkGHt168TEQtuECkCwRNe6J
6jEFHD7wxwFlkTq22OFlVYU7SWWsFLDrx0qzYRIoDlBvBwLTMlJeWNnI7H/TFLgN
T4jrpD2LXiLUoUqvl7rbmJeq7xActqGfQGTaWMR+UT+SebUDQt9vagB6FcCyW3cC
EinrwDp29X6YrjKsTYVWwo6KV57gxsqYXS4r6JtYC6PjKQdoT3qmUsmu/YZGY8eN
WCmOTaj6UuCbeFAESVXl78umTQ89UZj9PogkJXgTHjPWx1U3Xw0t+cz7EA/lAyim
mxLUniMh4zVuJHY2a9KThPpghZb3cVE7u+jW4lVIm0GhfJgE9E3RHz5YJiZOOgku
RMf4bfihDdP18zGBCkG4kYpbSkAAY4fRyNwKPu3uzqX8fJV5uQ5cvUFN8Al/zyjX
CSXrL8pQ/umbdivMUCsQyoaLxN1NWYWls1edAqite/187JgJtsGUkU93NIKSitbg
DeoBbecm37XGNn2zxTM05rhYylH0PAX7P3eqJ+MqhVfABXhOgPY/36YGH0u6ghqz
TSoiip/UJ0/QtyCtMdDi0lpxqyiK396irbL/ogN5rMgoq5YKQa3dtj1X0jy65etB
gvPCa61/PE8BHcQCR9Lnc0/VxsvNTj4OzCvi5JSEjzuR7n7PkV4NfxBB+OaEjprb
eUnJlCi7s2B/TDAcSOfaD8MT2yim/t/bosyPlu+0qSWXxJuVjoAaj0XuUUHH01w6
DTSV0nGn5fsCjSxNkUCh3xaFIrwVyppmFwWhC8D0aKcIXI0GTeGlWPKwaCQkGSDe
9d4VMWbTIfM/pJBvfMnPMqE3qT/KhKkQnttlnJG7RIjGG2vuD9BosECWCi6w54b6
4SXgstjcvgu4HDUo3sIutvX57HbviO9W84NiErjdMfA+qlHHw+jFAMRr7G+qgZmG
Al035kxc/3EKgi+QEGymoha0/6oRlTErTNrhzOMGuwgN0JQiQbzoQmy+RvPCVv2Y
qKduY07t7o3dSvJZ2U4sC79RUFksU4p/hKcbJ0VpxY3k26EqrhDzP2St04VqYTNR
8UW7th4CiVoEccU/bgPn54FiMIwXVejFzsHGsDzs/uMj+eNhpLbyF2mQsFSoaW27
C6FqWedwYicGbTeiJcGw1hdBx1mjEtcrWHM7pHvxFNJLfhAskEApCmPdM7SV1iKi
SIQPUuQFrbVky6fZG8R7hP73Td41N9JhKeYcEsiu64Pfcyv4xKJ6p0P3K/63qLAs
S4UiZ1EuppUDXfD7kR/sKfJrTJjzrWl+RIUwa0pb1niVNxdnRMGrcM6/QbnMh09b
kLh444w0JO2Z4mxsmvcRIBQJ3enpszNHTtrCe8dXI7GNW+VTqrqAs7KNYi1/eFp+
xY1tHaw6k8dQ6TLSl8nN5a7e2io0zOmynEzKgoucc2kKCiYfr+u+wzjlbU2sLnY5
Th/sE5Ee23x6EN/WQl5DhsyWU62098rlsWKemSQpAvhML+V6+c2Lb8r8nNBDJaCq
k2yb8ZKUsCSqBtfPg8IuRmkl16xqHKMx3Imewn2Z8Hr+DWfpxSU/iFeqmCuPTCRY
VgBk+Ky3LpHjT2SZx4twYu4pwtqR3yWPuPvY94CwBQTyIIBtKITlzxdfiBSmFgYw
0UlclCy6d88wo7TUpNc5l/Be8HJHis7HkEGh+IPEw2SF8nWvcekRdoQgUn8uPVBW
5JlSOYosdONpm2PRwJKgU9F96AJ9K4OWcJPmjUND72igAvRVnHcSDWjp+fwDpagM
WX8NmeR/OWvWlR8C88kxQX+ka/bNPXcQOTBpS9qBvRXkE8ZXC+QYHgHZ2vBYE58U
WWmeqGBtByQZ53d35LCrJ163r285HBuXgYsdVMXHdgNoyzowH964JeWNE30yoV4Y
lUHt7hZgfk1UPt5lPgkWHBNvZEXN7lxesbArn8+6q4DKZI6lSQ6DK1KTzx6meqvX
NAQi6SzvIxupX5i3rSs3YKoGHdsvEqpE75/pHv2pi2XMp9jCQ6x3EtG0XJhYGXah
ccEC9lBl3JK74i/7i1djWBgHaeZY68wQtFiNUxPPbYNqFCtLIDiGoPPZjP/H+8oE
3i56/AXBFoQIHCAoEC6zT184Bdab8us6EcL5uNWGozucYdCLnHnAhivemGiXKeZc
fziuIckra1gNj1q+kSHABS4H8DYiz78hYLb/hmylufc3+lAzz8AhCmE3myot1EzM
Pb+C1RG7FaZQjLwSTwSurwR1Wam7qEJ+1zSCN3viiyCwkjUVX/kNOlHo4x1NfVwe
PG4e6cDwGYdtMVmo7Gdl8VOeLiLupjyZaMhgNf2llycXV9N46K+g74fgnzL2abwi
V/PLdO7SYmwF3kKX7Vmenkp+iUhbfWV8LPV85MnxHWdNrAzjiWezipKAIu4AAd1o
/fYrCxTGRu36pTrdSt1b4AW/ISp0kFD20J2Y3QAajSZPUprW7Iv2r26UyGt/yrxz
pbCJJVLks+8bnLhLg8GEl6H2K6/CkS7d2Q2FZIc6sHKwcSA3Eb6bzuf3PzYtl6lN
Ng8dRzNf6ZjzGfnlqWVwNW+hwo5tTK3uMXEHv/jm8CNsuDoMHjJ/ob89Sjodrjdl
E1qijABdxHnTVKc0vtWvJbGB0y+wZSpIE5aTGDj9qaXyYY5Xcd45w9/qLkYoWVmm
cc6c3mHbEDplETdhyjVdeuEPEv5lYtoYW+YGZTB6A1vfIff6BWu81MiWq0HRJ8Hs
xZckj/JSg94liC6C0gdgFYxtk6t7JIDwbJb/KlsGuA1rP+rti1d0zpjTDYmQLaJ9
uxcYA+wXnNN6dKBFtQbRUDaihdtL1kZVzlUmP2hkM7Qnu/EszW9QFGOE2mTBi2eI
zWaFZG8p6CoGTFx+qmaN3KaAp1r/gWk6kMk9B1fyix0rPEk7ziTJQkNYKZt/MyE+
OoWusqpVX3xoY9odmSuPwXJS9CYuacvmKz5Sox2Q1s4o+Vpf/2RHdmazKb6Q9aN0
vsTEoslmsPjzpPvt91dXR4YT+1G0vCAROkV5eEA4CEa1yGbUygF6OidrAJR4Xn53
+QvXbyzNrBYtTxPh7pRjkGdkmjwvh2e3vfdJnaPH3kslS3+rFYC/YHgqhmoP3uui
WbSZlTldzkRPRUPx1I9uE078/gSiBHA9Mwf6sn7Ft22DjTAbL799XsEoPRsS1n9S
qoiHPXZVVxqVhvX/uOn+SE5gsJ5/KQ50xUqENE9TbO9L0iH+Uepzf/DI8K1xyp7Y
+cetZHqVx7VpOmJLVmq7sj3UP0aGPVrR9YT+/Hj50qOvzY/KG0YLnh4y94bMsYZ+
LOboQNOWEFA51/u67SFZyWbZ+Jk+HlJEBZgIx2HsXDAYrd8SlGu7Btompt7sBkua
22B66Ec0zsO/Thva78mg+HcPsnk4r45f+aejxKEfG/sBg6tlnArlaU2P34fmYaGo
H1+3egeL+z49QCSPxEAbJ6pUcwGQGPjPnIMfqxtTL4SBmnSrEr6uxtBxSb84en+V
CtUbrLgBKuy2pQHOBXukMLreTSWsTmySHsjQCCMxqSxJ+GmTA4EVbn0Q1h7QNeXi
MUarbk12IEsLxx0k7+fpsIfJBc4gu2+7TgiDsDTJx3oh7+dwm7HEs79tvjraRW/d
XPTCRdWelmemORkzJHNjwrwfL8thW13QB7O86lQeCVUvFwUIZqiiLa5ZKnky4td4
mbuB08YIH4cAMIE0/TkZym5MEeqpU37ioYd9KPuU2lJwBi2fQIsrSJ4iMJ8gMq5c
l2YYKGMgXsrTsyCewC7KxHuhH4R2srZNvHuKlx7psc0QfTFVkSifyLAGLQuZsK3b
2a0E5dS8dwUV768FeAhcJZEODmfbWUWtDU2EPVo0S0YF9bAQIVrJ4S1RK/++2c6u
j9CvcPVf8d6Vxh5KfQfOKsBre9M4cy0rXNIOpMr8owSwMmNBeHPW5RyWtxI561Mw
waIshArQcWk0ynra7ODw1Dd8M8wgBhWX1jUfnqaT2xh/bO1u/+gc6KeXbfQUqh1d
IYmCmHR5s2jlOpLgeaDCV3yrXQ0dGBFywDsT6JktJhiKZpcEUi+CVRtuoer9uPYH
wV4ulYZCK4dUKK3niYJxxH2G/Tx+087ehIZGh+RMcmRljzgYr9pUIlzR5SaAQmeS
g1/2Cldjufepiqu66xqPHhnOD+4KF7RZMNt4IdBeUbnhz1KWwb6d7xaU0EpcWqBa
5oCHYFJEAMMdUo5YmW2NjUUE6Q7GWElCprQMIKFK4g9k8eE/LXGO2uoEttv70M3n
L8mURdck+smWL7KAWgEvSWDEMumh2t5w0FS+yhWroMfEFWXdfm2VLmY1SHtx6V3f
1oLrcxzI0R3t2YqnAXyf44guyOqSuXUqJ9j2SjGYbu6qaq2VNy1xI8Yzeep2aVbH
LAn6Z9VL2aaxzYefcmD/1nrujsXCh6vDMS5qwTYskO6FKIuieckDIUo+cJahHK2G
/eGKUnElN7xFROcm8FbZF5S9qoFA4+LY1wGZC182bTOO/H5BzhYFHppj3VdRNofG
BHdNCDCItyALViFbdBFE+jYPSt0mlrrFElBqogjyNwbby9I0Mt/4IiMtQfkwFtY4
gpEdlI9h++BFNw1J3L/ipSJaqIRJU2euq8GeKjHu0tZGLlxX8AwxMGvduyLNme6/
qnOvA/M7H7ZosM2U4Qso3yM4tEfIssT2mAeLVGXFHyEH1aV/eD9xY99af+kVtiDE
HGMwbHzBhBtDh30UOI2wNvgMguU6o8N2U5xYsC4sjwxUwVkCH1NYh3FzEgkFNZJa
ckqgajuukFrZfDCblmvUXbzI+KRmhs9g/PmoWe9Ng+F8jzpW66rYbxTcpYSqYg3P
a7jGhQ5IoaHWUSUtEsMw/6x5kMYLbFTFKP0DR9eVaCRwgEruo3xtOJwuorJWTv2F
72uJ2PfaNtNJx5CsX7quMI9IvwMXln3LtTX3hfjHhavoyi7cf+hXhdCjxJVnCz3I
f6+YGAXfVAsYTqe2T8jDMpUf8cnKdaar89W7nGIlCSWejLuIL/Skb9NnkxTy5qo8
41Vsr6Kp4v5H+EPrQp9faqUqzR4VBUoouE3wX7cyHOjurcXYoh6Z4tPHj7xbofA9
7ZhLeKiG5XxX4nJJLT0OnY3yj+suus91fx0LzbCIfTSVWs//CenBQY3qq2H4I/Y8
zSHzgQZr55T9ONRYnXNe6OOfzzSmMVhqxcfSVDIvKRblPlKZ0JPljommQD0DwoRy
SLGPIrIVnlN8y+w1axmGwwGlOYjCa22tRVaXVBwsMCfQL1EHZpwmeBMqv7RKTaHt
tTTsXXmNelKv/dc8SMXksiDMlO28EfMZBfl+n2OzPgsvP3cDI2iG6SG+RtfQYJ/b
Gf3T0AeJ6IN0GfWjb5ey0Q0IZgtajt/iMbXJMLTHHASusQq9CwXPFNuUIIuEID9N
Kf9/CjYDyMgrJjyu3A26aeknJlwCh/yB1wgBTqWxt6kMvoBz1uiLNc181SRUGiiN
3IMCD2S7ELauxD0uQx3uL9okVa8y5wCfmyefqk6F1OJzIje1wuebS/auZABoDcFs
/yxroi0f4Xw3gc0MLqfKF4Xgggh+K+XIrOmRo5FboAiJLacsilL5v4uUPWboPbxj
raoic3oqD9IRyp9RHWCoaFPZHyc1/kiIj8bmDlKs5KjPthhErx61+Y2iytN9VyCZ
O8H0SBi7v67bt0LqnZ47MmbfnAd6iVVy6UdfaZt9LOjo9sialfpgyhlLfGwl3FAK
zzFBH7fnqkrIhVRGUjaOPFXl9EsfyxdbOJqqIW+sA8FLF0Ry6iv+jYPP6zjcifhC
PaUWj4fe4dP5uZz+TkfmZ0Xc61j1Aq6u5JlZFTO0rYG4UAjlibniIoCjtPrGT7XR
+hkzDc0BWYvAamWUzN4Oy8iEp8n4S7SeDTwoKsp+8IwiW7c7Wy9aBamJi9+gY4Ze
sBL5ici3AsiTO5ddXx4EBLhjFxKSS2PqyBC5qaEZTATRj+BQaksL8AYaicwitTNh
PN7DA+npC7IVoooySOCFBDeqLdg23Q9hSqae8Y8708qQ3AFbafsb69aarE3t0bLL
PieblxV9tSQBzSZDJORijx6fOM6TJf3MbOzifBvrypMcgt3oTchZ/PWM7JV+zmoj
jEoCptwgw7bd9AJG3JpPqkCojFVjGb1a3QDuyG8ipuyvkjCK3MR9V47B1RW7vmZq
ShxnAkS8K6M/k2oDV351AKxtPH6Z6xzL4NQZ0axWq/LQ7uKptYpBkcoPga2h9JRg
9c/UYFQ3agZ0jKpjL7zGL0HxlZ1WO2TR4jE9wgOfXVjQKw/dzfyakKVQ/cOr4LwQ
L3UtQsd8c1HYJvd9bzZNGse97e8ch0T5CYLNQJuJHUaIyqvrkp2BHMXTZKvMqpjZ
WlO0J10lRU+1dqe6i0kEhRSZql5yVjXDqicW95veHBBlc2Z9n9E6UQJECfRk7KQj
gTdQfyZu5+ZBcyiObDg7xxgFojz3LM24t0+23MSj3vYexHQ7t9V0J1LKshyGxH+1
tbqS71d//edlPLdz37C7Sj3UWFV8uMoHfM+D1ZOJa51YeSB7s1Hw7aLaSqcFcp3Y
bzTNZkuLn+8tNEBUrviNLahfeV4mTNByfLAkhEWtYnm+csjduwHfi9LiojOlH6Rd
a2084l7UqdCuJ18RL7fGEqJwyMW57jfJWOG77bEoygjbgn6MvZ/rCHY3hOZYJVmU
xwmfvm07cyImO1wo3btJ47e3yvn73cC9uhjWp90PAvtWGGZ3hGOSxlTVrWNeQXUL
JLmhkRkWa1MxRA9jlsP0uT1tfhcMaCraGpRpujUU/J6aA55Y53QJ+9xKNv6qZI8s
C1IMWHhMpalVn6JHMJPhTrEQojigLR6YIenMLCEEJIpxVlKkgSKh9ai1EQf5SDty
Z1nP8J3Y9qbTTo1spL2pc0r9Hmh51ea2lp0kFyriPpULFfZV1WesA6IsqOb3Y3m5
Sa/AAt55YZlVhx7mEQjggN78AR970OXRvALWW3zAOa6rpViUAEYSO4IUu5lwCCkg
osD3NFv0n3ZN9XUvvbak6kD3cYSgZMIlkYjVisSL/NrIey7rJLrYKKewIJPDTNXH
xEe2LeSwNpTvom1tJovaXc4dEhYg4sh+gvK6N6uTNfiQU3kylSAbOCyx9f8Vf/rS
B9kthupmhMSK9OGLDi3FPZNBsWCQ72727MLgrmimIIF6L3TsfpOhY2I6yi9qehBV
CF6Cpw0OF8LOS9Bjbu3FtN46DxE2TIkyvQ6QcHvVzz+KID7BeAiFFAw5nja1yR+G
Cq3phZOaSvA1LlQYFavD2cHnCuZTNR8PaEFDnPHwIylAMFFEO5lf79GdxoqVkdFL
3aS2pZi7LOljLmvlbDZQNffQC2WCus/PUHWpi4drIl4lKmulE5tUEE4+ISLgsz5O
s7n0qIztb94se9M1NHL5cyZpUuFf+OVMd5M4hVDajbCV915qLW9tHEXzEEGfBFHg
hq1O1JM0ZLbdO/tXzsCb0yZnzpFNXCwE/iDIrJDrej+kIjHozqWy8QjkBG/XKUbC
aytSoj0aHQ9QO+UyR+itW77cgJUY0kbqwt7qG6exTehZQ0XF7HM98CZhGf354Hd1
Lrby5WIX6Us7Jjdp1hdsv3/2/v+Fgm/OFril09Ooqx7AuHjHcrfvC/4thKIBUORv
GdUNVt+Yu9LM8QO5JLnDbTtj5/tr/gBcMFdLGdtr8P+/0RYb8GULY8MMZIdCQ8hW
Ig5PYuAwHTT9L3oT0TQZWMxVbZ+Q4r5T70EPM7UdOoy4GUpSDSuAcsQMIfr2veNv
W/kMBgbBcjt4EyjD5Z4i6FktoQ7Is97ZJD4ZfzqQ8aLZ+3pPP8dHdH0pCahTja8C
h25chmRhBARM8dN2z0cAPmKKhDCzHWB/Fagf3Etwulr+TiPnpc4bWXJwCeeKh+np
Zsrb9OxyD5dOKQ8S2tj3kkK0ZivHXXCA7FAvyVbKLsROimO9ibMOyIcOgJR++c7P
LryEgKcA5mKoDod+7PQxtCgAj9DtQIXj5xEtPpjhydqq4SGqwdrfabEDsu6gY2tI
xrqu1KcMbP7g1e8ZuvFV5k9Eqzd+8UusfrsnUG4HUgEojKj67CqJIByLZ8UwwaVE
TFTkLORUZHWq0GVcIEFMjkQ9oUWCdZXJ2uan7e4EdygxSdvs9GVvYVdC0w5iKMuS
94x+7j0EYRADPP5VRMVcftA/KG0EOmMLGH3QgZiEi+t5E3BeSZ1IlLH4FxTQtfDP
xBLJYgXKqqVfDQd+7Rpew9s7A5DZo/I71RMTvXhzHfXgK9CyCMbj9mc0l6ngt6Fu
ZQwYIm2dSGik4lqxKRQfDQdqEEdRFCp6gcsFKNQatJFb8Xcqhy+nP028Do8Go+nR
mwfECQpNovaWa+bdqpkvWIKe+G5Zj2E2DyY8uhDUa3AzYgQKdsVetuCE05s3y+ej
eUqRnz0hp347TdeiZFYHDQELn3zSvwgj+CE4yGzTKfsTPSjC+PzYWrqV1IMBuXqh
3fXvVa2nDLRjY5h+6+2WFgO9/3hpfsw2k4xCBPZsXQSnEsO7atXDzuyuMTs5VAdh
iSGOZDjWksMNg3/a9kHffZC27qL6YP7BuM3rqqoCkpcqRyHcjJpu1Ao9pKUR/shU
8u0rcGN6H4dFo3A/Zrir0EXHvPgHn1EF5NPnrhPNmtUTAGteEwt9AlhTkNpZt42M
eN+m/6frz4aq3f2kKTGtgioBFJ3YGxo+V5/VcwoAgpY09c7h335dwypFWCobwG+Z
Fn/OAnuUPuWjIaAvZbGxjYasFQcU/kqZ9MlSDtB72QTf8RxKZ/NymAINf8oE4mhO
PVALyofsZTg6jM6p6JQxeRqamfK/cEnC+sELL3WcPh+TSRfcQ12O0KVJVeciMdvD
TbzIRgSsk5GQRsVR27Hy9Ubsso0Fj6uIUm5w/y4Z12UdbhqOKwv3ikzrvXhHkNrO
aPWGK2o2nrOkHXBg/db9jloMlqRX79FgMIbZUU/p3ImxSgGMCk9zieod0ea4PSRK
g15SI87e8Fa37cPNmyPz2iSEd8qsbG99ZyLFPQoza+uxYxsomNg/UsYp2KPJnOwm
Nn/2HEcPB2YembtYfuECiAfBORBfUUUhcGnLi635tE93HHS27qjV2kEYhJO360Il
0vtCCvesE/DnAQWYPISS9DnqLVbndCJnFTyeB8ihR16MLDl+YThPTWDJUMlgAbQg
XnkIxCsw7iqqDx4bxQpuD7+MzSYaXeLKJxwmbyW+EXbkOgiTW993QeCf8XpoenRE
TK5FXpz1/0Ow4POPG9JbZ6OyfsV+Z4xEC5v7EZWkvQkZtIYyZaD1cVQu2+6pVIDg
tvC2O9wVj+LUovJUNqMQb0OG6zbrhOX3cM5wqizG2fV7P1YQMr+byEldoR5FVbI+
x420r6oWhzPUJbJxoVu9MWkIM7+EUeY2FGPw7rDef9DcNHAOf4dk9Rs3BENmU6WK
NYAVRg6Bss3wF8vPQ0T1rGMqS7JO/C5aQfRjrZ8dfn0MJjVDblVn9ryn5BPx5e+0
itC/3aj4HIib6krenwVVaV2/gPtbdIMKVia2mNMpoAs/mxK5YpwJdmv12vsuLg3w
zt4mrfrLYjcbqHejzpOC8+vNd4H1yps72qR7Pbj+T0QU6CzLYxSFIOaoSQq8Wasr
IATjuABxQOLWy1fa65rsiK3mCgsyEMwBEu5sBHDYtWpSnJrG2JYiCzxRygVR2lWA
18QXU0crRUF8sP7RoxcETfmsNSmaGXZ+j3T4IS8au8E5ziPPW7PSf5d7DgQCWrcg
UrI3NvTqJyS3HtY5yzR0NTVgI4AkD7irpl+xhs4Y+OZWMIQ/+6s9LAN2C+eDsJyi
DrKV0caheMFAGTAeC+oYZpomKlqHGODU4Kit8KF8q+KxDcK0Rrolx9xdKlSR+Zux
76TpKf9aLhr+rrhNsC6zYP2JRE06p2Qzkh/cTcvR19jBhxG3tIaPQEq3KPUHQ+Tm
P+qTU891j/0ecYEXgVAMpl1GqEbcx4o6yqbcPkGxhvmlP5PFlZA4pmN4EowIZHol
YrtFQMHmDXtnb8PQgdA2r/9KbUcaONhhzu4rfzi+FZXK+gx8CVd8/GkoJpZvbsoK
R5xkUrR+rWcVLEGkOy2EI7KV0DL1zHQf3T0D0LjN8bvpcfCuuuh2zunCvA31LdCT
wRYXxr4Z6fxAUF4Vf8OwBF17l3/jlmWIR0PeBhDJ815D7aB/ulPRATNt12+xXPRg
GahJuk8bpG2E7pQSDd50fWkNIlhfJogXiAMTgkFfEBkAOw2fAumYg+6ONxXI7kZY
262nOfhN/eW2JpUKdgpu1A4sRNFpqfT89yWIIgZ8tE61iIoaiauKqqVWVN72kLFp
pNeaLlzSfB/xRok73L0LZClSOieOu/cvUWwizmxZu9G40FMwuE8mUSYR3p9K1rgb
Yp9o6DBLk5zhafQtDzXLV/4hCrT6E95qfsStWfggt4wRGnuOne3woK4lAg3iZpIY
XZD4pOhOHV1HMgbeCZJitZqosaNhIheDz/w/2jD6zupxHwS2N5ZDI2PN42X4Oy2r
cX57NqaOZZsYGhRAixSHz3EGYLlYRM61wSTiwo0s75AdBLcFxd/2vepRsGwE4Wbv
o5O3kBN7ytPa1xzXYaHUg/aThKqT6xYTnQ/WLa/wSKTHahK5ae6iuuKXdQ4vIZY2
gmejRwKV6TjoVj5H5yZCkIzi9zFQTb4fTyOwJ38lQq+vpnmzVTh0nDucPzZsxtA6
fXVtb+68/z8IJc6RpHyY2W3Q5UbKnf3n8x3pUK0iCiUFff/VOuFpabiaZc2hBcgH
C/E4SYRr8shHwMBuK0k3XSlXHqAGpB75KXBG3MWF8RJ9kur0ZlT2BrOVAi7s+hkg
8rml2gVmXRuZ+yCl4DmO8pH12jyGtFtqFZV+UuvfIX6j/fSvsrvM68Krb4BcPIwZ
+C0H4I1iCHS+MXtes020xGvsa7aWXrN6o1/Fo1aFKxS3dL1sODunN2gf3HGEpUn8
PTqBs2C7MF4nSipe2dJrEhjg6R++UnRxov5/RaPD/umDZwV1O1R0LNKaMk0xQFom
sipJFhNxiENdcDYv0Dnc3phYEPHtBq2NPxo7UJSFtMW+OSNE3pe7peSVa6PMlX05
wgHIQzNkH8npT4sb7nWxFVYs9Qn4mASEI2kEITe7pI74kx1D5smgSkacQOaM0r9k
G3sPqaEG8IcVBZEJQp0nqYuwhyuNQGWXDpTBwjJwBVY7XKYViiHBU4JArABQ9wtJ
JFHXhzW7gOoXlZrPKWmr5gD7wgVa3Dp3UWDKMZg73XMd2S7PtHVDi6WAfY/q6OL3
j5HPm4HMNVf0ukxHLfS/TanR15cvP12oxZrI8nULr6lxpwtaxU3U3qtN4Z8KDXEO
f2AEkJ9r1P6j9FLcb651cd8BClzXpQL4rbuQRAeKbPXf6IZlgyMdWea2fccXqWIa
qjYVdiRU2r5FFqysR22FIlIq0zL1NbNG60r8B9pozelePie2d0AeZwUrbK/38pT+
ZmUMS8rltvUaaYYZ+QuOv27qDa6xOEutn5+ux2QT7HMOUk2Qqh9QPHexkQwiC9dK
G4Kd65EPlt5VnyiSQndoWHdOqvOOKa4L403bD+fLpz/ULWF8SOUTlJulq7NqxOG2
DBMxiE+0nBsPdyzPX2w3js12JrBaxDUsl1U5XhXH5tDXjpD+HHLAZebhoZUt8oEE
mHKv5GE5BScDpOqpDb51xPHtTUD6AubXxvBuwEglUjYC/zFI0atUXInaZ2U0c90D
Z3MTtQvSEH+IZOpqhWYrBeX1/wIJOL7hzw8x4FpLcOKGCYtSIeYdCsez/GDIxdhD
MKASTgAaVxTAxhSjDFXKQ/Kiq1e8nTdwCCObPRGvZqovjwcqmGu8the3qyosr/M+
PTA3tK7nW+qFBQaxHY80Gcpzs7jC0qlE+qjrIDKzwj6w1/USVx8+0QpJMGGtzjvw
P45oP6CKGulbWzg8iJS6AyXRxSZ/tGKr/lFVVexoKeXhoNHXlwMiRGM1JIoM3hEo
FCLxxRWPq8+OEuZTAA+B2+x5QbVWD/tQ8NqERq+Umnfvtun8lrmTxscmAa6JIzC2
JFIKn+w3oMiCdtcii+K46mQ1lE/jzO+Z4I8ej8iryNUM2wpKvVIk7a2C16Q8nme9
dXwh87N1RZ7Ng0IZxCX4xqOAWjBav3ukpkXBZQi8Yuwh+0meDvr/LqXixyNo4mw9
xduO09u4QB1/0lT1RD9VsSPkO6rQslgx+4+7tEylWChKWDhniNWfmxcWFzD5DNOo
bzsxS3n4y/VmQgY9m1sKhaAc4yIIUsAosVlIT9GUdOdn4q6LpDkpKkTfjtzzRE6/
YMf3e4FE9+c6s4GFdf6G8qpquKUnOFlUjzsfaiGwjnQbwtehzrkESFBUm+f19eHG
DHrVsdceFyBKdXP2o2W1tqDUlbnqb9BtVMmpz93nzTD26At21i2zG0KkgVNN7KnE
KfusWs/JHqBTKSHe4VAOaBUbTSHD1hgVOLq0awBRjbXlyA9+mON1CBcG+aYYprxb
fb5NW1AUCvI0qP/T5CdrW2t5obaxK5sDgU5Jd+lsh8hhpsi/UgJdaZqS0D/EYZbp
P1sbTSXunu/JHAPZymW+PD0z25cOLlGuk3NYPUuh7F+hNdvvDMntVhnNhWFk+l47
62TqJqQdKbRaCQk/DHNr/S5mdM01+GBvt26qtZ8PJLWascO5OufFU3DhZv5P9sJt
0g52onrSyCGEiCoMuCGHXuA/ynd4nr9FOHtvqLiAodv4pUIKzun2g9OerSEEknDC
TWaHHJIoST8Rp+QyINJdop4zXZrOSCXFpFSCCHWC3PM/H9ulOAGANBjMudDLlGwr
DCS4LzdfzsyRzoWLXmJ/xdtRKlxbMEyB3QOo72QCnyN0VGDZEmW9B4zQYe+DqVeu
Rk5S7MTuFsOKjAq++XyhUJ1VIcvk/ssHHGbly2iuK7kPjtIvIgWBBXj7cCG2UpfJ
nmUQmhdkszXSYrR8JRjMZa9fgrajcyWDocuPJaD5DZXzxUzTv1XO9SQ1s4JwMchJ
WmWQZkoOqj2rGG6Vw0qyJvwtc49R3KxyCdjdmtikAcwhasDgyBYyfQiNwBv4LVVd
EjxbeBnBXnXK8tTjuh6/Q0uB50dfelB3UeBBMBOJHeeVTlS8l51hWpt4Y6Jv0+d1
73fdW3DwixRU3wOrzTzh5oHqdQO9aBGUrE1mbl+331fneJG4UDnHfmSOswdUuaUr
v/FpHXDxGNyne1cjhyHcXMo/CBGm/NBUJ00A4lufTSRTsSXFLlSOtqqhv3dnoYIH
ODMRqCz4SzXgSzoNbs2AIVPNFFMr9UvEDhWTL4P+EHzwdo8y/9RiNeTLSPjBAKvH
aEVfJBMPgjVlGrjwwlqyi2dka74+18VB++1VjnUGZQvtIp55aNQR471lCEU+9171
Zxyhl/ppdxEc76FEXCXmMAxB0anr4D2DKrbCGWj11ucXrgn6mIlYbPiDDp17Dfuq
2yrpvj07aN2sUC1ItTOCD0viaDjQdQcS1vaMfqTW18VyFNmiVJEkBhAmMMyHzY5o
DMPks5Lx3oCQbp3Hr3BLVzMtvdAgyfHg3WY48xmdDm75bxtJt239eoh0FEmSn5Fi
ruBYW8baCIagrN4A7WP5rCOSiJCirMYFkklSpbBCWpQgvPodhzC29kXoztPj1G/w
A1i+6dip1tfCWBx9U8CphcX+NpMS7nvRXhx4lkYnj4zY3myrLigPndeaQA9F5k4/
wAL4S3xPKpz61ghTBflR+NutABwZaQguQ0aGGYZr7NyTNTTM92UTc5I+4hFQ2o3O
YRmf4suXly7sd1wiWzYXADdTSsfVv/vB0J7TEj8sZw3BhMGacHagA3rnzHFkANlF
8lzp5JK5g+Ot5VejY5kyDMcUg09MO/skORcrp3zSnlE=
`pragma protect end_protected
