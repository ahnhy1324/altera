// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
UNnBJZVFDJi42GPmqYebbbw7QLWQoLh2RWp8wAbd5UbRdFK4xPNb8KaYT+FmDX4hTlC89CI5pVy8
/KQ0Q+z20IOctGM0V+VxRYOQo9A1XLFj/PphuPjm3m88ExWt2k6GajxtUSa1DueajOqzl+YdoEM9
sgLvxHbjL2gZk1qATd/S3GQtnA2eCxQAEXAwvbXO1b1syZpBcnpAkCe+onstAtfKkjLzhdcPv239
JbW+rHolDWwIEUTJ/neZau5dk7fkqPabcLuytTYHS2f4u8v23Ufr4fwvczgQ2xz3tFoqB1yTTDxJ
4IFhlai2Oa8ZYB4bhncoxOx2r3wHI8HvT9YVyQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
yVv2//p5TQO6J91He4mihCrtOW1ydzeUgodQDhth6nRxr+CMKIDozPJlwLnSIzVc61Qnp/g/DwUE
WH/gZ/Tqs2SuRey+UwjRPQMnlNRU/Ue1w76o+hf9i+ysOXY0OkbC5kEyXxJEj+LEMhu+d+4NmtmF
UVO/CdAj4oixwSykmku9AH39N/2bEFuaRZjpL3Ter75OvdNnFPvk7tUbyxNZKFkqYHUL1duzHlLg
GkgYdusiGcIt1l3ixTDR5UR6Rq7SEe1gZxUZcIP92/Yhe+PcxqyroJbaJ87MWSiP7Tb1slnZc/Kh
4GiDqY2vJyPrrsJ8IZ3PqRCLVV4cY10ScKGFlMRWFQtFUddNZlXTyKT/42OL+GhB5VNemLuW/Yf6
Yn45sg4eCCilAEPUAXCMLshjeVhRvTWm2kQ+yuPrUees7fA+7WoQyNVfE5p+zEBxmjV3miO1dQuc
M9E+UZe0+VYimYSJQzM+SlfMED0nzfrp0nMqVBv0YtS3UX9oCRTCMcLjI+kQMeM4L8J9WFJvlxMW
juzjq9Dy+clGgQk2oS3dSUTyhC5Etr8W91jg6liUPx0NCWl0dHLQH6aSOcoL9sACw66mM+a5yVz/
zClvXFfYoZ9GcpXe5v0zMs0X0Q63zBgHgll7rQ3NxauTd7P3cfRLNpE1uiT+EYg1C8L2JfK/1jPU
3v2vHQcHvzUHU+rZxkw/kwle0JQ+K0Hff+5HZXhWnI/uftVArems0mU09fRyb+DzENbpZ2RTY9dD
YRQRaJ44tpnXEqW2YJevNxcIUVPD/ji4rsj9oKqRiXEkLTk1nRyZJKMjtoIfR0ASMY5cfFxvpX4z
3aWd7iW2oSP6nDq/JANcoikEtL8bfV8LOz4mKSaBYoC2Xx/vrvzjsH/uSQMyFqfpmxdd2okWCIrg
Sd5uSL13jkMy3SttX6w8YF7C0WOToRGV2SMDeGu9JJBtfBUAevRfuImiLL40mz+jN7UPeUdlTKGY
HpaMmM+26OmXYYTQs4jbSlf/Oktxct7SxfzSnMWSv8yngVB6+ZnnolMbcDb7nJliPhufXTqWk0vE
xtgjTAGuV3ay0nRgDMfRaK2bV3tM0EmPB1TyASK5tdDK2Znu+jSgj9oDvWUaRb/VBdb/qqry3DA/
th4QSuSjEhr6uVaWFEPLsZcoCcWK+NgiP11lChijGZyDF4UeoKoeEDOTqwuAxScWAbNoeuJaHuQ8
z6Ul7jYKk20aWIA8H/1xGAfU+kylLN79LGuAIHUt03dHEUk8PKKzTQYmwFj+SPvd0I0uyH/K+n2T
XMNwbRjOc837QWbfvqf3vX/Uu9cF0jRLqzTKj/mELAfBWfsKUELMXcB3sqjupsob1P/CrZPumPIC
Bo2cs4A8oIY+IagK1Mql8yOPLVuxwTnXs2XoWy1BxC6z//wNDiiQcepQNI1S+0ChdrPqzzmK+QO0
gxf8UUbMpZCueVKAv77DWTV5eAji/ASlo452j+A8XmbXGqdVFaZ5zy2kB7HyGOW53s571DVRRvxW
RZy3QQHQLRZYrGt7u1r/v6wxmJKqbjQDa0Rf0wlwbXhjyOnTRDafToAKDrlOeF5b1GLcQYbjV9np
+BDHjjJB4edpeI0ypTtvOY6o+iotnF23Jrvyj2+P/GNutQFcjP81/vxRfoWQo7EVJbmMVMmcigmg
GtARJ74yUz3o/c+R3d0M8TPl/TsTwuN7kes1SJ2lN3sxIqhwXAvbxpKigfD84RXcwifFNKraKZMp
+PFUK1AK5h4QflhJ3DVLxutTmnF0tWV8maJyB9/QOnNSyi6MSUPnhafMBGFcb3V+uSlD5582a2ij
eGHO8bVSt2VNB3q8NdC3Tu7OWGmt0tVQ05d0DjhNKhdP6DaZiuZVd/Vx1Ce9z/EgrtM5iMpz0GyG
GrQPnsKZxlc69Wu7oBrjm27WhOe32haFfVbBt8QOWZ94wQnXe8nvYj5a0CsqHpGfkC2yC+VuYD1n
odL9CPM983wzYnitnH72FLUeOIIKl0pzeYpaSvv0bTsut4/SBeN2WQp6Q2iQNRI/Ea3qnWl0oYLO
Do232pnwZqgfTnd9quOHCEJsoqsNyId/ZvGJ7ytEJRuDuI9inCK8mvJ+01Mp3IhwE4UtXBvJyDwB
HxtVTMwwBoCKklC11m+U/cLvxFmASw+ZMEjHUBzAYqNSx32mCnK2gujkjq1ZIS0fWREU/a9KtUcz
ODvEKkIASo7dkiLMe5Zw+KjdXsk5FXbwxwbaF0oH7/rO4rURS/xPfl4DbTVIw+4BOS9LYdfU7mFR
g6jTVHnl3QbcNgR2rQpZbEjvOXbjdhIBW9ES1hXXxE6C5gxJbQ3pNRYDINcDiun4zxQQAMoDl/0Q
PzVCrFUKI97Ov0iyWLFfC2x54dH6p7uRJQazsfdY82FfZ+GFBfAt+Ag/rxyEfoRkChtsLNsje3kh
Twl8U42XjgxL3Llzf+U5uR/+Sr1dnWgyX4n0TBjdR/nH8wNWuC63TXSt/naNFlEkUW6qqH+p1oyH
pYzoIRVlWQto83qwyPNO2Deh5C3Ic/gTdknz90SSRu1HbHb0hoZ2BTn6taKVWTTcERzcMNLquLXQ
eecUIZ9b6bynqnXNVxtstW5kqmynzhiLDqDgOmp4U2YjKWFBJWzx69k/dcIOV47pSpRZxXCvr2/G
BnPv1Jyh1xfarAY6hLpZsO6ydH783I14qZE5WwOJQ2fTDi88Dv670wjdeAA0Ez+3H/PucvTBoGvG
TRgh0GZ4X6SVqjYIt9fcaO9jfPNri3EvgwJ0r01jk581cgeewwUV0WaTl6jV0/fiPMMU+IQyl42l
HmMnuvUYw3mL2Ia93/io470yuMoE5jkY1ZSvpBX+wPXnGOpm99kMdI7aiGiN7QMfR2IyriVP9NeI
VnDnEu8SPRRd+zB14/i0Ujna4qnK/x1+yusIB0eF/FPsyvDXuCKzYzi1/z132741h9dvLzpFJR9k
ujDEGE7ZeKSOHfVn1f+IE7JL5NkRpKYAJ/Rjlm7/iBtGaF1PMY6/7pmt3a91TQECit1uDSO68L9a
0VZ2Ccj6dxornvJ8gtiT8RRe3vwV97mpeNStAdsWD1GQrLTfO8C42E2mDMcTba00UiuYfkVRcBv5
zDAnDGJ4wMA9muVgVCFLJOBGKfSyCzSBm713zrYq8mucfkjM1PUxQ7GiQ1uj4DVyppMCd/0ujMCE
Kgau5OdW6Y3QlrjctF+vRUrwsiZOGTiWxxE+piHa5d5oi3czvMGpE0WIT4g+T5z3q7Rf8/jGlVJG
eJJ8gYzKC/4uzo+BzHbGX7hxHKJ3MAGJeU7m7SNrMfR22pvbPF8Re++h699pxsYvie04TmLSrj9Z
58t/S+KiBYOgObVZTVW42+x2ArHBuUxkMHw9wQvGkKjriajC56mVIT0oYjj8SZNO3gVsQAHh1D/9
SKfbSlZ253f0px09+zMW9LtKADoEBqqsJBLEhb+as3N/aXzDFWfIANAK39OmnrH51e19qW2he4+6
EdDhP+DBB9NphZ5CdW4jVGmavKI2QZ6bMJz9W7d0FSm2VZ+dvTfVe8tksJAbyLQHCfabKglOBhqj
KDxlgCoqlTW2inuEhKLL9NTe5VoFgFGkUaMtaNm8aNX3HCuBqcAnN7MrT4xf5qm/TMJwTbk4FEP+
oPuaaIM9iwCi0h3TAe5GOzt8WnGo4N/ejcs8olsLWOtiFL290fL4hIFLuFSLjhc2r6XqgkY5ExQV
6HFR+Je0NcWqjIdVm+Uv/IgmmsWspMdBQci4wuhyX5l3FQzmmaqLhMW7aEvwfzb9QAq3wa//ZyNa
Br/0uPt2wbAEDu5pTqp07d0886T/Nr6eKa7fBeuNFD/daMIMaZ8ccPBs4zs5U53MAL53+TBAhecR
dj79voQtSAoD3td9cNSMNIDB3PGpG2H29Q7trKDfMYp3TSJSQbTWBIaIwjwTX/Zj5niyralUbXgS
ym4kmHbg0F8ECth22t40aLtz39p4i+atrI/bLACR25wopIyEz3WRcRPVGWBneRuVKXfwaohcdiVF
raoQjg87YRWA6OpWvWm/KcbdBEQHxMXbShY6XvmG9zshkrf5a/VHysr0syBuzSyllM6YMNZTWAJD
iihTvL07TYPqHNHa4iCfs7X/p5eZsPn/etHO+M3JKY7bKIDD4hw/pQX1f1A0niR1hv9UFynFvARm
5G7sAdc1DfyxBOEN1z/KWKQuaVhELK3zXptLqd2bLH9viEvqCqYT0VeZiuofaSOz9M7JWwUEdx2N
xkm+mQUJS55oITpdlBFlW8J1EYaS6RIjGUHaO+yzV5aWY1uk3oR+21Apij3Cyz2Wi5RKGGTYR3aD
JenfJPP+ViIGMnGAh8KUZyi8qP67e3zECqzhs6dz78M8+CNTVu3ivsu+O8C5YPAuJ/5KHLdPDS9j
/cPnrQA5OQL5FV2vNtT/Aiwrb1ebTubem+Yc/WgmR879lXRf/zGYzhhU1rff5hTaceVpBVd4Y9/H
8ty7yhgOYfxyFezoEjC/YRUZixgod1GCXkp16tBRk9fGP85auXrf1MXH4zF0PM6lUoQi3NfZqpFE
kxo/1dkEWQl9HG6EiOS5wRYfqvIdD1bn5DRIDtzH3T5SqSU74c20DxmHRs9lLsebtG/7+K5bTzJE
e8yvuMIopl8w9bNZt+xVhwgHvLeWEZpEhLM85d6uDqS0O98tl0nswqnwR6hrSuj5XQI+jh9w6/Y5
skHTJSAhjLSu05h/yvUu/ZmvXMBFAdJDDDs3rG7i97TIgM5g2DpHyu/402vsAah9Av3mYseMXpFH
tnfKldH/o+3s3sc9dmDWMHHTTpBPr4+Pj0lDSFW7RzWzfzGS/Rve67XiAjxmJe8DrEcIeGrq+nV9
9TkOUE8UAWRidsRIL31qzrMKmXOX8q5CAa5z73smJLPDKzTD8m8yKCm/2ApEDVqL4LWVcH1/iSWu
cHmURHPisLTJyTzC2QGDzf08b+dcnmNdmZ+dnvLS7b6erUlnAv+1Xe5vxNn6DkBzQde7rHLMLoAc
tkXS+Uodug6GZI1lQafDld5mYHQN8CBkvmOtUuOHmfMS2z/qqvoqGHX18yhXCxKz9wwJdrwKOndK
sfnp+Y0826+u13+ggVgUvcuUm1rBQSIW0ukYzdlqd8rvMWa9vtJuJFZX5i3rvv9sTv0SQci5+l27
cEzC/Qi+R2P8YmwhGkH6ueijaK9u6HFdkEk6KSmWn/KVyzEJ5vD4zrbclRJIrz5piBhpxK+1pv49
Oggpg2qbOcRWqOXpEKDWIijTGi4rHHtIKN5Ss5/zcrTLctz4ObwSVuBZxYEhi7pKVBRTcxtwVn0b
ScdJ7CsS7fsDTvwBtx/3JEMw6IqQ5DRJ+eEN7a0F4TbYHmKhrAm11Rg6cRxhU+8ePJ6fRSKw9iO6
ID0VN+XhPzkXhnM/R687lmQQJNPhNaaA1NVUJI79jetc/n9WuNu+GCU2weNLkIXFApHTqhYbXT6a
wFQOkQ692+V1/ijhLOh+S8BI194UllAKAXuv0qCfe3X7dUYj4XGiv7AyLAapVJbBzysPMNvWyF1v
fEiYdxd4PbhGlXdU0xm1QQBp0RSqQWHy0mKwLjvI9IdtXycFeZYagPwHRlYjkTIB25qW7OL6XPj0
1UdFuLnb89Zj4ggmDTbA9NKrNrfWVAVIy3oRakasxoG0RZXKLs9VVwKHsfTImGhkiAPf3SWWoTj9
COZCfG/hMsflmD0CdlwsnWfs6WQhOeTYqOVkOdnsEoU61LGlROzoY+7mBp+DNFjjZ3vZ0D7AtWPJ
v/dk59lsRCVY/n0IvEDl5pPHAxWAXD8IiqSJoKDUBaPbMW8cUb647oR8MVpvO0qwXtIdZtLDURNB
SylP6pPKbXI1IT0dsB7kQsjmybBfkiLcA6DMyebw3RDL4Sfoy/Xp8TlD0Un2coGUFvmev4NDS5LW
azKTa0KrI1vousnyFvobamWE+LZKIOA3AE6/TwKtAYkHUgfWuCD8/DNXSvrAY/RTa76GrdYjZvjm
4oHYHIsXlVPQlicXrWwMymu7jHj2Ou62mVEv+YB7oegBrspIMvzdgd3EpQNQwGntzyY6fWeUibuV
gJdeRRrW4jKSQT7HukZ2vJI/TZQCvf/sMIkbqcRvz1DBYow2LCpbUQY/QN4C4o72xdQ+hXzNpdMo
5L+M2PrLpXyyxwQ1ut/tY9NucOj3TrcZEgZQnIgFAKY520oOYZQNUiZTAAOP0O8Ca2uSTFH3pzP9
dsIkb82bfcnzoIv1TDne5nPFSmQOwMBvLnmjSJ6LG3ltPV0m/ub3HQlyg721iIt3sXdwaZSUDFxb
Iwsy6zlQKug2qWwFzV9K9AjJq7VNW0MXFp/UqAyg2FumkO8h3/W24jce/wMIDykYJyp/PMMzGmaY
/xMvJplVcBCheAxjjQNqN4eN5ErSoiOBzvutCa4Z9Yz4GLCjRcZSHveSaEjYIFXQ9fbCYHfOxasb
Pe1heYHMpZhW20gTxobYGzZWqNJckzStGCWrKQCbp+MkCzwjH5lkyZOK5nnftDkMyhx8Pk3vZsSY
DKILx9XBc9uA+JhJZnNMyb2VSxX7a3lqRnIY5jg1pbxahLh3gBdaGxbixbsql0RfxFy7OjC1kad2
7hqJN79ugHpgTHVJvC60Q9XXZuVnKcxUbHjxRPuTUji7AE/DipKSIfziLP6A9c8WIGD/pCfbbC7k
+1f4Z0e8fy8HeB7qJ8y+UfXJZxDgPJ6UglkYETrboK5+Mog+pRgA1tqLF8HjAFAfthabjPFVZMv4
e7eM/OErLrJQ6CFjSBcDliPP9QAL0Vb10pENmPWgDa1kkJyyvC3ZjFAIwxXHx7eQjfHe5EwRWHvt
qHaiHKRn/SKUNZ1iTCFHgVd18/u0O1JK9YxG9IzmccKxLQU5naZrroFQ9xDyPR9Y4HXoBICIVTaY
a2AqX2FiBc1qwaR1EFRkZ8KXWhHf8006NStj23VhsDfxeW1wMj6+MuzwHvhdboBO5K8R1U4t3AK4
QvdU5zyoZuXHL2zBs0vmd9brBs/T+nPRkIqxUFitI8P+Q/Vh/CV+qRjO9U+jl3mAQBeu77OEM+YX
c6m6QVm48BQOa6p6cve9Eqh26C/mExsFpdO2sgYS9YAi4Wq10L7e8QzC8O+7iT1+CFhGpyF48T/G
0ayfWG89ja/Tu6X90AHX2oNaC0doV5RdDtOmQz+nHmzuDuK3WZzMaE/jdo6LSl9ZTGqd0KpDRJee
7RBKM7yPwWaC8aSiI8ZnmWQKs7G6YYJOMqwFMzLPpjchYPE/V4kRStQone9bdaA+OyBBKhvTqvIP
GRRjwgOEn9zJOuizPxXBALgmgw3ErQVBO2+ZFsrsWYEBmGPaLGeDdGBRc3PdBoOh0LirGoOzeVMQ
uSYB2hcFOcJZzaewS/F8WYQ/gaOo19ORN3rhwTXiCoTsqzybU100lu6ICf6KpxxMckgQtGFutRFA
MbmFXeYBjd08GO6cS7Mg92gZSKJuGVBJnQjqL+e72IgqgP4GmRZK8kFruAWy55KTyCLBA60VuLHJ
fxJKOcmMA5vFZH1CVyWe9B7PfKty5oGjmp/+FZRYvCZI2QzsfzrgYDCFF6nhbyqGLUny/zmW/DkJ
1mwHiu4MGBU2J5VLDycjRuAjrPXey0U+vU5Lejl8KWU+AgMGJ4PgcVwFEHHT9dPLBtJw89hIuarh
kY/t/wB1WRPRdGyiqVCt9dQjIRsIjT8Zs9iubK6pdcs+scvzIMYdUZmcMVF02f9/VQVev6xgRylt
RGclhUxcN0PDGdx4RW0sUrwJwrbYcTmkbrXyRhrr4OSIWPq6VQNGwqr1yv6e0n0oAvi+mbZiJnhf
rb4kjf5FyBp0e/TP0JJ4trQavDMXt2lq5gZWsuCuIHqt1HHEKGMVykq9lz7oqOTEAj6zjQ244u1r
3BLZl+/wfGxB1uZNySAlTaPUpW4VY7GgTC9QnEXd+jj6vfItTw1Vx7sWm5ZtBlQ8dF6FfzGST0q9
ilZUU54DGYr/tCIT93vv4AitP73wX7urafr7WMSFHh4bHvq/zviM2E3AgBkDjdrrhMTD9sF299GQ
Ph6ASL6q9apYuIsZch6M3sDRyN6RwgU31aD6gh14zeV0+51T3LmXHUNwSlfotNBJkQJGBVAcT3td
28ay6up32OYaEpBc1w==
`pragma protect end_protected
