// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:45 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
s/dVtgdHPTYIsusxDUyZL3B20syIwNZ36HBmWKKeVy9Vi2ikGykL5I4nFbu5Vc/F
fzgrsdO+NYkthU8uhSPKX7blh1LzXZvY9adES0q/g/rYpUmdtNpg40+MecWrK10a
ZNPzYjA6p2QoJb+4edcEpkDdz7O9clMgzs5n/hVl+Nw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10544)
51QBBvyWMXJbLhmJk3K/db6wVKFCVBZyKL74/byFHFqTAizULYYv/R6MQ8y2G4jz
mzBH6Bn6LuzZpTUX63Nrd1HGmiXghhDyhZf2f1opw2AouHI4XBB0iacJmnAnoWn5
UVl9fuaudpX3BCgxNHI5dDNcUdsg4bbr9dUow4qBfA8UCbH/hdd8S2llIqtHfG88
zmuipgnsqu1qeQOe0DJHJl0okf82vB5q5dWx+TfI+7/sJrUggPILHKuXrpGRdCIX
IZLdCuv6K9AwULxpR+jJZy59tguhxL8/W4224zMPtDjMUGUWlAHQVgz9UjZqDABd
I+3RHuzLR804zIgSYZwzkEYYKsSfe4Ih2crmBug4Urc6wk8Qm46maUzzEJG7Lc85
adQUvus5sT/FzPPDqEkQ1EBAgsuQ3VYTPgNwMSWoMsx+LyMzCl4EDtpeSFaEnS7f
h/2MN+iQdvkagB6DeJ9ldzlLUEhIoiop+ITcyURsNULG47W5hxYqcBm7sSb1l4ln
DF/ILAQUQvVcIBWDdpd1YnKGHUqOUU7gk7wVV68PMOYyp54LJg9EFpc+Iozczv0D
ubli4dy4tkybXJClPXZ3tuyuCfW2e6xRNT2oj/nPUQi15zA5bb0/f6ZWUvO7gJ2i
Xr6DWrEkA8qqYxws4s0h/hMGASlbf1NCL/g0rq0xw6jDHcCzwKGAYRrt0ZxaKYSv
X+oDLs9iF/WZiJyFsOW/7ui5ozE2yi1cZzfkNVWnHKG5hk2kYvAXdpseUtBArugM
UXgZbX1YPsAhLg9tOhozqWwYNHk6KoBtVqDqWc4qS6rEzB2r+6oUBVGNfgRJ0fom
xL+6uZmq2fIjAwrmWEIz8/f3ufciSb76VAFv2r+8TEvpN9Uurtn1O1PV5DN6ig77
Pwy2c/weL9ypL4WrBt8mx5QjZYW16iGyQmxgwX35afrVRoFxugVDl3+pyqAHAdi5
thfIgNe6vZpGqI/OVOU6DieXq2Z3ljrosk8kSd1iT78JwsIfDEu18e3lMKGXmln+
zdhTkgIEc7rmt3oubKHZAzI2GAz+BM5GW0rfTdh4mensiK3twKX809j3Z7erZP/w
GrOXgZ76ITLnKB8lofSPQp6Ce+zNs5OY3YYxWvWiUWN5h6bSw4UkHfl29oR8eYo1
IuxFy1x5vnqq99MSFksAlnw8TARdsQRZr6162UXKVIDLfWSU27VE4LPsZFBp9Xeb
8PvvbAyQfTNSWeFCUrRy61Tgj8hnVsGmNy1sY47ZDq74cqcmebZojhIwd6an9dMa
fTyK6DnQHACkySH9GzY16tiTRWCmU4Rntvfv/94Q+6qnRmm4aatkImh4O6eh7EJv
oKGS3UgLfcQ+Dx1ceDBucsg/9Izl5X+socjN/1DAQeN6hRgWQKdK38j/0PcC5z2x
bDxl+FmGjOBrddemg2LGpXZjgERDTmmmJjlfih39ckP9dSBpvBTZgUXrzgyHYMWm
sA5oYO7+r0acZYImTs6e/dZ/ccDI0/R6pn5LVbHtTOX7x26k0sP+JbuI4mxeXInW
YfRc4N+QlDXQKaZetUAfEZcRdBsaeganWG2g2xkK7KL9sRwBhuPADh2ATm9vJD2S
Elm6RN8YC41aPbLxo1Gnd1VgsisCNmuuPedTz1dhl44zCZuD8jpgZ8VI63uOY55k
yvRI2nLFRFFCDrypUbPoSFOrAywcr3bJzQ2xLCHcdia80G8i54m8NSBn7mkPnRoE
2Hgd1ggN8xJ0yhybGII6m0iM6cZQrAuGRaoWJCSrQ+Sjdq693rNo8ls2zsoSGIDp
t5XHV7aeCcN6xQ+SSWb/9DYM94t3iXTHG3D9fh6jq/OmZjpVeySGVRCnIfxY2vyc
pxWKgISpZKEFE+rO1pCMGOrFGn0/lA+ufxnD8+X+AcsjpzWOVa8bexZsRD98a5DI
En8C84MmpA3qUdEO5irjj8s1yNHbUxjZPRZRHKzi2uvKcfuWiW8aw8Z7QOPBDVej
9XA6g1RskWy+H+OnQLEDteMWrtU8j+uPVrcJmG1kbRI6ivUlFOnnMpDAy2wynKvq
DKfGI/xpsaAs+fcCg72aojC9DY8nFSCmNb2jE5vxv9sJ+zne7SsR39CmXe0qKYcB
dLVM8X6tZQeBG/yE13wScVawy10hkHv/rp3Odvk7kMiL8iBZsIHztjinaxm4w7i1
cV1eO4hrFjl7UZ5lJAriAuPMyJ9AdxsZLNyVsZBAqnT9Fd088uZ+xjD/fuaM9ve2
vZBhKHICne+Hn3j2XN5NtRFb5K6/KdyOdzgdQ5t4dtJglFhVFqF6L0aS7KW9a4o/
9u9r0lJzsH1DNyiizPN2AEjIW9zrznIFMluZoAno2gVqL4U+/YyZaXc+SmpiZZif
VcimLMQod2C74t75rxz05966GfdeWRPXIGdKXa5a/8blvAfAesUelGD0ubQsTena
lkNvUZbo+64cGdc4DgNsI/ut+ugS49GOP2o4EHxLS97jCMQkg/BrWkgaJb0cQmG5
Y/zXeW8uJyNipLix+2FdnCCcyKosHHwA5WmrnWbEwkurPcz0QGbn0NQn8cBUBaBc
IXGTJttR1w/JGpQj3EU+BK2qTQu7XJADHq7HKIPCmRi4ZoBUnF1D0/FCo6A4S0c0
u+dTFwoJdnb3DP2ulw2aXxg9NliNS549A8R+girCn4LxVgCrQaocyY8QhJ0RQYh9
c59qFtzMZVa5AwzwR+TuALuHd8v5NZoBBsiTVA0fX/NsJyYU16IzK6abeWcWuJ5c
iMrExHyeclF0ZE1jjZw2uikkuHCEQq/w+UbkUWnSqIOtScuHKyItdPjkst15KJh0
yFsNcTXtVCZJIjgNJNExByDPEBvkb2c4C3NlCu7oc/3OssJivKWy16cLZrr8Hw9K
Xz1IkvhBaoVrdV5KCx0AbLus3+uHgrvVQ85BWKsKzxERbnPbt+Vwu2OxUY7rgB/N
2OcdWCnFwASLyd3ZQnYr9MxZxOouoGWH6c99/nEWuaJJhdh7KvAbvFv0M0rqyg7R
j1hPH4c/Dac87zGk5HXCnZD7U2f91rmX3Nw02HdFYQPL0Zn1/I2fSMBWmhhtPlo8
gHkEj3mH7pj3x/mdAKt24w/MqfpfcabzW7as6VDj5M/7Unr+3elnpripe/Rbkrt8
ycxH4Eu+JyVblZvqr2ZcRBhcakVxe7puFkkjHfxExmxX3tLFkQ4yFd1l00RGVLz4
r+qsmfJHd4zZAB/dcmxDuQB1RZyvGAux+0AIegZDiUcbVvYFL5RuPiXYA0+ChJAB
AfFvAq/k1RF61U0ctiqnonfy6sxNGVYMRUJrUocgtngZ8Jv+23/mrjjWo7k2ODsH
P4YMG3f2uw2g+hCB2297OYQLyY7yGjpx0gRxsy8m7U52tnH2hzN32RLVO8oXMUcy
hp0NgV+4GCIQ4UOl9wlegF5iGeGK83A+TJibvTM1p9Dz1lnfXbrR4THGKslJLjm4
woh6hKkuVDReYpdUyJmzSvqiW4+LMhPrNaYbMg8sh69W97v8sGVn5J3LsLn0GmJb
hDPpexFAiIdEdC/dSnrSz7vz3PB+52UTx7X0D1Tvkl+TQTaAbVS3NwWjFXyDszEr
/op7Ju3Auyf9Pm8zSzEqfVMKneCC/efRSBk2CWlPCV0VrSv1TVTdz1nwdjx8m3oZ
2+98XHvaysGy4P1Vft70/QEi2SthURM3axb75aVp+nvduYcNqM2GvwUcamHj8u8l
KBnMzYSdxL16BOCVEMojjEwLXIdXHtFowDfWEOjPcjPvA10+xZ3vz5//Qzl/UtX2
SIoR6kyRUWC9LVY4sMsaSt+Zw82pa8DJzARBWdtT8hpQgRauu7Oz9WBXxUFO4ATi
sDxLwuZx8z6dsafkaneE+htYS6c4MJGir6VH/sSiu5sSzFjKXaT9pUVrylnbaq98
cVKt2aVWG5tL8QzCIz/xUbfOT9U7QCCek3sOQ0rTxXivxTUS2vIvShBU96m3jTUH
HL1TQIzdO7L99bpfvgRoSqgrtGGtcevneaPFnlwma1i7I/5P7NOY8hmlJu4PB7CS
ihJM8y+OEh/uaqbmyXfwIeE8YbXNrfTpaywmeuVBC39StKT4Y40J+S39GMNxCaqV
P3Abm0qwAJzdD6H9IT9jFF5VEbAGu5nMEZK/gHP+eMnK9atJbtMH5VoAPwQcYMfx
WuGDROd2SV1PPd4ijt4gQ4zDofP+aJh5CRbXHzpvM9vfU6AKLjFh65Z3kbT3ye6K
UMkafCfV2mqcbc97miU6Bm9PazXr8evVw3pKJ7zF+4yuxACva+UGdHIkV6cOqI7V
YsgX6Dwa7syfX1PzfnlfOrJ85nAu1Nu/92BB4Gy16ZjOcJjkeTt5C2cdWn2ZsCz6
o8pDFQnWAMD31RYnQS1cZds9GjIE188yX6KenqlozCJY41xHEsqUnfaYuUpIFl+D
MFsHrtnbcBq0gvR7+Y3Eo5rrCW7txB1sgQ5tWc5sbO9kz/xNkEypcOLL6IFlxuFR
rZcQDSj+5GNIA0344pMipRhGfjhHR/vWiOvxu0i2IEkmqTHix61VHLQ4nlBqV1Ev
JmbozhFHYiSxQFOMhxu7326UtXnuQTa88Vf5DlrYZ7UNLKflh/psUK3573k9YB6q
1v2XHcK7YvuyaTQ2S7irO3P+v21oQPUKznzOW7NayUMWcEof27vS2xKWCtYxxPhl
4CTILYe56dXm20U8uo+65/r5UHAE5UW6g0Jb+mYUfDnUWoBHYPcO3WYfB73TnZOG
H3ITqLxFuxZxW49zg1qQwFTu0bczqvwF01lMPFNq3Hbo2qVyL5YoY87N1o95MwOM
zpH/eGe+sP8Wzlobswg3nsshRH4M+yaBYdMc4hdc5ma2Kj7HSPzmjKZglkmwxwjE
e5VxOKnykZe5wMOJuFjKcc7ybUb0UZB5E5/I/V6pWyn+gfL8rbFLYZux423vkOz6
s5JSY010DIb9PxeaJb2IEzS5Pwnx1MsZOBjy78FTmQ0iw0LUubX7fO7uUtE39IMK
9Mzh0LQp9bprwgIVCKW4rLowvfyuP6t7fVM/9WN7zRRqhF82autTfvIT6LZRBejW
NIsWSndLvaN2j67kBiG1tMYNXRLtyYzL3khkS7XrGMTOD5wFvfZczs1mvFrKFJKD
zPGKk3Wk5X4wHWKEcI/LchczjWoBHmCWSIBQIgvwiub7tAlVE9YWfbwZgANCR+Js
EDJNSXnXE+WcZTk/p97daC2QaLrRbIQi3IfJixGk/rwynBzbjo8vVFy/wAQIWg76
Uojyjytbt91GCMP/gR7qFbUpa//+ZXAE4tP3ztAMwj+RiQF52323FgAJuJKpjRNr
9wq5nHiT/pxFqySNxBU5JeODVN06EfMy7iRbv1B9KcdgkbmhtVwNGYx5XOxhS1Ic
ugE6Ajoh8N9nHTb5hPSMtk53tz0RgXw7RMpmDv53aqgcEsUqYLDUXgOcb3e+kg9J
hzibh1XAWo0rqcgx8UnX3E6U+atro2gmQfoL0rbaklf5sLisLSXJGkly1x690Z2I
Rru8YDd2J2XGHctvqcZG5wnEeDR5ZQydvZoBEVcQMupvvyrrFwdHr6GOypeL4Jge
sIsecdb9AlTMr4JUGmVVhNLwUFD2k27Ul5hYOFvbbqkSrJP+Wtub9WOgKHw6JVMF
7dzAxuLpDurIzgi8WJBrfLRWYpvVpWilALr4bIIG0rSh0hIw53NQQMnHyc5Dnum1
uGcKWMrmLnF5XFh6aXtvBz2NeeCWvi/9TVJU2/h49Zz6fAcaJ6XFwBKMOnoizcY6
WbcFaIv7tpEI2Rlg6nia64/CflBVyOM0hv/KDuXWYMcroDNxPOt7ahXlde4un/0w
oS+/tyViT8RBYARCXGXx0/+IdzuRazttkRXDc1vJ3OmCz/yHJu2UlDMwUJxxjMNF
APZSuBs0cKOm59reNoQg/NDH+0MLtWapx9Lz6ezYU1iZKLeNjX3+SukLF/NzfV4K
TOkhhHB4sbfX2Pvy3unNYz35TumsFZAMRMpDt1FtP0m28UKbD+FghAlNC1JHgFx8
q6bv4ulFTwaFxOOHiFFIqyH+xyVFmumEqy1WfwRr1/SjRkLs13UoW836PQS5Z9s4
z4NGeVaNantuz0Cd+YppY3ihngknexw4suDWyq4QTiVYME7BDYZc0oQdfy3DrzL2
AcNrm4G+cbmB91P7Vm4TtQZRA4mQqXfPX6q7h8bKKITjzVE3NBDANoyLdf8pFppu
TDnXre75PRUeX0ZXyyz9a3DJgu14d/SkaaUx01lz77z9uA/BRQO/XOMle62bT6/a
ONUcnpYSrFh7Bi1M1CGQdaJwvR1jgScoLu15IU2yFWeEM0X2WXlnPBdzkRsUTBoE
z0xIJAwZk7eXpvbIBPRkl+9IdmTQ0beTjD2wo+oi5tPNDu6kG0Kgoxd9AurI831o
mz2NDC5RBiROQxUwyZ/pKBdwekD3h0iFvg/+UfubD+/8eWpH+e2cp+OxNOSohYIm
IvPlG1CY3Amnwyw7xmERV4+3IuIXELlK3IyxsXhrphY3hVancpRAHEpdptKOW3w4
oPmVDpPS55rNj+JWg97a+V35VzgsEDYJ5m8agNKSbZpHbHhewyC5p6NWe+A8i482
3nayPz6AVmrSGudpMEr7MeYydYDnwDYFb6kZ+X33b+9801u4DXPhOSN/h+6wR2iQ
YgsZ7yZADSh7Q8GIoDngli/23YSgwZED4hn0yTSVDfXggLZYuIO5GqKwa9yNHozG
iKVLyLmwlZIv8dAexvQQvQnYrs7Mo/q0y0OA1wwqyaZMhVAaMEQccKbnSg/kckpE
UDh96dLfanhiV0Fy/tI1cRJhfyihRpG8lyp6uzf7HRWADNHxqg9YLH1/6zewbopq
rdqpXN3KBQlhsqWcJpJfjP9U3dl837elENfKnlillDNGuQ4ZZRaL0JYRNPrvW4BP
oJxk8AoqxZ3nVQgX6XgnxZq0HRKEg2tH6FpbalckXziudtW3S3IzZQlb5+uxd+Ay
xHyLJXYuQ0cp+p2hpH1t9Nr3CdllJ7Jo3r3j1HxMCGpELW6TebEPy4cqA0aqDzq/
M+jIBBRitpPYvI71ZwgNNqp7WzyvnCrwcgvwaYaopqj3WX8DTMzoMkni85pILh6B
OOspsEJzqQWQmtU0QB43YW7maktA1z4hfupiklX5ANcOJyyc2b67yCm0Ou/Hkrve
Ii1STTSL4FY/xErvnp8HC/qdy0Tj2S+CW3SFhflVJYJgNahzJWBEz465W/cYSuEn
6D3zDuI1unKjMK4cGhooGMX67ghtpAz+Ntdd8AzLSuyBemzR0IFadjmCInk9Knah
D9GNPJESLc404g2Kc86sPjUY1lZY75sEDNQvgSFqDu1hsvdhGWiCYcb5F481pEhI
26ddzATn08/TurzdEvIN3zB1G4dYnjmRJqIHOpMcIFrfcJiUo2KkkhkgnPMBYu+C
f4w6cBBVM5nHZ1bmYd4tiJOkKqiFq47n5yxzpL6PrALUzGFw2u7cQF4vPT3EEOTU
Eyx0puZ4nsGP5hdwKOJ8Kzc1HFgsftjTpcwTnTXiJNHnHb/SSie6QO0O1gz4vf+c
aMrG4LSDfa/qkyeGYKtbK4xHddTmUTiXgA7efg3W1gkcdi58y3lfb9GPxjkFudvj
CexwutYVn47WjPNlRv4Nak8maVLHVokiWiocM3qIWGqFUv20TW6vBzWk3ys0L9XQ
/K5/BqXeXzui0OUSwZ3ti/FHlMaOXS95MaErNodcFgHW/fCaIrHoSmjkNl+ePSzU
vIUn3MGPdo4ZKcD1PSTzfiQEewi5KkxrP/yFGuMeuEavFXkO8ZUhjgulUEd06/hB
23n9XxVaAsXonn9Zj9baPlx6g0r96cl/0a1BdYHCGoc4PxSYpAY82ft8eKxGtEUs
0OofCYz68e0rqPNka9vp4A+xodCS5dH7HvgZnqlHBLqceC+N4yVaiC7Zxey5Zhlw
NdB+PWQfDRPC/f2EIWryvyTjJFxJDssPSIA5U+XyYBA73mWk+DWBksvaOr099XNK
KN5EH2pA/TI9IVZeUQaUIw52tLGP0b2NGsbrG13Rkcgku0bfhKzW9oPY6ocpEY8d
oL75HLrsm2pkGxVs2zzsfg4ApeRokqBBnv1iRdU9zoFP9PJihTZlZ/iyZP8QCXr1
/hyQiv015VKE9ZkobD1JjU2Usi1S2VOnF8HGSOrHvsK+WDwFaIhCOolj217v3u8Y
Pz+1dwh753hgWiaFlqu3Sb/CCeC0VHrVTPBD+Mia3Z2kXnQxy5InnPsZhpTN/45t
bb51RiKPpIxHGrk9JfZtArQchfzyb9mqoW9/u8zs2YypMnlLltdZsBOL0ugGOM+D
WV9hUeA9JNjVGVUU5KdM+01Vi3vOagFbesXtaKaGmvvUJ/pSud+aeqyx9JVtfaqT
VG8d/21TDOcWYfnHdCoWtC8EAUkUpKmL2uu48F/z5bLYL45idLVjK61sTwB86crX
IUCDOwrX4exRiADW6Z62ZPRcA30eeqjwL/+pgm3KDhHUaOFQ7fHrWHU6KFCwTrml
dWD8RlGUPwsPIdK1/NFX4BiwNsaYmR3+wdCmkzE2xFIGd31hGb4OCKnFM587r3kO
/aZL9CPIPTyeTkUPYmTGx3rUP8UxSTnIbwvUAVSG6caLylcvPAzsa9w/tD1G4/xx
qxR9lqgmtbI9cw/gzZysX+cgRGUSMdzMNQkLy2+syYajDJIciwtnpEk3Zg3uLBDw
HzeTfO/zmyWtwTAgMGikFGSqgJQ5JnHqMDvHqmuxs+hV0hn2bSWM1G54a2Nbzvng
bIPqve/7gmhl7TtXYgm7z0dFZJ8Fo5DlaZEes0QaOsu469NCfJbsmjsba6AEiuV8
gNyqHkPblA41vVA3YNNPj9wsqJtCliViuKH4B37RadnqaLFrspJiVFVjF9mGCImO
irjlulk8pMRmZhBqVhM+78yItWvBhBrvccA2KT4n6gp0plh6KaWuHcusO4Toj/TZ
7q1+mmWdIEuregGJ/Kxu5Abgg66xlmlxBVvAxQW/ZvHeatxTiBuz2KNYaDsScw2/
+2Q3vkZh+v8B8QcumCK2qrMKpzxMGvzuzt0JtTfxh+k4ovRXffRxwDmqqoeIZ3rM
9TtCsPgxWozclu2jgOwGq2FoeZqpfjHZUtHiCDnyp764R8mjQVlaz72hMclz5kfS
t30uuIHwDoL44+1A8DiIoKpowZmqujpX0IVvAwlgh5SAgXPLb5u33ni4j8JL9uPv
Ppo2q6nPw/QG6nckhCy84ZpBvBl8FiYm7LBPFcOuOaaAXywuoGTbCYEH5rkd9JI3
GE31dr2QkC9Mf6qjNwPZjXVk1jJ7g8hNDQuLFRKIGYzPEZtfmq+jUmcinZsZG3dD
8rPyjsPsBkGbE2Azckx7BkdoIRXe2UuaOcNhPdPB+9ddOvXbJ/9gw7wksAr+oIBH
CmZz3sKzFpvQh6HMqxZppA69sJ9m7m/wvXXP+1xwzUKbIR5rXQTr31wYFczAKdmd
uuBXGgOeE4QC8K21Matyjl+Fhg7JCq54aWs50HSeoJehyzFdq+jnhdnevjQhuJnB
61MdfeKweiR1aw+L53nKuAzBuHZE1dD9I/r9vLkLKFN2qhPzEiZp/aUkUC/hzmmL
7sViyQClEFldv4MCPRGgDwz6sa605CvVTWesYJDCu2V9NOPta6dOUBX2PZzBIuSw
esNzxXKqdTTW5URR3VVlzfJuwFGM9I+VTLeyMMOcqxsvREkqDSfXM7txT27jQ97n
9lmmT5nKN0/DCCP+JRBxEbRzrHCJxUYiY/bDvfokQj2qZkKeUV+MzuQwNwy/KcGb
bSZbvS3MBltqQGZzCYBIhbk3E0lF+LM6zUAJnB22rVI29N5KGrMrOaOdY1zlYTNq
tFAW0KQkxPE2jbOLACkk7xkvOMGjTWJO+ie6lPvtpj2C5DokeZt3BKj0HGttMNsV
0kmLynSVupzM/Bgarwreyvxq/iOZYy1SS3O80lI/SPMUMTklLMUpLpZutFMhSxYl
8wErOLP7sC8p6sr7L0CoKzhdNI/6a5V/gkaNzefbyPnNumie6a5MNKwP3sju+j/y
Lqj54rjIAhvSKMDReWjath4Q6+66davJ1LKG/sNzZsnuuAfZQDPmaTGqB83k0IqI
iw39U7/+L9hT3W98vsElNMnw5eh+tD7QfROjVtg0NHZGtiXpIziJxfBR1/Wiwfw7
HMVjfjvJO1wdcgCG1c0mL+rt01XR7Oylzpk4VDz0GKtNsTgvG3xoeokeQEP/OepE
cpmrFhkBaOaP+4RjyCW8xqagEjsjxrIxBhg0two3SQETjBR3rAfsAabDl32/f+k0
5GtJkI9pvjWoJXy393sAhN8Snfo1KmUJtI58ii0L+Eo++dxbnG0mvuVg86gOBwZr
+LcSO0diC+K2UZWfDrlzxef/X2SRgwXamiXYRmIWqU/C+EKCDQoyLGD0p9gte/A9
Y2CN7CGzENIHpK2tpG74fDdtMj872hFDW8H1zjFtlX6U8OEuzkDCYpl0QdoPupkh
dFnTOS0EmrMZOI5PQhopT2RkpPbMPvVeJVUWUcE9ck739grfu78IqwYZFIZMsvba
LMK/arQe1448FtPw0Yp8CEtLW4tleuBQjO/Wl08o1lEMmgseJg/rMxztftMztlrH
0D4kE4BMsXAYFCZAyu3b1r4RcMco8b/9B7WyrML1bHZ8kcvdO7218yLWg7jPxC8E
VigL56Wpk/ZojDX8Sm8KaTr4+LpAyODagKtVRuKWbyrDrJs+uncDrMVDk4sPirwE
3mtUub/OWTzRI+wQUE5VBxX6P0FQvnZb0l5NcZlIZ+ROr7HIVrRgLiif1hrxf/5K
PVmyRfqCQ8w+dx0PNYND05MPG34KduvynxU/Od3j7AMx2xY6MFrM4rZdJFKNTntC
aflwAL9UfiFRqmG9TnbGvubT+aMHD1ameeN1J115M3qsIIGDWo+LjGj/TZet6RRg
FinJdsnligs7tLi3Tu4nlhCAoh8L4k9FABo4mf1Mvt9aMaqiAwrTklMecVqThisD
JRjPSgWcAJKIoRM1dKpbOulzGGZUPZS6ZU+cBEF+xzBKT1+55up/gwKx29NBhAM6
6StnCflaCk5hldsFWODKfB2qUcDHyO5iQLeDH/NZxuS6e9/48BaZ5Eh5mbvPtz7G
DTAU7ha3ToQk20tzgYccNKuR1+PYLx9PYPTnKfXGeUXCgoj8y0BsClCVEB5Lz+cy
Jm7Famtk8xEnQfS4geWnjRBb/T4duOcQo6dcmKHutJx4nyE9H2OItIBGOPX7jPf2
8DH1tkXENIow1ZL19ZYhVLAD70wi5pI1j8+VkGRQ1NipDZ8GelyOuMt1hqNNX3NC
iU8YvcE2tarV3MZwbCIM8bmeCtF6DD27wm0cJPO/5GG2dDMlAAX9OCvINxaiHZ8L
lffdrFmF5FhAIXMCCLW1goVh9j90VVSx0hvAaGWoO9xxno+5bbwWnO0ge0TIIia1
i2qN9tPNWGmsaDqtu/N7NfTJfUUoKB8FjsjcIZjoOmnTkwfgWuBABui/zlgPnEZa
/rLWtVk24ixpMQrgvZG7Vc7+eTiBe7bcGLjjsfXbSDMK2zgHKDtxbFYTShAydJh6
si2SX7AfvMssIgbO3ipl4imwH0X1aRY9r2q7DCFcMVlcYz0HsDhhNmaf3iPOLgdm
3NYij+XX2diGoof/EIlmEwI3ZdXTol/RJqMcbzkgroxx7VmMxigHGP+nE7kTwFnt
+F4XWaT6y4dSWU7HKf3frxFCLeU61dz6Hcciu6HqH2sIytwfpVjUpMLjLfnHQe5v
0CX2++48FOX0IrqJ25PUAT5aKWbtYETRxXDXQDysm7RiCDPhieOr/N9ClmtdV4nX
k29iSEWaaYB4KfF16NccwRgJCgoWCDm+hYdDmCM7lDjzZGb8g+PQ7m5Yap7ynqeH
oYVD7vo78HJAiWOWapjdJ24XIIJv2QMMM6HbxSvxZHOhd/3RO9+uC1EX30ffbvy2
n/viyEmCejwK1bbHxamky5O51Ehk7vW4Hf2IhiTvfG3+mqbKwGLRJIzbfuj+NES2
B1AVfMW+2/tKqTGG+avRZGwYPEGsLL6Nmc6Lpgz+4ote0gCM57oyrDm4b4VhbPyN
6sgz5OTUcBCItHzp4qSIY+GGMxPXbIqktJy6TYAw5C/h1QtXO5p3EY3qXxYtdWdx
8062VYMD+NlE9BLEe/Rv5BwQQGqiRlsna7fI8ydbmyfh9btyVq7ajk0xBEFxH0fZ
aE5+tsZMojl1yMEX9Tacjv+/VSXsfSSEC8RAtPE27mOSfPfQUDePYON9p+VSoXvi
1FJo5rpXLDoMGD2m5+oiYxZBII5vmsQ59A0r2VJiLSVHFQ4pnhz1G46NJp+PvvVA
9if8009zPi8zwN2VDT4WQefD7JNIqXNTrPRnG4bqZK6WRyPap3UWWqpFFF4V4UJ5
P7oMMCO7jvZfcxAg1U0sKe8yWuuEC5qsSjhrEsJk0GxGYCzTnXjtEJB5WvLcu93r
ZIYzZR4243QVMymAAF9SQVRO9vrd3n6gVLA0b4zI+4xRgjfhbor4RJROB/VF7eNf
aEh5d+JFNNXAAorKGGIQq8dbbAvdrjpGIBDSIVcJC+tdcnajSWsDANFXS3qLgeut
5X4dYndpsj/0NbDcPLU4QwCVr9MBkRDe3x3nBxaV3qkCutMrsKueowaMsmF1QpaV
VFr925RE0jU4+dmiaNDqrV9awUsLWHOXr0DK+nH5RzHgrF+qPy+ko9LpPdUzFYRv
/SPN9I2xajmlxWu+61AmbLHX00RqcI0mSJno/j0Ct81fORg5nHYaURBPscvR5MUu
EhRVCGGkh+djipre6AP32GrH60z0Y+3E9viLFpTAHSzGCIUMgwEMniomN784GGWQ
ng1oa+howVa7HlpysijNenNz+4+Qc6Qn8I5xiK3x8nMjwM4BiIOfsuPNeCQxybso
zTePixlSxNg/6hhXMaem3bcr0S3zTSt4UeD1/neoJ8wIL8l6WLpp2EQPpDCaGUmS
XlpHe+XuNVOSCcYmlLbrEKOQ76R8D9D+kqdv0bAlILCjdsS6bVXQngDPUXwCyNwS
ju3x6FoesZFx69Al6vtzgCTMlnYuOMCpQh8eosLNvNKsWvVG+e/JoUsazUr0aPi6
jZ2Fa1n+7A999dORwl9WlphYTBr0qs52gm6WFpcMip6KmpPqtpV1ISNNt6ZBXJ44
yzQGwCKrso/HU3Ch9mvcId2zjF/W4Qm9TDUXoxH8Wrj33flA2lXPFovD5i0R9spZ
gPdm1p/rTHig1yoOlObsPoA+EFHuT3/wD0SXTvQxsUSSTxf06s9/vl+mbOmOovXB
ZW+iEB6w9YjWXBFSQH0Gc/+Yizx9BeA33qgh0zq9hXwbRRe/6ajPm54/3kvuXfNj
GTnY49DnsSQrmT+GSsA16TcD1Apdr0hgo5sKlGtU5iN/mmFMQYoKwBjyp9R7AP7p
1gGK5AHkf1W5Kp88KPnDZcXETE/M6VSU6PIekhTVRBFrS4H0wLJ0Q4ta374XIHUv
iLMvDVN1/sZr+IKwYT9H0QHUMxDsMdRGu8Yt4vzjMkNk2EvKaEVJvKLEZM0fGG9H
dttHV36uZ6e464VRh0L8s5W9Mw3UJusZMNt3zhjUL5eLaZeMmxrf/aKnwaHa1q6Q
WnvdNdjoD4n4mILsCRi4dWFUGO6PGM6qeieelRzoBJb5QM8wbmcwkCfweTxaS0sE
tCmDEg5qMaCxvpnBgbYGSfvdDL1KUP48cerRMUy6oYG1KDbjO48911vl4qwA56tG
2O88VMBfjmGZ35SJ0+i6J3cC/vGihGE0UN2sOwimNW+b/YFJM8xZV/aqt3szAlX0
ZKgTXTAZZ3c2zxP5vngUHEd+ixandmrQyz9An1/ckaDaeOUHIVnnM4xcqmK29lFh
5eo6JDah2F5P/wYIAeSe9PxEzubXmxL0Zg6XfZwZ0a2e8aHEsgLE0oSRgocuOTOR
8XcBFI9ajJUMc5hDWJTmIj1lmqZImvJzxaCUkDLBr284oVU3ilIij/6uez3Xkl1F
dtgOFHO7tvhKlIF8CGD4X5zjEWm0mg9ydwqR4fzLatc=
`pragma protect end_protected
