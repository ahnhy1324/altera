// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GWP+2APa1u4jSqUB5xSMlIlhZcPPWJ31FVooOsTY5+U1FONKHBH6BFhBpE6z8iSb
vUIcVZpPi6Wfk2joWAp2PUnLhS3AE9OlGwWxZw9PX/+NnIEeIFSYgJMZH4aj7W5E
Xa1GOsCZp6tP3AiR9hZTDh5oOlPCMiol0S5SPG2qgmc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9808)
xUwp+Ch6tIyb4EkesyP/eLcVA912lMQPgmTPkVdwkBfrsHOg54klvI8R4ewbn3zL
sSHX0VtUBhOMBmNwCwaJrZFS19YCMi7O/O5Sxkeg7irUBT3w9bkt2urCW21QqnjA
jwv73oe88eu34Tx8dUMXtthW96a24pXePS8pgr8lDo2l/JrUFwsJxaySmjCKGwwG
IHGasQ9+vtK7JUZvp8ge2DDYjIdACnzL0Ok8bnefyZ9ezYRG3E08NPpHZNVeRnMd
2F0tz4jabMrCfO4OptXYfRD/b8vFkTCJAydzsO+D8EuAT+9sCH1CGlr57OiTTlo5
KwSGfxXRQD8Qzovi53Peb0PHDiwbbnTh45AMNJsqVYwZP7MzpvAEgheYXerBL69i
TLJpXKzgILdUDAKolno+kVftesbKl6Gu+ln2zvtIDIEZWRsMskX3tp1Jsk7dEXD1
EpoPt4Go/R/qkn+2VDl2sfUcvURGiB3OB1Fqc/A31B+CcEEROUk5Je9W3PPcQs4R
3XBhY2dZQ9g5c4l+XQngAmvxgX9vcAhl2/lH6X4JkwqKxWMBJDkpO0+IUeGBZLK4
dzT5wba9UsQrf1VqY/3GKU4f0Wc1gz607ggX74gpDLWQ/qJwg6dB1S2ZuHhgBWER
rb8g5xaJCJ0qq92bqLYd0Q1nkvMPC+xlTleOR+H+bjXMBqzZYOnlnLfGPPGqwsq9
Sbb1Nscr/lY2FIF/v8VMR52LIdbxU+ND4xUCGknFnSNlVlFuY1ddnGmGwbFFP+qY
aPoGlGFJ0JBVouiAcTxEeP3LqtRW8l3v4XZgrgAO9GW25YMAj3pI2VKOD553Z1/k
A2bE4AWyzGEIx5nVjjA+b+QhaUdfQ+dqLE5KHKd9pAEB19NKdX+O4i/POvOGmLhG
hMG1RXhQ1i6CYoM6B/fvvIpOqZQ2qchrtg29JFLdb5TxtoUAplX5xx0eGVlLeJAI
qyf2fK4s3E9IVSEMpIxwLrUL2KXBfKAeMmGHBj0Joz6+3Z7/oWUTVrIr1ZOv2FFa
jIlxfRey9M1hAVL2e1JWDLSJs4qbpZ3dcrudW3d4diolR/ZRDIYpNi27UXXjoEl7
AEb3rYK/JfoQqRWursDqbztqEzMz3q1/983oux9YzM27M/rl0gF+rWAqlrZ8xJfK
mLfRH/4oh8QUOMDFYiqnpJuzCnoxoIcWLaC6Fs604YyCuvalRRqsTmiPQhHI7vUI
otC53TtT20Gxg7zbEhvjH6W76D7zlT49Q7n9mf4fvwJn1Ak8C8gx+jNNWo/epBHc
6+7rm0ujMDyBExYVZ3hlT15DzsNC+E7eDIPHJtLIIatTlRLNVyvTySUSvZII1zM4
OiyR1ng3Cv3SYlumrhCbPQ4lIDgtPiH02c3Bh6+KA7pz6SSSGKFfID6FrDyWAYip
tuowu39GfcqrWrHbyk4cOBMxcyam0T+wzNTdsRkBRlEPW8x+DOzeWy6Ib0AeZ0eI
N+Th0xKUTrlMos2Dd8CnNtbRzGJWog1tRha5BAZ2ZH+GHpF+29ZY/SqI9wunvWmW
A0LIz8FGy8F0w+foTnioTVAvHQb2sMZIoxQCq0Eowkocdd/bleWsCUr20VMveHqX
x3dxrztY+o0rZNu55arg/0yKYX3TIFjP3D3q/3dLKNz87BmoWCPd97gbhBFHU51+
OnHUokqj0BF8Da97qXbrL/xNZeXJ5BLaCUatEEScXmIDPpgY90wSs8r7AqTUzL0+
CzWnOzqt6cy23LhKp8TkLS8Ng5D/FG9WgfPBZA7R1REHVv/E4W0PmFhYK+gLf89e
8pE3NWUEcsnKCG6sHCQ8wHHU/S8lRfR+RgEXjavgSeD2l6DQG7n1rur9sijVmHOx
5s2NxCbZM0zsG5eVALQ1lMC59xtBZffrPckrIfJIIk/SgEIWRqFIDapxEyz12ScR
kPOotcb73XbPw11EPVmk4vXhnH+PHCPzi4G3bl7jQQAC4FRrYaJ6ptNYq3ZIoTA/
p0iQWM61dA0FFLTotIana3+hDXq3oXayBbNDol0ToRN7GXHbZ3c/rcD1hTXhHvn9
JGfsW3gjaCJ3DsFS9RjvD2J3ItoAB6OuxL/Il47Ni26+hT6q1yYH1v6p4Azf5umj
T42m/P+xDTpMi3r3voWjj+4bPjQ8yh4ZQdlXUgMBbwgK3UCInSp4YYOJmhZvT0A/
T3RQbdbYuD+TOoz9PSMBfnGaEBDkv9U/t9b4kgQa1/38ImcjmNF3DqzxNGF8XN3m
g65crBUmxZbC6MJG6UKNidOssCAzPYg/1iEZ0pW9XB5m4KRc64G7KeowULlmqZX4
QRHZJA4e2rLQ/KHrnDP6M2br3X+XWtoH8Kh6Y3gI5hWItpRJo8onzEvoRbNMiU/S
WRxE7dos069JJfSu+KoV1iSf43EyqYc+gL5eGEiTvHyLQyXRRIb5WHSHFScsCmLh
ZIZhKqCUDsriINMdW5bFKW7PkyA3YgocOaDzxRKRa/KJ1Y0lhcNuJGqlww2hhcaC
fThgHlZ9zzJUvxgvW8gGdl/uEHDGdDkT9PvJicblpruQyv2iY/JsHO8fKO7zGSjk
T9gNbiE58eMlqwpCun7SZp233cqq9BEjOYVGQx5OaKpfisFzPF020FnUEDgHOC53
ygCV6a1wzJB8EKhshsx9nggFEuWAEyQtUG/PGxD/kMSiYkJfttOxb4dYy55Fu3a8
UvVxM4f2qbwAbqQ+y/3fKpkTs2TEwCqTJrXN4KWZ6taYES+xVSamoma0pHaMSc5X
ir/FRypZzQvr0E25GnUjGkV5RSFPvX+ctqDT1Own2MIyihjCfQ/lIcNm0nNNOvcC
bwQXYEPeCJFQ/cA1T/RPkJO+GmXvuRPNcoO/WS0D+gdDjVcpCqcASwpHp93L8X6i
XqmpeMcHhme8WSgiqjaNbzs4T6nDO5oPvPzue/YoOds3SkehHSiTYxQcUW58Hl34
t+H7dinfKhoBXzRh7Yk+feUMwThmf3AsTdl8JA6fmyRLf8uB5jTrJOEXQZBJUZkm
Glpk1UA4LBAFaJH2d9eJjEZHN6ul6G8riccILRG8Jd0rjANVIgblp58lXfGFniYn
cDGjtl0Ia3oVy4YNtYkMhKFqxfGrXwwluq3G0CmL4szTGmOWb2cxhl4aga4HjQBq
HosINhDHqJP+K8iqYLR9DozmKOFzpHeaC+Ewvs2AsGGdu+iE5h3yG2ZfbomqhPcq
v6oSI6Nc53FKxAXXdqEam/Vr9B2SQJj5Dnr4GHnHK87qhPZ6NtkV8yRYEucnpFSg
xaFlbuq5geBdxWSgh6WtixZKIUzTNJ7jux6YcxyqCfOSlBaMVvN+Zb39Lago40EW
jTeSzdZKZ9RBrcyd2tcuAWR6KpUa/3G+TKJp/XvZ2A15x00rTvaw3CgcvUA/B4Pb
3eGgTeDIsRytWP4tWnDEqH/RDGZ92NpQsiaw/FtZPLDra5C/forUOKOmO5HQtDPV
J3q/ddonJRG0n0KmUz6MLabT0nGQD/D1Fo/folZtu1D4f19X/c8P4ahFM5ATreiK
Fvjo83uY69pTVCyl4azLtUV0lYLvVNTQq7zpok/Xv/u9ScRM5Ua7QjQu+QF8hwqS
dW/EhCViSMuDc9s1eOUTOf6OUGCsp9+wQHoUDEACFALb64sO2kMBlALKwcD8Mh2a
pVj1t55OYH9sZDcuI/hKr2wip50lGHWmx6yAsuu7MkPFflhF1FVQAUNsKpbAvlau
uxCgE8oD3XQZXxKgXA5OGJ3M7q0lrAGTB/D7o8Apgn/Xk8my4HlYPBPgjtGocYGe
LUHCVHlbfNg3xP1IUcx6kzi2AVA7t1Bb2+0StKDTorGGPO7RSsRjxcVs7N1Mdmng
ZP9s3dx0taEFC532pe1OV2QtcDNCzJ9A1O17p8aOAQWsGGDReHBe3xaiztvbJH+H
GhR0lg7zPn/SkuoGnndc0xG8bgFkGiwjj0aj7uazEd8UCD336Gt5TqB8xQ+mfR1z
H5JgMxii7PW9BXiKd6XsTEUH8zSiOszy3tuQ+zIasjb63NnoYQEYWI/xOtg0Vkss
hKdqAEkETnARvpr7B8JOICvKoTIZVvvpGRumKuFzMsUqLUy/SHrfHHW+cUTVKyuC
UaMTDsrpkGGWZpR5JXirmXQLvpEKR0QBxZfC+AJ/MX9ZRS5f8UnkgfF2vJhsxxmS
+qFMZQDwOLART9Li3uKpqZZtJwAnVoPWncmds5bI0c6ZY4AqX7UUGDdX41TVYNif
GE8m9Taj0FK5hqDdHMEIzI1zKk9aBc9lpAPBAj8I9WDBshYwMG8TpLY+jMTIzq4j
4FWIvbj3EeNUI00ygBZQZBsAKVGImuP+bSu6tIqBv/2aslGmAiK+e5PZO4jbPyzV
tFiWA5W89DKBBvyp6eeoc4ISs+tHvfaYrIEyMQjt0qQdihGfifCBfsdtIL5ciZCq
CidsU5eYFN/dEdFCFm2XsEuc+6v1kHYfwzkaETXQwhSm34kq9Sp9OeWJETdOtgnG
J9e9FgW7is561IM13ul7VB7FVyiMmpTu+KThmM0oT/teTrtwYjfMwtYXCS4Y10XK
gF3dt1LMoy5wT/MvpaFhrCIlP6NKa5n829W9a1syY87EKk1kbrEtQWhMYiEs2Msr
3H7+xFm/PP9WHimeUMGnmf/O80Qx2e2S6ms+SGb/hrC3ZjuSJHuTJDjYlbjAFWo5
QBW6axlzZlor7V1pg34y8EV2LLs/33f0STxOCS+83aH/X6PqvZPapL6Bd/30face
EiaQlVlbP8dJD6/seeUUWX6QnrdbuWDghasQFSzPvk6hQlxLR4Eq0WmHaIu0JgqP
kr7tAdjls6wfPaLKenpzHXkkfoeT/JiMyWBJhXWo3lZ/eZJF9gNRl1nRA6txXCUs
GFpvKpJM57qr/8rFi65AJu01sjeqYZIyarc7bA8IC9UCXk02vKNKRpiqw65Em0/o
AQCPu3PmcyutLcM7IB3AgjcQZK318h58Rv2a07QO5wUL2trK2ecSQqB/pKA1fis0
Xhe6STzJVCEvd7uJnlCJEqHHPDKD0HElphWeNRNw7q7eqcHkELEcoqwEaORMkJCh
36BA8nRjM2Qhss4YtatkTqLhnW1wxf3nDjTAiTafUOCDGY0VlpFT2ohFCFPxMQIO
s2rF1G6TmdFvWwL0ll1jJgcoR3UQers3/0rEz7cyWJ28v9N0mCOd13mdw8res5Kl
Ofp61AKnusbr1i/h5odzNTNFOxz765z5CTX2HCFNBDpnn33FG56qQdy56PtsJCi8
LwEePrgwHJvQhxEuvWxhzWEbaYwxekwpCSzXq9+tuCLwClMtzxzWRiOtd5C2dcSu
+kHi7TToR5MeSdykqAhg3duZQ11fHYFOpwtT9JTGydlQwuy8q4M+4Q6YRTjA+mlF
Kqnmk9MjrLm8ACXSD2gIZ8tEMqUPrar9U/Fmkffpd3s5b5WGeDx65FRUkii28wgK
bTTXJv/JieeDnOMhQc26ZLL9o76x6/o988qXm7UJYLsZh6jmAO72RRxN1IkFzkmR
k2APqSkuL9Pz9FymfF+xujqoWdRkM6SGZ5T/eivOha/M32GudSvwx1DLdKiFocv5
FYdao8JP2CDHUjq/6pXP4jWVZBfbnTRQX962TKvBwPJrGfoaBjcXpCmVxS3SBFxI
96FoBEamDmWYxQSQf+6sgnNQUhUBUBTzDj8PBj/5c1/ljKW6MwoZotX/L/Z/VUXq
iLLJFY7G47hs9nWgeLy8Gsi2Ikk1nhAw+zwzOCEaXCuXvSdkwu9fmHZ97qPnGiLX
xKinUUZzxs3ZCC1aWQS2yV+hctEQAdGdmYpYZEx7dCucMS0f5d9CwMZp1S7x0DlF
Fab8LEO4tB1+LD5QVP9LAMAt0mbVRUpmFZd2lbTuJzg39CI3oN1KzEEsiLNowSWx
ifrOBFSPII9A8MeTct67fro8raJEYlm98kX0zAGSFPNU3zx3sOhSn2JeMMAfsts2
PmeLP8PoGXq1znl6vDitSVy1ft9tGp4wYDxRU84Bn2+yX+VQvnVFWibKpcrh4KST
UGheNCmadCI0d9PwANFVABKkDJv3cl3xP/4XsE0GgqxfF07FTLdKxcajgqDnSpgn
AoFRyBq47krxPmdzEYN9A4rNbjN/cQJy18Gd2Zy8drfnkkgdymo7k+ITBO+0eeNY
aSzOUxVZMJV9fpy5aYcLGIEfoHONW/lTSBD/buOtPX7mCKQzEONLywdgvKwGKs5x
RxSGarlt2Gne/P1zjrhkpR3jJhkok52pgLFca+jRGSwyxSO/v1RMFzrofPm6REGv
vwCqvs7ryfTazDrFP14aZdCp6V8HadJdCRGNXpWrcRwKzvZTfoJd6oJ9NL0EqzVz
KPSHCp2JHUzwjHeM/xr9zc2T92doxPLXv5MLijlGAWNhqsK2hn1zo/W+zxR7VAnQ
gfi8VS6oT9lPUPUBMBw53KgFRTtwNF8qlSwuxU2YIZ1COXP9sHDZeBopjKWa82NO
shsxxcxj0NsbkeGGtiLkH9mVehDUsgArQ52MUkPLndW3X3HWv1ly7vaAhV0Cnu2F
nkRcjHzufKLgECf/KF60yWqnMhJXnTk6phmdMK2uhS5KwyG/3qfVFJvi7pV7ufFi
rG440D0w/BJuOg8FGBvH3XgLhVpbQ5KJP5drGVAw/wKIs83iN22T3+0MTln2d87E
aiRBn1sU+w118jwxK5MK77UuC+tIZBAh1gKjxKFt862hARRmkb4FpgSMXO6E8XXr
sJ/Bud+l1jzT6LD6MWp2Rc1MbGEglNDjNArhd4BCTMewjA6cxS+IHCEOeKilrEoP
zheMuxfikTnxckAl7vt1z57SOQdf0w2T9xdIfL+aaSR/TPajXs2eczcPJjWEUXFZ
ZdihOA3KvpQ2NsLr6v+tuQ9ZQmZnuxQpJXBzUykir8bPEKJ5ltPdTqU+nijiGVLc
8eLnO/U+ZduisSyvrPodAPUTuy/4ZbeRiGD3RFgH8N6BfUsPLlTg4465OUq5Em2H
H3+pl6uH+7JP7YOL6FwWrBLzdnsMBzcuTOPM/6/zqFWKi9QqSOYH0y1WThewchKi
4vrDwoUAatq+LNdQGtiE0GFqAM++qH7ISSIT6yQC8ib10RBQ7kQipX0fGPImWSZS
hx4e0BhG6xJdxBheVV9cGqZjetSlnG/V1IMj7hLL7UR0VZzGzoFri1jKq2O55XNk
f8E1qjN3YyXqPLVMTaFk8OiqCLmuuMMtPYB2fg0b4J7nIVpLo2yYnvS9hUWmcUGE
YFaITvsuGgU9clHlvlPhwNYDO6fKjEGKa3zPBmrdR+GNmwWC7z4lbUa5Fu9IKivo
AhZ6oQN01RlMWpBI+n0J0YKJUPHCKCuatpwGC6pceAy5AP3LpvZjCwQcqytwDxrU
9ntamHj36ZYqXEv7RQuN0qbm1iPbbPhgYa2A4wxOeno0kmVq087mbXfwt5K7Flmp
ByoMnNJUguYv5DVX1Egv9XjhIeThks1zazS93UItMPiVSwRh10+zLsGsdwa819nv
66a3ZaU4iCLIxv4tsVcougp60Xd2Sr6dDuOVWfidQbLCmihc2eBVmbnBDkh5k10a
w7GzSmPQzeFV3QE6NKTAHTYl3efdzk2sVrf8e6aJgYV6PWHWhPGqLY1lTMi9Tn3n
ubxVKIotO1OLTqpB3F+9TW1kl39qnxE/Jv/jM8xlhWwYErN9apVU1XaYiN3qw9QZ
U74kaZCxzOJ5+2jsvzTfQSjG3WzYpQWz7njKC7PSxfpJtkylEzpie0Xo82AuzTIF
F3rpYrOdK8PojxCrcCnci1iVLy1oHXwYQTLAlAXEm46QtH3QYO4iryPteAfdMWjr
S0kxSNur891vxk5Er0b2EL6FUceSHLNOnP4Njo+EB+ksY/1pyYvGUgBKg1S6ryuF
2HsUWou8hupjWECc2AwVvYPe/v0Wv/lWZn3qnC5aqRdQ3GndR13rNVoOCG31yaz2
tzobIU4k5DgI5dhB/7ZCbdbaFv4Ommd+4HLgle/av3VJiMOYUlyMfOcMcQXTnmwd
EDFh1Lm1rgNNXSAsVo8tf6kVAtMHyqTV+G0ctZj8bJSuV50x9fx6+Y59AhUFObkx
ailIF/9OtYII2Ui/zfVNsnU+LbQBcPDlewy/Kv3GyGGPGVk8nobbw+6jNYBSjPGT
H9Dw8qifQHZKCR47IxQrMCzw0r3hR0KkycGZe73FFGltjh1HMYkwvwKW2L1OPD9y
mgpq70F9th/MfJlzaSZ0tMTPsi8YbVBxVe+QXoSdIPAeIDvIQ3wbSU9v4mURvqqh
a16QN2hzWqmNVXpLQ+byTcYACOVDiCVLMQBjKvvAP7MABoOS4B/+uFeKbvvXQPNM
2f8hnVlELgAWY71PMReUoZBTpbVWg2jFrmAEsNlrfJYcWSgxBl9aHJrM8mZbz08c
bpaE4Sh5n6LYOT/t5eTB7QZgsnUpau8Eb54rGIG2xg2NNUa8hzNcjl4AyrVGPUKK
TEDDe1um1HWSIP/r22ega0zM9F4GbZgiddEJiOJpzEZEWNtTS1wUyG81sNuEyYLR
cq1Ql2+G/WDbdYUiTJnOZlgSKEYpYmPQpsUqhMgcUhhcXqsH7Ea5VdHha628Xiqz
Ckc7qss6lSxIlhJGPf+SLdQD9XGuWXgD/k9BQHUO3Pn04skHcuNooJWwXbHnFRRV
zGdoLrPWizVCQxrT3+CN98OUTNLgfXHb4ayGtJDXUOl885mxQ0CLEm/zkPIxpsM3
DtqXlj/io0ggiSIWbn5XjdBrs70kEocQdbbgONj3wiEHoaed1+QQaXvPcMBshm0F
0HNuNJY/bhDin+rZi3+jl+knGmi44TvJ0J8aTqRNZ0AQEfnwq1iPDeb2FZDZvUS2
Z4/HuZqTb7t2elcqyZIEiaRl1gIApp9GoUHpH8mSbA6UopUx3mBhb+ifXWPHpL29
hXU5IMhBlRCCeBuDVWM4KD4iKCqLkGht7+rJp0lhABWhxpFCMHTJUwfACd/l9q1s
o9SIKmLl6rlpTBnApSA0qhQ5NE/+Om+rBTG0eH2cvOZs4lFH2jy29eSMw0XUZrYP
ZijBQMDjDs6o+GzFgwc7BpkzKkvmMSCto8F7/5vP0QkGieUQ8nILNX4i8gs2cgUD
NGbMv6zjDK0E74MAfWBP42HXzbG5OmO7XqhUsXKwADWPh61HT9JZXhkT5IDJBL63
HtKSsILSqB/WSt5AQkvDdZCZmMIIedHqkkPwXJEyJxvLQWmGwC9Io3irksxCYtRh
qljKuIaJtsH0FUtA+wzkW1ZcXa69Axs1g0nMomeaVYq6CrTrZIvuqjgasfMDOBHs
7IDe3D5kqlPZjNU/OTozyqZUyM/rKZb9OiMhJlF+27E5cwKSqb2v9e2sZK2qOqYl
SHgOJCFGVJfqlBRU1YnhjPiId4C+cpBb1jM6DWR9qaeHdZRGIa/RbcaCzZov/47T
OFx56E8yvppMfxoXnUMmTj+9ldIcC9kJjPlZbrdv06+w9W0LmIt8mhvrHk0f7L1t
yQltlWCNri7AYmaTAePoMwM7gYEZpHfWIx5p1v6GxZckj/7Qi1ZcY5qGurWjYuQ+
AH6RvU4QHHaW5A0DvyGT68ustugKNJxgnVbarITuF5nH/nOlsDOJughLtLgOqTT1
kl8Xhzb73BYjbRm3Frzx+T15zg6ZGIcPA4COKqAfe3Hlwn0XwxX/qvlmKg/uBi37
qJHZnH0TweNRycczthfRNmCPKGeWPpkUNPyvbg+uWTpKZ5IDft42CyFPFC5Q0ono
NJy0eKFU6r1aYzQTQxLCbFwJM+RajvAr+ENRW0ipRW6qcjNW8FHEu+FNIDxlNwGv
LM+symBvUA7L5cCv83gh5XuEoI6Ef3bImyEa/jeK1HwrsQKyCHT+Dh1+yi82c0Bh
j3oKvXIZ0H4ZI1/olVcA21hLGlGciY8hMeMiKYXUHGfBQbLk7OMT3pSBsie6LgKV
j66hP+VF307tl3Q4nZ964Vb+qDG+eHoYpk7Q8eOAgYaYAEiCbDrraILpENDSKg8C
zojrav9aIF4XrRsg9icLVB4hYW9lTyYoX9+wJHmy4mCP+NI7+evJN2U+RZIBnI5J
PGp0NI0dhk/nXkFzovzS1Tap839UZQmSsIDDZRRcuiaSl583eDuLzav2xUN9DTKi
NVZ5QgNns0UT3PZ36vyDpYfewWqUN9thTy7c+23u7BAn1tzQm20YTM0PFS/8cSc+
2/gDkgbew3wcSXa5Wk7HqrMK+voHlbCBHN+W2OxEeqMzyLKRna+1PVhSMN4UViir
4c4e4zoY9jdpUV+4kjnPGXDgoGA9dZ0dHN3IfVFaXtNAi4tN+vspxOwJCsPA9vTZ
x/pTqr0Iwq6r76C3UuajsNK/spUN0PM6QGFb5aNAQc/JVhu0RQSFAdpeKoA6TnfK
ckBUpFU1pTP7MDKyrxwV2R6aLsjLe80xvNXYyxLoZedfAFSot5789/GdzoHWWkaT
LIYXRDlrflKZdP7EBMc0wWH+QyF85GBBZ7DVasAvjQ5EeoPkEfnDPRIhVasKEr1t
EyxZKqHm4G7spH0tyCNU8rlBmDNIVUCmAf91yQLt1dxVnGj5JZUblyWrBy5lwcDp
NNrbzAZOM9yNe7MCG2HnPdXqnucrR3mvCgVnWZ2uQ9JKsvunIIPfMDEKc19R6puY
JHeyO3SCmG4NbgvLjJsdmVAlXGA+tnbQZJnbGgWCF5zq/ZDBRm2NlzAHxrzSHwEz
XMcnRK8MPm2irNqcrA8+7YYNyI4BwD68TiK+Ei1qgW3URRJLkR3Bv3UnDXuqoE2I
ideWQRYjf0lOOeV7S2m3968v40qtDh/2TEMGXiP5c9hvlp75pOrBY/0cOqeRvgNH
V0ts7uiRzbKnLVi0sBxK2K2+oDWW8qN6XSRCPUodeKat+kDRAuqz37o+Zo/ZZi8A
MIIJnAjdvJOUiSxIpKh0XqYx4nKMqdk9U3o85PSm/ceW0awNdVdKgjiZabvL7HsV
lXThY8BnhyuqvYSdpPGE4a/Rg22+VQbSBXOREn3oGcl4OafhtixoFecI7TjP1Bft
kWSOZHaOj08m/yjyoBT6KisaBBjvnTdFUP3yLT1H2u9NMJEQkuwsWidWAJjgtV8I
1bt0Tl2piZgZ4w5oENH23s2bZtEU6TaSTmoprRwP40ISjQZkq2VO3shC/wvPQsDg
sFYVd59FDngwxLu987SHfvYLg3wgxJ4jUoOSlI4C1BXwuR5saeeji3M/49osqXzI
x+uswY8gyM5iwBfjQqcTCPQrDukZRn5wHrr1CthnCqhIgkveWWXAAl7MuVivFusI
jT/LhOFyC4JcNGVh4p2BUAJZmOuUNMZiuCJtjhzNH2WOcXWMZfE7re8SIHxuordK
ht+aCDDF0taTKri3Q2SkSeAPBzPukC/R4IApdhitNaY6+XsHGacMrh4ZgDI8t7M1
gQLmtQ6PXHIdUzwYeruBbtXg/F5hQVX55pDVtr1thoE5YsfscAuoaKMicMHJpZMa
rayt8QTz8GntowzDvUtcQTtJcLidiX0MuBPg+MvJYvQ6b9mHRp3Fd0Ac0xX7OCz+
u4dQ+2rQfcokBo1mF+rfORMTrbhXj31ZECrvzV2eH64VNmboDqrOKNur7460wWT7
BEYXGCd83uN2S5SZQajyOAFhAiN4zG98qDLIN5c415ZAMXmcRNT3WIXql2B5B5XG
mtuzpnjah87Ohm40nteAJZ3/z4jdvTc3i+IfZZA1GGAFOLaYBVlhWujD3g6tqR5J
lMzLevszeYjiFoeVWeJ3YvssUJRGaHNrgucjbhT65mVjp89T1T7t2n3C0Q78mkgq
wm2raD+R8lwiox5H0cnB+bU/aV9IAt2Tn8vUdd0HD+WtdLCl3/8Y2iQKV3IK6/GK
I+0qnYK3C92VKCMXSS0SVZZgUodCm7XdN1BZ0ped3ZY+cd+tpx989MxXxi/CXIlD
azbGTl3com6WLPeL3GPGfF1Q3Bsj9lxA6HCioWpuym/GQIozouERW/euc3sOHz1U
2ZB/UVIdysr5aKYKpYJlC8L1YwlrnF0jZXUcIld+fwf7c2TqXjFuy2eIR1ROaH9s
DHbNp5umA5Bsbz9BrWeBxWDq+yFDLCBxKl2Z5JMLAb9xOEm86lFW32FWTXrPOcKi
na764dAcLJiA/6YUJZ/MzL6+I4nPPkwWsCI3JZl9nRmKjpAXa6Uxr9daqvARo41j
peXjv08Wn0UcY0/DfZZVL4AWrY5jqL0JUd+Ue/iD3WB+sp2YPkzmL1M/iIAYfdgA
l/VMFjQyhrbZmxpv35QOoexsUK2tRlTIZYym9EPMPAI60Q/TUtA4z42TczJCQJap
xZQIoE4sGyEMr9G4/HndLOcJ8IO79Jcgm1brLa0ipNfUd77U+qJVsl2yGcGK3hDw
8Epgieb88FAm/+t1lE4OuNGAbaixtprKvZ7Fve7zZLfTVkPmdgjQYZsDq2RwwZcD
c49afGbELzX0fLQ7dclObVk8AXIAIJLAsT4X2Osyqo0ofVgP7Ca40iK953CfX0rZ
qqHbPc52X/4bkn1ztYkJ6L+4/iCYOeX9tya3ewxw+WE1VntLVW9XcObNoEvNwQLQ
jzEpwqtNiA/OKDmF2yq5HwJHg2fcXb9K+zyP81QwGI6xhOczOAvXgvambeBfS7YC
cGEIMD7FExo6twTAqsIceOlJ4PhVtkaGOJ6gMn7wZGKl/ls+dZbN3NizKIGqa/RY
S/ja9iIHM5NLflPfaCCa2eW3cyVAdYvUh1k90AO0Nx4R0z/kDoyey3gio8KkxieB
kSrKj6uTHS0dun9A6b6CiflMn4o9JUU4d9H9tFtW0bgs+4fzihufrxJz8PW2H+n0
vTmZwdgpSqTBrxFs8ZeuOC0ZHOVtHdMIBvjZ5g+64IqXt6hljDxgZpODWo9Y3Vo/
JbTtvI/NhpT7MQDqXE65V9kq/VFndtyncaN8Psewatz8CmUoVgJVFS4Zp2JNo49c
etQLemKwEH1QMeKhem+5px3ht54d5FzQbgBb8Vov2XAGf3uvSP5ddwTrpbsMihw0
gF8Cyzv6xEfa1rYpzZTayIMGYgo3zl9jB69SUgwlFfCU6wxzC3l+m6ZfUOx0nSWe
Nsmn5YeSgskHzTHaek9r2A==
`pragma protect end_protected
