// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:46 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WAigC+7qEVw2ez3Vr2NRv0OXq0omN5enPgKvMwVepVeyonzuDh75x0dEw8zas1f0
bDfj99K83P/GEPXeoVjroB2fZ8g/hGIkMQddTh8fXAJS5ttCUWORwh5sIQpy3Z9c
gHvFswttRdkwUDwN6WFlvY1SS2tGmRFX1Z9RGviHq9s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8624)
vdKy8sHHAjiVfRudumxnB/TQcowY2UG2h4ULg3xg5Q/JHa0I1UommZOwNwjHz1j6
FJ+kXygKgTGiBZXvn0j1NcGMlrnkBiV+sEhRK8iae4yjsSWwTcWKt8QT194ZkUfm
MlsO7LNE7sxo7IHnUFH8gaK6rI3TWq3AGOctPSd8d1Leb16VWTGRDfDUtweDQNYa
XBBw7Q7uPiFsoILHkVOO9uiG2mg6QBGVOUCYzOgjaOENP1bhSWNS3sxRpOokAMYC
dGdUTf1rpMyJBA4Zj5hbDG2ZV8D7OLPSpNNbuZ/tRpepXcQqeoIb2l7AQ48YM/WM
BSFkIqjuf8r4uXu1lYSBntrkBvVnRi/b/5GDCwQ4u3DkQfJRU+T2u2TuQVKmIjEM
d44NvOTE2L0QXycsHontrPt+nK/Zqq9YZCQWCjcgqUSJeeVFmFjKiz1AqMukD89p
Wt8X2Va4lWq6qcAZqFc1LaC2h8KLLctnQK1pWqOcwOw3pLFYMkwl4M8DG3sOHFKu
UMpGZvEEjfaly/weMxGSYZecFCVjNafVEnP+CGFMfccAUo84AiTGfbw1l8kaXk15
CEi1DR6o5O7BsalDczVyTe3IbfiAglGnMukAWrHuCpXZFdreNkEaV7/GEwOZWFtH
3w2yJnME1T+3E9IixCvhUxOVpPP2ZDNa4GhadDe1E8Wv1TaKtlZ4LUueh1VnfABA
h/59t07LRX+xrdWpb5q0BJc++MKsEsnhxDbrbAB33mJxHoEWCoAg599qByzfeu0f
VKOsPNvJ59vg7xwLiwJTYhjSb+wYPBUdVMaN65gOSqSwRPgNG3O2gMZQf3BzgY0J
ZFQk7/YB3sF1UGklTq4T/lU4QtsOTRVRY2/QyKL1uTuxJjtIjOok7x4b+90PTmQN
xySwcmmqUtwAf5N0ZslOyWWNgu6iPLmU4D9ghOgYIIFA3T0N6lNqpkfUhyGcKfv9
Ddb9eyYw/6NcMzSgHkj5UHh4oky5SwfTixYcNr+Xk2gxMCjqGMQ1CHdAduyFvF74
4sd6wBzSp8yVpEAKWMpfCQTBen/0dZuACsOtsJ+IyhX9KCY94d4or/olXrWU1Gyi
jzB9C609rvyIM/i0WCpb1Gjr92+2lqFCewJLe7fInrW5hm1iU89FFB/qmu5pTIyH
bTpMzKgwetXTu3Aad9QxQbgvQtGB4apTr1h4zSXtttkHzQfEKkoXfZdAy9MYJZwP
qlqS2STe9MQTR9SH8KtYkHQP48mNm8fc+3RmPE48Yec/1b2zi/yYXHEbS1a/hDpF
3/1rStALBs/mIOZZELOP03nOmELW9WaN/c3YSBzpwtrb4XI5L4lw+NVlNNU89P33
9LkCl3pKauwt6tdXmSt0Vn+hTPDT3wyO6GQJkPOZbOWFk7FNkpygC8C5hMns8XTz
GgNCy2rHnCY2NXL+AKhO3nn4DpT0AAGxMPawVhHy35f2GMGPAts3u9qk8rIPAD5d
/Y22NUO2GQpgjwwgl87lK9aSXOa5gwk0aJBt0feR4kstULft2SaOR5UNxPHoUGPQ
X908LrKUKJDb3eyEiO4VfLeMVZfjUinIBgdtD+13134RNxA3GMldH4aa6U5pZYTl
Wmkb1orO6OJAmrv7czScDEkiiwiyUkM00qkkpHv1bNUdeXYudMlddue1BOQZAGga
H7dzgNaSa5m/WRqWk9B+3Kg2tSu/JYO/KY4szRBD6QKA4otq4fIZUVLz6nRLhzL9
WHdpkk07wNfMOMdpf7eLZ8+IZdBSeCWVl0ipGw4ijNKfYVCLYok+D7v1ou2EoAlH
FCHrciTemu7pJ7qnm2VXrVoVS5NgECbHJSYQcvLB3VTEfmQIi295byyoMS6tLIv9
m99St4vASRehTcBEWP1hL1dNLjH+20F7am4se+q9hYaWx7nk7GrqlKQkj4izsMvh
rah8H2GK9vdwOLxVInJtMxDbrY16BNVSY4IH+RopQQEI1tXMcMxdZBxNnexRv5HO
2LlTxNFIhicBtNHOUhaSRnmAhbB4X4qbLQG9t+hhXALHdcgZwd3mAHKsTaaXA4JT
xtVx4DddzWhh0DLcVP+t3j1NHy43JyYK1IwKYo7fXdppCc0n2jodNK3bTv8Z9dKm
Z74U4wHtrprnPqNzy6Eap4UVZ1qCJqSxEfMeuJEj6j/eC35AmQ5M0q2oWTISfg3i
oBJSiWOufgxrrLclEnIHx2V2MbNc2nr4fMkhSNBrL03yTfiKUB0F4Aclpdmoj5rN
FyZ+MQDmDXHJq1NWcOu9O8HETpfr/5yKwJFVs8CopZH2WKuuhQNjUFccx8WQOUxB
GDQz3SBiN3US/XFmUldMVZ52PvB/3lzi5HApIQ9yg2FzDEQutTdf4BhKoaT0+nuF
k2hpzFDPq1NIxqR6fatVtBfsqHIBXVaWjTZUZXhBpEDHNL9a2PjvMY/gbc72gYLm
8d7YOHd5wqmNlczrU4boyIrytKxj11JTjgLLNn1sK98Sx0IJz+bItInO6goDSY6w
GHNbl8f9xTrSYxhTShOwFm6j3g57FDAxWW0/87rM7Bu2AlXuKSqAdlqwqrWvh2Uh
0D5VLdZJjytF+p4U7GQLaSK8IqmPaoI/cVLYsneiPV3QKi/QJDL2DaWQeM8ryAFE
Th28tDoo9FMuA0ped1D2nLajS/akVz8Z56WKxCK8qk//2GBN1JBAhpc8dbP5rQGC
HN1zFXF4vCsdcgW1rJDWxCrK5awr5ORaAZA6bkCjPBc462Z4U/3pz8nDrGqSO0NX
vBht76Ty+Ft+qvoty90V6ZiISS4KkA5RpPJoP9ZAphIqPcoknEgPuoefMq4/SaPX
0B1k5Ec/vBwLtw7iFTKWVYBA3ZK0L+cv7TXRmEdS0lZqjHMcl2pwaHoFhHbtHfWX
JANaWQK38U4FXesN79C4JJYb+Uc8dl+Hzr8+nFJtiBhkxTrOQcOsnkSFTeZs5pyk
76YzTk516onYgY6+Jb4L4Cee9xnLBd2EcQMW/moAXHJfh/UvbD1FMeZ8e3qUpSio
visLcuUCntwIAuANYVdCddNrY1w4WWGRpdgLXvIvCzK0kk+dZdm30hcq+2iLDKax
3Gb2KMTfBubbqsrUujnGA2w12ryU32sqsRwE4ccrTb3NvgpOENXN/7AQqL5exWT2
bBfo3kXz36EiszqWyVzxPwYPPYADROizFeLTHYbt0GoYu0cAukmwgPPwAB7PnOCd
svncUU7KxO3tWn8t6qWN2NdWjCfUdk2+xCQH7/E9pr65KU8vALqEEm6WDp7mDMig
1btqtJJwYhQM/IryHVdMUUC9Awi+zsmivL3uVbDB8gzcVdRXtuVg9rMysV2jGtSP
miXpJcFAJvIQCU7LMM55jD3n7D4K7VaX+kqViio3sem3c9cH/jfN+hs60fZ1SshO
/Bd3rXJy3BAKm7QGLj9DD2JyGZ927ZVAdnW4xovTTiHzxG+552eeZzRiJ7mFNWcU
ZGRaxuaXCKcaZ4E8alk6cf+ALwNLzcVRfrHb5WzL2H2zKTqe534WIodbmZZ0ARu/
rZGbeYvatJs8pv+Y4P4+fQIVj5SGB8ux98cVkrb5E8/O2ex9PHcALuqeI9HaQKjD
zhsiDze63Koy2ozBTyDYi3sm914XwJivAHMWSE4sYEn8du6J9tlbAxOpuMaF7npw
TaR9IhoFbloEHbhsxiKDOJer04RcqyTPRAG4viTx4qC+J6fjW73QjEr8Q0kxqJfj
+pdYCY10llmQHjO92HuJ+rC3+UnChUjOT1dEfwTKtC9eW/eCkcKudoMCV+uxkwS3
OMRH6sqf0QmwFXDQroouVxnjQDdASp+mhh/C9RnYPgWfD3szsAo39vfg62NcKict
rTiFV93FFQh15USJKVY6Vdbcc/y4jOvjBfYvfZNUFLvJwchC/At7UfGKjOv0ePhe
4QFaGdsh4N3El3zJ5YGD16cyQaXgfO1KpB8fb+yV73NS4OeftK4simg4UdLaysK1
DQnXBpqwWCpFOFDT9SHQ+QFh3+OcpVui3YhNqYMaTNzJ6GuAG3jXal25QiC0tMqh
wKlwW+GltzBvxNP3/5Cql4xUzW5dCCWOtysqsewk5ONSa5h3zpqupIJ1uReNqiiz
ddsGzbJ9huHCDBosTawxanapnvSa1G/swYuCcitry6zmFKS7s+4yDRkaLz+fUjst
dv+z5a/1swyHflVrfgMtKpzn9ITA8SGfRb9T2x6l3ekSfbOKLvungzZUkOgfgMJD
mFMNdChyhux6tMDjd7PNcL/HcwOOtKOt+xydYR2ypZroNBXu+2ccyDoOlTmbA2cY
woXpdeUeBqkHheILUWzgIFq0p73c4qKreVqux+ZzkJq2DLva1mZi8+8dvIuDvlY6
lXn6bYU9doPnZcjiZcWwvV8I10yU35tlTPNpsoVVQpYoDCRmaNbrlJjaT0QPxZug
R75EmY57M/h2WTVq/0pzWTsvkkncKfllhRqm9D7aiN9pBqd4tJn23pj4TT6Wo3ex
Qr5RBbEyFEaF6hScZ6n9PGy4iM/Kgu5rLUvtYALMfg8EPZKwNnE009oc4kn9AqJf
zzFi5TUVuKS+2N43tWwJenxaL+8w0Cxh204u8mZ/6NJdxHEJ3xgb6wy+x0VvGxuY
Ayb6EhPrZwWLEyV9bMNms9hT+RLn9IhygnxOJxo8+oihqfzReijpQyJCd7UIV7KK
H1TrUibgWusa3s36Hb6iht8OjFZdHWpLP7agqA+V7TjlxrJ8jOr4t8cEma+LwOdh
o/NK4o3a36oUsk0WlHFOgmg/ixEpGsxhUKmn8QLUXtLxY3rJAU1vsZKPs/BClpey
CCkZKtjzTBKagDuEiw/nvZPQWyCK//Zt+nC+f28GackWPG97/S6omgeflJO92N9a
geMqxeXcv/KrPi4yNGjlNYllejkUwQVlL3SileFEoZQP2qzdEEuq/W8Me6H+xvzJ
EWbx5Da/OG0KtgVajh9nyrMDitXPkV8dbKF2ImDFQ+RLRCDk7MwuAhPg3cVypDJM
5Ywi+Z1srrQm17zZm5pv/HayY9YwvdzhgSj0elRPI3h8yQumdsXBdEjYKN88qCEd
iIMfwwhf+T2Ifava0dU9UwQ85YrDynn8BtvEswmCqJloRnZXYEK/jtRIEryGV2fA
pHbAs1n893hiYrqipWBN9SmYVyO5oddWO0sUIQkdmTJsOB53fhmNexU9QiWX21+E
sdF5K+qv2X85d4+Jg/ofeKBZXYDUi3vG9NxFaVt4WodpCKhEClZ9K7IwziJyLHcn
kbR3uhCo7pXE3rK9c/JmD3w2WG2WP0fXEOk76oeMYvgcs3uX0tFLuYPQDumaJy3o
Iaf8xtcpdWTojN25hBlYt+4MsIwLYuqv1KsLNLhWALUBcGfLoJZynN8laEEzqN4s
PdHbaYG6kHwE18IZYo3+hvhrUM//FnzjtmvfyQSEDu5Ru72x5Kjy7iBpJf5UaD8S
iNDu+biwr0EQCY/knsWNRVG+mUPIK+smlTCFjxcYR0bYEIxT+Hs2KxObM7zsXN5b
WHV9LSYjANu+jcHDcEM6evcXsGtOtz5uz992zlOlM5+0xo2nZeJpyCZtAGPgwnxX
fpH285hBuy/Gl8gPkXrLDU5/ohLmBAEuOwOV/i1WrlsHDFgfR2ESaGH01bEswzMO
0S9uH7aVs4d+AjEwrdaPJ9SdLGTrDNqmZluKsLAlNSC2rveoKWxkXQTHLAZU2gac
xotuQeZKyuVmFY8m+vqTsuTujGihWlfqBhfsjy4/ZPSkAA0qPlW45WgX111w8fgv
TffcsT3z9wHugx87ijibFIBvrVRMmEfmLanhBRPzJf8YFnsrI/Ks4DKJSK/3R6wf
1g2O0SZqOfH93z5sQTaXEwJgyTg2susONWZ/sd069DRBufNg8Btrq9of7Z6TV3Pg
JXUJ6Y0qcDUgsXCJ6CbOzCsqhQIlDpXIR0fw5O4XRi8jE67qpxwFMurlj6MyuEPR
+yxGTIcWhuYs+aHLvm/I0ai881ADilY2njg9B2ElOCjbi7FVXk0GFmlSLYQm6dU3
8S82x3ywbu3LdoT3IChiw0Db3lCCCDkx3pnrXr2Mzge7gx+YCY8cwDzhNIw/cX9y
qcruEN7DdKJHY5EzbMpN4/IjpI73ZwgnUiDKhVhFvOFzn1O5D6+l8ow+OGflWiPL
lSgZwFzcY3TfcTSPWwaI8jq/KJk4ndqOTnN3PhhmYk6YUzNrp1WoDfwZ5fMbiO5A
hwRb1VBz5NrnZT9jFpTftiZBsXAyvv2VyVVRTmGVyS60ZGbIOogm0Rb0kbo7gb/h
XYsUvyaTc1p3fsrTI4jzz+2fY8DwCY732XmRggqJEokisGncY8EpQ1DHnUrtQVCK
uQ3aZn5gEucC6aWboQT6kBYPqk0NOpaKsOHI0EXgFfip6/sZKu3Dh61seIACWsj/
Y7l5+qrO21XA+Skl+Ly1lc7ARoHmuXqbAUc2rAVV6n003IgFvYahIxCobeL1YWSf
jXLY+A8zjDxTot3Ja5NM8HE0rIotJbAHrIBTQxha+GdGN6jH2GqwfJa5wDzX2XjV
keqv3SoVgW465g3kCD+vsrdcij7dpJ1YfQAQvoAF1MMKJOzKojfLsAkttAbjyZp0
DH7WyogDG7PYVQdy8QFJ6OXckYN/ECCNyyPGuqdr542++3Iag5GYIt2ot9L4RakD
3nAiH3Ku70ji+NhJQBO5d4vZQ2qa/FcpRQCp/OZksjBtdxLSHk9IwKr5iNgq/2aR
u4j8i1drQbU9pJDtwLOzXSyryZiK6yKhX5/RgylatKiEGdAz2f5Yw5A4cdbw1Xxm
JRAg9ykMcEJLKJy0EMR2d0q30Tw4LZwP+AjA3/tGDOIdNQmoZ3og5t79MJhuUvPd
xr+S/eWtq1VpRoUUJHUnIICosXl2/IcO8Z5yrpLbHrGJBMuMq+hzIKCv5jieZN96
2C8qrPh2Yrmke4/9NRZ199pRUSr2FYZ1v7l9CBqm2MO/OGylBK6/cGArCHgWbo6Q
vppexXz8Rt+1jJ+ySKHZNg0GzuBVa/cOeppKe6rXfP+GhqiUHUst/sWLXq1SW1lN
kJCdQHBWrE+c7FxeMYCG3p7+cr/nsnMbPEVRVIvgqMBLEvfH772Glq9zQ92tkEvQ
YM95eN1VPNje5pORbjeYEY5lJX4jw/OGxf0VTfmHu6LXJu5s0H664TlIjP+ZP58z
oCW0TrtbaX1bNKB8BeezV75AQ1LDzozuQpFGXnutcYsHsr+3yYGX5T5yOSTEntx9
jB5r1rEfIn2zxNzH4QKr2A4JyCaV7MdO0G+kiIvC04pi1hfSxID3OYuLo5sBv9yB
JGfp5Zqf+fxg8NaaUIvfp0QvTAyK+hE68x+XAQ4LAMZvmycVUgfNnCYAfq5V/VjM
kVvv612mU3A01rH72B8OF0WbBOvv4FQYO+kFYavAcbB+IXUO5ZBESIJarAD8ibe/
0LHPizhlo/1e33DjLtUc403SBpJ//UVFUt9ckYWfhbPGbrhyk+oUuXLvrFjf+tlG
np7rqY5RxYvJnr79szRmVIFuWhVLbV5tCyPK82lzVzyhjbYrHc58WVsC0wMMiPs1
1LjLdShVqBp+429u5NDVnIKk+T52jx91Gassf4EksLm1VI2lv26ko936xz1GkAGV
MLAaqxT8LSSThbPOvQVmRoyyJiXcG0/bot8PmQP7Xbpu6aIXAOp82NVkuC8r+sjG
ZFKwBUDMtBvjZKZux/W4XTyKljNENh6xgtjwkzEEB4WlycN8h1OYUd1UDuCRNpUe
il9WL1tMy5dY1BJ/DdUYpHbIM/jGA3shYs/xZpL0tR2VJW2oImjACSzqGoH59iZ1
ghO36Fc8EzYee235XMefimOHua2RGS/ubBdAcWrBlvWSuHwTi18ZNFfwFlgqDs26
PXNYNzKhbDfGMNQ1Fa+qgpFhU82copeM6iyvFeZKARcegpgwTKdICt+2uMkWdVPh
BWz5CqjdmE8CVBUt10AkKfGN7dr1Ygl1JvuCRNXuSVF31hUgfwh1Km6JCsIf3iSa
ukXIYJVfpM4HOlQE8XF/DueGBeFwUyPPG0n1HhNFNt/1AMWDX1Hhibscb/RUg0L1
yL7HyKRsQvi0yHXfmdbn/BGINwnKBGm8JWcibp6OxPpbSEeYd5ZkmMumapa6sSfR
eEXNB2WrkvC0t6fpL58sigKMsq6R9n0s6/Kj6/ktQ5OnAtdcXuUwwEprR1f9hCw2
yQWRWwoDWxsTdgQsijv7AxBhrr/s7ueHAW9mqLiDtMKczaroxEUqsUjrh4N73YYb
rzu1OQVQE5lTuJwP7C2U03JRu33whN97ixl9Te9YFxhEsSIboNBQTd662omueg95
xSJgpV8eAvtkL23fTJpVEnwpn5p7BE75AVa0njAkKO1kWvR3qLNtYPSJHN34EGKG
pq9cqZ8TUjh+kvBI7dl8Z1r1stFH7rRtErlmBC+ezcAtobueUM/a/ecX/md43kaR
a8cOKWmtd7aayNph8s+O2h1KEPqUujPxa0CPFU2xKJNYvjj1afLIISVGC6YwV040
CGuNV/5SB6WdozFQ9hGdbJ44yOd4kbMA2dfgyb9mNq0TyQRw4QyIogXfu2u1JSCf
Zs/foCfH30QuHjOZbDRUFrqOXxxpgpBGsSj05UOy92fxylna+RjamVO3ca5K1El0
NAqoGyaIp6RQxQWiQOX7Ruzqz3toTOMa9nuYo4Nj1EqYLt6GGgM/UnvDqbJurzaL
NR0P6LoL3rbihFPg5kUu+3o+8sTaS6C8hdJ/hertGyW4ffrCmUKEt4E42VINGLVe
4I3cGrjdFRv7LeVexHHFBuZcVTdzWEoMKQk2VQ0sRnYetWR5RnKdtufjI3D1sFIL
bQ8kiRL25j9CgLdAUbTnkj+Eru+UkoLBTrOji9Mhfhyk+cs42S36F0qVuEiSmPuC
BSiu6FTpwUId9LjV1iy/l+FjYJxklFTXcMkSIzagJ8zExQjaf1feyXU8090Iu6xe
V499u2sWDIqDC9ahDExWEkFMS8ecM9/gepxcKlY1T6ux2EHYX6+cHyn0kg6BAdWS
mJuK3ME5A0Gvpxdp5tseFyOmUgvg9jAkSNk2o2NO994wht4AnmBHivk4qRZj5KuS
N2HzW5OwOSsUEwjZWyKSAff+oUTncPUQibsFagzQWvENujCMIOq9wipGbYnJmHjs
dMBaHnvd6dRm5R6cKp7tc2K7YEYGdvM1Sm2a7AQsnT1X/c+Pl0nWC6E1vQshe7uf
CgtfN9p13DTUIXdu4oNG/lIgA5JjMQu2YCSreUG5ZojojPErWDHGu92evThV1vQJ
kXmKDM+AklZvwgmsrUYMwF82Q9IMOHIP5mJeVqSGMimSV//E+0P6YoWr/t8NNOhW
CI19rdnLnT+400E83KrpCEGT8ATLzBupo+vICcNPMThcOsFzuY5zZaHS13FYjuv+
h+xuEbIWdgnx56M1VdfDcskz7jyCmIyPJ06DW4J/6AInZmlh32Sz2fqI/Bjrex5l
uyiluh0tnhQCp8hTcT+qSnqWF1/zUfizgM3r1igkik0ceoXQ3c7bZx3sAzfEmct4
v09atl08F9cDV89jRRd+si0vHHN4k7DB1u7pu5q/Yq6qVC9+5SBKX1SpyWgVFtRM
n+g0y/J9rQsjZjI/9ObecwMaeq024AQF+9zqVKQ2LSJMgzLJtranxCxeRBfzJLwT
Q9GZjU4eEkW8t6jzZ3p28PPSRZZhznw3SYpxUqbHuimKPPVZEPOdqCBfnGpqfCc4
Lbu6N2lSHEOLNK6qv+y5vXVtc1lotazJJNN5N+hIGF4soLzyXEyI+Izoe1isLzKi
kYqAmkTmWjom/iqOaY3xD3I/SbOC+ExrgntR5ykpnf3soNIxlMvIK4FigUBqPLG5
vvR0Kls5x3rkalMZWkhauWm15gH0V8P3hgrGFhRPmlAM8QL6uUxSUGJOIlSYrSLQ
u3XkQqGMgfZbCTX8ylAVP9XyizZ0CNjkUjKDHw+D5XYAvzkH2Qj22pyUSmLPa0VY
tnJf9M3RIuRGUyJhMUtHb+ZvjG3WYYVo0bDYbcN2ml2dCoaRP3Cjlu/45yoy6VLr
sVMY9ATs5uH/H/HuHSfKHsH854ZNrArqmlaMe/GYgTs6DLTnpQIV1Yc1NNcT3eek
sF29dmCJkzpHA+J8flzkYqSpfod7nUlzPxoDrQWSQAY3p/6yfYFHURY/caSxW2L0
SaTSMsdYSVAQv+IIX7FgNISwWjL9XhjR54ZjOSl9G2ZGsi0Ysj/AhdxVakTVAccK
vxrTQlq8SsF0e3Lm26MXE8phES1byqy/Wqm+7qFqHs1yOmnd0ZG944XRfUak6qR0
9OI8dkfjiKajmrESElExVbP0YFOucgqYho0AQkFz8erJ8h7JfcmKlM5yN/818+I+
NVkMXLsnCSO7DPMVY2ILNPxle7zG64Pl7u7hd8ITaYQT9XV2kSyA8nda/RVwqRGW
hZ8lgw9J95ceqM9gg0CW5QJqjq5d6aDwZWRgCYe5m8p3mnvU5EusTpBfC5i0LRMD
wRMthOF1cHtAb+jwOUKUG2+5rbSEMZXOJE86fmoGI1uAuRCbCj8pNTIxeejBF70F
/zVbUZS1zmVOXRYfo0YUsPQCOOofRNNHUta2C4QDH4ftlD/WAA+gV29OqrQdzfPy
hxIlZDobs5ydAMNw1VtnpqBClVkYc9swVhllePf0VaT3lLDRnLyBtLIzvuP4Qgea
VjD1Uoh6+Pmy7riqV8yT472g8YrfxPfS8fWTjdI/g3IBBb5utFLLSrHZQttqPdVg
Th228smGt1Ais45q1JtT6ge62G2MmjQxCr3C3B7KetPB5WFSVwDTeA2+x9r6DKqX
a7o24en6RrX0rqymetbBSxHbDyxwD1ZI9vlFmOg5RnvI1nbEkMyafrtQW1sp37bq
2rdPgAm/NAtpdn/ZpRU6JDU/Lf0c5Qu2xhr8tIGE1XtPfWE3licPiqhBS8Sp7Z51
+a8rlXqAxGm594uizhncTCOYnKppnEIrUsj8sBt7LWCbY4vEgoRKYee3jCaYkm1H
ZiF04eeen1GuOxkgyaLkx8oG9B719OyPBaHPCfjKbgRMNCzEFMs/GyYwzoQbyINQ
RcQTMgGOuuS3pN8egZ06tzugsW/6MgTh8DuRuW/4izAmKOv8KVkcEq9p7WL65zlV
B864lPjK9FRDXiThKIuuB+OH9Q80Rnp27l1z9D4e9fjazv+cSs3UHHmvFkmUmrWq
W7e0apVWogcIryU+I9eo2LGcfQ2KBvCS3V1LS8vejNYBBUEVu8Vjtv8zTu1k6mPP
wD7sHn3onDi9FMKxZz2NjyW3raowF7pubxSXZG47nY1vkk7z+yMx/zNX7AEiXFyE
erF0TMt0rfVSPPhKC1tIYt1aZsef+1TYzlpPtgzyC3yFPoac0n48M7vLsdH+tElG
CW4jGHLTBM4bHT96ApoMmLTqn0fbfYkt4GuYgM+HyZxBoSW0mBLXow1z8Y2Pm2SF
PhF/MT51+CiuxKz3kZ7cCL/u5iZ1XpyeNcz0RXkiU5I=
`pragma protect end_protected
