library verilog;
use verilog.vl_types.all;
entity clk1hz_vlg_vec_tst is
end clk1hz_vlg_vec_tst;
