// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NqAEAbpcq3vMM0UlnQU5KxKhNJzUMW0U+383OG+MxM9+xBCpMLCAJ3Sfhw6TfJvc
gx//AAZCyWBUajQXm4laV8hn4XVd7QOpLPQoiQTS2+NAG7fe21SJpNs4168bLd18
PdxwMeRXK2yeu4AR5lgtZDr+dNYNHk/i+KlZX+jXbCE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 85952)
gC3D01yu99e1023YVgHSDf5lbBnUQUYHayK/0iSMoxb/2VD7z56GL2PGWAb6qK3N
OVsT6rcNq+fIEAwYHGdjR9GtVK5xfs+EBwJVG13akHGTmJbvQxuAQl5QyzD7YstX
RYlUluD/+vB4Di0RR7ZBeCTW9fGbSOOnb7fAXEY5w3g11X3mCVHSIdEQflkS5mFP
AMH1nYn21ditSlRkNbUZFquRZblkVBqIX3Gx3Edpn1TKzu4DZko9DcZR7phe+Mz1
r5/5SagglrXHJ7dMKYZkb6GMl+XgtDDi+laC6ZA0Q7OeyoOf7ZR/veOKzpFAERZs
bI2eDFQjYttultvMgRg80e+Krd+uGo1d5aKetgReovnRoRG4By6BOQk7oa+BYgwW
uidhbGSfgIaVptzJUmNirUI2zy3RwLgoaTB7NtEx1X9KG2tG7wgbiNSX2lrKR5Re
3ECLMvg2lI2f+aWHpeePbzELgZitbJWHxF0ZCaTUz0LtOCAwIHc1yiRDEfLQvk+a
k107+dSIheSaFDA9pxo4q6EOqPqaa1PHEbQlk558FUBz6tBH8k8a/pUOxnAb7uk7
P9sswU4klPb3Z72XtLmyp9wIyMjoDbmi1ep2fQpYcJzhtJuAuJHDdq/3rwhmJ2OB
SVRr8ToySKxopNRhz+KFEXc8iSKOTm8xynqrR/6VgyScGxzigCcMkiSejwmCDXJj
3yaq+BQaowc6A1lR7hgUC6FJWa3rqknqIbrlvSEkgl7BN2bkAh/ZBBrrAlP9SA90
lf1KreZTaunPAjsQF3F1irpWOezMa4ApRbcoMDY4ADySfEwbv936R4WXtcHDw9i3
ikoL7iSyL8puKcsyZBhKOraMMytUojfrYOzOrMwcxMy/nfcFOPjdMjxkE1twxuo1
MpmCFKyQ0GtuBeoEHi5Szdkdx9xqL0vXCaqIhfDHti3XAPs1w5j1yDYtsbQVVsWW
QqZ1X6BKycOR7CzjEkow8cghjHaDZIq4wd+FuH6+FS2Cu6IogJh/GU0eIy4k/jei
Zhw1MGgNVsZVa2Wt0s/aQpO8QiV3QJXOaU+U8IaYx9Rpf3L1OpYUJ+d+ApurnjnW
DUIZ8oOuRhErB81aJooij69LSgJsQx1W/n3iAaCc7pmavQA1a+fzukcdYoakQOed
gRa10GSEz8A88BIZZYl7VDP8TOkTLzoyOZvkCdGlnidJSwiq3wMRjRAWZpyggAjE
rpa6h0xDa2R2+ztvMD9motpycRCL6ptlXuKEZyBxRwx/uCVhakeTtljXdR6q6kt6
/1X5yMBqrXaXKOv/4s47DvaidNbaEiFuhBHGUjocRtNZRdqTD1mMWXPDUwrAiGTC
SCnEPvG2fWb8vTZbnm0XgZ1yNPGnQeIpddhTz5pB7NxC2oaTpQ0PlFwO4pdOVBED
ZPwalbcdjm8xx2Q04bQLkn96j7cx6CcSDHB03GCgWaF/FEt4DCuk7nu7qch2Ksb3
L+bzNVesghFx5I33+hKsyd1skmlrCAhJvb/BXMAgcNh2ohlchtGckAo7VRKl6NkT
v4wtbTZJ+DjlwJ+aOzPepXSNb3wg+xda1F0TlX+hVHIp5JrI8A68k/tmWkIPvuCL
rgrktYzje15NzbwRBdYYgFZzxAXyO0S2Ddq19x7Om8gnIfibfcZHLa7AZPusfIt0
cqLTWWj7KpFgBtxeUwEcagw1ObXfFb1Z8hTmxKBBvxpJ3CIF2jOMgcXTeU7RedtA
bHEjXsZayz4Qw211DKI/YziG0xMuoz18R1p0mPtQlZc5ntHylpHq0IQ8GiLZg9e6
YCwteUPCeFigHS9Pgj2tiji6w3JVUzagt0Kb7gBDsH7b16Fr920nlstpYT9GhQVs
yi7IcGClrcwfSlHkixHPJKQvOkejT6mt/5haLEN7xfTErAkD8moK0NO+EMn8k03Q
uQrf4HSWJwgGGqY5BuZa4iH1mdCSpDAKGn6L7rJqMfPuIRVaGxT1PCch2LXT5w31
BtIdSM+hEQi6KBIjdjXvv0P8pp6AIym5m3Pd4h0klfVdQT/QzZ6ZTChSg0+i7Wpr
3MnSlqWrZizw345CYkESvERXzllm3VD8P3EoFIp5xrRulojJiNxARtZ9+QufGOtQ
LjBQVDJyr8ZXyIEf+VDXZRkw87LUt1c4aPOzXFvJ+pcDKXWInsJG2lPglmdt+C19
1Z99aL4cjBeiziUXuFjTUwWtTPgK+5hbiP++AySf3XAzw9CcnHbfso6Mo5Kuu9Yt
AGZsTJi9Xa3l70DBIjpoB1YJay0xqxzeYh+lkcPMOp5PYPxQLH1TpLYl1iJY/x4f
KqOA8VpyX3d8LcNVnaHmQrwRuec1i09xzRZg57vcDfhmMHvlxwoEuX8WAprU4Q+3
sfsDsubfHrPdKbVCvhae31SoZhM2wrOvpQTyakgxK6lST2jsgxYvRniKpHUkmoUQ
wUAxBWVO4wNlaSSzqoFZAjR781Q255086jbbnaPWdpmgD4Tz0UswDV1UsBLYcZU/
HqQcci0F+OXyJKU6PEYMaGOSOxZ4GQfbeAXZsNbnizT/mx5ZCO/qCtUeeMaVnTzB
iFcXaHblb/NiF2em75nWPv/rGKPwjAVxh4U2Q4g7ncqEYDDIsMWqGrfpeN0nNvDs
g607fDLFhnxEIF18hnkXF2xOIr2Oq5e80yCr1QagIu727kX5OkDSwKyJfp35eSse
IqKy6I53HOI9661zQwYujxYxxtcG3fMJ9KsJ4Xsx8aduHZE6hNc274AQF4ZA2zf4
GwfIArBGBCZbe/lPBhjjjA6Gpq81FhWTPPqqjPrT7AL0ObCfpnPObsHXo+gmLGij
FMo4kHyDQHooWWXJEr+Ug40bXb9OQYrFX5shuJ3YKsnsVwsYyCq74TWMBBDqKSsu
RN7XNNuWRVI3qOTyRVXI95y43cN1Bp7iMyHnfm8/OQtFWM47XZjQzRmVJV7AdOCO
aI86WCxmCsd2+zXMAWY/14Vmg/olGnMSXtb0C0Tb0KuaeRW5WqNMQMfM80d1oBm6
4GfMss9SNA1p536oVoiF+KvKguem5xyzFCXaKkbuUs1VEdSSei02iv6oxc1HwEpC
89VVfxbbq1pXSVkS7Lqkuu/LGWMPdXJ5iV/uYUDr9jUEv72+VYLLk3J6Kuch7Aul
JFQQk9SWIF0EN0umzWPn0h7Qs9+j+P8Q7XaXfCKh8sG8sBwc17z6M7mP510oX+LL
k/mxzrlRRDtxNQI5F7Ercc7MuYFrxmOZDEqG1jLnY+08kJKSj9KPH39UDAPFu48r
GVjM5zTODo3qX3Y4zp7zPYtRVBu/o7tFia39aFdQ1rejt/lp/lAaDIB2qIBqNysb
j5lz+9t8Ek93SztpVPaKiuRrGNVKneG2ZGyNuZy/ef9/oiVOSuFnmeTSuA/U/Zx3
dJSsLnFq60NQvPvP4mzmo/t4PvqdUH0Qen2omtdem0CU4iqkXyNW4o5ZWmt6xGip
6qt8YOQq+7OSN/17teUt86t3ZhGRRIONtKkuLCvjqhEsVCO86v7D+tWnQbNivEry
lh7tuI/QrMil2ffuyW9cCVxlhZEFFzurM/B+W31RYK18JgL7ROC5+z9kIUO8szs1
Q5dGd1chM92tIsPKfqwkDc8vSqyLy8XrHHFCQIrg7QY9jETEK4uZirEAcgzBc9yZ
+Tkqja8Rd/K4XzgRe9INRSMo1NtKZ+0+x2F1HTu1U3G0kjDtgd8h4n/z/LdcZ6yZ
/mSB6oOGEOm8uqnGTqUXKROfAgzyaMgrm0ESZumZmt6MkPQfY8/glnNqNuYbAHlA
7c0QS3PK0F6Hy2rAG1VifUCefd6s7caxJYDqh0MFi5qA//yJofhnv/6kkh2K3oH5
vrFUy+cNvYDdRdtwqV1x/o1RUbZhOMKLudBd88YDRz+sTTSSKRuTECFYpyTeCt0l
gLBRWnNa/9K3qtraNgCn7mIZvPyoIBee9PJ36ukmLWefoAQbREKmEZ0szLt5oHRy
As4Cuvv3FBp4UCvJ4EmF87viJx6YL1h7BR6CDsevQOWUFT7bi8CEndzvN2Z90Ez9
LGcomDL05Agua6dpRA0pWiLlfJu0edT2tAHfm1YgjxIdoThknFGHryO8JqRkkiNZ
aj4AcJmYQU6zd4yQLPrN6M7KdYhCCEVP6jehH1mo2/rDl2T8uuk8Sj7NMfGjamWT
TyzAcSp5eJxotUouh0TPdchjYFWyJbqC2QrQKkOz1SKW5J5516PJFcSMTyAyA2Fd
5F5NDq/BPfDn4Wg2RxsJuPBqUOjKs4dMPWi/slz29D7RwRpRChSI8l/ExAnDo9C8
Cl3V7Ep1bh1rQBaD4h6xPaSTwygxNtdxUP1RybKCe0vgSBxcAFeYCf+GM9NCv8Tf
dPvUR+9G4i4sQGX/4x4GXFc+dXCZk2iU2LsGjcr/VPa9kVTKv47sR9bFZuY/dCz5
qeA9soIrnj7qODzfb+OtXvjPeP0PS4IQmIjaObPzEY2pfyZsf46ZmG31Ijh5SEyQ
v3HWUb78LhOQjxL8hINfUk5QUqzsZ1jdaph5AQQv918Iunbbpy0AQ1WHnOJj5joy
KKOpNJ+2hzPUSAvcuo+bnAQaaChFLT8+wjV0p7BA5o1Xcx0Wu238mMnbNz3ARxmk
s5LuN2xsFUcQcuQr/Bu75G5wLGeRglstNhLS5SLEkaiU/3GR8nQ1WnhKSAuEDxSA
CDY8/Uy3+4/FoP1WLGM9acLZJv6bNFrLYY3asj6ha6y1c7mNQDgnTUc0Eafrn+vO
JHKowvWI+CNAxRDj/7KGoip8Ny6AVSaYH8RjxRAVFnPf/tgYOWMq5J6jjP06LOxb
FemCu9WPz0PGtjDdzrBTrb+TuwP29CShjCLklP2+KrwaaVN8JDLL8cok4w8LHC0M
GJXuzgGYKU7FKlE2c8TY6UQJLyQMe+zWdBfb6O7lI/0Pg7L2DCvqk3wyN6tQPHeC
1sg13BKWeAsaF8a2olTiyK0NYR8/AbJYewTJf7eZuHbkm8KSgSM3urom+IphvmsT
RGNRVT7gbHNEEFzECNAZvrf4ljCjzXbZqOmm6hTHhhHe8pZ5gyxJAPrK5kqPy540
gP4GpN/ddYOBXnt3mGDLOlTHW/K9fXrDaezQOWSsLV1+jmurmlODUjG1fWyie5rS
6YhQJJ0+cWi+1IJI6us1wTCc+XxYgW+GhIwZVSYcrYLuxBS5AH8urfygV1/dIfjW
2YStG7gjBOH2K/Upph4V+pP5LXiqOEbbKY94+psmcMAvrxzqdx3COwZ7buF/ebcD
+zsmgRcT5Dof+CAo17OBBMkghIWkvDdcUvBrbfWsJ6NyZqndUhn78HmD3hxLumag
VCwCld/Nah9TjykWjyRwMsUZI2xUuu8hQJZSFK/+S26n58jTkH+ykN81isRdET8J
Ngiqjv1mbLpo/w0dknMXkDvQ0lEM1T7d8QULKbMDOQ/h/qb1W013mq3EHVgZTYhW
bpiouRqAH4IZBd+EEMxNuVSSURV5JT7UYprQn/SPt6xvHLtDRpXMaP6CIxB+1ZZu
nycFl/vPT4EzALrlprhJ6uRF9+MMWjWjU1eC9UbMpIeC54sRwmblI0XHfnLr66bq
J+MYPzDWKcKVFPF8uMTnDTQd/Be3MkTeS08FOm5m7twnUqOjf1vq9uuhSmHe4rn6
HsauF7iPcIuC9iuTVKpTmTk+vpCbEenQTCymCNjt4qzPV8WRoq5JUa9Kz0R0GfPO
98/+BUWFv5Gu2pEc1O5u8vaXKMVFdUVofbrKWA1W5+DAZaZIYn+Xo0KV/NR9ob7w
r/6/rcWsjeSmw7RbinPSDDDTpm+uyOEVFUrVi6NPYGwOxMGCHUW9LyR27ca7gai4
leAK5zK6teaB1WRCpPkMP7Ema3oBKlorYDXrI+3lZWsPzpSMDJS9YUw9IMY74h3m
uZCKbjQt9WREpHMeC1urg01lOOJlKQxPOlaUU2i+WJJ8ZmRhqKTNDBapKvtNSyPT
WFLPytzzm+kt2WPTJT3ZNBKe1sgu6Jla06CVF75eDPljeBKbZuiqilfdwT9ipAnw
HsVpAGCqyVA7z+6tf1L5QtQCi6Ij78CsfeDtj64k7C5Zj/nqrYKtnwZSZnx+bLcn
Y+rXo2FrvbgMIW+I6BiqwqyspuShyRDAVY6Zj4vzq7CMvID5LMIlxGBkTEF5Ar8u
IaXfCy/i0c0OK+bnaYMqOnBqTWl76xnYfVC+Wxtu2zajQs9JIK+b9zYtW6AQVbuC
5wFXH0zTU4vz+tBnTA30Jzzl7yGxj8Dx7BEvFsid6e4PUGz+o8VaO8KtjprDqI11
PIctAM3P3c+vbpek7NtzNxiBewFw1/VFGeJ0GXylFce3+cjymb5L92DyjMHv5MUd
0h8DaEw/2IJbVxKt87AyxuPwHv+6n86GbGxvChqCUb/IM7lQGmneSEMfAwa4pPmg
aGXl8JR6MbYsor3FJOA81Z9iWwv/sbMGh2S+tQ7Ifnf2c0AE7hO8LFbtTFcoegij
yhTvsOG6RoO17OL9kK0S58AMM5Gm8xUrF5gWyvDxych8sf8qksg3/YDBs9f45EOQ
THXPDjg+Ywm+2ZyvqOQH9sx8Oci6DT+F6qnzJkcTdeTbGwQAu8Kk4XRRZ3eJVCgD
hX2ddTo6bx4uILm/Rh0OxdCcchoz7qGXfsQt4glTmYPv+7Z3ePCEv8lrZrCIfH6W
GzXcJPqJw26+GVjWvL8ygbQlyQPoAvOcj3DmdrFpIM8LG3jAPR1UxgMTmNG0EeGf
av1XZs7ReUwpSG6SM2BMSLY71PvyhzmmE/jyp2CMFrYifwTU0N3UmpxiJPShcI6R
AFQHHCF43xIbwPr664iz3s8V3LjauvIY8CWE/wNzTXjsIyDFc2Zx026s8G1Fst66
i9chSf9cN9c2FrxmrJomZuw9TSZdWRlYutAwSl9zxREirnEnMrWmIoOY4NT4fYq5
5dEjW3A1TGVH7teLFo4NzljQbToZMzUcsG3RCYjUlNmNXtvd8CvMcEeHnxaS/b5L
JMGNBSmJYGTfF8dg+iRqoMySuMaiLsnTrYxC0ltp94Uzyv6+SD0admHBJW/UD4az
KOsyZOKfIBSK4I39mZrx5bxtQrEUNzAg8lGXJ4SGidQx32Nw5L61IMi3Mf6vnWfk
j/t/+fEVAoqhOkDVyWBq7t+tJ2F4JQ9EGOQQUKBiWP2aN+LGz6YccHV6OxDSXrx7
kw2ZJpPI8j9Ebw1UJmnJyqm4tpuXItpZeUVp1JMpx04a24NwVF8VwpNyJBL1KrSf
Uu2valux7Aqe3zY5ZOjG0Il15VoV9BjHHAJE4knhwKuoOj32DU7ZZZcK9znqDtW1
yEP5x7nV9ECmGRXJOA7qdBVODQORhE+SKVscE3CL/HYai+YcZZL4SbgCw6RQl5g7
xzEzIECYYA5or3qZePEVdOxrBkDuNN+VYAoqSg/PdVzuwEcgf2rAQlqsvrmZ2gor
v3LpeloX9x5qZajEfNgAmbtGGslzbMkRgE1XweNHbicJ5RQRIYnQ4QqRszIlbQim
efmOoU5pQhLxT2lw9cEqLikokikwCDaLfO7VyLAhPnQPdGwJfF7bsMRKaQCRdMwe
f3eozKPbZ8CEAgwu7Jaz8YS9Fh8yGkqNdUeVI0XVsZt3k+krIeCrimOJgF3PGA+K
zV/L8ojuXxDyfQ/VYqKI0YoYkt3QvdPXrdlpGWN1UZtOp77jnJUMdPYhw5hG+7o1
IQmvTycdo+oLgu+fvpSwWdVoXDxFjdCvVgminK+qjqRmc8Ua66z1+ZuSFnAmLjXs
ePTk7kDVrr/vOKwVWROdXyxTyJSyivvpYMp3Sq1JnFKT59i+Hh7umqU3B8SSyuD4
fQkSjtJHysn/zTgOwQNPxvsb6oLttZQ7xst3pT88BS575ddoS5rimQD+KL63eLGQ
f3IY6G0mQdhz1rEEckPTNqOn7XAkrbMikJGqztKmBcs3OkH5WWq7Ba+lOP1t7QND
1G5uKsqL85nOBng4krufa1mLBlSH/fMIyiw3ggvV7gAIlrqLHxR0ZWarKj3Dv/a8
RTZAcb5rwrtwrJ8V08Fd445H9vVKul/SDOY0Wezu3Joly0qbWOx0dbVciqAms53t
5mL7sF10Zy76ZIHnE/0WiQZQT7tELzXC0BTuSDfCQddt4FfDHm4jJaf0NBzQISbw
6suPeWxEiEo9Pn9H5biLE0jdBIv9foA0+oRA8PRZRHI7Kmh4WkdcCA1Sxq7jmxdU
DBldwFP4aa16JI+ejEAM0OZVE/xqN9RUC1aKuqh1WfBm8NStDIc4Qt7Q3x6STaf4
xe8vsBNCcbSKknElZDDWJrAob3l60h05SWclIPe2vED0A8005GjXg+FzuTZ25shY
gmhVygCotX4Kcm7aNNDeZVUnkTkA/8aVcfmiEClj51sXDyMJi+DK5MIxxeyenokw
DVCUT4PM5LZ6MOmiXbxZU/aUSptkiIHJ2VTi2PXdvpmlTX0Kk50BGur7+S+zhJTp
wvCWFS7jrnVhIeJKgE4aTf6NP4y8+tseEwK3KmMdOGN2a44U+O4bMXpbk49Hcv03
fbYFx1w0TezJSF1+7TQwUGA0kM91evZEt/0+L40SjqeQLRD4OwoQesuI4uW5ivP1
SXKS375bvF0hn5FiOJLfnRUeqDTFHLrYeEJ4D7JIjBgOaLRBwioz7fAIfnlQpwaI
WQvGV0OZM7yPmV2BXp5nuFbR1Wi6e6LYYex0VL7Av+rKom/9RXP3oLopjNcHbvVs
9TTCYfjXm2FwjUhwqCXRt/zMcqr0EfiUQ5yVyVgDIBoS6zLeFm24FNA54F0/7GSt
/RaOC2bkrjgH7x1ZSuDWmg4is0xJdxq3hG3qV3QszUqmJAApcfAqbJSisVX/9wNB
DRIt6ZiYEZphJazXJD6Ta1BmXvKIpnNwyRbrBuhuPysmPc7sTDmECCV3EhiDrF0n
+429yA7GtvkiigEsPnOTbDgNFKiAqa+2wAaoAzAsRMg/NxvehOi0kCsmouC3R+7+
qcp0w1kKbjHW+Lrl5cLkoGrZMHOLauD3mDm1CH6O79VezdsXIteRHKJhjIlQY7Y3
p8BzABIPwWslHBqOH5zKi/Y1rPugbcDg8csSTAg2f/VO372o67nHS86SEGI7MCkT
5n4GmNfVLISm0HGJHe1WW4EqFlCn3jpyhGjYhZpKtImVdRHzas/72PYjERkr/Pav
nMmkeUVVyBl144pBtXUiSRYcqOiGqMMQePb9vHk8u81wypxtoErzXwex8EnP0YXr
W5soEMZ+6Gdd0fZkmqeyfq1vOIGx7CuQp6Z4y/Bn+TcCWOSPkWR1LqsWND/GjDi8
zWlEFv5di+IC9x0T2B+bshHXA0zEHS0Spt6drmoOO+dxZOfv6083oRK+D831oLKB
+NkwglLZ/th4h0Tk/4n0G/5xLVDU9DeHleRCjmx3ZmBt2zJ7gdbhRkDkUgsEugy/
3E8StI//jZ4SiLpSnpvSq+f5vR780/Q1rdzB0c93v4R1kd1SyVvBt3P58am9BcMY
gJLhV9JlmlUfshaL66Kboa39ldvU1Fr59/nv9W6lsyJXwlHp0E+KtBxpQg2WKHWm
kUvH87o3wYJLokDQTaGtNBPk1njo1u+J09iRamXatm96KfXKvUHFTNj5hM7YU1Fy
Qu6yC71//7B4d4otxiXMwBkc7lFRpNLQmIVOQyoRRcRDEgiLi6088lY7iO/IClhy
YdMBhDDM+JZFr2PoOY5EMGLP0p1M83ffhX3uG5SaiB+d1ehH43gMYf5Hu4da59TO
hUb32GemXYPNCmt6MWPKoh3BYbBslwYV7WdflGZpfKtQWSmPw2QJVXo/UcZRyvRS
t1MuZXNEr6RZeD7QER/VaPtVSlrDwzj2yoL7rxvTOs9EiJMlslR+dchb36mH64vr
CGOyvZyvstS5gkCCy4X0H5EhEbp4rUimFfTPz7dT5a9bIEK1oY26RkobmD8m1JKi
7IJ+eRkBgs6sZFOypZtpwoD8Zxvg+9ZzCfGsc7Q9T4nvZF1ubJjIAcXl0SGI2Dj1
qKjQShGK7YSTpO26E7kebceMx78Jb0e8wXwhMClpYsGqai+wxuooAAuLBzl+zR+8
txixVm3IZyJXHXSC/32ARdkXC6njS49PpmTYAT8z0orOIFimeKMdqTiSu2ZjVEp6
l5VHmsOqTkOn5+72kPak28ttCFFjn3f+XhZBy+AJw8eang/FbH8pg9239+O//lLw
XNhMKxge4ud+Eq/Cgz2QRT8WebxxNI5Lbn3WLkS3je9QpNTLQ6h2kPZE0OtLNyTi
mcAfvLvoCHmbGwKBmZAt5RfuDkk8c5F7zJgejTKoP0UcSTFloCTCyULuy2Ce8mpP
i3Jjb2MLgMia0Pah/pHa6Ke6892RkCusUk/APDB/NZk+/IYQ3zRbVuxEpSDPEKuf
x2zRA6xqsclDXX7WUQTRDrpU+YlHDl5TUMoM+FZcW0Wcv5jM/ATEpLGj0gLM+01v
6BKWIuUZ8EZB7rUhAs9QD5+zqIFEjNLyQhLTSuuLeNL3jtJUDz6mSpl54KyvF0L1
mQ0H1GasQisKqbUksGwTKB0/3/q8C3sDZ+A3eUWW5PnsWWoRnnveZi7lyDzcSXc7
UTLeIg5aOf1R0MdTylaD9cIiaHzvWTI/xQEDSKpK+Y+eBDgxIgHveN+ma3ayvlmL
Yp0uIYIld8Cv6VIeRzn7NosScH1tXTng+HroiSC/wKwvMYe2IWuB7Pys38FLkG9R
C4Xjp91PEuCme+N6RWh649mJCQ5Kx8uoU3NnKEG++B3tf/wkxi2rwI8lF95GsrLX
qKU8JfakIk1Gn6YPbfWLikFB4WB1iICJuTyu7Lc3V+7foMHrwu0xOwSRhl5GKSRJ
2yWi+GAoPDF+oWeLx1AWeYUqedYuyllshd7Yd3YMW61q9YhLZAeysvdX6twaxCdZ
osSBSk3vIC3un8l3CpqWJT38vz5E/OX92gHMIu7vwvIb49WnQYmlyFD6pw0P2bFf
TjDMMwcPgWEDek3UqGxNzk6KbpyVXqbX5GBGSl8XcB8M1jxVZRGQXXHuAgF1w+eQ
k3BmaiQ3LSxKES1IG0AlHMkyrZHbnkcZ/Ch44z/MTeTco6LKy6gkS6c7q+AomxKD
RxmrXiVKd7YlhAUVlUaKVMk/TnKK2Ktsasw+q3I72/udQE14IfdboKzdawkAMYks
s5nq1kkWKQXrOjbfVqfj9WboOt38zxh+KhP++4xsbgy4R/uh2FqoBGqfXa5sp+ps
wH/oEQyrRUJ/r2fhtimhsCyynu+AZAyuMxQekGwJL82zVB7v2vnATUfRvZAx6Mz9
9OSnnWN069RVYuNXljEaFb5b5OuRWnmtzScOlmyfRYPldv82PfsIyHENly8x9S9C
AqKziaXljAgZ7+IWsMLcqjbRYs5Gv8Iz7/tCmpFYedF2gymoPqHG41jNQIGPvrAp
oB03TxnpBcrTx+RksM7CPopM3vwP4UHWY2aa0FwZbZEsiceaFmZ02hK/Mi7Mi9E5
XBQUlRPJZTSqfQfYM+IWcr9Anv1I4HKl5rmGGHqnZ9eccL5/paOz0vurvXNcVyZZ
m+DyWs8jc/d6jAkHIj7rGbyfcMLYhWkWcSE2Ohh1kvFFsJ742PqVPfuNPaTK/oOZ
Gd+7KUZmfYTv0z8ER9UL5Hx+mraD0mASaoRAnD00rFXX0Ic8HxJPU2HkaMUdkkzj
ZfenxIF8boMc/1KHr7BT5yO7YQe1njXcM574N/zBzthTH10wnvX9Hqph5MJxiR0K
jFebxPl2uJVVL63pAyA+okDiK7qt0H60G9Xqn9QWWlVEwX6lkwwXqrTln4wWz6eX
PYDeQH2DIO48iPAHz8KMP3AVFBmzDxsxSPw7eBC3qwoXGCe+QKnyWyIE3qQUeWV1
lQz18Nu6KEteLsggnpcPgkmmgxMXyRoOGJzbcD0TElR6RsSCrjrHXYdYqAgkL3qs
Aygwv+KxTARL0alBjYkMGSGElyZ3suMQANDgp2b9BqTjtrY00zTgQUu8PfxG0OZp
4/N4U1fdZYvdXl8La457T5i4S/vLJI432x3kWUXvKFe9C6HLgTCOZtujKMWSjTZ3
Uesy+WfsXMjJUvWNsX6p6BY6vpad6mztAtYHFbotR9K2kx8lsP5CJOolkt/q4spH
7mdnCGYTGfgZS0mFenyJQ2W1FzPHvQAeAYeoDufDdvUHYKTSWJkSLsmii5lZqxv+
BoEFBb1hl0ri5VJ9hHyh8xs22RsSvttkv3J1ILCI4QLLNSIvEwOvAglfVTYUUVzO
jEPZpW7Mw+Tgk3uIgXlR1ZhBzZTwajQXhxv7WAzMiQhnw7BNFxFNQ272wrzlUkj4
8GNHmJ30VjRCo3SJJCchq+QPRF9+48xVYbIc+hW4WQiIUxx1GfL4wv6arJW5a+Kk
co7WvoLUcZBkWa9EZJAw5femXs/9e5gZgdqy3br7T9coo3ZkqX/Z9hzr8OFIbTiQ
OJnUvmylDqvvIdbPm+DMWwoHZ+kkKfvrgJ3mZr+P8R3FvuDTZzSRYk7egYtVi5V7
w4i/d1ycIdl17mUi8uGh6xyfnLGit7WzYHnRxgV6vJhGQ8y+PCoY31oQKI28q776
gXpnFmGq7p781w/Q470N4vmxQqF/4TCNyoMEtedxwVeWi7OXhOwWilnGIcQq2+ES
e/RD/+12PNer4Z3qPuZoNebCsEikxEqeVqO/iN/zDWLNqoMINHGo/wPt8gr5FdAb
c7mb/LeXi7s0EzTXGPkYdww+a0Dmd2Qkao1xbFxc7MkSueLZzFPeT+4Fri4hDhmm
4MRJV/62VOrwMwGlXkSmEBHlSPkaqgyn2/0m752nWPBDQMeLmR/BsA2p8R3UPMNy
4T8NazOQcLlcnlAEE24JId0v/3iNg4+YFV8CVW7Q363Ku2tNrY6PaCy6ucwNEiqW
a4f5PVRT8wt7A4pGAxxY6/6dhhwrSvpQ0KYeWZ9JfqQFSGT7pRqDaAlgNMoC7+VE
kOHbGXLArJNljv0ieerguOFvgGvfBJrXHUuv2vIdPCece19FjK9G7tQynlI3VSbe
3BWEl4ZaYVhEw6xSGny1mygus+sMNP26dHiyuBL67gahB7aLa9K/Co3ozctvcrva
Z9Dpg2T+VRT+WguZuai/mOOM1gYSj3PlEWu3geNB+tmbThf+NsXSaxgWKtDG7Zjp
OlQ/kyJmXtnF3asv6txHg/tAivw6PBbQMQQM73yMRwYQ+bx05YK4VWD0O93wubJo
ID8T4Aq1gp4jGuZtiKRaxt4eLTPoDFWukRZuLpojCNp5FnK0BFMtXHWkQ+UjymYN
Ztqhqg19vgk0mCDctXSD/BGfSRw4uuUZGbDmhs289gogxztHprF+PYrW52fQPf1i
T05w++DAGI5q/qctUbRBWy/Lv1GU3kY/Fwtmge2cMhvpYDGA0ur8gvY4FOF8i4eO
EyGn2oS4TbiznYJyjyUmPIUBE7oJi+ua7ZO9RiY0Ot8LtINuOoJHcFNGwy162mTU
eFaqktRB4Pvu/8x3P5NteA3lolb7DwDVs1Jx67S6l5CiBt4wNafoDB8HOxn07cC/
Hz8FJL5ETlTDOen6QMtf23qGezS0SDh/20P64mLvNx9AjSutJFuhTckSHJZlOTkL
bge51fZXLg3oNXDoAyFuwdMTY3PRwn3vRga5SEVXQFFjcc8lIEHsoASlQWJ+HrhH
3isJ+JaoskNbx/AGI8BkwpVxIRQEMW6fUZ+8GULtXsyXzgXvNZaua2shfuyKGho0
A0f9LOJYBQ2baESIAVh+ja2ON+OkFDbKD/6L+wITIcIc76tg9arqNn6eGbU283fO
u2lCXTtE5SA1bZiF+NTDXXXjKlerc3qZIoBfhWVyLU5hPoJhDbdp6DJOcDDet/05
doGwwMyWaMC4zVdi7eJ5hQue4eLsUEJLWq5ae2sC5fl4oEIlM3AHpxYyKXY2gGRN
FzbA8FLkY2T4pIz9LtVlQXIrNC05trrX0O4q5myT5vNXFJZfwMNqj9e4+9xpbVDv
KywEdozcOLEo4HN3UiR0cqXJ13rouFYdPoONr6SUeSYynsCHPlFVxtF+uXo/98/Y
ue6z1tswnZfYSyV5I98SSpcorgmRHVxagP3aHR5gfQZrgH+iD0Qh4X5Cdx5KWWJx
HlafTQfWzvqihD68GHB1yVZBD/J29dl9xWRixzBB4ayuGJpTUKpUtIbHjuMvVqBr
BN+WiaSjtxKA1DcrxUSwDw6rSCuMwmUrCxjr9LMH7IJyDBy8j7rIKKBmeWpX6Is8
RK0KIQPY8NAJUgA7Vm9xJe1+6C3hMVBz8716dfpk4FPJzSCvMbMJUF+Zg+nNh9Jy
Npbanb4FowXaD0kpdMWWVZpEdBb+aj0ID40/XXkHuUecO/HR6uHUSYcEMkf4bVu0
ui94IzDwG8SdnLq0af+wtPy+je3O838ONfIX3RC++s7JRAw58AQrRMXW7IxWAZoR
LrQ9J2AHZVNTDXlOLrdxRPKSgFsfOt2OTferiHFe4y3AvHcUPhSbB93jEBuxYR60
ZaVmmqCu8eJVP8G3FS4xAHztm2LSNlQ5uTGmSIAz3OsVf0NsanvtqFzWCvB1Hrdf
IX56+c08cpBQ+rAkhxYMhc8js7ktEQQDT0j6GwnE3PKLT9/UyIizwbnidPTojRYb
RZLfq5VtgnP15W3BKABO5JOwrjOqeJvAVt1jb80sTXRal+REH6VhEzcWz0LGHw+y
xrHEtx+cxS1B4ECynpMicvHgpuFRK50gEYZfqQR2WVoPxNCRPE4JR9Tz53bzfsJz
o1SgMqCt6RQwZ4qiOt9iVSEO1skoYIPjKC+/nlDvVwLV9h0l4c8XVXadSlu8308r
7xi3vH29mqMjfY9yrHOkABGymVl5feIRVOnjMZ8SVIK3xCmC9zZtUCsY3vzT5Iwy
70U7CgiCSzu1ekVnKXX5TWMhOMKHyE4psUlBUN++W1pcMroVtuyr6LnKcc8LwIjB
DE1d3GqdYIv0SK+tw2F/2HA0w+iC+jnBfuvtHg8+QesooVUAC1100km5jgVz0KwA
3ram9Hfn0bPlPUGVGQnQi/3P6jT4pSNa6IYg+w0lSlECkwg+fmnLfIUmgHlYhmzb
VscUDVah+hq/c/cjqCc//Lqci0uwgAjBS525vdTTG2nsFP8HimHalpLEahdGNQkO
maaJl4+MfmviPRdThKI9m6zG09D3/myf4BRQfLqQho9oLehcdM0WlqCr0YL59hKW
EXrOlWX6Kso5dZQQnzdUCMMnVXZCWygqDrJXJu0HonFAFtXSuAA3JNDqtXX2tVER
Tllef5BLRdGMV3wknMc0xHVPSJ9FzQKALQ+TjB4C/jy4jr+G8TTAulr3YEdQq9+r
JwbLW9eSetd5BD6YTTIo2IHPC+culvUMhkH61WO6WT42rzvC0KZIP0/JzBNH7RpN
4yeOIdDcAjTi7pfqjuV7dIaFebmweuycI57ren/Je9vyxP7UjJ6QfM8xYvAgq+9X
Nc5AMvvzCaro4b7fx1IwO/xBAVG421+/rYyiGZA3djOWiPooboEaOAtZKxkDL19Z
XD3NgACSs6meMtiXub130KU36m0DADTpUEnz7O3RnMYLzWZjtQshcHhNTc1gTCFT
4tuYm/PR1/Qwv5cR4bv7vhJTGaLryjdz7YS85R/jEq94jbDFSvjjYo556gPoLQ4z
a15vPf9zXOr66Ixxz5OBc2p7HzXhe2u1Mc7BioxUBSPPheN+BqrFGMfDi2wnI1bM
ACRQ1EG25VJnVMGdZ8tgLZ1yMSvQ8gylragP/GeKQPNTSiofyQqqdmF4qBgD5i1Z
BcbdLs90UQ0uytYK4fxru7W8vDnW/chOfyGB10+URWBshGXwHQT4aAam/O78gLfS
Hzfkw2y/dVipVe5qy/vCEIQ9S7hkm9YZgOvvgZrsfrFUgLHdBZMN1D/1Y81UJDZ5
TQ1+JQZB6SSgcCAfJfeNLQj6LCzxAb2e61hD8p0yFi01kFHpOqXSfLqdE1tnP3xo
boescod3JMc+WPWlZ/nuz/0d1o/O19njpp00DdflIsFEerYjQ1ep/Y2a98iDcm82
6GJx4d8Z+T9ZKN681EocieBj4ALpRAoIuYhUkDJxMLW57Moy4JOx2gNQ1D2R/4RN
XUcoB6V73+nCBCo9fh9iGIwHflOjrflxi0XR13iJ7gNDlbqQA88PPPcvbjZ688Qu
0X8L+QL9Andm/mNY5tJdkEGmb1IERX3sPrN1f3bIgmtid4JMADX5sXTmn9JOcEyp
wNtZQ2tu5ajSsuJpowObRKEzuL905w6cq1V+ZXlmsGurl8QFXU4myItVNQQP7SEC
HDKXjgMMOWQ72MKqkBVnbe/44iaTWWIhyj/6F6CidT9bW5kG/Hd0mAjo9yz7vBxR
1D0V4Wuyp1P/ZLrbOHPTZV7brnts+V3Gl5qh+6wTITqAemSIy6T6pSU+ZU1XQSP0
u4roJfamId6xRj0bfyiMXxceoatiFxMaCQxEzYdrrDlA2sKiVsU3s25NeFdOCFDN
a2qmCCgj6QEbS9Xdwl61lqaldAWk6TrR8tkO5AZmY/AFIvM8v5YGSZ1/kMGgS5Sj
GHgoCoUY5Grhb/mzA5STn370WPt+KF+2yjHCcpSA1CctMyfZcg9lQZUlyExwME+f
mgaqxFRnRW8mQ6eo3jKhmLX3OT2HnZdTrv+96cGWd884UXytr2AhxfDHRLuPauIX
LDvEMn5n9Y1L4si7m5bXkIxtEYaC0pqYXHxQgZax/9WzauE3gQkl8WRLV7wSBIx5
97E6onCeg8ueVDicvrFyVqOwqJ0NQoln0cr3nopndH6Go2WDeU+cJvyucvi93f9c
nMXVQVg9qTdNl46SHhXxTFLPlQFPcHJKnW3Mv/PWedITY4BnxqPqJ1q+bqYwEnnZ
14Te+6TDtk+ipHLrB5t4g04iZPuj3Rc1KZRRM7T62xgIEJpIohlQsoqQz4RE0Y6i
EZUZKWUWFA0Nw2TkFc1r00i3BJWdWGdVzgTMwiBYGTviZoMFOU6f5B1TcxxqiOU/
d/ctRfpS+OQizYYcrX0vxGDX1xfwyc522Hw8z4ZJNMwkEzKA6io9F1jG90rPB3JF
KgFqz8rOOgr71/L3Z6IpVHG7anCV7gTlkp2oeMK1mVu6V6TuXOAtyIVrBQiAdvxa
lSOt7nL2ViYTAFWZsGO307QpnN01053VUOlQ9IY9O/AHLrdc7syVKL0O/11hbljD
hjpB49rKV1ogfFsOV5AlUE9eAzVGVhEw/U5Hf6Xmtm/MoLcKloc2lKTAwQb3adH2
sxvfiyv1rWDTzYWi6U26hm5HWnGCuNQTrIJdE4V296OPBfHh8c+2zYu3TBAWQRAf
Wp8IiCIHymOWzQuMNoIvVIWOjVhqmOrAnOkE+/fYpHaWg0GOFUK99BrOIxB6RReL
bPyeQ6eR1fQNikfv3Q/GE9wRs+RcAgFjH0BbL9Kr3Dx1lxqJUwKYqU09MSltKyA4
wgblyNWsetyNRonVi55WugbScZ2fxjBPmHjK5FctbKmQl8tUmAw1QHdxU1MdAUFi
WfCng7RV9ekv1/0ajJOaoy0Z7t40Ck0kHvigmaX1kdlRVgXYHimOc+myq2eEI0Oa
EHecibxo40so7vl3yuDqB0YggMjPJvkQXM9m6JUCV2UEBqurZ0Ec2gr62fewbLur
abcJldeShVMg0wLpNwLXGNJKCoIJoWX5Z5Eu5TyrPeIAlXy+BaB0DQqhAa6U6X3v
rzvqgIkf6njWXIULIxYgVrhXBc3ASMOWQvKz9V57rOX9t6u39LkYCeVvrSGXKWT0
09RMdSpQVPtXWuTN9SPr2gu6IJDXvoU5R0T2U3S/01PUJgniS4/hNBBLhw5YtS5k
wxbmsoDPtrEpb/vuuExuNxuR/HH4Tye35Bf92agLb3svLUXp9NxUOesO/upK8NHM
p6dKICLYEPOi0+FyqQm5YClA4SPz7llLSpwxvcw/bad0iNqrPM94feEOGV/wtRq+
74e85uyvfodY4vAyPHvukgQZCJQZ5oq0vY/h26qTVAkw+ym28ypaazNuVSkQ8tXE
TDbdJrLzLR0sJDxqXElzqQg3sgbOuv/PAGwrF3CQYOek0HwU3X3WCqgLnuf+seWR
cIVt7uEFtkgpT4y/da8LfaeO+OoZ5wLW+wh0ummhKjZCSSFpi8g4aXv8B5HAM9pk
7cJA1aDRzumvysd9DuO7K/DRqbvImal2kw1Si/0lQz+rXyQbzzJXPaO7QnGiB4us
bRLAGogeMWq45sF+OE+rXen7BXBNzPxMcFydXZBlPmnz2IF0Yy9v1jCahrHAWuLM
i8YBpu0PMVH0zU1HgiFzNF3vvC+n0aQCh5/W7l6Ftm0DjoxJH9uT/TDOB5roZED/
JXwC6g3BwlEF+NRXNv6JmvttUvO5tXmwV4+pTDEnP1vCf7Y1c6zwKjMVtVAYEXxW
i1lMsAte17KrI/cHTvXKDCtAlSxijqup3diQbc06uYtsMmjG/1Nmb4XL+ao7pwuu
Xtwz6WZulDhnWw7y4urOedFBesqJZupBl0ydU0bW5NoRleXkVJLw4ck9cVH6+LTj
gW5CIT5djP8oiTP2GR/KOQBXDjWhdcnshqLWROQobd/apgipVwlv31mS9OtRARHA
zeJRwNR1CnSQATpJxGFPXd5xMu45LqIlEwTX854S5OEdqWmHSd4QBTB54ZeLCpVJ
EJroBKZkXofFxub58POdwYN6H4596O/V0LHEgZumR4AGRJFBHRHxM1IqPu38Bud6
re3kuTrkua3opx0jlE8mTPhKLGV5P9UIO3fG56yvX4Q9XYTQzv33V6b3FiYfTZ+7
Fu9udTeBQ2fXW0oHAbrx1j3hQpsOy1U00i6oJ80fKChqYxtLYvRD1cvkDdlfCArY
J4as2cogaCpAjqJNOaHCr/BWZ0+KjXaxrpu4TCRIj1OKUw2jGVsyKfobGZFQE0W7
DXAWqdER6LQUT9c6JFQXF+8r7HRbwxUXRlkqCtf+ppiLclBbLiYdKHZ4FLv+B1KS
Aumvkn2XkLT/me4r3bG9hoFe8we83L8I+jonh6ce/BF96zPpKUOCa9c+rwtqjlWp
f36kYxvQgsVQJMKficzxReJf3d4n6LFl2QbGQlARVwiRyBvEsY5kAsKIN5sbQTju
AhysJq5TdrjW7yzU+bu3wLXxQxpc7oeWEpXFrlYu1NJoCHd3L+yOo1ZPisDnGa95
cSek3VbM/AgIkXf3YTUIHTkn0yJ+uKfU6L1Xz+aS/Y+emZ57SC900NPsH0kzDpae
zSL6sTb6xRt32Bf/oATfIrcw/Kt8j3ma5nSMSyX+KVabeCV3tGPhACi9IscfVNXc
WTXcZrMsBphOvEOjnbaee3lCHmoPPNMSbGT1wfa2MbCTphaXbywlAVzdXjRlTYQc
wX1BRbQ7KwSttaRgSX8uhknQB+f5pY1F/ai9Tez4EAvZRdr6P23+6j/GX7lpkuLF
de4p83xFYQic8bp3vFhrwrcJvmOHkwzEladCV60e5uMQ0gynO4P2liHBe+ibQIso
JUM2O3K3K7InydgKgTD2mXJu7c8+TP7LAZVJvkhCL5hjA4aD8t2oG2ZZe/xuedKB
XK/ZHKm9FKI1fe5Q5/LrJ9RQQlarZ0CbsVPL+F0GISPuDHYeKPT8Q0852PrNEFXC
twvauerGgLkfYleK2BQ5cs+nNBMkpHKWAq1T/fmeVAuybDI+2+u4lby2Qc3D6wA2
NXzaTeymppYc+fBCUkospRjgz6gQjw91Ga7b/jBlix+sO6H7zmpY0qKaO2vnbyZD
A6GcVMg69mIhPRFHqTlgtsRopkF+WiQpCDv7Q3Uc3vXalRp10X5L2hvAAD/gsr1L
uvJWptN+/Pq6HeRMgkBausZC59htAPX+kBrRYhpBtLlhNHCten8sbJjRLHTknZDA
uA2REqP5uTPbud3olGxjIH1nwpQz7QL+9j7VXZYPkVdZfxdbUFlkAXsuMJ9wtye+
28r+es7Ar7DePWEUOPrD45xkH9EBa7JDcLHZhgypsJqi7BrRDH5GXBWIujIJi0J3
zbOAv9cj55p/E3tHu4oggb97z/8BhbNdfHTSTQDZuRMrhqkTOy03jdHgHXPQ9xri
NVkqlUGe8FlMKjKWNqu1HFfZtzO5M4fbHQCSu2Y4CAtQjb578pWZ5U+PC/mAtXgu
o1a1y2s0MNdEQAJOev/YfYSOHgb1tw8A3xOnf5fPLr8MZfTTSIuRVtWrX9Jz158J
M/vFoikAFAWzqfddiAf4jVpH6job8d94IvFJbiFBEOxBlg7BlPRnEjTTKkKnOqic
2Zd7d6dzZ+3ZOqbHX9beyQG2GGTttnEi1CQehKSqtqmAbVpyOYNh03BpytwrLMRt
kHfThsQ90++ZY/Q3DioRHq7iNw9fAP1xoIaDbfcdsc6ww6kAs+PJN39sFaS6M09j
rvyGFGAp5V5Q3zvSmyjdbiln/hrYcuZlrhK97W41VpASK1JxlNM0wGc8YXNrysDq
7IWjqof/f1tMaJM7xvgGzoEK/U07q1vHU3lKa8Y/rpCakx3v1HsTsY8wKnYycWEL
LsFBJSbW0dcTLykPJOzzEg/KEDq6qYaHfei+WirS4Cg8dnkfYvisxAU7pwu+LDsq
wE8EIgX14zP5XHW1htdnguvQrBZ4iAHNQsfNHnVYXWYzYAgjaSnzLLRNn2j3DCXl
8gX/YDrZXTmud3aprVq7QbHd+Jd5XOvneuWiP99Eoy9/oyVFB4p+ujWqP3C7R/Kh
iNMlM+aCYemdq0bLUVAjt7cbiGeIE3MJKtDCcMYERQlT8BtER9vKXlDV2+jm8Dm+
h1H4LqIVDrMGE+XuCFNF5jW5jAoYrJqtr4UMOxVIjxRRrWgB0+xqK1K2DEfZnZRU
Mx6d3DYn2/RPstU9XgKcNz2KVtYE/5WPow5XgXxEOtG8d4PAX50XCAMl1I5+c86e
PwNkdhVnBS/G/SDj1RWv7WZPUdekljtIzlUQ+9dgNYsZxzF5Ycm0jl11+SObC1O6
W7kbdo4WaybEOSmBMGF8MgwLh0c3dHJN1Kv/A82nZTKc4gdyQDzTtVMHEyGXMDyR
4Q+xNE/Ucn3Z0o47tivApAS+YwfmpyR4K5BYe9TZxkHeeyAOpsN1uLUx2+vWNfVH
vY14TxRQzP7G17FroryklZhVTq65ABnLse0BjzU7MxkOdpPCsUJOe5FMhMct9x5k
hae/GEGI9xI7uA9T39ga5vMEf+Vb+rmcYYNbRrr60H34AoYarhnade/Uc0//0DIO
mbqcCsdrGNac2xmxzCaZxUonRRyll5JKPdnRLgcpDjEGBunv7kaA4O3Dzy7q8Co3
O5fZ1e1XNLn/8CRhcao+hePHfIokW8IIpZTgNbAH5os31MemEAXwlgOuox5Eqdab
hZWlc27mD+teoqp7XW3DKXuN3/ITe0LrFVAgkLwQeGcA8DHk5voH3Sbm4T6W6BMr
ubkPwJlJ2g+Ziyufsarsx4SO5hiQtjN1vtDawBiTcKbiQFywvyoxhzIm6pgsrOrY
SWM/7kbmie7zt19qv9r9i1/9cMEg737kb+5sryZ+vb4KUSia4OFZiJOtBoLGhJqQ
GPOKDHkUu8wGgaA330ztjWLFL9SNofgYKp1oyTQf39rkyjh6Bjl+BHeYKnlDuT8F
l+Tymbb7TSdJd486pMC78G69qP4C93u04uQn7/h2NdNscJwRha79PPJ0kTG9k6Ot
AD44GxZZp7YVDVEwXJJzz3+UM1BeO0sathd1/1zUa2nt2VI8pQgTEQdiWPPlRG3/
eQkx+HYtzjZpBRJyxiZWgguMuS5l73n7yNiZk97JTnG3rAavcEwin4X7ZbviAcRz
zHdlRcLgwElga+1AoahuwVvYo5NhHoCglIpYGedOAEUAvNXtpoO9gyuEcZlmRxRT
fQrqJ2Ej8RjIBPRKN9qOp+QUZBfoud3zQByJd2vbYaDCffCH5y6EmgOxmUu3E1N5
vzVvN0BsXWT+1Yqw9zH9soQtmnPmSdkfw8yD2D5MHCtMbNVnvSDKU8FF5RluHS2M
zF8o3iIl08IWNXoM9ooz36yjQ6lar083AGDkl+Rw9xDRupbKL1dZN2KIuBum/N82
Mf/wGmQMABa7r6B66aKGMFZrU4Q03T5sQKMuRYouBNRkFbpoKafFLlAURlCN+xMo
d5F0mgb7Nj8ZpEg8x1jCWm9OPvdWwCZwkaOEzWhm5hwPGkd1Gq0Ii70NSNn5TT9T
DV8jmHYKKZlWQ02LdTECcDiOiqTEgbMIZsOnv6pMcnXKsKDtXXO1+zrIy6EzxFX0
qsLMebDWmwsnfkpgv6ffc2yf8kouI5Dl0kPNiFEmOvOyN7WIdYoDzdYQcK3l6uSN
7lIf/spWKZdQNMqYZMJ/8nwcVqUylTc/EUvCT8TF1jJYwITurfXnqx/YCs8E2OU/
uLpk1g7pT59nccwx9ZEnzh3HwoqrL7WwTEUx2mLTZ4IsvAXuB0KVHKDr7H2D4SSh
PJqwjjot3kAwphSrVnlcA8zBonkLFapcpZnOMLPEwBbYdcRaTJn7Y4La0wwNbtSh
ReMZIivBkkJdKj0FrNFiaA83wM1n83J3pQfMFITxYq4MZKCPrDjz+WthnKVLSlnM
nlaoP3nFHKI+4PrNl3DTyDRKIQ18h/xZkMEyjy8dASeOhmwgOQoT5lz6S6tmUURu
4Ig8VzPr3z573uDHHOmHjwkPL7RXLOBnQd7+lJvwvTIhCiAPCZQnP3WvXMVcs8wX
C+yBbjDJ/0KdwSXTHY6lQvbXuzdjN9oxICMrsZFXa3F1UPbbSn22byQHHjFFxCXI
KLkGKdrxYam8liOzvB3QJuCZJyNDfYmwrR+yiTA8f67pbkmq2HhPgQuE7jcoEVxv
Jv2UsK4pgcYjgymVsaiE6J/4tiVZCXmm/nGyuEZGSq5ln42hXzXVKeBfikfBWokz
hN2WI1aLjqut10e2fiVnosagUUcItjfM7J68D3kOHhcYOhwmu9bHKbZ49Z7RoCvY
zYYGxUi8kkBtujYloC550wzo+Hbo9pjEzzU0zoklwc8ohD+GLDEfBlYO9MjiGAHl
hExkwJUz5vewKKSVzCfI9bdW/12D7SQ9gaGT7WBuBUM54a2BLB5N2h1GRuAbRSL4
tcg7wVL2P1GBnsViP6zW/TMI0vkQck6NskYChHyms14CUHFinBX+zPZk/mSVRkzp
0fCbJh4HsjvoIR6sGoMYVmYuBgrhrgOuITW9fb9i5LmxDAp1Met1um8ZRKIbT+4X
R7AtgGmPQix4YG5A7RAzbZfZh4NWw4VXV3g8Lx4evKU3trCWdj2y6qC5hfSlgb9j
daU3C/dY8TUN+rNsyGTRW4w53EPuZn2AqGljJZu9Kihj/O4LusKEL8HwkqHDWk35
b809eogUGHrptqbfKN1lHMy5R8pmlOSBtHHdA8wWLPxQ1nV1ekUgR3jTLUM7koFA
l9bjbKjQiMDwBCDzCuuzmh6AoPlRzAs7sp1jQgMbvRIBdZtBfrL5V5px9k3vzWif
0ZaQQJDQ7ijCu2BEhHDYIByyAKZu3+YmBHWaTeHWkWdpkOzVDlYZsNnbHqj1j0hv
o+GosJehshOqvcQTydxQh9np8hUxwGuWIycGYgkTWdclK9eV8dtwIEQ1Xhvp5WBH
R2lM92ZawHeOrx+oPUUz1HYMozwwszcNWhtW6QH6E/rHzd3weVehPQSzQoOP2SuS
ZuHgcL2D/KRnmjz3DgzBKwXlfvrV6WQ1NRekCyINs0BT5QF9UiilzSGkrK1UdWbr
GJuvI9hMnhN9FClyr6QcqVF/HoMplQGgi8FIdDhwPWOWU4jxzHdf9wPy0NivqGfl
UP2sqn8+E14pUSKSx7R9pIaTvniES+eoMMqglLnO+OP8c4IkJUq+nKmXn7umrC86
lA4RpJ5Fnpy0dkBSz9Xe0M4oNxHENc68mqrSATx2JnViijNim4hseAAB87vGTL7o
nsxHUvERwvwCq/taFsn2jImvOEVP1VX4IaH6juXJoTmbSuY3XsdoZVwhR3BjTrea
pHPaO1GOq+4YBuQ0V9H9SH+6edkvM0axVFeDqaCKcUuO9i8tAzPDMyRlRYBssOK5
jRBJnD1ZZeMFCUPtk4YLwbeYeNASgMiwx0q/PcibEBV1JKxh311Q/mjIQ+rteOTD
t594Qf+fC1BzFHvhb+2p56UMalgI/KRNQug6gPAoRhS+aZd1+vw2Bq2aijGddc3V
18TcH2xF6ySFLn6upSYyLYXlJX1m/Unxb54k6h0H+7Jr+CxTLtWNd4/GPo7x5XVC
3eUzE2Zr10FjjKhAWXZiMfu/VZm0SpIn4v21GjN+8AShLrFsxk3GRIz1lwG6FZFL
HPb1cALCpVCmdespU52poz1xUe8uqdpzV4NlqGW3C73JhGBUVZqZZ89B7NymckXK
LglaYVsKuck0PeL4tVnCmZqowYL1g+VRJzvCxZ9wotUPijPG/34IfnKWVz3oyILV
sLPEJAWKICbNh5OJqg+Au372CWdnZlEvmG/j0RdnZSxAgTTKOZj4POInhZwGwagK
5gdWDpmKoeSfZ90ufUXnYhFsKqMaLSonaPiiZRkrgxyC3pANhh/rSfmD7F2ozpbc
zchJ7Bsv0bmy5BSHJMFJtT7nMP5+bxx9Sm4yIeiK4ky9Y9cqvcNXcMe3mXbGjFXV
u7niEYKXI+a6FIInlpwSUkDisEckHh7i3ApHVbbQJop30T6N1xUnN1Ek1mzJRT6J
1HOCX3z/DmLW+MDnLKvHtfNLhEUHfq+IS2865qTVCY6dWotJdjA6jH+aABfUwsXo
KrjN0WvWPtOvejot2FMSOyHlHhconjHDoCp9EhAWhzZQokKZvdRsIrG36GvFT4Ba
sqO8SKg4fvZ/KUsXo6JjxdAqyd5Qjuqu5Iyy0BCsoRvefnb+dBw4gP3n2PxTTncd
aBNxnoUoHXkrHmCgdF8sNggVKr6ugzOnsfTmaDxpxEd8DiyXS6AuiqFbFEnhWp+A
3b0doQ8nAeM0xhWVzv/ALvRcU01rZ904L44by4nvD/aCZ0lCr81Vjcq5iOmMMXZa
fSFFQ1riSf6a0kG7h6CR4VLm4lANy7etlSZ22QuZSUS9/NBKr06FWmLNFyj7USAW
mbjaEoLrJHreXg8WsLxmO0YBvzCSwW6IndaJDu1seq6Kml0jUOZwSelzjiIm51ab
PSpm+q+up+ggJWh7o1UUzaumjq3Lwi0MxpK6PyjqqcI56dH8RKdCyWFNkhsx2R0V
Bt+tTu4uX0/F1TOp2ITY4oDdrEbUPt8mQKVyps73cuUeaweqYS5jNgDEjVfIMZEM
5ezjCxTHOO+Ih/GjR4dd+DYRTSDcinBOAgpYZMyl/dYVMgROkQRTCsD5YS+mcAdI
gJmORw9B9CRZMzvlisFMoT73EXp3egJUqFHjQQCsCjBum6qSQoTcL9blSiJtbA6B
QwWyQQZXD4yfPpfbdVii71AvGLvZQL2FEmexmC9k+eJ2JdBdX7h++BRuJGdsWNPb
y/sSzVXOpoAo8LwZyPJ/NpB1mDpn1LMzVH0nw5QELPe73BIpZXIThtSFiDSKtgWr
7lAA3TfSm1o6syJ9EijWgGU0YPLrDKUuZqwRhjZWjPAPKXOGrflJy7cOrRUtDT6K
CHLZPO+azvPMALZdVuto5UxtzM5UoMdA8eN1C3E+21CdNAMkF7aJYd9Pgjh5sg/k
RZrfjt3FAFhI2SSZ+EvbedhbDt/xC0GFUOJKzHkPkCcJAPdAJmZlv3fXkThE41NZ
faaNUhmDVER91Ew1N+6BvEVOzqQFkGHZE3/MoZsABlfzYbkO3TxTNSGMr1aJwBCB
zf36ykWKBlpO6zMw3iA7GCxrVkLTtTOj1x4vc+nEWycRfXUOIv7kQhx6/5v5CTKL
oqMB7hZwN4FT8VUHaXrmsUII818PTOBcdkMDTBE+Yl0dAKO1JsA9ig8CWdae4Moo
Fb4puaM25RrmNQaELTBRs9LNvygeGG9p0HdhLvkydtAeUAIVuazSHvP2p9r7IPhV
rV7eNyASvxFGeFl35gMdTFsGyo+blxq/wpBHdq/HPdtNWIgqIk9Gqc34vcINRrap
WfHVX1Faen9V8DS3IUSI+rw/VXawbqYwL48EO3M55N0U6b8nXz+ho/w+SqLVjGvg
NQLUEBBrtG5RGbh/JuhH+Ts5g+u16YZKkvnALx00xgK1Pf4o4xKGGXqkBkbedede
EOIZIznw4GD/uCvD0KV/Z7S+CuPhYyAVWwa8uUln37ycjfj9cmuZYINS/bsJVA9j
RFWshWeT/OtmTMOTS4OLh4WjdrgUwNt9q4DFXDhtg2XhFWTjfaDJa/4hNfqcqT80
IqPGt8+9N7QWoz61ljBWAcZ3LDn+ImBxaEXtdwKcUC0KoEHSJkr77+zmKKzv2jCI
G8w1PhM4L9cG/oEQhMWa85byLjmgDZwoEG/6McenKc1KJF2JzcJLpN3T4yDBSK4c
Zo9g6XpcujLHdgy1GF3Ze64SKzf1ooTclYX/VACfaFjgk/z7yyvYLLFUKeCc/XF6
N+OERQ1IqC1RoajLhWdoVKuleP/oAXsjoS0B6Hv7/oqHpIetNpvreYGEGsc7MZoO
mDUzui54hwou5H1tYZLvHrZdU/WGCSc4SRx9Dt6niZN+MGZTAGDv8LoT9FezBXZ7
1SYEfpRAL7SjfW7n0HpGOOKg2tb7JLaMdHFMOsTDf5S10nET1Hgx9K/MrqvWBLJW
yNt/nbsySBJEyvIJlFP8AVVbEhfS230lLZW8bFevE5lq6PIn476wdMcYfp0Cruwj
F6xr2qBWHFcSltBAjOxHc+XhG4IxHys6MWPlfXLGVqBlAU6g5A4jrFB/xLXHwIFn
lJ4n+xhS9VJI0xXRkyPh+QiuRUXlev0pdygniQ/8Zm63rfYlZqNTNEy1X2zC5gEw
o74qz5h9nA0t24qAezSmZ0x3tYFVCZ99Jo63zFQwZHEBIGQTp5RaVJ80ChffSbtw
ipQJ2WSZk1hNuI86WTq7fr0HQsoAhl/7XlwKJDSS0CjVKsmdnJ9zF364Yb+f2k+g
vqdnFrbcO4WKUsWpXdvdcM1Cq0IPc1docPueexNq8Y6uANo9J77ZtuR1mXslhYlm
JxjMYaT3gEGq9eYD27bFHInHo4017khBo7BeBkJPobeXiHbtgxBlD+75weZpoBmn
zePDJFpm+fQyIS4ug528ss2Fkw/16KjKJX4ar40YiffFnHCNEP8LhzTUXPUFqiDu
o+k1WMUNSY2D7KlBMUe6oTKU2tIphvjobA0PPJjEh1PJDe40bL7rzv9xosIUQe0K
7ISXW0DAs7+bAfVUpASwixKT0+PxxZKB33LGrzv2G7ZaR4j3Xz2qcwbmOmruw+wQ
nmkZeHwNgQU8lHDNTvQGylo31vMS4UFpmvNtw+Qmz4J1q6sM90kXTXn0j2Jo2x2O
CZHVMtFCexXBy2D4qExxz+wSiLQ7iAiHLlmN+MmOSZig79p7xMFMiJZ5sgJcjAUN
qnOcpC+uYU34fmpoL51KNyBjeVxlIAnS/YGs0zii4jTspRsW3FIx4Btz6Jq1lZtx
eIPSvFRrDBMSS5YyWQtLghr9O4MW0nfWhBPHPxZxQq23NIZYVF17083A6RTSzqvH
6R/jO1vIKb70E28pPEv6ZecXTV1b/w/nwJfZCOHDdYk+tdrUPwC9aGSWEzymZkrX
gkvzpyoWZcVcIPUKz2bRtqfoRtr1v7G/g/uaDAsZfUwU9jnSzmml6c7W3011y9OX
DlhvPdgMlxCXsG5S78fs0WgMaQBD1o8vRRKswLrukM8Ql/eqVTPh3ZmvtxMbcUcM
VsPhwOOrXvb3snqI2Sx+Yqa+v2urreIATAdJd+tTdr8+MrDyr+P+RR1XIygrLJYK
qwxDO7/Ak6iuqmAxIbimOD+HbM1I71eOkRGVPoMPZ6CEAy+pok5j3subGo1No6uI
/qIYN0h4zctUAC/UI9l9TE6DhLN0/XtqXhrWHok1pLO1jxeNHvnRzoSlk5C8eryt
jxudoDg0fqzDm9zHgebhmRNRLJztBMNi2p9r0HTo5KO/GCWyTIdyH3LQFHY7J3LJ
Qo6Rb/6vsBAh5/VDkP1ZI0pm2z3QjTYQUuawI9lJU1uiDN2yMXpC2oct4PkCX8i0
Rx5duKlVXTXNdBNjBz3P2aZ9WXZqfRY9MQLPsuUj/YEMQdfvrExohGGaSuWbdo1t
p8iryhg/4UIIWgzrwJaoqXDIYR7uytNRDGsR8I2hrXsTc0u4FFXHjnbzmHGNLHCA
nhfx4gSEvz3U2zaI2Tiyp9sDSVFlZ+5kD/I9cZVaaO/v4COZK62jWFHxz5wlqDlD
P6ud2ecybb8V+1sBC5vUpAkn2m8+LChI0OK5mHC3Gk9f5x4fvPP1odvbDZUlbNWj
trwGdKWY93/Zf8TymnRixMzA1H4R1A0jj3TkxOLacyfTjsyO4gj8qx0UNFYLBfoC
H+es2+sXOciecOI5svIi02LA7QWiMXZhHHjzRU7NcQk6eKaFuLwDeDQj0TX97USb
2sNa9kclrJDKY5rlnkvoP70VUx9G5u5gO4eUOi1F4tbar54sDTD3Ton20DlOWOxo
2wd+3qvvZbCjNw4cgZMacUgaxxT7G/iujXUY+Oeq4P99ERCciKCCPLFSunGvdUuA
Oq1w2mtIVAH17Pc67SpjmuvT5/EkzqwJ+QIHDXqacM1UF6JbyrJQRKDqLw55VBhc
6QeXvtYAL7OMmE+F62QPu0qzzaXvtiAqdYL//sTSEPazkBmYPr90DItBwxhRwgn1
vP6u0CTnA7vnlj19Tp41SvMTvUazG1GwqJQ0cMSujFRFtinuGEcIIgHl3HG28Xr1
ZOpYnVFjt5fLavNogsHZdI91PmTrWwX1VWAZCLX1+a6WEj3OZ01Fq50w8BlmfqeZ
pWJTCSwB2EtU6d7cjdWJwdFhn4eyDJY75ce/67pRXXA7i6RN6a2i1hnYbQnLl6V3
eM2Qr1UJVukhuot+pihQ9vSuTOTIDYOWrGKX5zfV6K1WNCBkVaWolInSqjIDse69
cy1kvmIxgHkyRW+ozp8B4H6P0cbC/xrwdWedCyYs+kTmEuVMLd4/i3OvrnuXUkBY
IfQCjFLDL9eHYIi9JyV82gyE60wOG4ffw1xm5IjSMKv25656H1C3GAQlYwxEU9vq
fhQ7zDEstzvBN4IQf03V8gXNVpDa9ieFk9Kyabwc6UcY8pePDq3/f/69tsyd/TFQ
Nz+hLc2vawv1WRU4BLE0j8vUw/i2WookOE6Eu2On7NJfABshaG5MGELzto7Eei8D
S4c0aFbUO7EHufFicDEjjEzzV225m+u2e9qN5UD/sLt0r8ZK7NEJNN6Kw86Roswa
GfDTcvYaOkmrzOCGxpffFfS8CPW/4TaO9LAldQU/cAKbowFKSmpawbYnxNulHM8K
bvgdNtqEozadVJdIEFBkXKx9DPq4ILemYRTibm7Znh7X+vs8iLHbbEnyyKTo7XFz
raqMoLh/GxC0hodNLRlUkogkShrHq1K30gfdgY71PsghxwvhwumqLOWK8ejkyNXV
vhMfrcw5/IwLI9tHTOSQLchgvafUxHzobJ9Pu3U0xBct0Xts23b8zfRmDnP/tN06
CL4jOjlitOYENOW358voDpqy0Yvc3Pz9/tIgCyWkFvfTBTy5viTZ8TnRc9Qsx94K
Cc5Mlg6WR6ON67X1rXDvlc7wrTW0S9hKkHwmZeyCuffAeI7jBqRoLbuEDhflHUrx
umUQw0riNOcaRawX/W9igZKk2koWM8E2elnhjCU+4o0IWLvRdHfCkmdZKjz2qLLP
0AY2JTgnyRydgdk0zsBZlrJ2NthotHZ/9EDS6faOzPAQqSPdkjpFpG8F2mq43OXm
v6BcC4t+DHt6VvQs9zZnP260QI3WE/KxqfxiPAFGqRw4M5sp/2gKildsrskRJsaG
3QWxvZhmOkuhkW2dW98xQkcipVAur8Oolv7Tfx3UBZndBXN640VHms50xy1kJkk5
1fLCRt2AIB0aXV6PslyR0NlKfEtm0ocz8fdwPYbsv6WJoI1fZBmbri5m0XDqSphn
IT668+KQGDbQ+xiESIw0juf5iZP2GTTBa8viASimsomR447huakeJzfsXvEMBXu+
Z5E9HFtvW+U7J+YYBwjOHx5eQsH6VwpNd4OXA99yH5V9/pf9Tz5WhZpTUIbfNsbH
g5MzXhNZhyt4rweESZNqf4bvWw3W/Km3z2VnCS21bSjapsBYAMVY4qdh2haCqHph
sZhGpTqOrDyF8U2ZqGZ995U0HlK3vX4JbsbmqO/INQcN+0/dgMayfngtVrr6a0uE
9bdZLIBUA+gxF0hXCFFw3eRurcNUEiHCIhh8/CJmOTeV2XBsAgYhEL+0ueyr2FxY
f3s8HZcJU51vOW8t/PXf7vVdT5xeDMeXBucgeqz/Zmmh06dnbhMH1ry6GaI81spY
zLzqQYegvcTYY2/yy1kfug7Qwv5zMCUooKAc6DbONOYNUkXrlGKEWEvz7cYcgVEr
zUmzENXn+9gl0oIIn1t2yXWB6+0fxQuyS4kjNhjKl6rfjXPJvx437iKYNac68dEy
MSECb27j3/DRcDDnV8nd9IRC1okf+v5AYYfD69xTsGUfOEwgIA4mCWHYbw5JEHUR
5iw9o3ZoA5MpqRoish4WNB9PQzTAvimVaRz9rabIHVejhK2z/M4FpsufcZExzcH8
NdMnmO8dt+G6MsrrnIvgqWqlAdrXpX6AR6+d+ODwPaNQZagmItREd4F+3MdToQr/
YT0+ljz+kJGaTroZPFsoB9CU9qxY3UuX6FNnuyDBCCrJ8tQTdWUknz++B9AnO9Un
PsXDM+S/5m6xq6QYvXK0akoxH5fsnpwSY5tJ+Jw1fzbgLAFHUmAl4G2cSoew5Snb
YEWFygf+NDDiSmfYkEAUNvjMXE2inUQNS2XzUALikT9tilO//+604Uf/5JH2Yp0d
9qr7XfEKGtZweFahuA9Br3IbvepitWEAltHxWboDisA+44Z287h3Xh+yWYZJGFSC
6WDIht5KEGTlHGQp2pLkW8u90sxyissTtTekJJ9HBqFMlEgvYsNhTdi/en1kdHU8
8qQFM8Qg00Lnq2RqyVXqTte53ngGI9H0AUrFFTZl/9zDgXTKYbSDu3fjRxDorr8J
G5eGH7tduTXDBv9NdXtyddTK+CoxpJQQDQTOzrph+RvC6EN2yDvQHM5spU0JnKRD
ePVDZllcayNBGY0v9sS+k8z58+FCY0s4vV93M+XmkCRJr+hUlxTkD1OjCIJfjL08
sZuvMnpU2moA4qtebSrcw+K2yT6XmLszn//fTvr5S0x1zQbMbIi7LLK01LpbncwH
hlz7QGgJ59TC5fO29c7EgHQMH3DXdB8iGvcffiW7Q1evs0oyCKwBmozFEJcxvuWS
pV3ihEICA0qF9hN8BOlJpJpw0jMQ8WuKZioNRTEmZUqU4RzhD5ro5Dx/noJLnbEm
wnU5st/D6b4OITnDX/MlpGr8KC8EwGAdC4WZmSKM+9aQBkd8aS90ojAWDa9ra5WC
nuYcKBdVt1z49aVGJHGyK+jidqbfvpQJL7ulMv1glxZ9qfNtIvRBlHvXbOmji4fz
cOAiBP1rERaERnlBEvE/KfNGjYKXcbP5cFWYN4sDsJB9Ul1xL87jnZlaLYTr6anJ
pFRUFjyXqb7x5lHXwgTokVYC9ovXOZYL9xTBOTdy3VO7wD6agEah88B1YrP4hcD5
UsGX48yKbOj1HU+mmaMoEqEwOjh0hHwo5pCHntEFCKRA2NarRnI/LKQxs723A8O1
o+bQ9AwZ27ZRQBV3Xc6ffXGkIT9w2vGaWyhGPLlUpR8dqwlwuvVp+LQBKiNeUNbw
QAE0YIf2qqBcMKE2ewlZ+nywbS/4bfl51Bmk/5tCOJJ6CJREMlRbav6ay/QwgjIu
R48skjjC588VnWessBGN36YTb+p2BJ/fiiMdsnpwQg+s9XUY3K6GVlB6RqAZMYaV
/pkz/5t5FpVoPiT2Ivhv2HOAtVNzdmMx8HcmgRM6YqKEdZxLHC3TA5eKqkq2CzCa
fQzoJeWtVJPEazlRq5mPBribphcVPEQBF/gdIyIsntN/5iGg2pEVrs2ogOMf3abE
OO/ZQPK/gaAWfR+/q1A2RwDpCI4trsqBlYRtLwsLYeIlwCy2+XspvtJWkTl5XGcB
4nKywzn+9rCa1cWnJVQ0kKBqhUfxtiI07BfgVsDajh3RDsuFX+1sfouC2ZFNYpgt
WcqdyQTU0mU+dBNL7CnVQt3vO+DzVNzy5HnxBDDJ6q5y5h5PkhN3OdoWGqA+evvH
n0SREj5mcsNq501VffqOp07zKvdpgLhI/uKWh70NF26sVDQ2qXg8K51ythQdg2Ni
XmqSizHlYzc8L1ANCTFqNIwdDQhgvuNWtpLGT2xdun9J/ZyPPJ45dsPGbHsNrYlB
N7O9a72Qle6C2HqqLNjgDWcKvwrluDAfEF22s/cglBbq7fqiI4v+gqcsq/tuMRey
Rkzq8KnvzbWUvQEyhZj9KavjPBJ0sOdypP6g5xJ+O4jt4EDAyr4pDhDheg9mg8bM
pmVCy3vBPD7WVtwc+FzXLYkekpiSpLgorVCrnbUVM3nPBqenRDxBMGsDeD0xeqal
OxVbkUsIG/sRO3orm0LjKvpVvKVAQfjb8Hl7R9oeHb95EKqWdmMXnHaGfi7yI6EV
OIGzyOCPYIOD2M8APdpk8RJrk57jpbHWyvEC5rm+HFX7s2dh0LJRyczvEDFJ3hGY
psKiFYSV7+bvFawPYR7eI3N6gr9CO5VVxPvwMYGX60N5zBIqp8Wd6w+KynA1Rrki
kuf/T+ReLc1qFrvX5kl2wpII5q5YQd8r+LXHfB85CN6bgNofKbrDu5Kf60wYqH9W
f2FlZRuhoYYnFMWKh5tlczaN24W+ojZuVXGMcnesRX80Ld/8XHFM3ZQKH6I5rnH8
W+eNOnGZF55uFmdASu26rghGOL+KANIvTxPCPebszqdJItT4EVVUJg9n2POnfzH5
wSUhzOV4B+4mrkYbIN5OTHrW7fFHIJPQ5UolT2y9fduxeCaOMRmrQoY3kAqbIH72
ZZeiQ88ohvwoc1227Q91Y/VHof/TkAmoOY/ksEKjZZdJiKonSOdGOa9y1xYiK+aT
89BEPXot7RfS+/6Jte3JMw+u5AiuYtiVP/p0Wj7VSD7dy1O/qa09hzO7jkDyWPWS
X+nKr2hrJEeRxRzgGzRl2h0v1ElXGHz02TZJyUWtP3thyv0tq5xzRU1ZY5Dy9yRv
sF+WDIOekkJH8xUQgXplSkW9zB2dR8D31QBJctGmSVWHK6IUG8HkQMl917kcreOW
kLnexndfA40nHl4H5InrIk73AP9CZchVuxHbrayVq5SXR8QaCL4wA9JqI8BzKWv2
PjK8qLstYtF8KSYg5/QaDyRD7DDUgFd00X3dDrlFP+CsOXM+uehHZ9jWwuShstLZ
HElVQ5eTXaRc+j2Jags1OUYv8f66VW4wbwR63XjfIwuvEAlfcSJ8dJY9bZEGCGS9
EVwCQch55IUF/Egazv4t58XrJySvE7/VD2frA6zoqBE571Z8Uj951mcykBCRgC1g
+kPSI0Mlr60VKHJbtMJsEU36JKl43TsGbB9X63CIcxbwyefvbJgslko4R476Aqxl
qUDWYnI9jldygZi9DZV+PbRog32+ACqAn4mvnY9+pTPVaUvLepGAuFjMJ+Aiz4nR
SzuuLprAj0Bts5Vz1KJ4XhFcIm8hc11AoUe18wUp1zJxlo12R0GPhGJT7VB2h8QA
lofip+3dH6QUq6TstO6CtKoKeyiydxplfJA0MGLhBB31uA7RCZJZeUx3yEpLOnwV
+F7EiFc1gGZlLLN5Rt5D5xok1c5yhQcwy0oZMGQGh7c5PLu2Q4SFjXYE3OhiUqNK
pOrkK+6qETqacwKBkH8k0AxlzQjWtiUAOB3Jg/vrCM0/lzgXjxXYESKPV5sOxKzh
obPY0u9bFiheBgfkww3SFVzYVWnPdA8Xau3F4ABB7CAM9C+FSV6K1alKZr1DsJ+5
JkG8GpHcBGGiR3u+/LF5wZr6pkvA4rotJ/wHE7sQOe0Nh+rF6pwiyidOFJPlhHbj
3TBa1AAWOzXpeCScl+DF9ZFR3/1rXKwnw7FEpnjNyYHV6bOIbW70B6kfTEATx0sE
wd5E4TWQCTJ3AIPBioYUBE00RwuwTLU6qHBrbKMFaxMDmOoMQ+xoBWbbT4jTOOQP
2IxdkAfYehu2gdMCsPMBwS2sB5/GrXp/MmYwyq6QQjklZp9k74sJNDlsa3vdD+TR
PsOJL/LmgvSORMa4tVkbuJ3He/nxIDX6Ti6CxTliuSWaoNzu1ZGXn8trgFQMegN6
ecYGbvV8uUhaO6PpGOwDjqrnhOYOyQ3RKEdduY0aysAUTO1dwf5B0R/WPjMOKcsU
EjvXhztK8bqF6oIdAWl69xvqKGVGCuzQSTaw+EqMoJ+0BT2lgXG5emhXgs8tgOS1
9HLdoplopGbWtTFQRtepanLgrrZtOqFdYIZ5hvhBZY+VuERtHl8iBQZVal++K47M
gMyawHgit4LKAM/PEL0ZsI4C6L6HSo2ov/IoaZtgIr+hDErEVCHO0zMinrtlIw/c
PX+3R3JOrLxz4aaX9xuzWXQupXze/baz+X5TH03i0zcPkvJP0gVHCtzJANxZsJjL
R7jMgTgO2hGH5SILoZ4g/WEYxHzgt3nP+Rk9tzeWFFSYE2pdL3J0Sp86t3OcuRBZ
RTf0oOT9Y29ZZwYWKDkFqbJZpzb5GaOGp870gmMdArOP1qaVhFwCgLceDHA5FzCB
SNpV2tTtvAJzlXFLNsqIf8zDz3Utca/Y+EPsPNuU/Wko9J9JS8Ydjeb/6VsR5Ixo
PjNA65ighSO318n7mcZmloIJHTQkRzGeuJegOK09INMf7dOKBN+tpUm3YfDDoLLT
l4L1ryVK4UXuQUtAmWQeDLeKZ89akD/o0scL0mbHqBfouT3q+iwfqdcfb5SKSN27
cilbPDL5bsrImavCxLzFsW0meexZbRfhUZPK76VBbpjzZrrPnym4sZpguTZYlV0m
nQmqH+oXRSkZNSbsxOaeBhwR0uEBrq6f6fyVZZ+OWrQlBjsuC/K+vh9VdGgxHA14
dZVZtd+WWvyjhDLUqqtAPOsrCIOpuFz6TPreibCxR2XGSwN8OPg70AWFw+kY68y6
i5HzafjORqeX1I9u4sOSK+C64P3J+sP/6/vKJ8+WjmsIzScMjynx0U2CDG+6maB8
Nzy0IQ/TpxWRP2M+SJyCtGso6LtSMX3Y/u5k6x/blK8N/U8t4iSb5N8F98TUYwc5
IpJpuGr0fNYZ2MNVKE7gBKYKkFG3MSsuzFk5/oT3+Tk7G3G/2RC1tkoiM3t0iSS2
MhAHAhFD8bQL4LgCW15AOTpoeDqCZJBi/3Em93MzjN23gqCbJB9dlFGC0HWc39dN
IHKp8g3xzJM69Nyd4R9kRmZ9vMaNZAYLypU2DUS+FNkdQj8oKTJ6abj/xhNVeFOT
bmsWazZMJl3asv6kkKaq/4YRcm8rPR8dmO6168mMz8xdDUcOrdw0a3TTWvBmjM/K
yZ+HnXSUBQDBjJ8MIn83ghj3LIfjXxZRWmJYImlI2Wuk/2p7ob62qkVAetsDLsyN
I+krGnT6eLfAJn3mwt05Tsm6xDt6A68AS8BB5z4eRmNZxRKAE31MLaoITuYmbMro
tYeS6pZtSWgKVKPJEL/z6RaS1ACCrT1JX8NC2mSyfXMgm2BQQ8gfn8rUB0Ys3nuM
GV2vFp9fuwsoYWqfO4CR80aO8itwJL5MRzh7hcytruPZBDRCGfs+8wrQ4fMOiOOr
ZR6y8rG5goy+/VH6aUOGXbHLHDu4g6sO9BqPnr/I7kem65Zbi0+sBZf5MPg3kbki
yDmhcOn5t+HBpCQWON1DMyOB0fDNqVH158cQWCrVX/WIG03q8ahC8DIDW6gURb3U
TyaK5ZaafUjPK8KggCfOQK1xh5/gkmuRSw3cEbZYQJKKMNUMGeEDbS8piwVW5q2Q
TVsXTa1II4X5eAjAeUpER8AP+kU72ZWipvNDXdmQuhze60483eXmTj6kFf5d/fSZ
HRB+q0Q73qCZyV9aZ1EzKvoWDL4VYmoyyPZBl8f7DG7IhSD7KBGkH+4ZXChpr6TH
IDiRTpaZCDR+FYb2gbFOaUWgRRnJoDIM5hbFRn+FDaY3dq4/xsOIo0faj6rLmklh
LGTwHEw7PIiX6BTaV8AuYz4qNYOwBzjYKreNRz1RkZaCcfzspX+b66HmtOYdiXpy
fp4nim6r1BXEPA7hTap9mXVz7mh6SyDt2xxkb1MJUduEDvjPjTdpvGqR5U/ahXMb
9o9qcgCQKlC4oFduXmDYMd4RCp1R+YDvuGsglIcSDB1KqsaMkU9aMAjszmYakhpF
tsu22fr5Bbo7guewTiT/f/0JPmgxhUwVwDFlQBpvC7kfDLuxyWSUnn1+pGqK7x2K
6ZTMBM5cCqvQRjExdDqyE3UGcuSBHHRh3fqvPFUAcdqpZSeNu3fjZWi3aZXeV0tv
OVI0Qjr4BoRWk+O91kQndU2NePLibkMg8OsG2mtUcATM9M5sRbajF3reW9rPjPGB
yf42t0AnJqV4PPnIr2948JlMUHsLszOj+AyAIgs3D5Zj4bPpC5hzM9gQCr6Z19DD
DLVlYv9NIHqDNXq0idSC9CZVXb18nNfAu8oOCTYr55mD6eXthGTEjjE9c00BYkRG
dGh2kKr4a0cAT2AIbLQBid3qxPk+Voxg4VAsHkSBi7Bcu46Ju/o9kmxAwYlrTlvA
h72BGkgkNpn68GHuDjbf+L+9qMjZraYICmAoFCx8gA1wb/XZBsc0PO7DFpW71W6F
9YZ4e7KutVUetFc1oUK96jd1dajeThHIQ6FBeEdDnEbhQSOHnxnzq0Yzz2Y/l3HZ
2hEAQZiKYF8F97scsez4coqbCkfHv1vlwxzFLIuCn88SRBrPBeBygwatE9jNEmmw
MymFZxWtvZVtyjU1D6ko3jcZ0DBjyRTaHgK1YwZuI+SJDc0gPTeNqW3TlAzRobGG
gI76Mbfz/kYCqF4MeyuxWqElNH6Y77aoLZVtaBbH93GJ+XlYF4lUbBJypRYEEMKW
f2xUEbH1pCB+/xA482C8Q7FrSjomU2YTUuhOPCPDPWV/KnQnNH5lhSdQlWiV1Xez
JuMoN+9txbiGjf6irGfXh291bW+YYwYgwRVgIg/MG4SQqEDcpL5+dwh5MQcFUXF4
rkRSCH+zr5NkbFuCv5eEJ9jnvwl0+2n8XVm0m9eK+c2A9Q3iJAs/83fWPZNOoTKK
h36oGydPLjKgDEkngPpUkYuhMTb/Ream27CdxsoJs2o/TbHZU2GvfxFWeFlCnsAo
HDlt5pE5cFT9kTINXaK+YROG3X9G2gApjm/5sB7r53XZjGS9ky3zbdxobkhmhcTD
8ZjUe+X3Fj8HTzfmH+62w3Wx2rOeElIDZqf3YxcytSdwJoJLh2cuxXAiqwtDwub+
IHplqf0oaDhAPq2qodJSeiUeoeBerSKdJO/wcmMMU3+qGkWahZtwwCCHGxmYsYsG
iYX2qq8HzYo2u90wl6WBdPZFtR0cnZdbR3c56rYnO9jIlT3rYhRKLxvbUK/4/7Li
l3B8/9EDebYPiCfHZRf5VmgJSVnfynkC8JtNqP80sAoKEHNg/sRteGNfwb2dpeNl
dqKPpf3SOvNAGBxjHmDoh8XpMOB/Ac3uNCsJkOgpvOfchsc/8P4ppbRwHKgVe4yw
VzrSaND6Egbu9dOFBP0q0ByE39XNat1GBwLI4IU88+vB7HxAs5pOSWsd+AxVQ50S
xribHiLHpwSLWVUdThIk2OoVau4DMBHR/Om9KVft8MFqtPR6RQQRfAmWWHyXqcKH
LvNWns5HodpT4AHxdF+xu6RCBcm00+T6JoDJp5B7LHkzmBzRJa/mJGwaCd+6tVGk
pFOk2lZRc2H/Q6xNa3o09js74mmBokjI1PJSUhWu9+yPm2NKDoI2nNzU2kMOVH1B
SpiDuLNyhX4VKA38r5LqKBSbNPd6svOOapw35Z7xOHTVfdEKjgvzR++zgQdQv2Ig
GIc4DeHuwFCsmSnvKB1j/JPO4VCpffVm3/doWZSobhDsXY5WNc45feVOuQKg6c5Y
xEua9D50GwYG39f9w5aSbZvhmpf7INT0esGz44WgqvNu320PY5sjwh75CLax0jXV
BVzMQPnSsguYnu6Rsri3Zkw1rlhHJab+QSfyUlmoY5rTrA+jAcIt0kmdfhYF6BeE
cIXCKUm9RRj7//Rxr+dj8HpUenk+9rIa0PErZxsF0c8X25uzadT1VTcNujYmjBOP
WKrkNm0Ek7J/lR2LY6gBFvIfPIybH4EzVr6JnZjlDIBk5jO8IlYrZqZlfnPxnCUp
ZcMPhScnjMZoXEvjLzJmhahfFI7xhDoxs+Hb+MRCL1dsSt4ysp8a70z4k1cS2KZZ
87gOj65xhIqI1JFJz3h+wrJnDHG5rak+CGGUqFYAWmLo77WvRTJ3l8sYhpWnXKGF
7N1yEz9MNFtVT6M/1sok7hQxIb6FkNjGDJGQW901H/0TT8zFmOLMxE6SrOVD83Il
56T4v8Hb0fwThY6DjzCiITxk661iON9Exy7iJx9cQ1hR6SKZ7tNj5sxoX3bjOr7G
fBrTIotcxZYqyGhrnj0+t22jI+bofY3FxIwGys8aKv7daX2bQ0PtqDql8wUz2oZB
00Yuc+NXAxxlyshKwBTL6G10Z5NucjW1vwVH9DtXrd/iSFgPgyS6m8+q/0uj3SvH
OxUHlJGATd53MQydBvaUz0R5ympIhakR2u2Gbal1k7jHMhMKS/iIN1H3b5J6VMiS
oMG0f2wc3lHzvhjZ8+qxz0XWdWFl2YPm1J9tIG8pyfmTwrd1gCynh+Luh7qwTCPZ
hiTunWzmSNVjC7trOm8pQFC/5miVNfPlVf+4La7d8Tfhfxpgkto8NYvDpB1GVtOs
pSEipDbpdB7uGKbkG9oxsqRBXJDE9TKAPaeJZRBmfqdCrpy7OPwPrnJz5deHDf75
ALGeML3r7n0Q3Z1M/oDuHaSPvNfT0dDAPu96dfJnF3qRrHlHzgHdc0M/8prNQqho
K+CnmmcNUoi0EqtDoVHnb26t8Kgam9J2hq+SWsDZMaFRgIqxlxQTvRtUvoHuU4BR
J+dbQmRVMq1Qqu49A6dJiHSsdVfQHX7hIIX+8cFjSniQFToRHHH02AZRCF+k3Wuq
Hcz95LZZtQY4gmJsY6bMXXChZj64E5WIONzEK+EJhySzTUER7/NBQN/y/3kSKbC4
rr9jMi6i5kypszNDKMRdQw6ahCg2S5BAhovw7TOiSj5OZlwhl5Txr/LsyISjd3Hm
vvNaJEx1ZWPOKKbtvP92O+ZKAtkMfV/DY3eDHQPODLMaTzENGElbLitpP80FuYq+
avJ+bGu1CiIDYB7AYRGc2Lm+4kaqScUv3CFANUfv5zlMceeT4OBVbhxvdLLZQs2a
B3PIgDxq6npC/12qB6VWlXxby0551ifkLUhrppMeNKUUlUUfhGFY+YYng0v8W3vS
xdFmoxhk7oYDGNoW5R36+H5EOMZT1UNvZUIzBSSj0CI1/ULczxDTUoMyiPhg8jU9
Trae8JO2DUgFvq19Q+t1LDv6Ajjn84sofbpSCKubUkfZuP6kvG7YLLI81V+eQ01n
2hYGcS8qrPOwaFk+s0uRFrcQfr8Ko1/YCloaPh/igKAamzPvHE4qrHwhutzaclU9
zzDmKf7X1YmcaiMM8WJgpn64WQDIHpWel2bxbyCx+riJos4LvlpvTxCOIMGu1Dj+
KmVKOP0BuKhMSYxT3FYLEGG+kE7j+Uf871pX791MRFi92kg/rWydX+G2yUtYw8r6
G+RncSmyS93gcidpv0NiSlFw/fpk9FOlZfFIvRsHFV0W3rZJAbDRA2F5AB1Lpby/
z9tsd88N47LqFYYa3ZwA8d9eQbAsFcyWJY25Pmvi7pERQoetyuDmCodBJ7tFBPUN
oOPuukH0WzEd+ri9299QkQulMZwgKSnhfv9FRsQ8Cs/kxAIxcpVonO9FrmjK+2H1
OJikKO2iSlw14ybHG7ln4svJc5KdnJYxEnzmJAYJ8FnLOb9A0y1SuB7zFscA6lEc
3lxUXyFIjYiZ966VfVdCBdCrid0WcmRaOLkIXvi7td4ob0W9pFhTS55dWanL4L3m
taKRVug8vXBV/agRW9mL1JgKKk0jW7lh91o4Eec8QXRQWNOmsRmhH39Mtk0nVSGC
uztdQg+2OgtIHbx68mb1u00mpFI4XwrYfGmKl31Ss0MU/vcCLxc0pKGsEkk3DMxM
3pIPOu2YBHB4jYZl4w5HIdQDJbuyDbb0IfNeNwEV9XJzwRbu3B4pRD6dvKIIQMXl
sbEFb7vZx9Q2Var7h7qp44yvZ3vzV/ihZEdphnXxCwGAm3c8qDeosKcoPtJMx2G4
cGFmIIl580lB6tafBw7nrhPt9xLrh56tPsIGgm28yVuibVhDBzkF41Z6+1dsDKvy
//6mjesUAcVU6QPmPOWTCpqxHhKoliFYc8SIt9Ef6H2b3BS/pzuf6GvX3zp7m58r
qp3MwiXliIR0smiFySkTrrD2XQJ7jT7VnotTZBP7yoQ+RdL3y+ypaOYxb+tj0P8F
7XqnwLiUDpyC+6XUIkL5PnYgM9a11U8JXDHDjWpn5+0MrqcLN4ZMt0r7dr4xwJxT
oDgzs4MKOKUoFHMfIiFh/+mcd8fteGwDchROo0ifliMjip01gZK3OoAU1Tgyk7Xk
kAAr66MHJioDocaUspYuK2/aklSPO3U+mGsA/wY3kL80aSt011DH9UZ5pYdRBN4p
fRv9g+dzSQp0/455UK0MZHWirid8OzaI329/F0rfaT+RKTyGMzPCph0LSCl3dnna
7/BXPBX8X2XakRWlMuuXrP2KQbfuh3WC7pCqI83UKW8F1uizp8FIpLqBUQYcCkIy
p0LB4G3yY/T6dQqVC/tsDEfirwRGWRyfyNMXc9PJZsYSClDbsUxHNiVLCcWAg5CA
MR+v+wXTXyiwV+lXrQTM/MYic5Qn7BR5Fk/Gj2hTXKMoz5He/rtunQdYTI8dViGt
nfy0pmaksV2pi8SVK7TJOhIPst1Xz1MwDubOGwAgU+UDbbW2pINk5QQKxNwcrsK0
1H2kG1iAkeypVEO526kNLcceZFWAI+3xu9bnZOp+su30E3wJvLTd5XSr5P3/HlLx
od/esOvWnk9WtUisAF1VUwf7J1SF9TRTKlwcjeCRUQMn5HvdaOSa4th2UNQih2dx
U7z72fc3E+yxHv6h/42h6PzLvyZr1eQ11gFLyWVbFXKkgZYdQCXYZ2UN/q+EtyNU
vI0fIMjZXI9uJSzIVxeL1+qPnZqkje4AvVsz/h9yBM3W5kx+W1WAqZQGBFCwAgbG
9QaixpTuc3z6qsiTs7bbfEPIXGhRJ8S8Z7ZS7zw4LSfGQCv7lQUpIN9Exa4gmN/2
7faYzg99WeBwzqxwIF6+TRY1r1VCvj3bAPokPF11gSuTNS/DAypGLgJLU3Q9x4nG
BG1psZFaBPPPTsrmJT0iQl/lt7Pti97mv/WEgKcMzK66tZ6dKZWgd4l28oLkpYjf
QpFaHCOIBCZyFtR1eQottMDT6aDqyOSvchxxwcW3tJATFrWCR+fJGgI4gTJPfUR5
CBJtpKmMY33D9yVmr+VPa7GnR3VrK2xg0TYwrqEJU7jskoGvpcwJxQW8uEjcNmSe
xxxqtcxqSoXzU2uPwKnmbZ2+zc5bjal5s6w9jdb1UOVlYsaeD5kbn4IdXw3JB/Bz
JgTfsbzTNTG0SY+2MqmWD0GGjLdXubwrMp6vk0fpA5fSdNrXsVtEMWgIKSxFQxVE
JzkPZI2MsFK+Vi13/IOtTGP6vTryqpKvyXRJT4Dd3Nv2UVcfF987UO5LHfuljgU8
bwv5OeVU+vWgzJSHDDygMr4N6Lb5WA51HpL964rF9TOh3d2vS269Ni6YGpjm8mIj
qHWdAl/jjMYzXkgC4glzyoJgU98ldXMbhSpvEBiM/B4G0a0X/HduBRkpVHJaeQSe
LxO+qLzmLGAKSQch/3bibonRKUF0oCUUlMgEmC9M7lziupdxHlKSJKwequh/g2UG
wh7j+JwT+qcZhnlMqPggEgnLSBw+2aDtH3VGvqKgHM2Hf74mWTTDny8vVQ2QPggy
q+urMUKXsRPWeYIEXB3dbcbiOjFn5fA2Nfv+xXS84mn+8r2V58Oa6q4d1OsvLZNA
nP3Y8S5kWPkjR4qEeA0NKC0IuJAUmCWoDai9Bndf191wwkZKoRWbQiui7aZT6Ziw
6Kyr8nhjJkbFe9+R9Rthr1p0aGeXY/AgkKAfkRMypj6nQ3IcfEPkmBibRuXb/NvY
duh3UT6R40HLWiws5r7HGS+aSjzyLI3Suc1r4H9BPmuGsvj0Z8QIFY8Va3BPrmvd
xsRf7xFSOTyOgwic6/UM9fJ8oSosdfKM9xswnmKVxqwBNINT/hT30EmpkwfDFi2a
YIyE6kgJUkCTiFmjGqYbvNKe7tnuq6mS2DbQRwYVC8Sy62Q/OEyUOR7ALivJOkn7
fUIcz4eYeeDSc3i8zKSkhFaf5MtERdGVsbQdjw5S12P9QUru7LSKSmnYGG779rd6
b4GuZmDLmiWfGmU+aRkqRA0dmjTYYjReFEeL8W7/aiWKefwj5ALT99i0HRg9VQcA
eZOjlAttfHd/pENl+IqTIPG327a+1DpO4CYyqAhQSeSI9t3unIgimO0pZ71VBiuJ
VYiN2P+xy9Te3Yw8I5/x4l13MxrOrxZGaBhKsRZhTmHdraMkaCuFtMxxTi1oZ8qL
AwhTf6k8gYH2UTZp+OGzUzua7B4ivMk2YtwwESx1Yof+JEdh/0IBk1pUKyjaNqBJ
bkwqZLauitZP2pO5V+VUmELkSS2u5spse4EpKQ9Ld9SsPOr/oQRStI4ODbJEtQSA
MYizRS2cgpMRLFH+tIcktv7FoRUtIPV6qXY+de45znOqLZFQ9wVdf1svOIhDXrfs
mRBtTuzf0T8s1C++upJFEuvHmTTvVINvshBbxR1STNaWbwkpEklNFdpqoSYvW/oE
015E6NsgN6DB2T2HLlwYGD9k6zHZZvAWrxca3+1NdjYCJUpLEYrUp580qQqHsbQr
AyswzMx/bkcaGq50Rur9n3Wwa3fkME6dKS0d+R5T9/dcAlzM7cVNy30Y9rzIs5gp
sW7vQhY+myjWuXviN3FX/h1nlnhB38flI1XozeGYjXwECD5SVs65psKCpIEJ28JM
7uqtqM5SJofRmWHHF+Sf9NYskO6XS337vUNyEVm2v2dTlCiJIAqCnBq7nIaeUT8b
XHaegTG91C3qTHrn2h7qobKGN52+wJLMjhHHCGkQKBFVoTZ7Z8wkrkesXOf2ROSX
2pWG6Pc7iI3/T6cpNGY7jXWnXhov+UMIemKDOYPeyG71ZrrAtGG9gxBiTkQODlsE
OELYDwCldK3cGM29fq8ExTvYDtC5B7vATvsZ+lGYohxS7yYXp5MtV+jQJlRRHEoy
CG5/HgF8lj5TLO/xLcZFAhhSATPJglB+3fgkZz7q2DftMjTyuaHSMfX3wUNcXgIG
1BkrXPHwo3q3KSZmiLTT1of2iHED+zoIhFs9shUhW3jIMV8zJawpFnFPTZq6TYZE
t97c5hyfEoJuuQSmVJkJPGB3x66Nj1sJaeSgIGtsaJ9NApuagdfY2ZjaE/6HsZKz
cwTIrwyYOMPdVwzIBvlwnspNxWE/IfLXyFUedDESn1BCBc4wOL0+FhD+geFSR29A
qh3NZVSUNSzjuxYIdD5m0Sx5E3Rt1YjBVtAhloh+z6kYC2g5lNhso5/ohBdzEjm1
Gb9+JNJWCKK3Dom2RpqLJIuAYJxS1pM/DtXHp+M/19cpzUR0FUW4CFI2d3DvgRov
Du9ry4ni1vyhbrPm5AcSk+m4U+pcUT6mGQcmhMoyNuUqW8KtzpNnnKjn0F8n1jLt
HmwapSu0z15fx3CLHDGyUWJbSiub5e54iD/1FHLWhPYxcB2Ol79mjjvHBh+O6OZ5
RroivDuPTkEbMbnee2Y1D0iUeOI++CEeoJsIuUv9j+aX5ns27cpuxDsml+Jn1NLj
LKZ6ucg7bUlvYz+EsMyLKClkerKjTV2DwQhjeJRD6WWF5hye8pUJ9oLyk2w2wgLT
Ub3PILXCK37+cmzhwAeDrEqFvBW9zrWTPFiWe+owlX0rpjJmOxGvuqtaOOfcS8u0
xhOfQu3Go4QDWbonCArqZw55OpGjAIgT0aoj5+gt1VHwCpb76RwiBttBdQVpUDa8
xAb/OApcriceMKec8uTD4KK6tw4fmompFcM+kTkftYwMkYbKBdmCP35vp/g/HMfg
670v/by+jklvFu/dO8CG8/TvXHooRul60/DhVrk4Ob0bsRyh4VFHEp9Jj75cLbAK
EkHxETcgcLhMYqUVd8EWEgpZ1I8hkYKe3MTWBEpLBm4rpGJjBFE0F9GGiY6TC+DF
BGlShUqM2RId+iV3NFqCMbvwRbskYoECkn/6HN8s4Gn+UYoVrEfoENwB4cqseSwq
9qHCmo7rfjHnPlYfm3mzf9/8wSKV+eg0ISMFxz9jkRmXWqWtyPJevq8tZ1ffhJdD
rUObbT7KkUTsjcCz6h+0+JIb7fr3WZatVZDom4o0WlSk28djltUWUy8LD5KRT8Ba
x/WMQRp0oD/mAuI4cwREM7Rlhs9tbGVpnn4xQL0myC/svqUIvXzZQMv3pPLl6lzw
iySiy5dANsIUtxxsB/toEr60MmseMJ6lqnAOEJM6SGzfrsaRSrEyyj9EffCw4wQJ
NRccNmYHiuhKpHr7KoF7zLphINL0ukzXWby0eginscij4nyA2MxTjlTtKoGAsg0a
3BY0Thxv1T9uLzk1QBU6bzBfGMnIoDsbxgeGMfn0L/dytg7Uen/HsFJl/CtWpTZz
Lq/wa+DmTEWrQ8fw6A9hHmccZWEd5jcxweUCL4ZQ5nx8N3qeLfYE1wqncVwrsZHI
zuwiP6aTXPucx4K5HunWDEbWifOO3a5gHTshhCoh2p4oKSStDSSWbTrAkxc1/2tT
GBTeRX+10XacheyZDVF+mPnZGWQnQlcf3eOxIndVLOeeLD81vqlPp54n/MSb4SxL
ZbAxNiM78Js48eLGA2LzFdsEm1uW/CTBR/dO/rR825UOfV3sHXqi7DFaAZs6r9KC
eLYuCHIrXakpoy0xntwZMSeH+TFoVUmJyicjXqSwoI/l0Ul/s9BGbqEgXy0R2z7V
8doKDy+e5WVecaDblWH/uEf4DA1nO67tZXurVGH5+3oM4CK0JyGMYrAoG2IDnTkJ
kSeklXhpJKKZ4jio5M/YksCd0jUdTNWUjJUL30sZHxrRRISm2rtEIRE7GlErFHKJ
MK98zsu6XQT+xK0dJ5fnZB6KkvyfMdAZV2xrrFS7MT1Wl71Wz2UCOY7eTtB6xE8S
9lKGQ8SqW2c1QOP6Z/rbTgAqsjGQk2qjCss98hUOgvOz6lGMe2sw2R3iANO+cjwC
bZ4wAyX8FGS9ZVkoTHsFEsRH/Pm5MWVn+xssYLAnJ3ll8+X42VY//FyyHHx567A0
FD40tHHdR5HHOadwqOhxw+Bo8dzmEt/FZPZQ33pTEAiVTCR2Jba6mmgkhV/zxSsv
9VjzHKswikc40GrosDJI1QpYfzxxAkJsfoV3ZEcX1G8zrwFPStE07MJrLZrPuhNT
9qrKUy1pBozf/zmLMrX+6CzkUij25iBrPGQhiyR63ME4ed2w/JbTpfOHTWzcJGs0
hQrF5uPFO/NHGd7mkBWp+bDAQ/v8TpgDbhPA8dEtYQ1YeD9I0zlWP/UMckYaaqA9
9s9Rp5y569mGc32LBbCNfO1w6zmQDDx7x4+S8NfqbIlv6UIPDudne40damK1Ow94
OxG5G+DREbSovtPy6AIG+8/9oiK6VmlAV16/3AOq6EKo5GJFXxYfgSaRzzCJH0wj
LSb8UiMeLPtbUboFuKh0OXmQ8tDCN8dfsBB11pI61ouyezuwTRpki/K6I3VPUFjx
Co4YsiiS71M2G0yNMYQBe3HW4+IxBz0PxcOWyd5dBvyAUJL3FMOYxEqPoqGQKwqV
1yKeemgKV1899Jyt0vinN7w+JUo6wHlIDEA7ry+e68m+DP0K6fGZSdEtJMAy1nJL
hqKAb0VQ9GOy3hpqN6LtX00yaDsHFOaUZnpvFbK7fq3AVh5d2ER/PM1Yz2tJPlnK
omXW9xHUHp3u44yZ0X3+iaFgZmKcmRZyfSdOCXohU/N6/PBnXR7YAOy/jnbcnj2S
wDZwHgmrt75XzI+syfyqIZjJnOn2wVInmdT+pTV+ihraDLmv8M/GAKOw7r4rwutA
AHp0bYTUaD0GIgMPyBalrpTA7LSl0PNQRQjCDfebZ8hskRMWq1d02dJB3m1bil0F
klC+eC9iKkk5uRQdgGR/o8Q5Iy1n6Bpa/4y+mqikLCylUP1TM890qXD8SCE2iUD5
ttW9mX+U9IKlxspVNxYc6t3y1XDPpnoqVtX/aRY1ujqdePg7mSLqbfK2KO2zSZkO
O9Q/IHYnEZu9m4dJpLB7xU9Ygx+trkUjYSmPLBwmxGxE+iB/6MYWzyItnwT3ewSf
u+3fR5al84xQwcgvo1/YMZ8RvcD/+Fl/nCLqq9pYG2DUNs40am2rmOsbTLXIsP3I
tJm/4X/0OfJPWKm3R6KZjKY423oVT3G8ThHckNSnGcRWQyVCAbCEbkctrigTavGv
0Sc4klclLpOdRI2V6xr2rkzOenaJyVC1JkJp4hefiZrzely0S8TngltNTK4rzrXw
3VfAUIulwQ/Y4SGdl0hVviHJXNNZAzy2dS5j8kKUqGJh8oUxI8AN+o/O22fN+bSe
o9RB0ZM2sRg4kz/6+0aAfov9fRFvZdQHVgcA9CHK6j1ek4WM7/7LBMx45+Q69lcq
hkKgpUOqB3z5j59qiESX2xrpRjLnlNGT5lWr1KBr3WkBzT2ALik/zbNgsLtgEznX
THuAlqTJDHbotFLkZfbOsUe0b9HjS0AwU6jY5KOAl1cDRaC2lKy8HxHv3JjFk/UW
cb0i4AouuH/t56k3ybJF7/Tb9emPB6CPdlov7ornYPmmkXgTmCeGGKPKEUG+hmL8
T1evjXg35EbF2WmjMD+qKb5E7Han51F/RzNDPwLITxhUMbcqvN8lLD37N/NlrjyK
P5HlBM1Wc5y/3IukVw3ThVCL2gNcm49Kh8g5leXzuYpiGTKeEfobmfAbY6shLYtP
gPebYnXNPMZW25rlW5fFP5KVINXThiARKXu3zt1dfhZMkZRo/SMdl1o9gw4yMK/q
qb5UGYrWPQINhPt5Xw4t3qjhW6ZCriF8zT5ocs1J5Owww/JJn3r1q/kP9Vai33jn
lF+odnQlJOXw7/AlKYNise2Rlxv64M2TSxSllOvm0tsL/UWXzM99y85EFiwk/8zg
URWNaCxG6kkdntUVqA5Q02mg6wTybv9j8V/+RE8bvT1rf4f8b4DbYpRoEgSfbejN
iltAsxDEjaBqtfQZMKOJrJWfBW9I2vf1tQKtr0Q3wugThZeaFGwhY0lvrmvmrHxk
30PfWL20GbZwHZK5lpqfxs8Bu8R4I2Pn+dVGJovbOE6MpHKIBEFPslzwa5Xm3DE/
vRUXGKS3B5EkaNthRY6eaP3X8CrAjpPJKQKpcbpvXMhNFXK4yqulUcJMMabgmSHL
LKi4YmsuZ+7ddxm4iA5da0acCnQzq0q3DOSkXz6DAZSIbAl6Y0AxMbCMbaPBAyOD
4gesARK7Nd7Kd2wmAbFdpNg7BveNfSjI/q79I/snGf3+8LrSpaEJojT8Gvm7dhJF
nXR92GULfyhlRFpP1VoG/NIZ20WEaKpAKHpq65TLDt7KKGekMbrcFpS+TLVWCiHI
o2coKwmAwii9unGzgd1ZkpWBz+F5yHwnwBvUnckMq6jp+tae0AswpAQx2Irb6kEL
KOF5K6UKiR35mAKb2JSaIB2kmy7NX/dtw+vmAnctxIP1OgSmBS1YVWudzJvgY/ot
gXgs2kMeKa0fWd3b9dd7UnnSY62eRfpnLUC+2MAfp6rfB81MyX0Hx6VRCKdVx0pg
+8gb7O9KfyFzqcwc8IOR0+Jf6vCM6HLQ85H+HsGHU5/Zqsn/6pKlyqDdmCnvIxos
caR/shVy+7Z805/yuXPccg+AjovIGLzxWf4T4jgieP1GhF9JV2QLdqWdfQhBx5HB
S42NDOWWcC7Pt31A5trT2cFwAxoiRtoSDjxcPm5k0SOW9tQUjFcnGB0Yt7rbTzRf
/cw7RDolYR3OE8C87EwAz31N2SExM7YngGnHtURnb8JlJFkzWzggmINzmy+7J+T2
z6q4+xRSGUo2U0PxC3gpP2QdHdA98c+i0h7rCq/vi6eaZ89qAtgffIcy84ClQg4Z
OfIvXYG6VVW+tdPnNiuSaFmWa9zUlo+JPydx23CIQ1kld4cEifgu+bH61eZnaSD2
A/yO/wF3hj3PB2nboeZ0/qiRhuCo6OL1uUpYl/FNsSijblewu2jTOsCI57CYJWUO
/siHe+w6/MHeunB6XHmtL3H31mfFyKM3epGqXbEaonaCFN88u/qdXKQo96z2oVZa
ylhEhr7AxfrPBvNUsbONQ4CvmC6OY5kgqpsM54Bpirohbd16HbGVQHKXy/2fC98z
tWvDsx8UCqBC7uVRWk/ILuhZdbPKVMkSQDMVZIjfUnHHCjJChc+MUKaNcB8vcDZV
unISj3j6jM58vEYgDa5NNmEdTBIx4Ql3VzkKDsuLILHQ8Ui4v6q0YyZUmcf2dbr7
Q8/97dPvlp0ng6JyREjTWC/eFE/7wi3NG98tgHqzQ8mWZNvQYrwqeHP2Tn/u1GmV
cxOjFAWE8VGoz6RoGrKglW4YuItsLwo5Zr/oh7VB3W0GcWVB/ef7+S5EhnmYCWsz
Tbjx5qEP6qTgiw+FuZtHIch9a/VYq6bKeJCCpofJ6iK0hT+tJ10pfAupH0LYbFG+
vrUXd67KQ6XjvA+m5/qyF5wqPVCR7w04hXLVOZCnq5lY3rCpjS61ghnk2u3HMrLW
kWk17dUSJ0jeZWaElmS2O1OIPZPUt+p3ndnCqjkluOIw5F1tBVSQhFbpIlyzdV7G
a9sTEegVlsReoyGGkObbKyeKEx45SsmQgm95FzBWqApxJoFbmFUrbZeLVcSWNN+F
JrU1UNP9L0ZKZ/M75aKM1TonYCZhYOcu2dCQgjdqnDk0c6ND6Az3HwV9hSHzoWtG
bZeJnoxjJ85huvyrfmDYMEsQUTpa3EAR3cIhnnGYI4AQ/8tERO7Jxv7T30HdZ9Gm
EcWFBlCnOws45E4f1vyePXZv/O5IBvAbiX9gKwvZm045njFKtvYNvSuKitJLYMps
Oh6NkYL6xETfTqONU34wtPPMxPxSpDPnwxl0QYXYW/3iuhLTuWoKzurlXpSRHBbZ
m/Pt3XKxDZRCBvoc48Kbk/5oFhCWMikUIjpj/dA7/LoNS9EnB+vThWKJUbJRfXka
h80TYetCDpP+5SnENtKoku9TrLNsg5eMJLY4nSD1u0hUHN7W76bQlK6e32OPhRRR
botJU2+pkn65gKy8t6aPDF7jsfHLHfhtIQnc/afXdEMlrz2I4gUpP0+7QHgRydyJ
05M3HdNMGnjuCYByiJByJG/WW67wYk4i1MbMvTGjlN+K1TirzlmTJIzzTwFILuyD
z/EHbddOLAYj8NlQYKyK5RQ4mJK5bGwbHGdxX2NGJn7i+hNwBigamE13xiXVBGjQ
91KPRSK2H2wvjgoLV8r3DPmU8I7Y2KwKGN8CiF4xMOjhEdCTA/NdObqSExuVaxx3
Y0AqkrZrrmrz41TtPchhhaQpX+Er6ARAzuGbGpzB4QU5eDCepBQAij+981JWCIl5
HZJH4rgyr6EHoEA/RWXNlnhqvAQGxNPxs96iZoc0NysufLYk+937wObMOXj5a5/5
nd5Hsbm1ZF9DIIpBqhR+9YZ0T8y4M/MlNcaVaIbpYMQHvHJ9f67JSRvx9Ytvfi+R
PVArfkVDLPBtJgEHSbkRo6FBfmoxhcZaoKre6uA3zGnhFznqagb/cHSCqTXfolJZ
LH6DVR8NTr93ju8h701UUSDsqqteki06qozA2RMSl1tG2W10HSo38Tfn0qjBB9EZ
27amnNrqqOUShLaxjeL6K/xo9dthb2ttZvA9AnKWNyndSIvsyHAeESpt5QyS/I9q
RWa1ubOaQ3LIb/Cs10XPgVoDZaE3jkBhrCPpecZnAzNpOJzYCTdSZokVLEVC6sVe
CU/QwOYBhA3odBFcvaZrFx1ibe9LPxK5Z84EBo0qaKkS8BOquTOLuzoVo5VIcGCS
U0WuyZ2lzgbl4lzVb/XHMwZlSjLxUZhPIyk5IoYuVqclMp4W7MSH2uBLwjLFZ2XJ
TXLzAb5bKlzGXozi7wbDhKWLk7ZbHZDXulT0a4j8Q7Ipi5ArvJIxH9ZwOijOhmnu
FQhOlUQfvnBWBTV6eYdVIe2qYm0hjyZIvPcn+SLPZ8xbA0WcYnfeWwVHgyLVt8jD
EGoobuzruJRc2rcnFIy90kTF36HyRpNgIMrK+P46P0c09ah3IhiUV9ODHdEmuj7s
C+k9z3/WeyRRHA7KpxM+m9t8xhB3bBHrqAuf6bYooV/Xpf6VwOR1Em5xFXlTxtpT
Q6ahsEZXLKO00wq0Tb+O5iU0WgX/I/QSR4SQZ2XGkIGrDUbge4n8Wn2zcGrQOffg
iKp25na19BLZs61rWjA7PVlYBiESTOVBjyTrXp2WiNNSKeczzCdUpPBZxlterOc6
RAREkAbdJq3Rjgg3ML4ZPl++zGvVa1GI0aYt6nSsrp1bEyTckYQwCF3Q6gmJeSg5
4dsELjn0j15+dRWgSJFx+WhLg8abvDFSBjJLGKDQuVaIR1RPVy1TBYcU0G3Geppm
EYdRqBs6bpGqearEdFDeSXe1/lOCaQEUWlRTvgJlREa7BcTZCbpt3t6CSBCZdOXm
tivdbSXr22zAOnNUjK4NQ83z30Iu7MU7kxFT3ansXEUyt8tbDBtoioSm6Z3ECPyc
3fIiNE9os9Il83iN48QtyqjOgqBI0sPAOM7mw07zGXVu+UveFEgBVfnpG8LnrOop
kJ0YhsnTCH1oGLxVftPYxp4qZgMSRL8pb8KLlqlDq5Mf1sOSpcj24EAZ9D+PsaYh
kGXyQoEqd8SPLecSg8X41femUZjTtQ07GwUvOZ+VnTO21iooPBNfN9eEZKIVw5mp
wtvwo6et7AVpdP4LIHkLMRWMIE44aib2ydby53JmAlM0MPryMgtXeEkcVnSppORw
pAvc5ka9xal4l+NCEoqSSLgcuzkAv0T4y58ZkYvRnIAs/g1imowuJIseKYs3Oa1p
aHui11L9e++VHfwahV1QyLav2zfMhTvlAYEYtsCFG+M+5oTojUet0v+qCaOKVmsZ
dlRlE7mpiwnqOwtssPMqHH3Vg95orEG8yToXF6nCqvY+uzxvKdccXhUsawJs5yeM
iux4ANPW90wk2C8182IuyK3TNRc4zxk+3wFJBXRyBqtg51VN939rQ3nBI+XkcL8Q
chh3+Bd3zMtksSXOz09iT0vLyv1ijM+XKwHvCqFWqqLswcyMCIbhVIyjBLv7jh71
zL4AekPcF4aYpra4Bu+7X8JEocneNKmDNt/yNWBJwZ+obMiuttnedMDnNbvU+RXs
r5BDJBsiXket9uJGQfArNEMSqRseiAWk529mwP0ABD2XQtUR+iUCaxbqf6YfVTwG
bwQYyxzQqAvncPrru+J8XLQpb+pyoykbHyhTS+4VZywzOO12nYCD++615jMc0mrR
MdYiO6KxiKBzW92RsQRq/mqpZta/BUWsJrF65j0QDk0gpR6OIoXGkR6zdSKkzFUL
O21oTYuj7qT0kMrDn4V84tURs6rOQT22ABRR1kgDyapJMRFZlQFDkCQipyGT04u9
JReWaXb6C8Pg0ZMXKB1JlTc2m/T+Uyo/CZ3sbURPOSqKw1qtGlL0+RcsrVwmHOac
dc8z0UcG5MK8e16t2MvX6oZI6w91Ucu44hghZCHG+prQgtyDYLcRrPIZ7lXfRa8B
t6rKPAcUOTLDD2qxCxOGAQpMurfgW6V9MtG0jWowaU5CrLozwXb7lasl4J39dqHS
fLS8kwMtOcCTKhGVpiH1uWUY5LV7wujfFyIiClhT4WkfvnzFNnLRUlCKjxtc7xOT
thPxZnnwsHucBTirLeBW5vJy0RiX298HHGHwfQMRuxDxyyrjqhAhFTL/rbETJUcE
bQpaxHMjXHSXrqQcDL8q0wtNeMdG04wehbOEwKKv2jsGUFzJF7YBotcUdeTfwzOq
yrH0bLwxr18z7+7ri8bbFZQ+EzLblLppYd3b3yV1bmXeGBHEKI9HQnBrSJC0ghG/
IGOK193KG/+GLMpFp8jusggqT/8WkdL7U/+TA9lCmoS7IdCJhDB4uq4zowSqD2om
7oOaAJ8/wtlEJMCHeQvmJwJzXHsZYICIAxpvtGF6yANBgXINAu024L25BWv655Uk
JhY4q2L+GVizE+W29EdZimBj/GaZ1pjTdBI11g/tkT8pagCLaV3JLF8Ah5vy2g8y
UYEaxFMA//TxZNxKmLpX9sgh0zfajSMk/9/i/CodZ2qlcqqDKlKlW+HGQoO0UV/v
LxB7WE3jCIARpQR7oeK1NfhUQvzyHyUHVIDxWIio8V3aepZrkrG4vtu7q1SZGThG
BFNBpIKOMOc/x9lj4rn96yGw+KtdCABodFRL/AC4VtXrVed9KSj8cbiYM62PoeyH
IZMv2Gd2vJcfXnkXl0xt/3fScmsDelqChRpdas3uXjO8//qE1gndUGZZJgGjJupG
JsAw8PsM+0S5xwMfX0l+gHjy0JzxFhLhrb+gsQyNY8I2oRQQdoPBHRLqv/zO3gH/
TgcT0KUk7RBcHupRcFnnbltXrplVOjiX8fSVoRLa9CYl2QrVB/59Mrw6+vupXN07
XGuVjObf06GAw+X4+1tuqRSgUG0KNY6tnncoItrVIlAL/KR4cdG853/Pwi/EorL/
8To6X4bY+HoHsAV6B5duJKdHTZuNhmiLtikUV6aTrWcZ4IuEjRgWtUvikOfTezdb
EVs8aEQmOyctA68SDSg8QuExVr3CnB6VUKw95HK2H2J5RS1hZkOWYFZ8p5GGhqA2
EZsmMihoBIKjP2NsRnqhGywRhZ8Yqr0vhW1b3S4UDfdr/xmS/cK4SYluofUT1MGv
s4zksKZ8aSzNteSAFDUzrKFMVhbITx4SNzNH595tUlJHFPei+VxLt1M8NkapLuLn
xCcpKnUXq9q3bA6dHdEAWIKIPpek7GDzs4nRnqGFQnqxlRPx9jDdkHUD+teNWHiX
MXDE91emVzvGa9096IWN/U18C2gBBx/QEq++OTpUSoXhoqDGsXNiJcnuJhP0jHWo
fBITawtIFtM3y05TbSpavlRTF7G+eSH+kwmfGPwUSms614Kmeg/3nqfa18Xaq178
s0+yyEBrozcvq1OlCdZneFkrrnbhVypD0qZACoE85h3aj78FHqYqCGpRFRWAUCTp
vyzhwP+O27mNZoQO30pXq4uVo/Gn6xF7HSKCGnYQsKMvjGJmaeqybO0XA1WcuhAP
KdQ9p3g6QY6bAIbaOZVP0/tBIuCpiUW5nXjk011RN+8gr006n1Inb1blDe/awkr1
MsGji/qWd7aLGBexoNb4DxOZ7vVGu9srV+ms3HxMobLOKHnXkJ5Vye+IXBgBEEx5
Qjqy+2VXAq+pBc85ek6xlRI9Cn3HnWZRjmEKDZfkTRIeZwbSIhwuy7BWalMY1iHR
ihY4g3zHuwT+zwZmk0Q3a0dpHyaLYXTIHK8sMaUeISzH74w9H37pI/W76Tu0WzQB
r2tRpu3nZ67vXhVcCFITKsw5Tsj7dD/y/UuOFFExflm/dnTqv5PYz5yYrDaVZsyi
wtbDeDzSzWXgZdx1FG0R22fiJKxqvBjicogIhta3ZfaOGr9o0eF8s/0tYzoRE2Ot
QAQxi65RO6MeS8C+pATpPNQ1a+2onfjbTl2xZKXgB/+tjGzJ6shfmpm6YTCME6Rm
1UqtJm5SJLaA7Lv2R1Un/3+KtQYb5K1VXY9ftynDyGnRDILRHcoo85eRK/8Yvgx5
j7rhvJcz6vx/+l18Dkzb1xq6LHpz8nFEjYTPI5ssv2aV3PScwCEJEruGpXOoVTGD
/eg6VG6NQSrMkNlt262UhDWO/vsK6emPH/QRR1vox0eQmbigjyWz0LANEPqWf0kr
VkhKJRhXfhMbzd7pxPH4eHLHLPpe/Q9nI/rr4kKG/8QWMwgI7v6Um5UCRGibSJKL
qAXsASWtyvo2CAu7yFjqVDL5x8+Pk9x3qrcw7chBiludsXB0CLSbtMpZ0eiqwk0K
KLcGPS095UyHp9L/DZQgla/DCqP44IhvMfBhgenk7kK4a//eHMLSe49SiU2FDAf8
uyfU/XWgslh3OuhHbPl1oULgym2m1sTe7gMVNEJNC7z+ak3B+ds/gCWDnQdl6VMU
06DQ3ALrWzb/VA15ekqZgRU/jPwwMdeKU5BuovLlyse0yAMjBFtXmEC3U+n3ju8V
iUnXWtgv+oLWMTtTrjVkz+phidQRbKomvwzwQ051qom8d5bEtWzMQVZDXgf53+Pg
ajrrOTfEg3OMGoiXcEi/PCvcxQ9hFCC1eNA4edTfGkvqY/Y8LpCPMCV2wIycDhqF
7TDS/mMScnDrVAP3yUlDBbDILdMO4ReXvA5HkP3S9un7jR47nr9fFOrn+N59SIW5
UeQANpOZ9Ek9NDkQdjDooMEeACGLCl9pa4/gmtkkADXRedj47xcWkwukCunlPXpi
c3ZHv0AzQXdZOVNBO6t8WsJe3N/VGMR2qGA2Lfp1AWR357XhRNGKR7hp4DizXmHo
kCPcBi1F0RcZIGgQxJDKKOoCgnLDPQp4y9AByEWvMBrbz4G8zwSe7uSVQYQ0qdto
v7JqF8ArmfphTDO4xjwQRjQTlEOVvE5Hs4W5aE5rFiHpOMmz+eMOGfcMOZIg+idt
ejRE9JwmXV7iB42vreOUnVw8iuKXUFJxniZ3AEMJvO+R30KaEF4s3CWTEiZMMrBW
XL8OP4Y/SR34kI/sSe1b4YnOFS551YoDlQ3sZEEMepGl9BMGyaDg8tkkltg5Gom5
gej59lQa4v9iFEAzkv0jSaikfzuAlSvYNbxnMYsyDSwUoLoh+FFoxoyv4WJDqJvb
ZJRpbXyMTxIZGXSUUjMAyDD8MgKWl+ELOcveakOgyDkRHWzLRTB8UrfyhRD2K5IP
ox99a7Ikm2TH03FAbMjKBJQTSoEmeVrweOQoeCNRWbbPxunXemIKhYr+xan/e3+m
QEW9+M+qih+6W5qLAQI8WguOJlr4hcH8cQnPrnsL3zfuTWl1IwtMwH/gHL9N7BLA
GIjnllAXiWEFguyVmdCoxWa4GC12jy/zqV0N3Q5K5+U1yqbLOfqFO5t8suykTQ5I
bOC3FU/w8EdM9skUjnehA0+pvuJU8/hvGnFkNXuucbbtw6L3K3q+aE7YjdGnnGku
p2I0i3FsVst5p+OeAD2EyZJlStQth8J/GzKIdSStHUnVdZwUi13tZRtLCl/7fhjd
PQqAPDslnFI1oOeWYm3mIqw0pXoMxQfZhH8k0KnjkFPb9NbENOKArQvm2ewLlRaM
IZtIeEH5OqKgGgzaHoBPmdwnRbU6LpysDBe0vMJxTQ6aOFe4B+dY/3KKSKJDjm51
4iXnRXQNnPtLHQuyJn/jIx6UAXH+PfQ6JLTqeRRqV/xz2wzdLfwrjGnqh+D/0o0z
OtifQXA60vdwMizLajT+C2lGyY3ar3anQfHIBZqXDbT9I2ZJj7uigBbHZvMozwJC
9UsXS8zZiqgvX+ABX/pRlpCxsV0qLCuqxXYc6l9oIePeuMR1dc2wr7cjTrX60UGR
dVPTAgbd8S3ncsIUNvLYhVE1gQDFLqRdcifZxw309jIWpgiljrFNKpV/eZ7Uok7b
3HpsSZl2LRl6ltMbgnjMzEUBQZaxoy1wZg0Z+KIzvtEwCdWcfMb4d6IJQZX2dgaM
/X7vbCc2IxAM/KMrvm++j5GGQSEDeteEMcJxu6Hp7+XRDnEAffIYs62VesKPtFCU
3yTw0QaYshWf1Qw6Ik1/ssa5F7I6H/ubj4DGx7qRhCe/BO6gVcTZa/Kj1LSft31a
Ika8JmvAdhePZA94ut2EHeoNCAsE3mZBut3znj2xaXwiI/HcARa6d3CZiiS2iAFR
NhXziViNfV+bbjUNNdmmuMnwM4q5SuUetiBiN2+yZodfUmyGwZWbZXDwAHcduE16
MQAO8OWAqB8J7ijAH3i8hSsT/PLi0daD/6pR1r6HzDT2WFbPX/BleAm5kFvLpWrq
y35Ihgx12lRHQHz5bVvNsrGYdIDoQLEfg35XPFwupgKmYG9GV1kY7WRFX6YOqGja
6g1FJaA868Ki2rFLe4zGt+trPk8LpD+aqf8AgWH2tvalloWF23uAkJG+5vKKxPAs
eRXOwI3+Z5PfApvLc8Zk3QAx+KqFnv9sfBiTZFeNVTs9Ue7JtFp2V7X1JNjN+Zbh
Ybz9zX8hPmqUE2z+cMhvN1GskLp4/uNRPMbUTiMCk5aX+UeinEZu3iN8NpBmKx8n
qQsv2WrmS439Qf9vCl8DtElcO/VDVo0kE9qwlafbYAJ9lMVGgzJQfpWXTYOx5yrg
8t0SIYif5pbK4XIGqAsb1wkw3+aK25In5m3Qo20H5NSakD13OQU3gH2c7t3MGe1F
wss1MUoQhw/8s0K7ToTAqeg2YYrRap2/Q2ZqC6ic0wOFmdsa93AhIB7psaNzw7dD
bsF+yeEv9iCsrDWLj4fEIvxVxhdNDC8StRp0900+wEGLRDnqlmxFI0Vx5rPL0O9l
L45kFDalHs8QuGvXtTQRM377IIX5iQtJnLPoeVtlblCK7RBA74X5IaN2DojvwTjR
aV8MX1+rQ5hk41zGD8zMgDnhbz2sNgacu3W2YVAmBSuOAtXCXTtGDHc5NOOn7hqB
7/8Ng7T0bnS+6epZLCVEhtKn3cnZKhUtmDimizxsTAwSamCu9JMp16g1rEWnQypV
yb0ov6jreBCoAd3t/p0lZgogy7N47zrtKfXfysrHHF3A1W2H/OEMrqZek07f8Sd6
1ZcZxpuT2PHAYakkkpOIgBh3PUxVdpAKkarnwKD7YvXlR6QYwMPfO2VL1NwOF1Q4
LLUVXclH53dxxhs+zHWvM1dVZY7fXWR+1b2GqB6W3OidCsAYTUsb+awUIAjoo8Nb
A20KTl/h5wlIJk+csecpa0s75S2hsKlIqS8vNYghjIT9wRP+Yl08Gq+czrPTD78Q
P9MfZ4v7PtI0y6ixmRggBVXbsXNZQRyCBxibuV4/vJERHcsGFGw1aHK/vPTNsVia
7jcFAo1bkzdKUO5se5MhCxO0osTML7z570eruMEmmpul3iPzXUTmOVANn0sIusHL
FZ5uC4jmDdOPxvaAnV1mymKw+ADjqXFOa6F5y7bqd5zC0B7sPiPPM3QNnQ84AulR
Gmj4nwkcBE0yX2j0T1vVkyi1q9nMdTKD0bmH/xunWrinPCR4OYjFWecdNuhYJWEd
iDPZNxC/oie4E/s9xqhA6TLek3LwYC+HxA1ZtkNha8NIgY7PXJWkImsf/qP+ZURK
KNPr2o8aOn7ky3Pm6w5XfJ43xWmyHuflk61PZM3caKsOiGhE6V1xLq6nSfBofhDz
FFX7OQ1KxGAlAKx3SVXgNpE15aTzMvABNGi+nazZspn2CuFXwtX5yQCEgtBkrlkM
zlIOpp8UpbUj/fHhBWnw1ojY4u3EZdrj6tRmpDcFB/2/Y7KaaauZr57Fjaz6TDjW
4jD4VzV73ajMYNgIxWLfr8MWGzFnTXC6wweDFjLKoCOhT44wWvZGIK8sit6WSWSO
bc8pXnCHRI+QQ/SzhX+KFnPJWtRDy7TEzlLMT01ZsHdU6bTPhvgLn5ZwBoMNN9ce
q7FvprGxj9bj+83B4gnVeEImCb7JTH94CpXqsjFTas7Tf/XP3VmnB2LyNA5q2S9y
lQHm9Rsq9J3IEsvKo/v1uDjyeMG8tgNQ0DoF9g3KrPUD4xBY2bED2IwVdW81bElI
HYxhzEMA+BrasVRRlFuevFwe2AxbHLI2ANQh+wHPMY9A6MWvD7gAHerqQOEmpIr0
vx7qQvYhSsCHIqyhS/sNqxKzZoNJqLbKCLs51UeN+PedlnzTXs/WWXMxyoPwFhXH
X7XRAcGznttTDcUYWSWQGVIqDnaDm/evJM+neT1LhBZrrmXrFvfM4pD842pbCV0P
trQP/G2WogWqXBvBBIUTWAIrptcT776JgPJH2lJR6PUNd69Yp8xnArJ2Zdb9ytab
3pNWqmiSaXdbfA9WYpQ06Kjc0E6efg9fa2bPLCSoPX1BdcVGxkD3RmrIXXMDcZDl
L39aPSJJZJxmB2QJ2o65T/V7Lo0SnGSJ765GboyK/+UTrHg4qJnDAcXQCcP2vbRN
ziV+JcgHtGPPSz0eDX4kuCSX1IUBCX6MpFjkWGFKZ+yh0zM5fK4Dxne9WQUsAomS
hTU2ol63HGVYvByXqfHivyRmyaK2Sx4Be1w0RuzlxjgFJJXeMcje92U1QGN4oedc
e1dRaLErUAK4grVUdhMABSzR0C78KNpujJZlq5on9n9BusgGLVu/cPoAn6KbEAmA
g+V0clMlLXHkvBcQeCDiVv8RFZhNdX8zaalxW1JHp8PljAklWdi4TmwLXOg+UFfP
pdFc8rETkI9AXPv5DhdiR/daTP4QkrtB11dnnGoPAfMR7SEy1ng4nNbRsuX9OodJ
4gCv2V1sE03aaUubvdETgEt2nrTPVrx8+h759Xb+Y7rJMMRIoepaJBQFH/qXPJYC
SdY18dmaH/QkG0e7FYKjsw0JQPdH657h5oBjB9gs3Ugi+RfU3mNmwTXa8HbGCIIb
5KqpIXokR857P1gOgzrpl8mZffZ72pbNkEvU3TZj6eANKEzD+0xAyK0yBeccu4pX
HGLtXz6Kj2fIpA0tXoAr48gnX3kWVIUSsfn/g8/C+pBHqh1gH3yOlv4hbfn6vWIp
UCFsYHdbEaWxUMWMOT24sJASj15IDBu4zUMu+F9/NvhouhbmWJakURF9dLW/a2qz
B+dtZsU5h/IIzV66yi4Y9P2JsgtGRAoxl0XqFtVtTBRECeQWtzOserbn/VOS30ug
ObOhxJUm6PThnefrXLMIVdC5f5VQlHkHEJ2rMEFgDnT4s6q9vZzF5JN+NZN1zFp0
19N4jHj3dwfwxwMmyib8Yn58G91PX0MnhGrl/1NehIzlaWL/lGa62ztM8iWgbshq
DmROgxDc42+E1kse3LLRGFMPfcNSDeYQ94ALLE++T/boHIIhhWkfSBgMz38JMyF1
vOq6Re9AOlfxhruKUt2yqZ+5vtvqMe3fL2VthlCgL7OO88hdxmoiLHPhLDCio5DS
MXI6rhrs1X0io292zbT8d5e26s/OF+2X5Kqx/ovRx1wHRK7ZSoLof8XGYLoldKQb
RZpX99G1opgIUdEo4L6ftLsQupw9d3Dh5iSmI3Amw1GC6gOJOgdu8qRutL701V1s
L455riNBeONS143fJ/xJAxCM8ORIEDu0Pj3ddQvnLpgdkJPNtiCQjdX0SjizrZsn
Q16S3Mn9j8XPChj3kMPFe7LcmZmnQW3idi/AhehSePlpW7DvvWdi73ulCQH4rGWt
2SlHFawu4/dYZg8ySqiN4/XbPjfA808Eu8IMfn94QsS1mysjbeG99pk3s9++1UXV
rdwfXJb/QYQX3PkCKYR07AbZmQSJ8Yx8pZgfe7cMToGfUBw4pYh5bOd21sg/wsMl
lug5cI1Hry/dLUVqQiYNQrFIO2V0WaEYb6ibRnoNGysiASyboh/I+Y4CiiBbnPKD
z8jnhsKJXzmr7sP5ptEBXQeLaTse6gKX/cG/OFEAMStHi/HC3cpZtXRkkEI8s+hf
YKoifrgiy6j6LKvA1gqcNeu43Zuz3B08Dj+LJdQP+mWcvMtmuwjwF9Lb29e7ONF0
DsIShj3LA7kcwH5VveSM6JC0nYOZP9LvpTsShViv+l9PJbCxH/P8+zUpo8FkAwnf
3oQTte0nxAgXIagbOMyE7IW+lG4KWC+hfNXKOJ/pZTdAA4gC+LUf/+9Lg6i93Thv
qRfoJW6D2sJqiHq+/Gasba+xBFguoymuF3k5gmTKe9uB1XcKPKkGxvn8Bl2wM/Rj
dHUw9VNhn9W+Me6MAj2TqAKddkRRRVDatmjdWqQFVkZ2Cudp5Mm6lpBhnPhWF+TS
uAOq75qvC/ElfczQKoIscKiX+06fVL7I7JASMGF5bRN2+ivJR7oIlTwfpMI6JMwA
7IeAgwq9ReCcP0orhmfZ2hlH8qM6P9YTvoDu63yhgasVSiRky5vx+1P8H/spAbxB
MuP4I0c6TipRhsBuZSrBdEhoPxL+RaJ3ILFQJO6uQnZV6wlVeukniqVUOQhgCMxJ
fEmr3S4Ym1uKryOC0wW8ag6IVgph/PAocUWbm7QZg9JocQBkp9T6MJAdJ4obBwnc
p2mcU0FK7IKCWuBskWni2vVZE/lO0+AI1O6BMDT9unPwn8BWj1sgANa7/hASxE+0
hq+MsP2neMVN8Gc1vfS4EnzNyppNhRGm7ACW775ZHllG+BquRKsvJYiByL0KylK9
Ssxg+PWpZKiRqCEj+30OUE/kPp9tvmm8KBJywC1ar1TeqnVEkj6L8cZZqTFw72nG
KOr80ACvDhvfI7cJrMn0CRXZZPqZj9snE37tMGhzxnwfQG9XGPwYMSosqvk6WR6s
7FrLhffim88hsUzPSjBhlnT0w4J7hycnZY4P3XRtXG6q2K6VmzX39ctdTfX25nPL
kRjejjRtUZFuiXTKYMUpM7HTXvIDvJxdM9P5boCWvZTfDx9QQyWxEWFiOjjbkj+C
oup6fFer4/l8ng8doJ3en2lApWZQ/76iBSKY9puSOWVIf2dpwKGfS134JkCF622d
lqb7Yoyo1ZT+Ztr5XCXL0hnxAqVVceTPGAsO0SJ3ja4J/GjODrMplT2oc2K3cjqJ
Yuh1sTDGHQ//9tlIIqvKQI0CHi1OjrdgWtyMQl3X2Aileq9JfI/pCK2Hbqi6XQhg
MLXNz24WCP2KnBwORVk81oHaD5xZomifXpXXm8i0XfrezF9V40aYdAjs1Lo1GIpx
EQvKas30YQ9KCSd4HmRm5wXoEKD7MhtdbazsgtrhMI2J6cw4eR/lrSYqzK1+a8DK
O0hEtR+Pf7x43S18XDRRprIbkDbJdeIJtqXloD40gvvI84KYiKCeccwt4Yu/3JiR
nvTTRkKAddpNJkJK2weV7DQgn3QM6VthghrgWhA4Xu0/MUotBat+qTV0ITEoRBts
MpT4pmtnbGZ9YrQf2EbRPBbfwfVB5SoKDHvNfNhydFMzFRFQr4mpc/nh44ECrGjd
suCqWU9BzuXQa+Q3hYohj298h59Rr8lbsvVwijlbrpO1NsYwQ8KnocX5wwvMYbTL
ibhzDGkHQQersOxmbEB9wF9DXQsZnGRB4LJvoNukKr29qCjZ1ydXFB1m2foBsUri
cnirbooervuluSv9HZ9Bhk56dRFKNvdjeVLfO6+lWSvJDUF5o0TTuW8zsdQkqN3M
NU5OaURcYP8kzx674TQQalrYqYDCUywnAwAjjdWf1ZbK102yTbtOd6OoIiYTu6Ha
s+Aowm/nabtTLiMkrV5N2Q4XiBdBexSB1BvBJS12RdbZrlb6XqDoZyXXVsp2VKfP
GI6SujMjatL3PkIvtSsoRpc8/WBpFs7cAfCxmIrQGyha5IqKkxMp5NYc29jhtAsv
T9+44XT2TlrZYtr+UB/ITPQOXkbhk+VIAgDu5Th5+7ozdr5SjndkKZ/BdIXgppNW
XP1A9VcV3v6ECAq9C801eT7qucjBDlgIG17TUC3X42T89YE6JOgreG+vxFoL+Hrf
8qhlBzKt0DWaRskT4DwRVYOJRs/vI6Oi/qrSP6EnNaNH+KWY/1jIXhglTACCKDQz
hFErC0GvUqxIoTkliTAroboxrQ8V8tG3rysjtp7I1zSg7XKjYng7ACD8zomYH7/R
FPn8WqruiaO8Z4h5IUJRqjhklOyHH3ed4bljNs4k5vMM5eSSWJQYJrEyLcrY2bf7
h4aG/TYeIUfxSzDFf8BGyET02R7THgyJTr4gpbI/F0n7/A2AGU3uGyl8J/cxte4n
PANvNbjytm7EJVEX0IQ0yFwyeIZBDFEKqwdBZwwTJKmKrO21hYUHqD0CbcGScSo2
peyxiUIixcUFGKwWb7ATkp1UIGqHvaOMukBzbAl7W/OeJHw3IaKwcL+sXfgATwqR
PujMVqYqiY8VXkDaYeWqv1dDeFtwvhfElHOtPgHC2DiCOR1TmwCM/ufzEBuffMNz
yqZQY0IjP4lr4VlktqznDAPodZGuueUMqZ+2UUvkD0LvegfmdZXyFixhja8kOHg9
+I6KSRMrps8a4yVjTu1n6YenDYDyoAbvGNds/FBl2OPQRDWxSNh6VpRf/aWPk+kL
PJWEMvqr4FsMJsUM/RO041kJcQq27LnyXB/YqRSHAJiew9ymIujz9CyaRFUjS7io
tjvRSatTfi8Vuyfuu0mVjTKLpEcuhSRGRHHPkP6M7PV5f5oZ6sEgLqSDO7rlgdxf
v2MTSp/UvfO+tmJow5O+CVNTGEs99T6GHNrsVPIMiTM2qPCnNK0uSVpPWMEKebyl
+0AK2Hm8t6R5K7s/RAL4O7q3E2yJc+S9ToKPgYiqCQR+0+TURQwMWsVKw3oeaUV8
cAexmDDWbQ++W64KqKeWU14XCkAli2DEEfOsf70GbpfPzsXPgNiIq3qlTw1Kf2GG
iHkR2ezLdvT5jiH+5A8pNBp91wwT1VLcjEW7OsfubRH5ivRpbFTor5bSDYpiDhX0
WoHp/woAyItXL5rntPKXDKhNu6U3x2a/LA7eGxtqAFbLwWmjSjlquvQt3om0Sc1K
spzi+1MIqUG206LJNo3t9IbDvn3+/chtURdyeiqAW3yBwGbo9rMii07iKFCIIvSO
5AaRGf/CQNDMzIDgkWKk3ZEeHZhKtuUJvBwhFxbIixLLXr75qI1erq02ItPjHZ0i
iOihm4+7tVOnrzNlUgDAe+dflw5U/30YIDeiOrUPaJfuv6GZ3pJm6nNIjBBMLbsT
cc4NyaIwTFrarv0Tn6129G0vkVV3Lb4y2F7PlPnE30cIrto0QFLEFiMtp8dH82wm
nFnFYu60Qi1eFxajbwWjFZVRCjVJqlmOC2k8uPk3V9aEs0ZqzRos6J8AA7kxdBRI
dMfksn52mljbb1cWV8McIydnHfTZhCkQc8+2QiDXI8qBKLn34t6+uzbQ4ZoNInu2
4fnuf7m7b13IR/RqsgAedNWffmO004sEJYAE6tXQa/DIqaM+MBMTfUuHMqDp1Pho
AF1YGmuQlCzljORGc2WpDwVBkRHEL13XanA7L9yQpFPWbgFWhKNRS/ggKiaDhJ7a
dy9IAaB+AHJjs0/aYKX79SD8pIYlCTtjMT3gGJejQ5BtysYnJgi4O9Xto9nILXuV
zCNqsXsuqTQKeYGn/mFjAa0vpEPNMK6k4MOo8Q5cZ5UkdeNGz4tHP+P/rqiZyb4c
KEigpPwXPMVAkeK3jCqVr0KB0fCRe6eYQHEBhNO3pLb+osTDgkNc4RYJ+loNnBpP
ic2sVYwjD+8a+ng7CilRrskALv03iupSP2M6QRwCibqP+OdHK/EzMJ9cxOBhaCeL
YNcYthbKgh0rDjdfi7YlNB8dH310+ipkSeAuYu+Me/yla8izQzVyUdiJekJN4rvV
Btl6qmS0PMJ8Srv5SrKQcU7rGLUGiowhGNWKXxaixhRmRiiUvsZmx8LGpFCHVp6s
bhKLekXg+/9SjZgKqflu21DF7An7P6tTLD4Vytkj2m/YoI/nOfyqA63H4yQU9J44
Z6AEzjVX/8WCTogwksmZ69arRuD6JXyq1hY0a2INTPsepgpwW9Gx9ApIEXgoFaqq
KmuSZ03pkxXhArV+sfr5Mp9aJUdExiJ6rcWO71Aht47CY1z8ZdpAjSbKBfhq8uKl
k3bfxjJ5z9Oz2Pmm86F+fGJeVa8lwyJFSjiUI2Bo4+XCUlfF7W9fFCurqrw7x79/
N6qJCnhJTIrGMZhqiWylnDS4CK5W/0ZxhSVFX0sMMJxtySMZTkISti+TC5krGy15
aZIw/lPd6MuHrOEXv18+SGcXRlDyZKiJ9pgp+pXbm84bxiOb9YbJ3p58vlcpQffM
qh30Lb8Kl0KqXLiwN4FwQl3UdmeeiInjcJIO3SyAVolM9W9yvp2iAYg6k6zsi6cy
TUTd9TKwUdF+N/QnqugcP4nzWTeaoBqsCBeYEuQDGAi+1jEgNYzN/ZO9V2ZbQ0vM
XPaGf8w2AEip3Q8+QXKKbSZxIn1tksrLdlK/Lx3J5fU6RZSWwWIh5sshKKD+XORM
OUO46Mi9eGAN0hVj68UQ+8V1GuszdxvoksHL2J7uB1QlaJQG+gymLMiUI5i5pGRS
Xw0pZQ3u1qZoGGSKIZLGcHskSXqSKT+puyoHLU4gA5J7I62ns7rOoQVUO+iqSNjU
ZoRZMZ8bL/ctfPc1DJUtIF7GbvKddyqQugql+fE88Ij3ydnSuXNlNXUSWlOWaDLL
UfYJJPrT51O6T7MxoL+fzUGXH/GgTufiyhYq7sdmFY6nqa9l2bQ8gc+f9+YVfwqq
YRvRaI5Dpr8m6aLXzRHthRrSnkgJ4In8swdiupJLKXHS9HHI5h/d2PJdRb0SA71O
0LXE1g+Yarh3WtP9IzaFGw6u8+KvFlbQu8M7+ycIM+lZB3n91NZ/rwCXRZkd+KQz
PCmhkyilrlTPVEI32k9bRcGAI+F7sn9Rrv/irkSyKDbUNt9zJtl4dXdL3n8FjKCK
gsq6j8CH5Uy/9wflBkv2pEruCUtFkHM2SbJlBcaAzqA7Urepe+Y59cllwBt/jWwS
65ekT/+ec02ilv8RyQGT0+bbXRg0pq8NNPYyrbYQcvEHKUUk07unC0u1CNQ03qW7
SFeUTOK/9QuUMo/N4tcFYjR5Edb6I66zmPLjWu28RHcgeJaybHGhKe9kM2AjRrZ2
5MWY1OlyeGjkeSgt7/d1HYlISw0FQVRhiuqhRK8/Ai081SytRonU0/dnfuHBEdiN
xxdP9tAp5X271xFxvK0zTbtRB1Bfh6e6Xlt0lBDUeJvki5uBIjGgkomGcWVf7qLG
RZXM9SUcpOywnNjJUPFBftwGXmszfe0rDE6PNIaKwuaC7wTrHdRZ4LGyHNao4Euz
Gaz5ssDTRmstyMzJy0sXej9vN18EmeLxYZbu0+4UqK/TBQyMcg+nn4kq/ROXYVYp
9DnfTaMhZBOLFcP7JhUOmBsrLd8liQQmw9Qv+loEl8ZoEpZzeSmSGwp6Ev5ojcLH
gIFrfaVqbyk1HWrFIBI5Zj8nHpgczTqGzF6yK0Ioc4LnnAJS3kWy+iTkBq/nIu8l
eeWDnS/iN3WlogfTVVHNOF45dk8nRyxZ7io4HFcMfY9OaznnNiz28JKBJaOpY40M
lx4+MwPqJTscGen0sebZrrqvj7UlOjGc3iicT63CurzhkSqi30ClaPCJm5qIdiBj
Bj/ldIrYdjDSUUZac1C8CJhShDnLytne1fCwV1HQWi9fDBZxh1Bq6rE27GPk213d
dWYFg3k9hGIby6SQOyxeL0VUmTT18lrHT6oYpsin+VN4es121VIy2JwSCHk1uKF2
1hqvpsteSvDvbnD2DdtWraz65t3k3w+qmvzhMAa9rfSiOywTv8YQeePOZncvs7Q0
DuztPgcd7VdxwD6DS4sL/pNo1N4wtomjAidrJSll8dK1DsUnZHr2d0T3c7ScV2lo
wwnrBp3nLgweGqMtb8NU1+rvNLbjv4DZGwINeP2axihVAcrpXwcU87p/7SaTkOlZ
TYFZBtXCKhLWhYTAbKSQXTJJ3NNBh+DiCgcrhQJOatHib6bNmHJ4xsdpYoczZSdA
9PtdCgOUjehl7BtjWChSMfUD5laWk18ByW1EIzHDDQX7Flu4ZMP72HcOZ0wdz0ml
N/orxvxcr2cu2QFKtPg5wur1kN8CUzdRgsRPh18jzcXfa5tEjvMwhgF9cgGhLkzu
8pEofTmxvI+sbiIpq/uaBaBf+PAu/FzntozEaiyGEcwx0YTx+3JKe7TnVdeQFVcw
qw5zU6L1CtPV4mtlIGLfDVH3n1C3dcedzgpBi1HBB3+zXPIvAL5I0QOIpp2M3tLQ
wRx82LkByvt73d42GMdCNaNwbSA04h2g9OVWwmmdbVJJxh0CC+Nb4R88vT70+xOk
eRbuOF/SBQzeonpVgdRGXKrvwK4Gya0lNxVQl5TJpi4U/TpEnxeoKlb7Er79SiQv
Gm+pJ0UxqIS89gGBsn+ArlqEKVEMrCE7seAdaAV2pAV/d4KnWSwejURT05byaPdB
3yDDKh9At7s/lGQhdRVyTg6chPvEGksOGRAzZG4jwgcjeGacfUXGOb+otQ37sfV2
qHxylvi8n3nH5sdHPS8MLRCzWgi4SqVZEP8ilaAZNdcWbHrYu1YHxTJCupYxnMde
mCmYYdcaQDgW6SWJNTNmshJG2SKyMcV7hPRG0XNnaVVAzCyNqYrESts4Fpt32cfN
ObnSYSD38oEZBGQdJe9R05oaQmxqCH/5hUvdLPYvULyAul+aOjoGYn9r1y0Xi+9B
acMWEQMbbZBfEkavsml96m/AMVznpMt2hdWhBlI+OXMW27Nbjji2N1ZkV4RhqZNh
IPdroTfIU7/0Lr9epcdYH0/UWmhZhkBr1LYzPbot59GaRC3xO2CTsM+ZLW5YX2g+
+DkxBiWS7CY5XKb0Hh7H3znOnZb1tSs3nkmGqlcu81oRrUtYqZNjmG2osrZLXLu/
NgpjN3alOhaZn5lHkl/o1csqp1LbPAoOm5ZSd59zsyeCwykIf6qU6eHWeyoxrflO
9Lu+zlHZn7TmOnw0VCdjB1XnFHYRcMYULqimPDDiCOroF77QmbNBdm5yqee9lzXU
s3yZ6wK0f19cYVif9NJ7SZuTd6AB72f6k+HzSRT9K0w602fpZ2UkTkcxQm2rH0GP
2sA2RyCjA5RPa3sUgMAJgj5fDQ0dWZzjaAch0v9gBxyPTn+IJP+gpDO7K9ZCsa6C
s48uT1HFL2b+K0Gop2j3kKTsq2uiPivQkNQy9oLvwHIhVOYBiCcT3Id/gcrab4cF
oi6PfF0vQ02F4r1wowseR5FGyzJPMTmIsz3kDpXja3H9HiuyQfkrOi7nCud5wEfh
76hbTZHBNnIfI2AAbSE3qkEHnECsPk7ajs763O8+Isr/8VLdKQAf48WApj0puoqf
WUe2+yM8EyBg2RRMFxkQArDmDEbK2c43tUy/EsFPNyMKUOWfEb0Gg8YS/FokX8eX
1NOQrcmKe3efw0osPfZA3ZrEO/uR/ZLeTzLCvHRwNRRtmS1ibUuzfsM65dV5kAWF
emiIGjTY6D5p6t5VVBMpeY6ppP6EvcUunh566ycCHLBHkNNFljI+xsJzLWZO15wk
0WI6Nf0RSQfqqNyWRSUPkHEyE7ZkFZkvr8/v4czzYPSbBybAfRhMltivcyzGnZIB
BqCgki9N1yl5SPNpIGRuVmvxTVdFDjAlpG/LRtVnhmDFvPlz1C+E7qCHohwdLjQd
gUbCXC5jq9UFKJD+yz3yDtZE3Mlv4duvCD4xLhUpVOYvGJvImv6L0CTjfLGSpENh
aDZr6wJ+xhODpCFl9Rc7NF8OHj7ztaXby4GQFDCXB9f+z4WI+SwPllFiiMlszJfQ
WqHoSHyEPaZlsPeCK3wfRaaHwEI60dGWnh/QnODejKWF9tyKkl8jRlLkQu2SJ2rQ
2ZrZCQPHi+hSnvolEaYt6blt3rBIXx/AYfEZ7E3Bn7/0It1mdaem9EdhWaW0Kygc
KoU/3yAdkm/02cjuj7BS/zoJeIBkkH/GechHpalxGA+NzzlPijV+tWteG2zPVPNU
Jdrp3vaNSCK7DuevTAlmuwa9Or1Hj2IZU39eS8EBXRlluTGNSlZdVO3gLEFWKjsm
P9dAhKyXCu1A+2k7O6bNy1u2dXOX7OYRxZvc4oe6B/JzwWcvi5zgG+sRwIRWZGTn
67fKDQG0LrWU5tA2TA6VgSkjFqTymOpRTdiS3sPsKLZ0fjNRCJytDL/2jJcBAt/s
UlJ8tjxHQc9X5vL6zW8Qp2qAKY/cxuf1lfOiNbPLICFtHGtbUIWqaT/ciAa/CZV+
zyXFhYaiWNx8PIKouU+o5Wlqx3ptGGUo5rhw9tqcmSMgLIxtkUvEF2rLKim0BjDx
nRyqUUOY5OFv6N/gsPnfA4weIpPXccRS74OU6QTVKs8Fs6K8FLVmpyG3DLQDZj+s
pNUwtkwAajKUFKHU+Cc7SlxmSlunK+jcqosyaOMeDi6keIyIhLjwLFxV7QGPEwcY
fK15/OQ/ep3LQlAlLqNXicnFLZ4V1Fa8xLn5AJYFKz/xYndTHa9zN4Nu5HJBdYTP
POMd/h6EDg6IZLUcdq08t963JKF59728hXThTKYRV0xiPgXsy/uhTwo3pECTzy0r
1qYtC6mkodFCRR4ixLWBllvuzZMOJEKavIwcevlZnyCd+XXN66r9cqIZIvJMmTxM
M3vQsS/qSFXWChycMvyu6WdXlhuxMl56GoRhTLx5KocKFDo46B8ZhYqlp54pwLqO
UfyRx2Pbs8Jra+RWs6tNOHgJAnRBuWaKTzbwAldzwmzYgZ6jkk5iOTHztQpqQgSB
LhGm4PxEubjZCZ/oQ44KOmNMndpbjN6vSYOUkOa0DekOH6BQQVjSyRP2Qv+NrvFC
3dGqWfi0/EfqVGVctMn8bkmv3VZjMTmIR7GEI3rnkUi89E4wdJ8DMn5lE2W31su8
X8ydguEA6Fd62r5ZaUk5FmO5TpkEk/AqQTdqNdWg34A5GTh/V2x2MDvqt5hF6T0x
F5y4Coqc/omzOL601QfMrpe3mdlIsdgKVbj+KGFEtdq82jXX604LdMMgdZjigoTV
mN4ycQvmmfX0aN2wWFvGKBk77C70jUIR9OqHxK+ZZUB1UxhJEt/kalTdD7gjTICD
eEhMoVXj7wN2urUcSAKtJdvmoxEituxWXhYpLwLgjNlW39VQSLNApGz7fyxYugOn
GubTTPFXLgxf08eFmIf4E+jozCnGwS9sYP7uNmnHARBWRdxrcG3aMl/AJ4d8/iOL
toRufZBWZNS8DZ8XahV8Z1U/nvB+IIxtR7Ei539c44EFFG+gRefzBsN15qmBXzdE
zYEouL/QYfIrgLtONbB/Yh4pGH8pcHoSfMFwIt2h8OiRM6EmbBUA67GyqG8QAc3m
phtk32gMZ86irJX49Skx6d9F0YsDfnKQ+/mQLruGdmhowNT6RWudt/OWDCfR8uk6
jpJ8hDvK5nkTPzhg1GLER//iHM9TWa1dCZ6Ew6Y55ZeoTcUq6vn2eNwLz4/t/dRt
JoksRyv7Bhh/qczaJUUWq5LX/X9aE8gGmpnjRbB74ubTj0PFJH+z0zihqwS8O4sV
Mc5ocrR8neVMp8eeGoV2SwbUn16mjVnb6GG8JrcXpfdkiHt2+C6A4eqph+69e4Xc
CvzbBgTese3oC/nY+rcx5B4hQegk9BIgwVq2NWIh2i8dev2+M8l84KpCGW3yYVgo
NuS1JCb7IZsb2R3dbPEmKXqg5LFSX51IzsodTay7I4QZcxpiAP7vCCD7eC5lp1NT
dcIbgZ6t2Yncn/moihAVt2M1uB/HnjcHVy/mQCKMqw6tYueqhgncDiDmx53Zi8Tx
q3t+cp/m4lpUu3EYZ6AIyNYnvyfP9N3Zh0iAcVE3H6L87+4ETFxBpuIWS+W0ko8Q
RxuothmGqcWGnR7iYw3sKBP3Tn51YiXQHOvXqkvzZy1D2K8+nIGx08YU/9dbKREC
o5hYEV6wmqm4cPVNee3AN6lLUu8q2gd3Qkt9PWKh1HfCjjv4xDeJA5R16wb6fLlz
zRqzrefd9iGL4DuGzm4my2IKVXFmK1BK4MK7zg7O6rISZ/OcvTqd7T+0925nB7fh
Km5ZqLSfCim2jt7lx3c5A6TUcOnez+ueAzO4HrwKwXLKHIBs/R1YaQbevh2qtAuy
3qXol2b02Vc0lCaa2VSoywB2Ez3/PWjJI8h9TMEllhqn2rPTgMLE0gSGShxRZXvn
LdB64OfAwnv3Km1Ft605tSuvQl5gaf9RZR3n1g6W91YkzNdyPu2jGztWjYxAOaQQ
XZdAsmd0IyqtbSH14dq38s0uiIT/GlaZU8xmeqcthoH2z+9K1siE7NIN5skLc6fU
jOGoc7BXk+/ZY7v/szxrGLyuoihm1Y5u9T44XACN7jywWzBc4GDAd+AVkimzhFvQ
V5L+Dv8nWM++GGUVZil1sNQqMAs4DqaLcOM1b3o2O2dvMWFOYe5p2M6b2w5BKUof
8huJOCeHgiKVq13KRnbKPDXmQw2wGRedVv487ZU+9HgyiJzEpuoivRxomgV6691P
ING+dk//CjKodpKQhjLtzXFNi6h1yC5DXejlEYLEeZ3S3v5sTzxFvJQUcMnz7KGT
yt4lp5V9hiVvq74uYXiTGugtoF71kZhMGqdgyG43ZM038kPUhhuAVUYJmp6Kqy/H
/i19Uprjet8wkMWibUV8/JmOUsVqwVmK+yoemDwyp5j/CEVKdMIi0qwRy6Py4/kM
+HFz++GQ4Q2EoLXWV+6RE8O4EdlthmU+YPuaJ/tzSHJDRhe2oPpqS6KNNmNjJW+g
e9J4OJp/0G+CM6mMdN/TSzwieB8/PN5QlKSQGlg9Y+cI0WEY5PJy3pDw7F/IFb/O
SPX8CJkNYpgIWnVZM/GEQJ3akBJag8tThTLNAwT45hcHGE/FIcwyNb8NJvXRzz4p
XEw581aPqj4AblopHBesu5dqgIAiI0hWr0E2B5HPDp2nUfOYySpjCDjcCpSTJ26x
+/maHSIh/HMss4NKZvGz23V3enXbvrm1/2fg4iTTOO08AlSlLZrq06rJF/aAqPW7
C9wRiKVxIfHclNz4NMvBldnpHfaH3MW5yn9KKQYVp3PQvJTgKZC8iWNcmMu0dzVD
Tkc/gM0KNsEdMNdbLG1yspyYfxc0HJ1XbxHt1Fbq56Ph+xbyYTojj/tFkg1PvA8+
VYsGm9B5Czt1F/NCHqZFWm0lQQFDGJVsY3lDhUDCTP9B7mmcj1ELrfRt/gdKUyqJ
vnED2kAH0pklJjfQNu0aLePt9k4USBNlwMZigtiq9d4DhM3PHIWnILPavi2dG9Lo
zFGDLmAwXsmuqKtIGw11YcZoDF1pX+HAmqvKfw4haATgozkiIOURuiUocck8Um+5
UiBsbMflqA8l5ML8S3LuEALdf3FVM8lnoLCgsdMtMi6G+u2GmTVT8BxC9Kz/Ji5M
o+bgOhf/JcjDnn+5N7S/mx7xSpdCpS97s4VTOv1TFnQXIJz8F4xzkFdPM4DbeRcL
gnFoXxW3BFFqI6F0Ei4dL/fc/bKSy53BY6sQsuMdoJIpHi1p8Rk55G0FVMOwlBSO
mlZd8d9RzrBPEImRxOkbXLCWoiTmUQNW2JTtshnMRAXjjpchmvNZR6D8Br/cDUh3
lEc19yzKUcl+AYYt/Jb6pNzH/j60CyGo/iuNdy/C/EG04S4hip2tToLchfL2x7ap
VIC48KLgUMeI2Rf25jyPrLDmXN6dvaKK6ZaX1GoHyO0rF9PsyGlYSe56YlnM/40S
t/iCyHXhWQeTabCcauseXbw924hpZ5YMHn55OkoqErm5VJDGYodz4HVus0z8s1Cy
j28CMlmJ4pWpAlh9ReYZCvTxW9aJknX6FPM6l/Alzr+wZunuZJiMxtDrISsG88UK
pTWjeR9zHT4cCQrF5DnyPgSYFOZJfkzueXqj7+jP8L96xib3Rj6TBqMeGgkZrpDf
cXIJ0xMd71ZNepA86IWYKLMjMJiv69/ZBnlk2TZ8hSJNmWwpZyAHrww+agaClWs0
I3WIiaOhS7adHISMRnXb50XLJ9IuyHA3cEA7CxrC2B1kka7HQsidzQMcAL5W8baC
byFOPuJ0Tb0UzAuRM2CLf/mOEjoZyYbHmBuXFfA314D4RQ02+1RkVMJzA/depdeY
H9v5e2Mfmwvio1AsL9Ug3exe3lQ/uX1zudIOr04b6UblU9UdRHR8CzoBsuy3SYRU
aj2zvLw5iQ1WY9Te/oST5wgElX2G8+vrjWhtxItiR+sG6Ksv7fkkE1mMYh6+j+Et
0jDNqGo2L1IvKr+y6uXLgu7IJ16FgLOl6MLIr/B5prIYUcqO4BDN40rTV0lbxD/Q
NcvlpAUK9xOZntLyL/av/vwhoZ5V7l2/OorMP87otmppiLuexLM5cV/9DEZfapQs
y1V9PKs4MXUR1m6vDACB8+7KK5TmtP28eAhDp2ujrpwhqsc1DMs7aUEF3st3vGxk
cQh2WD561M4k5xoPof3aah5dyUqmYvNVDELJO5FWmbu71JrCk2hPWdQXfMmLTU0u
mcTtn7eigGEgE1A55A/N/+xM1VZ4eES16U0mcxPc1nQwLD4/EToW1BQF0vGBU5ne
X9ZCEizAcKy4DHjKViCTGJ4pqX/0DL4FK6fZrT5lqCPk8Z6nAWY4R8GmPD6dP7zO
sOrBiBBvLGxAquku/lgppWfhpLxKn+Ad5/TnAb55FCCHq0hzDb4yBvb9WCi8GVso
eVIWZE7zwiOBDrwol975lOloZaYus2r8SPzBuDJKCGp91Of1mm+aCnKotaq1Smpy
DTHNMG9M8mQt1gdYfWdJWGXgk66YlPKiLkhANl64t3KPax3+nsC4bq+34v3z4LMj
7bfmd17DfLzaJrscQhpH7fTHeOEXCcrJAnJfIXLkTyVZUD/3HFwuiDFiA1WZIWwB
oxMVnWCuvgKtyKnVoeSOP6Y7ZVQApaUw7t6BgGy4vTT31a8HpvBtiCugTpsfeRr2
qgXo5BoxAvFu3Ztm3TO9gCU1GtN/ocmi1s38ayzXoD9DDkcvWSX9WRFHG1xfiO/q
puxP11F3KNs/VfivnE7TSccYWRT7aWgy6dqbIOY4/bEcP/7fDKHO2pNpTTyuw2cp
ksrombQy5+5xDP90fVUWwfULgp0EDxAVKCSKULLwEpZmae74n5Amm9K5hFSE2kvB
HukA/jCcUmtMgqkS6r9d73OEr8EqiQ7NjvYpW4YgODKnx3pHYZZst3MWrwVQIzWj
QKOlF/Jfq1ctlmVR2TonnMkfHTG0TcSgcM0jMYAPdPWCPMThe9gwSrHWPrWfq9oW
VfKsJg4jC48rk/chKbGSOfU+erM9bU1mkH2bC3w+ph0KviqMZA9Te6OXwK86p66z
OoWcRDW2y+BfVDDA0ZzGA84kI8rpSlQSMmHhk2aXZQ0xx7ipJFJV4N5GUxmctRpi
ndSybI8v/loJPSG8ib8wsDH9vCfXjfvz9cZZuO8vNHkN44sW/n2gmgnbReGbvkxZ
kFHxvf2l0q3SIREdiw3BFFxikjyaIUPJXzQdsJgBOifK6+gCFbelq8PPLRX/iWF8
+cCdKCpANVDohnycv9uWnoFICG8IH2rLNSVgPx1b93kdFY3TIVDHm1KiVQBKTkVz
MqJglXk8y56Y8QNY1s8Cr7v2HeoVDU+wDeifpDio8kq55jsl2GgTiw5fQymJF10h
76bHZcRET1AS2qszT4HbcIOZslqUAiUVq13Jv1KNy5UzhYDEVtVw0u6gyL+t5/n4
Ah1JME4QBfouX/xCJABRCCi2SZmw3E1tKlURh7DD4ZCNCHzv94+A95FTSEMazws2
X5ogrZ9wt6269XUZEiw1gCcIqjU5IP2obqQkhtvXwjnDSmYh9OGcSp1CTo2cxFcB
008/Q2Jnx9j/EsemJeNd7Qb5zrqkoe0Nro0xBqx9NTYjK5x06BC/yrFfn/Mv8yoz
vQCUshfBTnnJ1qEWdJ9y87gT3waS8fzcXmgZZFrpoc8iA3ha1hB0snhwGr0IhjwP
7vObhayXTZUWecq9FAWR2jr8ClnUzXNTIzzTOcZU6uYEb/1XbHqDWWj3EZAewxHF
8d6jaIBwMco9jEwLRKR0X8mUOtNs7g9fLjzc48gF9a27ukBXKAk8ClMWLnH8Y7T+
R9xK/+N6vWB4WgcmZxuc8ScQw+kzp7aan4bRe8Pm6mtkfkiMw+RydJCs5irLeprk
uD9BuROuNvlzC0CGHHLGErFMcpa7zfN80ipHrglnEre5vs0b8AjQzNq0WQRK3Xxz
8l3zgvwebolmBDH0Xu3htzF/LysaGurZ+3btRiOUxieDylznPi3zH7GK8doK8CiK
JF0A0DHsd8aaD7A9teW9H+w1iF3hFzo2Wbpt/ycjALQyopEu3vpgHbbYipbvIlC3
MC+tSanOdXDZv0xig6hvLUc9pZ0BBNs9AjSKj3RS7H50nwpaQdegHq8fxpDHXL7q
YZB4XR7rmANJSk0e1dW4Y3VHrm5GDkjl2AWX43A0LL60idCtYayGwDQD7B/Ksffs
iA3mPRVaIRDYFbm4+FYsu2xqA0lVHFNZvN3If0XZx5Uwl4hnw0l2893dA36mX+p/
u1UduXJdmWlmq8Fkm5dRiLf23Bo95lyWt5cK0zZDED2pMWCFJnpoFpUqCoztvvfe
fd3uquj4PPChS0N3dvgALaHD2kzjJ5a8Mc5PD+j0Q7OHCJMZEe0LTY6piy+MUBRU
LqrqWemB/2Y0PrRcbgfGG9nDHteo+FmG8+DvnIgLz9kJHOvZ8gG+X//7tTbsvMx8
nImC6jhJ0v1fTfEFHzMaIM2pGD0dppMxQ92exze7OkwhxE9ouUCUnO8hTpZO5Cif
YQ4edj1JEnl8BPwMZLJmFqzKMaPwrbSMznWgoeJZDc3ONlvWYDWRD1Na6F7ve7lP
QfY/bBiJ2YfiX5ggOsjc/Q7JcCJuN6HcB18YFhb7PPdqYEFq9jL6wMKeHv6/QUfK
yegJTGWZpA7TsyeicSuawQyc+fIXMcwB24A98S44X0CbuD6dn3OIIcjTGqBs0/A/
SggTWejLGxPvMs6+VA7wg8zCl+GSSMhYMvOnwVAJ8GvH6NWc+BtJYxBjjttaiwP5
oxlBEHL2UpIapVgvH1J0N+huOBRmd1B/CImqZNDy3OciCbDkzs6j63YnYZLsj4YI
M5aTi82ZzZcZYPIQ3e0FW0fWQEKKSK4mUWFX2p8oQRFMzqVkzDJ9lhKp1va4zABn
X6uGtzRuGh5KMMMFxs41XEyZmQ9TolDFdBk8+1YLCTNn5yIWvPYb79o/zTDueZmd
MDlNgGM261Vgd/n0kbWvAw036oCohE51albeHMUv6ftJtKjbnVR00gGa3D6F21Fv
mFEdtcXADopMEIe6FlGQ4RjHBmOCaQy/PbD3Gx02eak0Y0XdNB7SJtheB6KAR5ZC
UJjqkGpwdLtILju6U6yxtH62oFiHcLDoJzQ0AGefM13XXDOTFfiZDCKJ3fYnyK5j
7rCgmkBpaojpLLgjnShDqrsBrMkE4xyrDtuMbquJadKW0xjcJ+TrV8ZjSEtHCYD7
am6/KWpv+6ej/med6HB/Mae6QhXAEvnnoEm4eCxAeIXBby2xysbrTHLxlKfOpnGM
FcxYai4NFdwtGdgzmDnsRdHlASpr4rQ+ChA7xkOTDszi2Vsm7qnWKN05CD9lya6o
e2Q70o3Wgh5KpV8ZhWiAHcR0RfkfulfmuDbwXIYM/S77BkmAUScL052qIYOHNbcZ
t8YlYtffqqYQQxjNds66d4girx/6+Isb6AjWzhA8/rJGEscTUMxl2oSzH70y/Z21
nR1wt8KomWyLKdkAxcsk5E2EFg+pWM55476O7f4BDKpihphNaRT+4JjBs0bQpzIr
vVisuhwwIzVGao7VYKTBUrl8FhfLhQHMYmcnyk4khvifymr41Aa/FXSfDsM8pwPX
jXXwSR2amx8RN6HlEp2axapudIDeKbt3+ynss941mWDT9cfTl1ewOQlYxMFlWhQi
OFDk2ua7lxaOOYJwjM334o6ak0+M37lQlZ1bUyE0HLDLEaZAAGfxOKboAB98eKy0
oJRupjDF9L6lExYX6/MR1XCNqjFmdnTFblzXnKxczkncCzCVC5cg+6400f8Kbeu1
oHwFkS9fVkm+0pAdPbxCxB+9h1mafK/ERATs3fX16RZKAd98+EWdvZNShaGsB12c
1zLqB/pvZWjtrQZTM0bO5VVNaBK9pjWsL0EQVNTG2dsGJimYwXZyIj1afZV8DhK9
piW9LDsfqxShdC8AoBA8vd0iIqRT0uU1zpzSXBAcUGXL40/1MRT+gFa/BNO/rQ+9
8nKa8Gbdq4pp0BbUXFgGDPOSWkO+BuUx5Us/rCjsHj05LC30Z8XMa7ZC32IO3LCK
9Z2DJKCzr5pt0DPwOscfiWUVccamZuhFfcu2zNi9GZVe4562tdoi7biSxM7D+Nrs
5DXDRi372GUjjcO7ir8a8bjXwT/qxXxPqjmEYiHWVyUmITjrRAcRhqclreGa3U2R
8kzUro8Yr75CaFEruGoX/mxwo33zAEf4WqYE1Z3vyDWanbMa1cSWCqyVR8Sl2V2j
P1m9A4Qq0/8nud73UPX/jgD5NzgC4k8Gjm3VYa0Plu8Rsuj/ZSGhSKGVjo8T/0Af
Rac9vUxY0/vEylu2ys34kr6fAuCH0qusFYz59FToDaAFccWuDFjOhmUz9bMm5FgN
vFzFhGwS9lSdRXGrmQspJLJ/uVg8qTfP1npauQajT1yZ/+trbJZZEGwYHxuDRUZG
/1Ai25DTsM1Emxh2Hixv8fsB/OJuLfHtJP4yognNxrmiHvu2ymGrbn0xQcWHzOFn
EEKc+YvanxAYKSwCTb9sJnUrZxPFQ3mL+VUikF9P0sVz3OY2oj1CqhLjj4I577y0
giYL05uBpsm44GQatAkpRL5AZeG5Poi7w2AK061CcsRjuYRj3sCxzhKOLJ7kNMx4
Vl7BMGx/+Fd1SRcTFDOuKFWsScfRvx8OaM+rVbWT+Ohy8caCbKluQfjrJZDAprFo
J3eax2TtB6lqkrItvpGiTsY5EIV/+MhagUBh+/I5DgNIWfkVAREC4hvbYFpd/jML
KC/ttQ3tHGPUGSPhD2ub68CE9Sa9fBxjNrjhVJvEnXXJeULOEa7qD1mKU0XAt0VA
Gja0hnEPCXifbSkBCmfQyVwHixahvXuh+elM1/bQ8U0O7EZ5iNrXk7RzBLoqb/kQ
QGZ96Ze/l+CJwTmwZjyI2w6/4YBUL66RUinQNbFJ020bITZjP2CMJcRK9wV/EZEv
XG4saFP49V6awjdK3WHl5YQypYNy98XAwxd82x+iAPT1oDPZbf5QqqCWn2UDzuuU
Ll0pSEQEJHB0aLBudZTdOyddzWyEVUyOPmM0GULye5LVS7+jTee1WJSah7HIIDad
0WdZDh64/4vibKIjq/KSxbrOcHYlvranfj1G1WmkkgFBlOdxKGXsauMl8gq99LXX
RinGDJi46a2ni4j2lsIwRyVsAUQ0UtQ6iCrY6NaEIOyv3gnltcPRj5QdDFMgZhyH
qaT8ivjeGKK4T0RvxMB14FqDn6Vhdjqe0jx1Eh6w4t9h+z6lpw4MKh5JfgAk1UyV
Fyh2KfZqQ579ZedP9dh5+Ffqm5c87G7Mkj5PEiiv3770wCxZMR+nYNWh2nzbwzGk
9BqhPDP6KNEb3Wb06iCXsOeAkAD382WtJDXUI8HHHNd4KtpA1xWJk3bUH2SfhRak
PaV1iAOxskIaFZOgf9FNpQDIYmTcyey1AdnnQ1gGV0xCf9kfX1kRaHVmyi0dPJ9G
EVsyWj8IIZ7/8+WtfLpw6GsUQOoDIhAzYowad7me9FIrXrQVvx/SpI+JXmebFxEb
TSe2Rv+BE5K3zv98vrAWFXo+BUKHB/MtQDtP7d2IkryhOuyH86v+7hdpm0LEAQgs
+r9hNUB9ogV7QGAbJNa76rM8l7XjXPUcS88AKhBYb0WwqJFbOwY//+EGDiEZaMq7
a50OUrJPy0vXgNS+0Ue9WbyfDrVyC5SShxGx/pW2ovRgF7nPIuBPEWS6LziUxMTG
vv2P89SgBnqqsoZukA5GCzipebnR1ofIenn0LZVQV4e8VJxdFfZvy6tgmyf57qRz
hom5NvzWlqMDJbI/DhrupLI+IgijSiHRZkq/bDt9mVH/IcnSIeBfl1mYwPokIJqY
cSm3EYHCQkzOPUPSrSc/pyJW5uMRPjYzha6tTCu6OkRs19szJ4AVyUpsK7/bihQp
OX3JSNKHWixklKC99wJ4XeySAA6y/cFCz3Qd7ZCdXvs2r3E+CU7ZwSKDFxJ3xMEJ
OWat1a0r9j8lsELxVtOB0emmHee5AyqRn1wr6guxkVqD3fz4Bn60DX//BtXPCEDc
oNOk5vqFmrrYKmSJSHfrl09j4rfen7MTXpZykdjQYi49U8MuQUfj/xu1O9AF4OiX
kpkb+k3rGOvC6iGtsODK/Hu3y838V6/vTR5ZJ5wDMhy/q1bopx7dXGObpScOit/b
y+gC9Ei2GD8ehW9Q4Lzo4UZqLHJ6uqMYiTvuhgwbZp5qa0o31RsLLRZexy4AOhFC
KycGyKBEgyQ8nNKBN1qWwOC9KXDOmGcerWWC3/QP6RIqRZYK8etWnls3r73g5Qt5
YRcAOEIv84hThjBUZXjpPDUQHa1PQLz5axGotU2yB+vIjkt5Oy9OW0IJx5iZIMCA
JGHLnjRNZTlE5UbRRM6Q5AcaCIdGBg8IF0rXYTp39PPprKYWVZQRKho3FWcyN2t6
oBy880oc3EHp35ZaefUycAV4gDhOA5l4zeMIj8n/Mzgz0Pb1ahbdsUeAEIAVTQZ9
FcIl8elyI6N4jfC/QK9I02hZUneBblDUKPy9X5ZIpgjTXlEJhPyjmWbclb+z5rxN
03vPISv57Bgkq1dphtDOFP8JpV2vFcKghD/A3hD41t0SwXutlsTsspKP0XfS5HgX
kAtNVX00bylr6uyG/xY4xbpce8cRFb5Bn5RAF4mgi1VdPnrpF+XYYVfnbPPDUNKS
Ju/ZWYhnqCmN+EVRfvOUtExfZeLLMhbdg15xZjUNak0aLc1gI3ycLdxOB5XIag6s
A3W3xleSKQXOlObuQ2kStUGQ/4j4bxoZ0BTEEo6wREt5sQqtjbRh0aKlbxoyc2nW
N+2or9cbb2XXr4NR+7lp8kOAh9mzUEBa4+7Ez5FPHBXq/p0xFVnYlS+OswiqfBUx
FvNSD0WiD0j/LISIwkNpwIR00XhpcuEl7GqcQMwoJdNiiSwnlhB00YgThGNuVRmh
D43to3PLu81imR+4gkULVhGo6xM6jc+uMQlun4Y1lxuH9FxVBgIEmWZmYExIJNtr
X7IRgfLK9MqnO9IlfDs5lYmWlYei1jczDMpOlfMmQ6Gri4/YT9IxTJYtE++uE+MD
OuHrVlvy1A55MD3qfBfsbG84ak/uG6amMTAemd31ddYMePUaYKaW3KPdfiWhqOOH
hgQInk5diOzmuAFZi1cKwTPnyymNTYZ+Jo97+Oi6zUOTBRiGmyIncnk4sIFXtj0Y
5HvxE3jTayiPG3oQTewVc4pzvfowx1iZ29dIGViURwTER3W1V++wCpiyyHyy4TyP
tbpRThrsUljrJ9j9faoe6VfIhUXES1Ce2vy5De3XdO8FowWpej1VQS5laeY8ZrxC
AJpIx7vmJe4fLUhCPsSgaCAGbfWE5d5Qqm/qFdOmOI+AM1/MvodaY8m650sxREQ5
mqMRf4MKOIlH8I3xllrmC+vEwd2QCdVX5+QKhuxDYgCow89xTTWXYQkJr5IsPAII
7Q33HgB3MJXxCn8+szfduXl9w2xDD7Tqe2ZdXz7wnxBGryGARVCN2gopE2oLR+98
lzbzufju277OP5F/ngqdUJpX27TcfFB0G5Z736ARCyEcuUJNM0SosUAyK17F8psv
0R4zTmWK2vCzg5/mKJgRgMokcEdBzg/7OJYV4pYkCcbeWp079TZ4kySjUjgHOQT8
0frERy7rYoWvPGM8HRt11st/Z898U81r1zaFz46ZZqPXi3L+y8xZvRTZtzz56EIv
k3XltgHh36FNt3Z230JwQjlLVxrtJwzKNpvp8yKMFzQZPJPbac0lMoClJSXaI6Va
jnIP/wCBYiYoYm2Gtmd4GX2SWtc0LZwAmPQgKXsr3ng4/FmADLzEyCysjwiFplCR
VLC5RVeFYtw9gAXMlbK3UssGW3QHEaP9sStyM5A510gBBsDYFdvHZYqJKuwLe7P8
RHElLbn1Wy7xFMmRxvpbEZBNPatgUG833WX2cj7ACIO3XgO7gygJtJ79i6tKGmgy
kK93CAHMKcpy2lM6k997oWN8yvKEUk2ofDXB1Zx92YpfyRqLRsMUKNwgg7ABPyH0
YgGWYQ8w94dxaPtxs9zPC5awHyfNTH++vRDQYilp27GSgMpuwRLN4rsAGezs81Q7
LK+yML0EttpKOGp2EZIr/L9fp5ADqQOCpBBbVQrxwVQB30Ab90l3vDgH0PBpSeqy
904Vq0H4HuOU4QNr8AbpxO0B2KGN/NhkoxkK/9u+2PsPyoIiIQGCjtB05z4ZSClS
Iuss8MwadT9J+wbyWGuaa8/4dIYkTQIRRo92ij4oOZQYQcMqy4jP0EqZHGNQv9OG
g7Q96kqIXcERrwcUs9pgiLAFYPjX2mCFR1N7ZJqth3eaqyC7JVbI4PwZSYo7Me/9
2HeROgqcLo5D/Ionup8W7YnRJSXLG1z2/u9msb79AKCA+p2yyrEZZRwNdb23Lris
1YSV6KWBgAiXcT2b3FR7KibZ71IHNr0u8T3jbeP/F5Lr8bOLUcqZf/Yg4M5968Rb
Y0f5QtXfonintWXsU1NkDOPtc2uukDftbDxFPSivf/Q2t5IavhjbGYFu3gOO35h+
Lx3eSIOQkV/W37Q3gCmdTfK9WOyNg7qnQtVJTohzRVWZUBbXh/3N+e9B3Bj8GgLb
hkFAIfYsXusIZIS6O8yIiTRPAk1N/LEhkVXdFIRlx65OKIRSOwfvPgu4p+GwEIi3
iIBqbkSIRMLMmyeyXFLbhkYoUXG3yd0CJ3kt1GgKKjKvKzvsNqGk9/I+dOjm4mJM
sfQajeiLi73D+L7naqQwifVIVAXzpFVHbSGgx6RNMYk1PC24gxfUJurzuM3jGDY/
cMd/gVTPhRoOTJ06Er+5qH0/AV7++MNbq5ySowG53jg+mblKRWSs9k6hrE5LDO4i
ZWFj0ZgzS0YuVLsqMev1AUFTdQEMTHu+PgmunNQIH85gvkUKggwPV3/D5QK9Rw+U
/MB6xfsqJSmBVJKKpcPT7nuWaJnXoxgL3yLr+xX1I1fZANGxFH+MDXK63sh8nbHO
uFY5dp9nNB3rh03txVp17eenbKSznmQzKdTZbutIsafgbWNXmb2PXER2xqFjRWEa
ITrF86jhJxH9ddzoHVCAs3cR0wUH10ZSLPMXsuZmnmYyKWkgIs1cGLpsJTw322vX
iC2rob75H5LSoNLO1+EQuKwjnJs7UMNa9c94QmfJGZEKo7c36ItNQvVOOtUW//Tm
0aPhzNEPKjlypJCbENNjUbe83O9+1Dh+Cf4RYokBHbeWfzJefcig0eNLQbJSxYpa
Vt9E38/6ryBKvqMTDVhOwiDdJ7mslUaIvDBlvmPxSbWaWH4dkhXaho7mvMtW4p4L
aCaRSc0DgDxU1DFSs+Z13y7/M2RvEauGwpNxVUMY7VSK2p9WPmnlUoczSY+I/3eh
yZxgfMetEzR5O/d8R+h0n591EgtyKYpfJJrBbmL53bdoWdzctHe65HdsNjhbDs6p
yWPoBleZG6Gc/QtEWSNHxmrLPpZNrk+YykH5utHls+yJmQzqW64kCOa+ypwZSURp
3lhtWl/jcCVp7EL1fnVBiEdqGKn/WcGUb8FEon82SNSyudyKFd1poilRR9M6982a
Q+EcOD1HF8Rqh0etRpF5bY3eikFKBajHyn6HvhQUoadOdpbOIfx0XRKIGToif3Cs
yjB8drsIQLuMB7UgEXCXxs82c1FOQtKwZFDkaoXArePKEzJJ7haJ1v7eQ9tSn6hp
1+shi5PWiQ+/5c31NJIT86kvO1zm6Az7pifP+o7k5FYKsgMOqLsMGxXHU0+ikjwM
VlpY+BGzDlcC0Oi5uH7Bu7ftsHYtNNuEFEfK0xDs+5gRHGRS4MjL4hrTfgreSLjE
DxMnCdwme/U2JyLQfONptic+IjLosdXixtzcxA+bNAyQkmegofFQqwUxKj5wT2Hu
B8KiS/0DGdqbd/E9JKtpZPVi6zTyQZWvItsFP9outnsnFpbbs9VKikbVUCdS6siX
66iBD5e4XsnJ7Eh62rcK/M6uJO93pU30EvCBymDWHb5NiZ9Vh8duoSNb8BRpTN34
yI9l6OM24ls3eSX5wynPp17/LVv/eWgnndR1djdgiQgm+teAFvNi83ws11QnilJJ
xMZlDpydILlXqdrimqRmtQ+m3N9Xb0gNQoa3ByEO3siQtStkWV1vvA8gl4jvPDu+
PT+WCyGYze9iN4AMX5NBxgZERm+IAfGuTHmcNWmvkppG/eraa96+40reUqwflkS1
95niDyvvNHvs2+7d9Vl73xiaC/6rSmYdU1gka1Iz8NOJ6cVyjiWk5ru1gbDbK6wQ
0UT0z8etJv5y0bjKM+taiE+zcp4bwhGsjg53FZ2FKAGX67ZvdjgCG9w+s7e5B9C8
/evCuhWWjgQIGQx364skEWEQHZ7M0NFf0lF2yT7+SZSTrTWDItTsGdcttWVKtwPf
SeAR6Sr6HGTKL4S0uAVv7IUGjrIl1ij7lYCt5peF1N33M5pQGjqGPzbiKffs1mhI
efpSbiJpz6eC/tVDuYXHgWvBdApCQZEbgeSOC+7JdReDo0MkCFpu5AeLUmSH2ORu
uroVIzhVLjS6L4BvuLcF5Io/X0bQxGGgzpaBNJFUDyEdC1r3JZ31wsfQ8sai1wVd
iPFFNWimZtBJL9JfAvMfRj4Fg8r7t4w/3NwzP0SpHRZHk6MvPR9HmRe2DBNHht5t
wAh5G2Uk3ZrhP4s0Jw8oDY6TYbpXvoww1lZX1Ty7cPOlBlNPJktmvZofnKqOFTK+
Mzsjll7WmMYbXvy2bSC030T8BPXx5vzuP6g20CzDdguYu/M6wgOggP6hu0MjqkQl
ydPVeLtaLZ6s5dwkco9fK/9oh8zrA083MF8lm3/234gsvtrkc9pg7lhBqQhDo88J
aykKynkDAmKgEHSIBdAngDmbvlrzBbslYZkKuK+R+ynBcTnKIb723djhJyzKW4kC
DxbrQ8fOgyhNFCPueuvDOVKg60vidujI5bMwkf/Vr+i6u1n8hesfMZGnZbs7ZRLu
ncRdkoUE0K5QwZ0fqOQTn0Af3ynqX2nmF6VWqhnfLRzg8m7YVxAE/tQ4kc3PQvW+
FkU0xIYPTUcEYp8Cb0DWEY9w7MOH6mEO7Mczso5CCEzOA7/GnJ60DP+JXbxFS1YY
5N4YUkSqUTqt1TJB6Al6lUPmrxsxjJ6Yfrlg41sGni4Utls564ayqmrTpckGVCcX
ZwR2cOtKWNAiN0EuZXrcz4BGUsIFu3t9cGMzliesO4VioUAzpSK0DCOdvYz+n6il
eJ1YgaYTTbzWCJc2ML27mYbDI+DMFG2RjcBSrcI67TadMXMJeVlMlZIY+L6d3wte
HDdj9kj6QD7srcSrVHY6FziVLt8d0WvDLwydm45ZB0Z8mAC+/iEFv7pjKN0GZ6U6
mFoE9a4DOwuD4NLSu/iMwUUaItwJPSa/g0tg9fMhfim3p0GxUFtFuaRc4FZVCgbM
1oIoR5JkBMVz7kXGnv0K3j02NpuxV0+wjulAUwY1PggI98+Tvn8zZ8uLIKoKHH2w
sGw/13aoBB2txI0v0uyHM8ukHHO0HCYrbn61916HZUn/hOqflLdjtONofnC/pNz6
2Cy+DcZf+rosF7HRuTuQt60smMuYFsRcHv4ft5FGWKu2Rf54EqGHJ+8uB7O5+JkD
j5FzVyM6Qb6oepmrBIb3296SUccBA87HKuERGy6TtddZyL+j9Rg1Nhs841SoF+HS
R5ptDYQn3Yu56ol8ubrjbMuVaA2EAqfxDGx2An4F3Zco2udhch0KcCfHCXmXwNF7
2zdzhhd9x5fPPD7YEzgcJVGRYzmvZ7RMLFW/5zWydIePa+ihRH23+y/8R1UK/KIO
Jzg8nPvqhhQHWUl6usvstl+n/i5arTkBPptGo/pluALG8ktoctDjeER2hrf2Lo3N
N2Ag/no1DfS1I54jTj3bgkDtaYJzy1sPx7d6qI6W3ksZQwlYnQ778eeOc6vqPEVR
PtJ6d9AbIcaNJFTU0LPDRO7rAPA3SG/FrfQV0SspU+XfMdiZ69cEnIEi7gvibaAM
tC+3T0IV0aSTkkbDJq/6zVI/CUkoNqEzM/Xn99xuSybFG1DZ0vQvIGwqaE5HLbe5
0VYNadqqz+6My13JNjxccVSIk45DDVmm9s9jlS04pxpc//DWXJOCQtYyJrT7m1Ru
7cGcf1Nnn2Uavgx+CGk16QCrj9srJjVujukhrefaM3CAorS14cFi5hH49mi80Mok
xqS6dRY8FDQzLFOJZ2q53IqxaC62Gw8uwZslKeIrXBZKJRscKjkJv4LXVeeRWIXd
MKhydXaU/WFhRpI4knf9ARxJbSVHgSdvz6gijRve7Qaxhph/sPYBqj62Y9QNhwlR
vXp3GAHUGKq/BC2L+FysbfkiFWhtweHQfV1EWo420p0kKKuduRl93TPob6WsUmwh
0wvWP9zxV612gAIAclSySC8B1njC/8Lq6nb1hWjeSVMWLvNSBa75/AmkjXHnESVO
zQENf2CDIlqO71MKrzuDIi9oQ9kGeVRsZVWwBTkvTnTTwHzJnyRFPg+xpishIdYE
Et8hOGJhk+qQ7a6VPtTHfW6jFuvhw9GRPGUN/97Og/HGZrvLmDVmk45CODAN+yk8
uoi1/aCaH0NmfnyrC4VPbceT0954/5V5aeWUUACSAPOn1gBQeJJLSBO6cu2hVUuM
/cyPMLMYl9weLWByCEm3xNz1l5HzTOmLyRKdcYsTvjSyP8eX2meaqGY1jgOtgvGu
Vq64XjT9EJcLPoaXHXr3dcnA4uxWsFUZfCM/Z/bcX4LMv0EyjC/0eqYZja1UC3hr
xtLnFcK8X+AQWyFUHN9QzWws5hk0AdsxfmC/OxXyiX7oqNcE9UO2v8lh2s4Kcega
jb8nSj9kz+bitKf16yvqdxQx2FDiTMoN/P3K+q4rGiHui8vePhv71g7mFxw+RdSj
YZ624Xi1+lihpwsvvPoNTlqm4wQ0uk56Y6IzcWSYxp5AG8ByiGKMD+n4fKTv7N9j
lxO3v+MaNaPpyft0rnTM7j6glOUpvWwI1eqbrn7Mjs2c+BarK0p9bAxcfIUbrF9Q
bmeE0sL59ZBkdxNkfjAU0Hs19SD/+DEbbU54vBatRVuTNnJT9W7vpNrBAEGHJC5g
HCUS8m7tgjOa0oXAhxkdjQx8O3yjMRYGwYIrgVx6ERC26cY5DzOwGgZxz0hsXNq0
39G+IjUT9SJM5e2DbGPv3FaCBm+DRNTx2f7cxYYG94kOHbh4nMZyJwMSTh/n4hpn
dsQcngQCc7GeOCRGCHYoRyR1QUG4hFsMumcD8HrbHLM+e0yRZZ2PvU7mb/7hJnd9
HeTI6qh7fLN0NtQFTulLjaUJyrI3yl/OoFjMLV396BrBQK3haOHsJ3la+6zzvuQ7
jO3WVoRjY/FsliJkfIm5TQoF3LJMIlRcRYUOUElmDEcObqSJyE7OaP1ZaBdSr2JV
8qmiIcDtg+26CIWAlikf9oSUG2KSLozh01+GoE5iGoWKjeHzgTrDbma0p+Enytbr
1uCEiCPrvrLSh1hTzSE2QlIP/eIkXM/iCW5qy+q9B5y283/SRi/Q1Gd5T8fZNH0h
vpaYCpAQtt1Ys/sTyYecBTkxpb7OlwI7/NdV/2Rg2VyHMzsbohpbBYLaVh3LV4vi
wIqy58XOOF2Zu96u1n4OZQ6/QhsMsWmBn9iDPeQWRleYYX9f7wGNGRDEQd6g3+kt
A8H6/bcX+sRdOg2Dz7DQv5+sLlhu5Izb2hf/JfgMHAAzbq/QeTpxfSsm69U4nOr/
Y62geemArmCKGif17WFzQw4vNChH+fGhdpTuHQ/efk7pBXz6emftPVH2HtLsCUmL
8uXeVTxBQVV4MD0LHdwcTsf+HPjfpmpO7SH5E8sHEx2ilzrt9hW6Zf+hoUOqMePR
S8yEbf0J4SZPBdNzpWQnvqprDxiyOo9MZj8bEddmPJC4l71QPmDH0qLkjA0ajvoC
PoLZg7sjpXlCK5unf2S/AlHcW2mTCaCsqRf+3TgIFZY4r7uSYn02kqN5cfuhN33e
RQFj8vXrnAQAx+i0U3BAsddRYwbrtqHA0zZvzgZzMt0ZWSxSA1y4oPbAiqqO01l4
Dmy2bBrxJab4R4xqb0Eg2MIak+tZj0Q7tNIXYffU7fbwyRzAFasVtlHCCgKH6lJM
k3H0ecjt2B/4/ePYHipQE01cpgKdNjROHwiqbTmUZFRWOXjPoKxeV+xIXGQfXO5I
WKOEZxREvlxZdH2VbLEtnPbaWRbdnxu87gpuDZSKGAjSylb7+FRxcGQxt5Iy25c9
/GyPIvrdrK37B5Kis4jCT0Y53lRCaPVcT4FdC8Lq7NPRtW2Vjc0cy3ziM0roQQ0W
/5n9AZ7pnNq+NGxtJXOB9obCX78uX6AO9AWpxKgvNNyaI4GlIfQFDXz7dCa4CO5b
NvwMBw9x2KgXKuYPQNAmpbcRHMkSFdtGLyvEh7tZAK53zB4Qb4/T0sstzbQg8zJy
aqCrWBUssQ+vxL75G4cQOfYcX/5UEaLzjYfdvRuWezeZc1BjoMXm5YhSVhfXMzvb
2VHYiTXI7NLr46CzLkCQcbXMbwAQWlkrEz3K3QzIULUJi4wECUF5T75I9zoe5VpK
0fcxMSPwHJIuTRdkcCTBJdrRHSs2YOMX8OYI3856BcqlplsEJ8WP+pD3TCjsIgIz
Bh7AcIdwIEltdmO0hBh+pP319DJweeN25LqBEE5581ACEV3s5MCjpHxDGoBgZVWx
BQ+xV6NoBIHvRougYbF5F1JzXJiYfL7ARCwYHEWb7O1wOZcH+oOq8RQaObzE4i3X
6igYxJUWYGSIEPBbhTvqX3e2YecUUAag1srkXY8QtkRMILM4pspGLVz7iok0LOSW
3/FojszWavC1KJPfYq2gs4zuOPt4b9l4E4oVCCGMrX5u3I/Yq1G1/kamZe9yffnV
Mab/XMDtxd+jwLKoh+tl6Wduw45OIcq6VKT8NCOn3fmVAIxlt5FHcN4GD6HdVwb8
9IoiQOtoNhZ0XjqicSAG4LnhwZtSCivmiWIbr2Ruql73m90BPRgRZ0igHWdl+2aC
i/FTRp1CljVoohRDaGnfrjkzHQBrh6nDFao1kTQA0ZzJ5KlqkSQfnCLAvzifqphE
RVaQJCvXnOlztBvkVy5PLRUpl5k8yupUNK/F2WDe73BzYvzDY1iYy+t6YEYHzrY4
NIJUKxL4if+eL+VXipPirU2Eb3fd55W7/l07+s4pUdC3FTM8FdD+W2ZYcqp5i61U
PwnyKmxkRNXZsA0kSrbK6C7q+8DnzbylOmetp5GAqwcO7FOdwdWlYzUSPKzYxUud
hkr4NEBriIYav0wuq6/ZN+eTjPwCHsUXndmnsLhR6kOHmBscDcTiKo5PNsqov8VX
pUoK/zSX1/qclmJXUroGt/dPAakXgvL8WXmHZ96l4ARKTQmfSdMgOqXzJW0bsZ1g
liaSisUizh/Amq+21KbpE4lxF5KIRCm6mA5lnS3xA2fgRv+Tro6uPk9Y/GhIp1By
AzLQyHigMK8v+j9kUz6Dqd6HxCk2E0zQQ4+fJ7QvaOLfh/5HX8TRBJIUw0WBSdfa
0q9nsJpmCGsYdefwHPaH5zq2jIOAjY/GQMxm5yi6IYjnvJoDJ1cjPaYrX+gnHXbS
OaPA2yNfFyTSz0/6rzVomTuthRQfPKeSMD7KXBo1AtFhiDU+AMs+IZnrmSOLfgL8
Ve0YKbW32Q7UsvuzIoaL+kN+OOWg9F1U5I56+3cmpKyMJXfiSAYJ6BWJZint1P06
27NQwAWAfVMTfsMqXHs33N8nsuwd+IrfShRGQfZhWauUbU6YC+3ARiwtyfeqv8UB
XtTGtsTIa5PKRQ0FOQN0uW5KHi08sEXtrjLN/F81PlK/wVj5IHCqfzTLYz8f4uGm
YdS7I1nSQPoyK1ge7WwmPxB0w8+Cxgr+nD+qSHlDy0ItdR81tKZoYjK5Qu4doGFV
XF6KUETLVPAei034uOpPBF4NZ+Rt9htGB5i2niDI2w63oUazBeTpEyBWbQ/+L6IZ
iGl1emoBAOjV+shhQvljnx5ypZEIzvVTYwd6FvvZ8xBms089yCjWFraJ6Uw0dONu
m94jit8L5SY6Ox/xtuC0EhKFw2yftBgVMxYirUgujGiG1/DsC6hDrCFanb6YrkL/
Xd9MV/JQotjTLl1NCdcJtHSl0uqbs65HbS+F+/9q900QX3RYRlF85Mg5xohtF59h
Uy6SPqPMz2thHhlhnX43MfbPt87FukI2VmPf6d3SEpsXPFpGI7rZ73nkN2YbFJks
VNzGRDeiOfjorD+HBlgunUmmpJ6D4+W/CPlKPKXiLSJLxAtWg6keh4mxwGvfGgsl
LkQ3qO/SDI8+P3BC/Eq94zucSTa16UzmHoUQbg5XkQ4UANoV561cWu3VvaxTxCop
1hJHCzQt8jzInstGrqeLh3kvOWzWbACYb0g/wIvEG9KIgwvbqsJe7rFpn+bsK9nN
gAOvMm7LMoc9tyg0omjHVOCaNFsrY5PR96aLdZhO4ZHmZRBow3WH64WdieinoL4U
ve4VAxXWD2+kZ/dM1qRXln1wnxcUB/5CvE49Q71kZA9GwOcnePveDDCc4rvl2JrW
E061v4e8dBMrfQgmSdrLcQL/KsK1DZaHo2/lFWdyAzZGPkVP47Q/UZCKO7YkZGXY
rjhK6I3YBlz42854Gwsdps+UtGelSBW5fU2JnZI9RNFFpB0EqaV3+gavG/j4xJe/
k2HrBELYiG64PnW6CPrU/QNoWL5h67j1Aj9FIvZdMcSLdk3Qm96nGAXhCDC9jzjI
5vBawi7V9sB3Nwp/WN2ehadFUupFEQUfH1xfjGa9Vh2ZgFQKJ0xT702KHg0U0jrl
X3gwAgo+I/JRhHsajvbrE8eHswEMusjN4Rltdd8llhHS2bgE1aEqNUdBpK4xIfml
b8CKgxhqBZSKHkg4uhfZDWbnhuaIrXleA2D8ChXt1BZ2vCcHg0kZagu/a2eOTgt6
F63pCX/Pv3h+6HHYmDkUqZP+cKxLS/T7M3j7A+KpY5OzjcNMYY3lwsHfeWWJju/i
MZkPmvHdLbBlhUZaU19k9Uetg088vFK7CzOp3M3OdcXdERWW5eOCABhrrfKRkjCp
aOmAWFS9djN+xzWHj6wIJ5XeZDWVMsoP1evVN6/7O5LvkvAZMSEl1zVpKusL6k3w
elw4eBrTf3AEfJYFBuzMTwxrgalxd/Iii58F5uDxWF/V8hxNfVABtCuZ1FUyL8IP
5z9bNxtttBTdm/XdFBk1isOU/6uOr+zJrkTq1Uyc13n2ydc/aA3MBxQqcBkADSMs
qdMNAwayFiY0A44Mz42brwIQybcvbqVAKD7Nc0XFtEkXVqPVp88ccCi50JewqaTg
3QtvyBsevp9EjfoFDjT+xGTcx40+dSR2XcmR+Yj5ewx4S8OatfxAY4QVi6XZz/Ca
AWBcY1YQM10hSflUgMkktck8a4lOpaaw3uYpGUqxLi/p1mvZLfqxV2k+KNPjMwt7
kVDqmlS8xGTOE0voWaxr1hjnaHfMvXVDG00eLRrSQV/BTG9+RbgU3iMdGQSFRBu1
honJ2atyamB+v6A0SWO5+yLTb+Wnqu6RjiFRg7AZ981TxJH2NACFJRPIIyg0DBxP
WDfQUnxyt0MHhVasTGdcGwv3G17pHrmjq6+H+0jmyAcuIgaMpR+D+GhOMyCStRw8
/a8YQjBcfCebjtVRwGzRCjQmbxmmY4ky4qX3jxSDPFkclMRMa/s9MqhEEAz+I9A8
P0Jf4RtY+ngw294UhcNKAl9QaUgaxseMItsSFGb/pbJM8vmT2QnVDzWuPcwxNcc6
8G3DW1rsG/F2an/qBSZ078AN2BHkWwX/fM3wnpiLqovvrFfgvGj5KIootQHaew2o
nrib4k1mdH1gNWAPqLslMi3x0OIckKk0DlL/kVsBz5fCpvZOQKpRPCCT4nCit6RE
l/GWeQEp89ccAdMGXgCeteolxzP4ltGlxuqwDU2ut/ss4OwINalB1SgQGUv3P9wo
uEwlEFi8mEinXgbspoYP7V/bOOAwrd4ZHuyalEl2DaUGcCrJJ5HVkMX6I9UoHw7c
PvMRX/1/TCSOiB60SXTpp5A1iRtwPXaB7c+p+fSAXq4MkGkrgzbZooOcQhIJu8qn
pt869ccYWlfPsnjNksVxdq/AaWYq50FsPM+As8tKPzeZCn7sOILMU8lsQapc9VVc
gj+aWSyq2HgcaX82858ogMoZ1co3y5GyMmAuXmANjWe7Vo+IvfHUq0i3FISmGSuZ
Npab3wttOf5+BH70got3ZVIHIrVxCyzCDX+2//KveFnLsRbWyPx+ZOxV2i2lVJuy
gfFxGSHIh9EATnPaD+Jva7KSqv0yFEGRhlKRh1lE4fmxCaE6CkzozRaOL6YO6gMF
2u4pCxNh7xk4LjtgS9pPSS9IqLtYB/ABPnaDu5NpRwHuSKEIsWH4YrdFk+s2di6I
rs8ZWx7Kwwa46nszQZA0KXiE30QV7OIbxaRKC0BLwZar4xifFwa6FUfnINKbQWsp
kVjiy+1s+TCBGDOuoqnYIoyP4v+/Xv8Cyt2YZX0hEhJWFlzY6+L6hGuXrraFcaM4
M7nqHKu/Q7m7+8JpTVHv6lbhEGgp4bKQabcng1as6qWcoE7JFLYoffpXKUK8Q3XD
Wv+2LdcOb2AdwavdyZ2+OH//Z75AucaCqI/Xm8JPv+QcDU+KODfqL9mZZrTNTKkk
5iM+YuF/4s7os4Befq1zUU6V1BTBSMcBAiOlUslpPeOqvx39XIz/pIbKcu+oooPT
YkVqAyqaGuFDqrbJXJNOWZys69hRaRRNhwNwO5i437avjZtaPhxpe9Kg4oic/m14
D/z1wZkpT4eIlsIrPblK9peBAJmfNjkOshuxCGi/vVOVXLl3S2cQvq47tZNQTEmN
8JB6lk65AHe5fLH7mIB5EYxvcc8/jneCT6N879TjZsRvJPJOiIVVdY5J3ahMUZ0b
hEfmNGoWsksvLrSLism10mSCat0S4wa+emDdUyk79BBiAHCrEJ040JTFN+UIjdgT
9LBKQJqUj2FcupLMgJ5K9PwS61QLYQ9jwt2E8Y8htwJNV4Bu4B0oQcyTopHWMsRG
faHCED0igRDzeNz3viq2L8WSWkVV56JYAVIv/PVQ4zCMN9vjLzYxH/TfkEuLhRs8
1yCJORfVemQoG0tGAakUjbZ+V9bpTzJrwNGpzUA03WprWQHncOQjZHhDy1RoEB45
9sA51fppwSFABbFYAYAf77y5YevNMB7AiVMEnJaRq45QyVVzvHzWNRkj11RDVtq/
XnDx0OtjlI8mGD8AGolClD7KMAj1pBsrG7VS3qjn2blW1KZvsdNaSKr2U/TFkhFl
iLUzgRJKYf2PTlNnvVNK2gIy1y39mQx1qTt1ZKqcJZB/2vTVWuhQqfOEiIShet1h
jgFkH1xgQe5MjIMYJfy9QdoGJglhD6WBkcsU85hazPrkqJ+tYD5WW8w9VULOFh6V
ySeMTRKsml0ILPPLW0y5qMRSISbe3op5gmMWDsYqeUFvHwZpLBHgGwyKYZckhGvK
s6ju6Di8KJA6QGPK4lg2XSHnR/t22sgnrp03T3ZppIgHJKaLLaF+ZI4SE0FVs8oR
OjAp3A7nZtbMwmCjAioMwKxbhvQneCw5LQHSUMdNRGF/Xc5ovcJEhAcqxR6zLlhe
ZKgT9d/cJp0UXTGPLrs0KCPah8a+S9DMu+OXENTdQCDyqOTKYBaI/Xr9awVDAp0u
FKO8qM1sK2yk4HcSSSZHlZCLEFMtmIvLsaa7bSNcLL70bd68IcQnAwV2bCu3CSkm
0rGmwayA+fjM1PahOlu7BhzjgfywBN58McesTEVobdRVXTk5wMocUMJv7pa4mz2H
ge1uLSzyhpp9pVgIlTf+/ZVFoNMGdMGGPJfcon2jw/mdqOPoOY0/PfJZG1uwApW1
+DiRWlpDCAME68H1o/2d5sbXjjQrKGQ4S+VMyq9RjEltWDrCYPj+nMzGgqRezEiP
5RvCx5HATUd7PsZl5LEtfpu76oTc5HRKJb2oOFuEmXiVGHqUgjc711VVVhtckRES
NEMzlmAIkUkVny4hTZk/Syu3Hq+wLnHwI4u7xfqenLVwYsGpJ717GaobnDyyFmD+
Bm5xonCKPxG2M7SP3535HmjPQEsRlTcW5w4Ox5k8yjA5cWJQv1vndcXar9PaOqMk
nkAYxGbUmP1j7BU9ia4mzk3RBxlH85hZm6ccuEPOJLbrkOtlD4i5rRcOxSNUONiF
MsNR9rbZZExFg4QfZgeBb3Zi0TYMfUJRU5oUX+G/mKgGNI1M64Zk/LbNSs7UR5hc
WIGpUHldY+gAkytV0agsbyt3ubaK9fI7z1eAfrXfhIQLklYTYd/l5bk++aC9xgDS
ynungMmijRorIw88PPxQCos1jLwjaLWUwuBgJhs3GycTPTob5N9HuqYfDWnjjp39
WF6dsp8Dib+66FY94YDbObbrWbe+TXQ19bcWsRKQGtwYdu/54NcdOsR47eFNl4rd
jbhgAGzwzQPY/4AxRJPu9exdFShSoVsefhr2hwE+mvOOAs1nsjyyUdWaMQ2j6i+B
q9/4uReKnMkuIhICXS11WTzGNdCioIDuvGyk+AwEYDYIuj1DhfYrLWN3DSiI1TrW
pv1eirrHJ1CJOTubjl5kxsU/9Xge/C0ZMVgnJf8975/vPZlodb/5q8Nz9Zt62EdY
l7g4EUzzBN2eHKTeZ3IyzeTFqt2VHhHukgLNBpttUssaMwt8THyKfB8mpBAnfkJL
fWvfbcYpcL/00w+hqxtteWD+DSfgNpC9VAt5+zp7TN1cEZIfZNJNzAcFanilKxmD
VqJBieuZ4KNLFxQHQFpgPCXpPrBDPBIkOQYmNq0smozwpsTbPpzQp2J3K4MU8nBm
mRbHV3MVC9BBnGmPWfxXmMfAqCagwpEFiycZF13r8OKQzYmIqBVjGFB8/0taRuIr
l2ldN9KwVXf/R4nSaWwleB2O//af+K/d6fbgJuMadHgVRNphbBuA44EY8OIG/TAq
JD2nd758yyMokz8DXaRdLodBgZCBv70GP9ihEbSXKazmpBYT8awlIuy5qrLKWcaR
OuQ0OctUDtbnTcGWI9RUkFYy3s+9xVCXhdS09yjBTJIUFnVBrkHj6yK12N7VZb0k
bGA3pC/jl3+sTtkL9MI9uTpKC+C6PiGUCp7dDRFgWx1+WgGlLBzytR1Gb3Rfehr8
edHyeDUnuvs23c1PyIWNVczMtm4Hvg6tmjo+VIo9GUPz7gIJwPGgnG5fgiEPz1Vx
uAolIdr0WXHyIgwoygMgnvHGzTh1G5vyx03qlE7RC9q0gG7KZWnM3pTT3VJ6waGj
M5udwmhBJ9hRYfgrEuO85EWzp/rtUZJ8WRaTtV8XFcsbmnOsAbC391Hq6Z1JAgBz
tHFR1IpIQ6k5LxUStEzGipCv3hXEqGjN+cCR1cAF+4QrpWdhInh3Ye9CJkI1wZrI
Hhf1qRCE7e7tnN2MQnsyS5LsJc+v9TmbPnEmVqERqmfumz4laFcyxIbSZbu60ua0
I16cRsJtm4kneQGLfrw1kpF3/2PK7s6V9VCQNNEBuuRumFhyc+1eqAC84bC/Kqb2
keBUxj79IFry/0ONlWbJCGh2rk16qYqEMUtNuPMs1/lkrnBy7RNkBpetYNyUrIxc
vnS73qxs2WSGnBNm9iFxZh+lYU6bL1C1L97h4Ex+iuyUEOQBeNJPHRkT3tvPS6Hd
AAfg2N2u3lPA/0OgX79zt84T6Z/U3qsEuXHq1gkkavTIVDeaxjyNDIUXE8LiOFtj
2O3CM8gFd+dtgmvOiAHXhJrditI9Zqn07aR/urlZvlIyqu8cFqmE66eMkoHT5R5M
YV9nCVGynDKEWN4tLdMSHP3WUvEXs761SK8RPhpVjBii0ElM618M54Aclq5maAnf
3lb//d02pb/9C07/J4RUeVSYqPvCryu29TAK/0Cmyq7XlLOXED5yEX1DZ5gB1JY7
jMhMCQA8hBuHFBei0u8VXVq5CWi4NEgjuKERWsD2r+F3yU5bpXvYuXHvI7A3NZNo
mGF8l9A3lPDnKRiNZ1BJFXkyeTYlXPC9q9aZ2PtsJ+iu/OvsWFXMaJlsJit+llMm
OcirxksAtgm89yipy9o6Fp3tDANzeLInsEdLQMXgP2FYvYmTZRYSTrNIsBtaaS/F
QxtE+PBwCSFsVgaDoa3pX+jRAJAgXdW1jUNyOVNwrkY8v7ruNqVun2GaQG4EPFca
saFwsDvA9VNLmTRxATdGhKCg6eO7WRJYlVG0aAvIpDNzJ+Jorg+jSU3LxgCHkQss
Hy36TslNDxDVtgZW4TFbnL9TMDx7yNtmRCSEGjnoKvY1u6Mo+7HTZKJ7I39wFSJM
w1QeVn9XAKKwqpbNj+KiiqBlcQLipLcYvbKdBoyG2+x5ztt51eyVtptlepC5KUZ6
D3CbNKL3BmVG0NRAkmzkExa+wihMqenHZrrFKTNFRx0F8zvK16xlaiZXLK6U09Nf
DGCtzm4yuEc3HT2/uKBNQU/6DXUatyGXzZ3Emu/zF5SFWiiji5+Z3lYCqJKZWaPk
0iuE2BlwNmI++KmjQ3Z521HW5cN8qcuFBhHLLyozL2MwZggi+wKyu0I/Zkung1pP
XFier4Y49BUB+8GjZ8t+iMFk83E9AoomeYlHIl7oDXl6WEbm8LeOOyrtalAQSqfN
a1eV7nZX6LRU0qdseOCCgb8MQQNHTiCjbf7ZMUg9Kryr4t52KWTnMSoWzraRUM3Q
Bth1y9HcG9yqc4URpJ5+cIgfP6qikJQQtCgvOilGLRhLsZpl29U5FJyp2hhL9oda
HLGtOKggbolAP0guGKbcKeiSsKtFwupmSazEoI/3V7l2Iv9UbPer4n6khaukpj88
ZBtBeoE+y8JOZUZ0HwAAWzjag70oUhdbpZghXjz2P7eocOrpO+2CSiwAaSwfH3rl
yI9dge6ki1KxsI01+OJXurEA7qRgMwJgccywbbH6aEaXfSWm2pYOLR9Gl/L5pInk
yWk3upAVVxauQip4b5RU9DENuiPXPfTnc1LfDIR+qohB4QN1idRFm0UnA0wTCy5z
Y+Xvo/8znQbq11yChut6EGnhhHKZsuCXgup2fGX3jC19ev9spmpgp/3B1sbn6xk+
hv0urCbCm7WYILU9CzsWXNYxiO1Cf8cf29GxrBwloqWY+1K28R7COsvoOmYBz8wD
pwhyIBRoFu1Eo4S2LePt+RNPiJfwPW1WtfCe39nNp62zsF1wyJTNp/JZ8aeE6G9x
2mEgHGhuxqX9K+VBastJE+dfOGVjtOle02bw+8+azceL7fWg2Vozleiq5C7h2K6j
zXjESRRQZL+s28mp9fC4+/dtdA43mEyPAU/sIx5rdLmt16ESVhmSNRq557ilwvzo
EURdUCePbsH2yg1ae+x4xV1JtMvLAOfiYaxv1NPPESjZTiIh95AONXmCygl9F4Oq
JQ6lWONPMnxC8rfHkXGnaYuYf22JXQ0OsWlTgjU/M/GQ1bvywCyXSnq7b5VZW2c8
ny/1xGVzwciym0O8QapxZltQHnjJtL9oIcUYhW5j+P1hxcX5BCmxyGt/Flys57Hl
YvjdwI//7iQRvHw9fYbSPB3i7XQ9bu9pQS3z/qFqAyK+0sm/rKsNa1u9xPBvmvd/
flZqN8kca6tvvZWmgrev+3w9Ug94TkmsQnJrBH7JCZaMe231re+/RMOpMG4hZm0y
evmiSavG8TCJ4MUWo8tasxSByqzsuJVnScYsUKuo8QJG8eFaG8Hxt9XjAWphk1bf
oy/zH+3Z6/Mz36uyh3sTQcK9B3sRq6LcZKnuBhD+KMyDXlvDn+PS1ek2n25V7jX6
dmaNrBbSGlFd1K7VCtYN5W9yk96VSsKGKOhQnVq+PJGmvndbK+hAwpcAfzi8RxDO
qMfI/4iq4FR8wG38VBzRf8oxpUBdYTVMnCL8xFHknHGS7TkTK9rpcK8EjetRdXeR
u02pacTSon9Z0hbTPVwVlws2KiadcuC14YCESd9t1hSd/gN6ecLFvPRJ6lbcyfwy
2ilsfE3qro1c8e91p+PfYZrXZoSykRl3w4Bk/2KnBaI4UzLCpAZrFMf3UiJHmNq/
VTCTJEp8rpSnSUej3Ceq5ggnSt0jp0lwrIBGMA8dKpcsW0BrGeoREtsLW/sAsWZk
XbPqJzoyuFhNdoAz2PKfg2ey953sApkj7JeoYgjGQ9HTzsfPWiRlglUAAwfwwIAr
s+xMFeyElUCZmwwM7uGqUeoxPakkC0poW+x7uGca6/Z3OuPCoO/qfkRujiLKhWvh
GT3j8tLGc0+/DClkymDKRMCqsGWZsaWVfMsnJ5WI+FlX7uSQHXil2SnVGaE2fNtS
k8tRMv/5CRBzxN4rA1CuYSswUH3TtQVwlekhGeVA4a/BqZDjxVk+DhVIoSQTfT5m
ZrVDaERJXsQEb+LW2We5wtRdytI1wf9KNVw1mZQq+iwrPMAy1mTMYdsjrSfKfCuU
zZvaLgQb5dh4TZ0Irjx3o9WD5tb2a2BxdqRzTimINE1c/D3DOEPGUYthLxGIZWFO
1eyIpZIT9xeIslGA4W5h8TejgLxFCU3vhE8zCCeeyouGY0/8TImARyoyj8sp4Cjg
Ub04T2zRJrYuCjShULC2xtk5gc4k5s/jKljHs960dHBgAaeX94iVlzsWgCKDzt3e
Rs0UD/SesQM2SuDOhsShst7rpCwTIygbb5I6pP8r3CWH4TDSAF2Oecnnshr++WMO
gtEdB1k5YEOF9sM4orvvVJmzT/001gnd9pqq5b5zEGNxnR3YlrNbVbEwp71MWDN5
H5uA1lxTQcbm8ccMyXO8erUdUj+zII3wcLetObKV4uB+pUi/dwfdtmdROHBtIOEE
FpBRSSQ1sQ1NVMYHWOtQi50mscz73h45y3k7OnepV4iRIGTeiEgEAl0GOXi3s+UW
xGnNZt9AxDRSkZVArBsJLU/h0i3IsbFo3ZlF7D4c1eZpmR+bQLyCNga40up9qdUv
dYPSN7ce5Uf3pWFJG9qsfqvf6QSocyGL4d3lWkxvrWLSaNr+3iA65VUvxpY5GPkE
KOnu3RpyKmfx62bUzdd7J8DoefRQfFhc7i/DsVwRwCXya2dwZJ5Tw9szOghFtOwh
px8O/c2UptJEk5ip0ZIdZdPgajS8NdPwkoGaAG1L5KVrszXjGOPXvnk8s6M4yE8F
DxBX3QY3jFGB27sgOSL+FeMzhZB4R8FGcsQPwTifLH6uMpgjZ0NPKlID83mCHRhH
j91S2hHTF5zBJt65fi6PG8C0l5rkCwi3kJh+KaaSkER1ZpVRVZNLPPh0YffCle/W
OAEqaS7UPJHwaFrlED8EEQPoRdRWKcVrZfg71jiCFrFdKGsk4JXDDQNeZoSLPJNG
Mk4UYsn9i/TdJ3PBDhskk2oS8o4S0K+7mVMwdA84eNdJdhyQRXFsQznJ2sc8XB4P
4g/XM/F95uklg3W6LL3O+rM/Fe3mGWwXrAPBuYe3x5rw6FywEmJzD1M7TKSEQSRa
aAyrB8wJ+7nPB8xxVi7Hj2qKSVpCgEpj4Ky6NRUd2Swz6ZOhHrXQyRn6Iwb/guvs
dTcqdXiplDFIQSfh0mmgtySiFbi6KUR8pmyRuHoSF9ELuqj0HMaFKMYqWOtzv0dM
kxhnd3RhM1xL/5txQ2ATfdxG/DW8WBnm5CHj5/HL+TS4ESYQ6p+A3X2GDgQoFu3W
p1QP8nY5D4zESCVpGzTufrRVEnICGmw6p+Klqy9HlfDiqxD6xLZwbULuDyJajTU3
8av8yAWLsVG7fTeKTHkotWlUIqA2TtYSCNUYnOq+kR4c8aabaJe/6NNgaTpsD7iG
Plxr5b7KL1Cjrt1xNpmtuTTbJIh4/ruStl8/m0jCHebhIARDmrbKsjTtAkQUeoXP
Lmugg1hI2yYWsBdEdIHQ8FnF87DEIzLbQIgdvGnxOA9Cxy471q66sboMArNoivTH
OrMhgJf1iO3ZOA6XeidYgisHRbAh+vkcGDA2CTmQk0B/prrGvtxdV0LI0oBmN/i8
wq04E1VeOLkHH2U8JKXOWx9YIB42MvstT2KKxTsytinZTPGt61OHWkQO7NBY0ZC4
cMBu8kKmWKwJn5eW7r1+8j9FNP6ypT2T1GwfXUqXcRaCiCplvtuDJia4jwoLKBUi
JYgnsH1T6Lx04AUaFFrKxUatldvMzkEOpoRu7rhb59IiNWX5FH/0cXV8B1Ah2obn
MP3bKN9NsZKHK+W3FM11YRi+oGdLcX6QDo3egSreF55eUAskviN/10dtLzKMOVNl
Ok92WmsTB+oEfAeTsqiWOGYwOb6UWF50dU4dRdmmIlQqrSGOcqedPLbE5vKDqKvP
m+YksMCVRck9ICicyiXE3pzjV7XeWPVbABBR/sP1P6SNI6ivYRZFBVGqMxHVaLD/
Pw8Ot0ZWAhvPO6Y4fcvuNhf0j7Y0eq5T2n5nKd4tQfzUs2qPD7hVhx4pO4gOymcz
o8vH3a0vU31POjl2S8oMRmysmpH2nI9fAjUAVZamyYoW6bg0w39dGOh1ECVCa30X
h9zsOk022XUdTPxWhphJeBNWAJytP3M7dyyaXTA86cw4sgRka2ZOKT4xE5mHYZIu
vKTx+JyLMFRMRcd5LB/py5BUK8cjEsQ4tSszqRj9TdenPzetaFZU52t02xKA3i7J
aOP55M0a9CdfRkhV5OKX+GPITuM75VU5jk2aEjLZQQbdfkFUK0OoGDkvE7sZK2Jq
mIQEGcKSurccCeM864nZ5T0VBNXsW+EnTml1KDbp+XtL5aRUVt4dILLiDsHzE9wh
PnGM1Q84XPY8AH6almexmKDNPrVszjc4CyA2fhd7dtxcODHjGZbIgianwBL0WDky
vCrgt22X2h/VJ4TJgTnjnM3C4pq1P1+s7k3IcV3f3wQR/nVro8aN1uLg0GKCKVJl
UJCcIovUQdLfsErlIfPBKVoe6PnpjyZsoykKl8EalPdtfDipmX8lTLiiGdp3Ase0
haE893Q5UhwwhHrTo+C3p0iQWq7LaAbxagkNG5LWVWP0fiTzBus5sy0ElRSQC5oU
aUMrspE38rScGGz1AUFmJCqnTBmVfL7Kw7WrL+FkIS3caU849DmNoxvgNC+1M/dd
0BtQ0EnnSFdp86iUW5R9O4rZsWZiuYBB3qh8Gu4Vwdi5fCxRCNjZql4TEMQyYsVe
nY8OQk1tVjoXJsU32crWPSwW2NgIDeK8qmXMn2wEVnmh3ohKwEP0BfQlDUYlccrK
x9VDfVvg4C5wnejMySTCtrZ0EI3uUiDXxQKrFxOlPa+PlRVtvAen9UNTfePuoN0h
XMaDevydQsGp2XhPOy0ROKAtEK7V6lt72g3bSJgFcXGwbQTE++D9zxjAvzHKBdy1
6XHUSUsbiEIDOvWW0oQCxHpnw3Nk8s9MgMSa6rF/ygyw6sKLH28FveLlCPz9U3NP
adp8ov1CEjAoYRaqD37Tl6hemTgf/fb8qoh0lE/ekJ+rhSRVcKfe9kXUGsYA68IA
l0PzQq06wFPaJqUlJOzku98VI79gqjLKEx7k2c6lqgpyX7tJzUvf++zhHGX9dmAV
qj+EZ8HhIMqtjdR5y0WSiOvcVP9QK08AUdPIUZ6UctPGufe1386chXCPrMFpW/Nk
oD14FyDvwAGQAqjrGtt4zAFq204xPL3njkwGsyhayikUsrLG1y/zd6ixC4lkoQgO
FViP+kx1cQH25pruh1JNl6MYQ6pODtz/aFuUKW3GVnyLQg2C6T+5ivOhJeLyOEG5
5D8yxEYyTFRUcVmlGlu3lxm+iWnOmCQG10LmEJBHN1fzsqrIwAsAZ+/cF5zh3sTk
ScBcTXvQFwSaRLbKF4v7sT7n8jB75F9so4DUjXgmMMbntUVRW/uYJUwY0T6PC1sh
tsMgHF5uGrZvfZfDEcydwCV7exvVZkOdcomgJfFC+uJOfrdm2/Ral6H22HNAzp2F
YSotSLW0fNKh1+w8GtmIu+gjpJ6s2f2P18Yvz+N005aFbI8NPduWCXNFUffnmjdy
W+azM2ijYwDjytyOHU+eE9f7n+o1637rZli/s1FJ+fuHBswoOkmDLXWZsBOUo14X
aye2up1Q3woN5GE8SR9y4wgVWRi6V1cQEiFNvzQqqyi5hTKx3qUYmmgtIN3pyQhQ
R2sCqKuofYb7yvdg/RyKrLtUopFdYXy599UpYcjORGuwOXrtZQhLa1JxD5yqcsW7
88eFwtV4A8nu/n/UP85rrvZ4U2DIX4X+0s+6jd1XLlsqZzIQVhRqXOz4cEo1Ks2i
9EGcghhVO8uLRGLS76oPkrVyQPCgfIbty8K7sEjmfbSg6GlR4QI01yNVVKR0N6MG
8nt+UMspvoffPCwwQ3aTgCWbMjs8zRKjlopCA10MHHUOc/LqVrlT3uc6hvXMmb5A
3Z0JCecXyfr83Fktg8pJTQeZwN1/NJ9lO1uTwvtud1NxH4j2mQkSMDdNRxDN/RPq
TKNVQVjZEx7DJ9qKzgif+LIEL1WDfIj8tMTYMmWTqATQKNZiFmMZ4Azv1QAvBJMu
55ygOGCVprC2S7f6rvMJKA547pX7oC2/i4Kpy88fjBPNZPnr5c3iTCbELMJSel+e
Bmac66XfMYl7/v7Th1uexzbD/7GoCSl+WJLEP4osVOgLabRVNt/f4InbzswBf/qG
ojiW3GR6BEd40QsxjGXg0FGpFECitlabURSMxTqwubjTj7SBA9ZyGMsOXs4k1z9J
TwuXBiAWnE9dTCRc3KsCz4zndwMER4+TeF9l3dHyFyQ9KJ1DbhxDcPh/A+ItD2vR
APxvebtiX3adSpY4slt8QUKbmcuhnBtmyQCZMybfNLExc3ZPvb4L3tT6ZOkKJQ3R
AaU9YFw9GvjTr+6wXwWr5+QsseWa7DQIC9lXDtJmtXNz0zvzzzZ2k5gM5fYm2tol
7Q3c8qw/ewmESDSlUGSQry3eLQ+6aJeOMmJpKCx8bflRTtR3rcE6e5A6tyFSHq6w
Dt353QIAz1QeNOCq64/uw65/L15WEGpexJbcqyas3NzyKwtyPB+nuI2E9xLHM+kh
ceBkiqjEz/OIDNvj7O1N1bNsl+hhTODIw+3ZSth0fvRDawGe7OIb1bmJ+rxUFlXF
BOVE4Yu5k8I2P7rPJwmtl4bQgyaZ0mUgX3E8Nptg1KD1AdeeZiJn1CFOQE7SFeaV
V5ZKOjKO24mFKCC3GGTBP0tjg10mT/2dF89VJAzDDUFaX2T/vEasd7UIwdrQMKpP
MB7Pdqzi275yL4vvk3UbhEwFbCjcyA6yGbvtmG4n0w2E/Ewrhrx1g96uatS33oiK
jiciZ/UBgbMoSeJ99BCf690mPDHkpNXE0yzvF0gti1fPW6Wfur4jvKmj3rEKcB5e
EedCkuvPahR1EGnuCwZ6fyhOeiutGKziUFKo9HWdNfajKuL+ZJV1M3yW2vdD87pp
zcVqjWVxKyWu7cvElakhozo17c7227OngD5cWnJY44XSlzb0roCN3Z8szYUNS5+d
u8AHJErGXIhjxYwD95FI/UqNCkx9uuoq0THAkc/JEH84JMyHnBAQQRhi59BzOfvN
GPFvoBkvOx3uL5tc7CDlhXMgolCsqE1VkVSSmIWbSQ3SNDZKv+tBUZG+x9PYIHvT
Q6CcqBjGqsgy5fNcsow8baJni4YYoKnv5UNNmORJ6CEPdalrYrlOGYuHG8DKeLqu
gbf1dHtU3VUWfTZOCod5CAOk0ZxOi+ylorq9LVAILIhWlt2tC0IebHXg1NtGnCG9
Yu56rkOA38a5YiGV3k4ssvNXICr3l4bmWliWrIrmnor717s+0826l0nHiQ4QQfdN
0fdBRSDzrhVOrPb6lhftTs/bkTk5WvWaI+vq+RObOIwk1L/mVQ5OJWZSv1++58L5
3JuyBHrKjrMCBA18125JmcOOVa20mWAtRzsOHZoCYGuPnvFqItNX6jILnCy+vXwk
8e85ZJBwLO5zI7b7xANDew8UJHH9WgkAhG3IwiWnKbasUQ/d6dcFgDTBI5QY9LiP
6pT/kIbf6tuhcg9qYM95UaZyxq2znSgxnyQn8FCt6cWDkOYvp0bwKHwCO5b9y2yk
77IcYhZgtWCZA+c9RmKXnMoOxgZiAM+Mm/1cRTCNDUGr2YDkgWLqHnxgzpBCbgbn
2zZyPMbTH+sWcCiwVDMGqCbphua0mY0A98WOJY2aKOQ+fluThxOvwDb776BL7KPR
tN3aMOZZr9YeEJrzXguISpRmJW0PT8csN2cGoG8PzfsinMlTsMvVxuLCppq+vQuy
pEto283zZafm+ZiLbbXcVxCOapc31lMSQKN7e/aUPdvTI/6h4hbinfVtOvqXZQrV
F7VDBPC8ttNfAWIyBkAuWMt7a3xYWurjZF5k5FuLDtg2f6FBAu6MCGsZ5ta9HmcT
K85FeIPWURU1K++LtSU4FnvJ9Rm5LF3tyxPGdGAk4eJAl9PWlS7r9Iw7TILJe2Zz
y5v8ILQJ1t28ciKCP97r62QgMgEP9Kfv/VHOvns4w9xDuyjXjqz005CIu57e74za
klViL/yny8c9zxNZ1s7+7EwZsC2I5mZdxEvfdWfs2qC47B84N1hTGNzjKVIvma5h
yuderVfHWufZV7p4G80UnsKqSLckbJ0P38t4ih7wUH/r4sAHTXxe4kGvjhVRTYuU
mM9M2vcQ/JOdlm4he11HYZjaTDvtDhX6VMlIaog9iKazvxGWcxNPfADQbRmk3fyZ
ADDsfAKA9rZWYhVVznKeU9egxLyqB7gUcFtnaXPRmsIlBTnsDvd5gyUaELRe4gc2
M0BWMd86Qbn7luq8tfMA/MOicz7LdZrg0Z8B1Krmx9AzkUi2pT8JvomaPyX2hwhV
6L56UxmyT9q5J9XFmsiENbhTLJqnFK3LhVNSlbc/iRY8PSedpfAxbj8SwSfwehqh
bSklK+Yttk59dSx22cFWGHWp8OQ2oe5HfE8v6APK5ApoKfcj4EkF3GwzAniZ6xli
Xoiz+Ubx5w5vxICS0wm3ZbkeMdapzfjRij/0vJtt7jzc3dZGpvnNgx6V3ZyDUaiB
HhS6pmBEp+BAHT6BnolczcJxzIQfaPHNUVFAH5lkjk8e9stz8zgsm7c42YFv6GJn
xmIXGSevHkkmcyu+L8F8IYtQImxmgHa+Dx7Df0G2+TZVsLO7UNdFJcRGi7SGNkwe
HUippBvRGox1gtosnpdZy7PA+fr1EyqVsvFEctyK2X5aAcAU5aaX09wY1i/TI0zD
zWMcIWKiZodlmW1xE8KZmu0U1MpMTdZ8Q9XdbSWJXN1aZiHtxip6mKet3Y12ZO90
TZfkMnOQu0kc5Hi2NhcdjK/YeZtSvKHK1e84zy1HBAebrvNmzR/4kdr47bpQLUSG
4Fi0UG1rzIkc0HiKd7vBakScPDZR6K5ISto6PZDHVukjjdjMrUYlx68HhqrRaUkM
vhnhTPmFJjgoBps8rc/U94Y6oQ92QPeacwvGkcNSyAeN5/OqisHKiwtJUKV5xp8O
s38Jbf6M9h99BMtpv5KZGGzaAg8E0LSxG5Rl3DkkokZsdZZ/4S49Vq1NNYyJZQG4
osyTwCmL/BTp4qpcOnET6B/x7h1XayRe5/NxSz4C+exIM9geZkihYQ2N3AETqhyf
nULQFft2bQHE3uebo2H+Tto9IqEQ3XnYz/Nx1JKp4KHxX+en7zi8/0SYVf5blhkV
QfvYQXIjNsJNDMpaoo4LAkUNthgYIF8lIh2RA/bOvYJuuusg741meYcCLGmUtH46
u1VTD19Az5COqbjYkpmLWzjJa6itvSDw8Q5TnCwCcVEdFfM15RaDlGO69ayimnuh
y05iTWHGAYWq90bhE40lkAWDOUpQ2616tFAdZQOG2g1IkHutdmsmNbLBQouhIoW+
Ftq6e2i1GnUyv1suBsWYpYrbOeuRLc/x/A1W9KM6gYGFeEr4PnyNYPgYiwuQDf7W
vGqKcA7UHgY/yEAYvHkIkdJQcG3Pz2OsC1agj2WFIHQtMUqRUqPCTjtlhtArq78S
LdgmK7NpVOQYLiC/3+tNklGGmksGyf/eZCOY8Q2KW+elzjVdc+BvAqyM64hvswAj
5lRprP3QAuL/ufA1BRxfmqGvU8sc0yTb12lb6eNIau3BhJlWjS1xWBw2/eq4YtDt
GNN11F8sWo8+LZkP3S8K/jJoPQId9IMsXnNOaco51GFKZ4IdmZxvaQmNUDRMWYQI
ZSSraD2a0/IfYGg26BOb3sZiCrCdwiCP2908/gRk4cAzKv2dWEIN7qNo1oD1t4sa
C/UhZQ3vOHOs9XWil769R3deZq2jKTX/+joQIEZsrMoxBTr1uxul3IXs/QJa4+rz
XpbC4tZrPMh+wOMo1mqiEQJA4123wi1G/4Xb6iK6Vix8DEPOhpkx234T3CpMHnv/
XkwnLmTaY9b/dlWwXuxMxveaVB11T/PczqDetmo0idESOss8gETKWA/z1qafexQf
Dxqbt+SwHtPZtrTaKAwsU0+wtILJmfipKXTqQOwjywjQH6uo9axLfBnrFDDONKmw
fKzQam9QbFCKMqQ08FJtZGMXJhokbC7Vz1gLbLqfTZV4HfKIX8J6pfuMOEheHgAD
KNvqv7Slg0grSYQDpLIr2YAwqJRhML8Jlaaiz0Fw+Z9tXqkcgDVuttnOaUJ9WfOU
wsIxuuNtZqz5DQCcWo0qC0lUkgjjztiCjosyzW6PLzUTX+rqK0AaTpzL0+9VYst5
luiPqqFPM2kszyQ2ofLW8KDlFtGTQWcAw+H1P+vSAVB1CGSQCnG3zRpX58qBF3ZW
f2URwk1AeFqI3ZW/EBssuJv5gC+iS91D+0uH369uuB+YCUqKpj0bGNdmrlKkEIrg
qgKLEM6h+Ti3M/SDuLlodK64PMSYRN0/Qn5SQjjfDSDbLwdZ2qtAVRaRVlOfxmbS
i9fE3RM7qWNCwk3Wmx81wTCMYWBbF4CcVAVlFKEuuqxvx1MDAXpI2Q6toiPWw0cE
hIy4f9goII5fG9sJynvT9MfHQsTy/SM1e8BBpVmEnnuJM6fIXxpcfoN5cnNRjLV7
J5NhfSU34nfvHiaOm7vBxJcxxeQ9chTyl9/A9FBcGftPz+5ZsySfkmdmaZDDXn7w
JzPzxsi68CXnFuvKXuXP/xGGIyPaH2S6yq+MsPQHAbGi9quAmeuAIcPs3KodX7a0
Qai5CfWutYw5vEcMhkc0za0e1QsIkeoCYBl+YV9MAPeYV2xDGnXI6QJcl9YlIK5u
sDjXydHxsd5scT5QSVT5zEdR2w7+34sFDt8AqT9j0v7iYYEHoWROBQPSfqr4WDCK
gqiZ0PJD/jcqaa94VU9CZx5Ts6K9w/RFPsm10yeruYOfN68+vYJ0BV16nTqtvp9l
nvtzK88IghlCG1OYMKqw8QT4dv+OMSNITiD94k4MZ6m43nJuo2wmBKOFT5/D2eR5
oSUePBpxd9VF9ucWby3TC9mE7RZuGUwHOTt0Hc3b7pw+mZsq0+rhLC5GmbfvGBnk
rhnupsZ75y9N/BIErj7F8ghaV21kWGjv0jyRwDUsxtdVDHYh88GacU3sr18Rmx5H
2/Rc2CjXFNfJCLJAOF4s1kdmx5KjP4Fgte5KqczOO6MfMWuhS9h2K0Llzfkm7hu4
0/S9Um0vnV39KY5xxvBGr4rT30dGeWWthpkzAnNnbBaBXcWWWuo9sRc7/vRL+A9N
mhB9Euo7bAPNb/3UUlfZblkAYBtI2uPp1SITUG8SLqsYmovUzD6gAuzbBhk7FN9+
T4C/NHSNCs9rM2WxmGvcSGjN8lxnGYr/muC48ZIu9cppNx2thAGCcJqswc6cR6sT
atk2c2XFwlqf+n5AXWUpmTLBrFnNqtxmtKZUTFZedDgXsd36zBu3LkZLUuPpss8J
aG6oeS6TYLxGQSXYyitc3cGNL7GX49Xd9AjSwtLny/Ezq10M0BS38kEZ9gjEeecG
+5ms0UtvVaMg5w+BzdkwMm3YuDZ+vK1VM1wImryEUy4q+nmbaFVhuZiKW0+dcVXR
ptai2dgLZiJtBVn03dtKU2h0QYqC0BRFI/q4YgoPWoacUD7Vq17JPjlJ/f7dh3D7
ShL5w//jMXphJZ2VePhVAN6eb2q4y47u2MVnCrvBGn4pAXnE7uVNvoA2gdKumWO3
sN82qPPpS48txLwdX/8M2mad3JbI+CBxmQbD8aLqcFnahiq0zd2WR7koZDVGpnwD
zyk3PgovvobnYDmgT44hgf7AcMNDNbWm8aqPahvbNRS15G8G8pAgJbHcfpFRxqHs
GmhJOTKBYeuxmAy0HjlqFUZRUyHmk8fEB+mRfy7m1IABPmM425ajmRzc8nkDozz+
lJ+jI9lZKJjEkoG7A35Vn3Q1G9YpnoANwxsiiKfWD6F0EvcDx2siHclpjsbZjwWA
Biiut2xkvagBAVe37ERzBgr73dlufTLN01Jzq7oWKTor25pzG8HT7pd1xkVXaMfj
IBzEs1lrBPjmdhxr0pL72deMnWytmmwPuGflFEbnNtLI5uDtxHwppm8Oe7f0ntn9
maAXm3qZ+rlyXAYLJxlpv6YecE6OfW5eeuR+cOhmd+kFXRwMvV2qgaxrKoUv4SFn
/MLR0DypQGzFiOS8aBkJsTtXGkzMQ+lm4Ov4xV4qr2nUOaU7J9+8F3gjFnW9dcQY
hKix0uwRkhzWkRo3uqhapwjb1kh3JWb/dw/nVjbseuWpq2IVpuf8on4c8Iz1OQJS
8ztMMXXRUtuFt4FkHylGyfjLc1PA8ci0vVNA+O+KaAkX2I4G/0uhHIgxIBKL0mTO
B36WJjgbgWC2LxlPT1EFbCaaUSDZSyCXXXUunpFmmI1mpS/WEmM4FELtlOfcu9pH
z4TBGv1SSiZKuJWDrDxAJq3t68f9+rMiK5ncFV3dx8S/HIyEW48m1cxzDowXOJHr
j/uDF/Yxz3wt8ACTZohAJ/s7FfeeXlVqI3rDqVLNoTqhIGYY5Pda5rBsUnAsISmJ
6UJa+Te9GYpihuf4roHsB2QdpslLLuO4ue+z9x5zUTLGoWuR5pYZjNHhn5P9IY51
drA4lnXUy/DdlNRxig6Fzui/Nr3qznno5rpINPvaxXH4fLgSvKorT91kseZ3u9Aw
XFd7U33jUQf6RAogdfQDrmDxGZ06YcKua+lbuifWzqa84hPge0ha1tN8//4jWEAG
/tLYqy2J8dtvFdcsnplj8F/qrUJHWnjyFkLWNg4quyvpJxc1Br8aA4kCh+OKFcsj
OvU5HHt0KmlMndw6EIE0tn4ww0vPfRaacCk/Bl9jyfQJHpsD0zDKoT7nxQ6zfBil
mw1Nty/XdKgauGs+DxGvdahI3Bf2fxYUIXmnen5g8ZWHf+VUmzfQBeaX79H5vUr8
oN5cx7X8ssrGTdEl3/JTpkUfUfpApdQmLki0vwM14eesrQ1sweCMpQ89IsqadTZj
3vQ+n3x7f7TB90j+CzGjUZO90+FszN1RHjKCyh0+jJxX5GzAqhjOBXDvy+ga/mW6
kZiGOx8hYLUUIU/U2FriLPk8EVFyQLkQbcTLP99K8siA5MOpqFoUaEKfM6O5ctc2
lCPTr+U7VAY3SZQNRKU9ONRTjpkFlxCiVduJnxJUFa5DQN3dnoyKfqRMkDB/+vqu
pi2XdCg1UGOjq7PFHjTh7x48uOGQ8QzP9W9G2elT7sLtEPvfMnqTpjPw7QHnbZK8
4GvzEMFhblnxcg9PmmNsqIFtE0T6Ll6azQbp2fcYIg8k4Fw77g+SJqISdBUet4Vg
pjCy0QI6hcvSRclga20lBhWEZoy5mbXFVlRhb0zb1rjvvRuCbDZPYBJyiX0dGOwy
JHaacieWB5Mdvz/5xluTNuCsLtd6Pm008/CdWHNj9ZeTBV4fiVoJA0p/qVKzqRFb
zzxZjEXKTaqEtlh7ohkbTlLxYcPfQxiAKgxLNaac/0xkR215xEXZ7a2iFusgoNBT
V3HGcPVieJI06pJoc10eCjiATzRcWYl2dBiU4UnNhFaNoferFFnpjPZPZS49mVsy
SPdU7+4xUA+BNwHqHs3cBDMbSPkO4jJ1rmx0WiikPKS8bHsVXeuYB0aRK33T7tzK
s3cOikR9wNGkaHIKlTfP50j83BfpU0jtSuBb0Sb7WkyCoXT6dc9/EcD4jKZbwnZQ
wzxKoiQKmp+pVv2oTL1H7KylguxLSg+i0q5aSUA0nORuxcuI7lX0+q+W/Sj60PGG
QZdJijVcQfaasNEcPFtHUTp9NShwTiXTGfhTOGgjWwjK1P8tGVLE0RXI1+iK3Qp6
8oV+nBD43TcZc7AipVXW4cinHHVFw/PGBG8CLcbKRCG9xLfKQkBIfWoNGeTX8jll
oHvwt+IFsh3uQq+ibXFyE0W2HM2Q5tPUE0ymy4lBPmk177ubplhoy6/NqDGoOOGt
8/C0kWvpQYE6goVMFJE9Q0EaK5nritneyrGilB5t0R2KPVprVUf7673fqWwQCN4g
yvg2B3sPEnlYD73DtQM3vGNz2kNwBVm9UWTUjYKsyOrn6BZi39GW6ls7AH8/sv54
M1eei9v/vRcN4/vQlDHFT5IrGWYbLTUrYs0TYiFwdACol5q38thMOiL6s+fy1F/8
oiVbTSd1az0xgE0QJYnZ58+NeWS2lWoT3jNjpq5KJ8tZLOa+4NuwcxMfHmbc/faQ
OKZBX+WWG73JWU08IAx+O/BsORwD36mq6djV8lofXK6HyZaHNydrOo6aji9GUAW7
1A7JUTxxWskicOWnV7wkijqrAfgMRnDRv+/HZ/8+eLuzU1tcg/anSV1MGQIb7WrV
AjS8OzvtRnxzhALJo4iFeHIA1Imb3Ac0QM/u7h4Wamk9eCIpPP+roqt3z6PpPXur
n6N1/JOcuKcABkLzckmvlRbnz71kIDSKKE1U3t3nqa8FIThRQOU0h6gaS3fNKbsi
OH0/mqa9Z87hlm3VZr+mM5/qcj+u0EegLO8ph03kyucSjvWBUtYzoqFv1B5K5EP1
Rqr+kYl0pJ0qnIHIQQ3jh1GRWALLF1BPezIc2KgyjolJNypPRkj2N1qZorQrWDnG
UNW7WKFFoPZR4HXkOTyrAozIXYFq0zBRcWjyejpQY9PGp4MOuSar/TkaDuquqAPw
6+mYEmHr696InJRwOsSNgxTS/1VlBzm2cBn7D8boIEGSies/63U6RL71a7+8DxUJ
ZKxFW8wv69BoKlXv5Re6sKS2ZG4XwX2Zw2XQQwYg3z1ytncR82+64bKC77T5wXH2
MpQcfXdIky1hHJttuu6E/huARQRiNCXYq2y6pMVJuWRVy2YXAuP10TjPvAABXuHj
4/4EtyvjZkfp40W7XIdKoANlxkuHQwWMN1Yb75SOesWHD1nBOEuFUcJ2YjjdUBzh
lNaBjBZTG/jx79iqKJ61iqckaOCxhev1MJqoYJEkbg3QDJ37CqPpAVOLcmyDs/I/
+DJmArdt1/Af34iNAqPC9tTgM7hZ5OspNysUfHeeevsgxigZ8e84XJepxMLxf3eb
9VA8v1JA/I0LKGpeZnRQOREbfejx5jLoN2FX4RVlBk/Vpl4GYYqLUr6r5UySgEuj
keTBTC4qFZHFYkMW9dscRoHNp2ovUEO5m7vBs5sXxrBeJNlsJMqFD6uXmk6E29B+
bDOmfU+S//ox/dpgYACeLdKveUoEpDEvV+T4kuACq9VuhcJbvCjfyiR04wDQZjLy
gur6l+mpX93lEhaqbQkLIxANfXxZwjZZH5F4mmWK4+KydRTWqvB/IcMjWAazsblx
5ZYHFrL8cQqXDgV708ZandCiIKSX41i4Gg6E2cTI0okmw+57olqifOpXC+fpvZX3
1BPvgB/tevGAdfpmtFI1PYIOvE0IWzRgyViejc7dL2ggRhS8tIxgWzRV7UOlO+CC
B7UU2KWPbAwP0ysHc6O7pdbv+vC51KE+abgxz5fIkgCJNhMwUCf2u2nny4KtysRo
vErRHGP/nyhR028E/jazL9AI8OLgJIYcxHL4+CzEFXcLUUu905uP5cy6br2JmB9M
pTa7ljK4G1fNnic/divNwFpsTi33dsVrDJXOUevAVdOveFEBXn4iOwxSgocs2iET
R8wfiLRD6JMSIASdyG5CjfYAQPMyNQI8bdwgAsf/jRUAi3yknSr2GF4Da/urbm9z
uio/ccdu1kBukEGLu5xQvN/bvUixRYKs3NaD22ofjSPLDFdcqGOU8uiZKFu/f32k
HMnCI8kC4O0ofPmUmr1GxmaBiO8Z0toHVCnBehh2KXJFj7vIz75uOyyg8zn2DIRR
tHEw/Yt9e8JHrfA/J83b3Vfc47aTZJ6vdnNFN2tfeNEVJbASZq8jrQC1pEp+q6HN
tx7lIrLyDtI7W+NUCtk08ojbrvCWGa6I3Q8DM9PQczhuKAOPkPJYt3OlkAuUomSj
RLhUMi743m/B47SY0d713IM1sRTwRmcApnJoWGPR+74a1gZPHSoynSHIuWJkxdxd
aBWig/WN/oEbK5hrQWTN7k7dmgs34gFgUH3Zyv6B8K7Qzwkq5cP70slNWEBFR7SK
UAQmbqAZAWI22qC0NWeN2RUrk5n8rC/WW7fNkKwKgV9me/nndM1hlXNcAMxxygq4
tWKX8zetIpnhscJvgofEBJ2THm7WJARbSzvm/0xasckkRmXzEnoOUoztXQO85hs4
xrexlBq8qTcXo6dNUV5gO8Gj7MfiooavvCfGh9OIZCO2hhBIxgvj6Qi5AM/xB+/s
ID1CXp7NGjxHwehvtXK3JcVqRXuYCS0WDWkD2OuTi/lIZ0hCtBDAHd7nMZ0hiFdC
fCEfWbf1HWS729nsBiJs4k3KRxxw0Z7qRre09BEhlBal1EEdNg+QtyfjfTiexh0S
DXxRX1/AlN7v9i6Rn5vLCNtAzNULTbdrmSThKpJ9j8tjCOW+biMulgePOK0iafJs
K9uDGdY5TMRc8niRlfOPwNFbg4qjnaPBXY4IOOdny8VuSKlNcZrav4adcmGmtovf
ijP6ls0f3k7rIM+3o/s6lW4VJQxf2KK8CVm6kbh8LH1z6OzLUdl8BkxpOcZyLckd
PZ238xsoknT1d1IVJTG18LU/IRqvmtfgp0yjqIA6xGHV1QGIJV6o/zBeHTUYRag6
jMiQb8T1WS0Vv4RJQi7dMqlYAPoZgEpGtQDtF1mBwF1xpkQjVzrmThbVeJ3G9Nce
9GhkHd0XMY8o/4n8Z1JwfXOjHOAajWwJmAKEhLJKQu6Y1vJWsneU7xYXIwRbj/SL
wuMVOad6pxK/3WhQDyQBDEcCnLiJJJesAxCNf8i2zDDLTv1L/FXTjV1fFbghkZCv
hnkXi6a74wC3Ay3QZtF/ffMZqa3fX2KOKtNNfFGWWDdFBzxvqCiscxziHgAt0nOR
OCXjz5kpWeaJI794PBOdn0ChDDBAOJB+bkyeEIJwWY0W2hguNCneJWgcLolFoHNi
kGtZtqRFsK9UEsG10F8ypBS7bPGZjJr89QNZ0MiE+h0LnMZzI04u60EPnwPW901C
ZXod5jUqFJdYhX2VwGkpGQOiOK0lMU2f4jNVbITl/kaPzSO4gbeaRS3WzIHCU94e
m9YHQn1MvC+R5M/9rO6eSwg+zBlchj6u2Pq7ZcbWS9/PXWP3UhJXNv6H/pdcrXT1
SNmYQWwGIOJUC2BBfT22t9ul7JMMCBlTdIKzzeUIiBn1zRAJqgflKgHbuzbjst8O
YmeVzJGV0am8NcKUHOJzO6Bk9uQlHVNhUtLJ95PisllpJfne9fwFZ42JKWK2H1Gp
8lShYum2uhw+OWXhqPjAtl5p4Zvti9V7ec06dhw0CQJUvj49AyXZMZrjz7tT1kc9
DpLTMqfONt9ppwtlHExbbpjH5e9yY7r/teZszygVoUZZI0R91He41asldVJRPnei
imMjEasjQhyjXYHJ3v59DvNoSPZEHX9QccMmHcdoQa7EUBxMRcFIcF0sD2YapcPC
hie/CKEiGJ6owppSW3qgYfP95OGfXDpl29XPvlHkAOns2f/rrQGhkh1qIK4C3JeG
Yi5DUnyVXBnuLachZJ4r9bqZlqgUnqze3KqdZ/FNH/gW+0VLCXTMU902R/8T59Co
qLiwwtORFmuyr8bBdePjyRutqdddYOsoIYuD/S5KrLPa+P+3cLHAGS6L9VMDNh9s
1ScqPci4SlUXSulQwKbnNmw2n591CrxZS3RipVB+HH4g5Zv+ZwvhnYwrOxpGRwj7
5FaEhBXOVvXiA5le2N3kS8TZKLk5hdO80eKIA/10II+i8jULgbPDFxQb4AvdzZ84
ODRzVQ3rlwVdo6/F2JC9cZHD++yBz5OmdBt6Nrxa4I0PVenEx50fG9WPBCe7Dgzp
nnLKzJDN3Cn2gSd79udd1u4irTz1phptX3MehJdkwt14atV12InD91BpXTGb/cKo
cQybyYGag41P2Pglp6GEocy9zaeC8a/ddAhklHXJ1QAed3mGhXIoVGEgmd/SjcrD
ob6b6nKbwAhqgVn+CVsK8eZpe0Bn3NVO9lzsgIkW/JCR0SCubpzWpEVjvxJ4X+eo
TXPIid52pIxUqKkU98rds4RgSaZMnlLkLM/AU0vFAyW/a/HpORODjJ8UllRcBl6o
Y8dpvrZnl9AaQzd15cqF1dHdHE9QrI7ttvUkyT7umzLExmIRHywSoLyoP6P0BJEO
dfVnvRjQGONf4h9TvhwQCtwgA/Swd8c0tcYMJUu80EWV2cV++pv12IUGeSzgaZTI
lBIPJERGLeBKuGSQXZlz9zVYrl22I7EA7Bng1BYAaSBIv0WCO/FfRRUpHtoXhpFC
RKMIsurAcX4J7NNHhW906kDtxVlwPiEpXbb8dCNo6hnu1F+nzgCdLm9Yqwtw6nSE
tuP9NNJxmYfNT2LaXGCrDcj5xjVxhBJN4v0mx8Tf7LH1SP+dadcpubGjfwNLEbBT
kusy9YMDXKHmuG0D4ukk01QFzJjDqon3W3MCkTKbr49/QjVwntkRvIrd9auqYBWj
z1WoSq9ox2Wl4TJDkTON8uxRIirpJDQWdRPRlO9FsezDRBhSg2akwZxhTLSFkOd2
9QyeuFvvT8XalEULDmoLsjQmHHFwwO03ZP6lfixW3iHyHhsnyr1GKElnHzwTLqRb
scz3AJHCXKiku1Gy7B+hk0GUV8BB3rcq5yKgnLMrcLcVSIbv2xg2FMv1ChvjYHdh
tGrKVJZvxI56PgcQwmdAeUXAMMfvgi5jnHXi99zap7RGHZVouOVJOWFXU99YLLjG
eaTjgWfI9D495DbIe4Z7KoD/AMP8C78J7lKatSxDMEA/MrNs79TreNwdzlxGRcQE
rp8IJZOHNx9yuSF4TNoC9hvOo2ykDyUisVmY7c1HTmhtObDUPlMK0kGUkvPqMRKE
cPjQp3BVQZmq+GROcRv8A3yeAhfZy+VccAgwnEOkb1JkIG0lvFMpYHSEMBuUkKni
SfZbSdKFWdlOO3GromZxgCBLhDcSAReqEVMU4akggq7y7JvwNIA/3ZJ6NjihMS1C
fWsTiCb9f/nhy/mjVtJGz+EYqGq218vbJiMz11uiGKn/fbsk3PtyRgkYXQgnEk98
jGx1s4pI/+iZuvvH9m01b1vr7c0J8B1oi8gQ9keduVGkxcqHFehXr4hEX5DwHi/K
8KwR+W1J5YguLVuwZSVUN5mhm0Kspj2ZkbutdWDBbiGWCirfr1F7rcWxcL4L/qY4
TDrDis2u440o8SxAdysVELql16svAJxlgvWy8DhlNo+ohzEgflm8Fa/4WIU+ATuG
+mrW6bc2EYrCdtdXJL3Q8H10PYGuqPQZVl15IJu2j9UmY5LTsNzq3fPr9JPDFEiv
odieJAN+GW5+uLq/kvvFypVjXz7h5h8RuSiTOO5psTENTD9AGn/t0RfViKPueAox
1/09tNBv62m0sHuBy+8RAlBd2yEZ0k/nt5gawsfjGC+ZZftGwk3L0LJh7IppDOe1
VuzwiBpn/CSa8Nz7sw+emYc7P9A7r3h87xSmSfzhl2Bg0da7HZgRdy/t0FkCWwkm
uvl6u6Aj3qJ/H4t6hrpous9/mrX8tSVrJizzxxHcLKYz3xJh6ddcyTb6FmbxsBNl
bY0ItAXARbXV3zQkfkV/1G34UMQmi/PS1e24xLX8LS8N2Skow4o/GQU2JZAiyqa4
4CmqZAoT1yFT6GsB7wKWSSZNIbc4iraMkSEOdqcnHdhd965Ws6NJ15szU7FEqt95
NjKUYUi/sTQ+N4D9FgbDIRECu/RrSdOtGJ/An9a3GNjHa7DFglGtVEWxNw8nomVb
SDsYSH3igwPIBGU0y5Z/wB3TQxQ77N/RPFwanDQMNi6JDomSi0JXpPfQXg99aSXI
HzrfUq/tqylQ1u5H/sAg+1MYSP4EgyS06X0D1DCpZDt5Eu+pDTbi5G3y7N4vaNQx
SYz2n5IR4wYy48votAW5Rf3C5KSrmlMTsbyuJ3BUtkb9HAw34yZR3FqDQybiDJXF
pVa6Qu0UEWmmr1chSNTg88n3TBSSAcBr9JTm6DfwIl89sx3O2qiKTtpvbzYuTby3
gzO8nvCAb7gOnhVnFaxz9cTOom7jMe9KTnOTyxN55V0GMd/Gk/exiyTFwxN6+KuD
VcDOxy39v6jFhgz5XW7fo37PdcXJg2UNQ1HTUGVTO42uGLUnrjbRLkFCpql7pN82
J1tQyLjAdBovSEXtAWfw+9S79aWn/LyQfe9bAo0WCv+2x+21ZM8hX8lBb4UnbmMj
AvOqh0RHg4r8+Zz87sR3TjWcdKCw/cJbGCdlD4QWT3U=
`pragma protect end_protected
