// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
QdUT7F8hQE3xsqjfCHYhHuDRZ+pCx7arin4gSc9Hm5jOKhr9kbKiEHxOlbmpCWGXcojhIPho0UNT
eHBTiIL17NDZLUyzJQPA+GzWInoWEvyat84Ro+r4XRn5CyPjm/FbAiidqAiSLerdhPC3tAIrd4qu
J2thFjKCk+aiG6kKUd/SMk+ZsacN9peDjl1MuN99OFYxteIkNmR0ua2k7SPkdLagvpwVYAI/Nci6
fTvBG40VGzTrx4flfhHwTOvIM38Zan5yRUKnuyptxXqS2/Yjsw95bb9+kT7QlRyMs3uVYmW6M/fL
nRcN8TXZi2Hny16Gr7G3gZ0NXKgfcp3/F27eYA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
QiT6euqfHHvNBuITgO33pjOIpgSIjPdEEenhHIIzV9mJwKJYQPnAUn/u8otf0xnodVLDpLefMk4V
/1VB9HRaR41Dj5srDgHccH/MX3Fcp+0YgHhWfCPgkRdne/lK98OWE6BAQYdQIi1zWElFq5f54xCm
38G+jCInabmytB4tkaKHZDD50F5kumlK6kn7vYDKwnls5JoxoSvhfQ3Bu/Je50zFwIi/0twUTuKB
cT8gR449DF71jIDu3LlgDHBm6Rz7vMb8CWmYYvUHIejyCJp1sKuIIlQqhRFOFrhxmC4OIFuyP3tk
6aRZLVx2FKPIZMx0CKSnlbAqq3anbyA/dI/kIwZKQo+u8sunUaUjeRJjYjuDyXbJQhJ42xoLF1Ah
0yCGnqxufW10AQVG6RwVOwE0w0eCb44/fYabHHDVoz4XlquMicSO1fNCtGkR2TyScEMi1lkt8Ad0
euqrr84Ex+vDCsNNJvpt/A8RsLX5f7gG08tw7fJpcBxpC6QOPrb3HS/j5GkFcEHFC8Ve6uXcHpYI
8qUxBREjDhdatKnZ3oqxmnv5NyyMeR6jCKvtOi4NfsAN9ZZ4C4iXmnmzhwo/F6smOWQLicX2rwCn
ImNMRQl8TGgRDDUdP9uBcrDuIurKMYJR9K9w65atgAhn7ZQhZVdHqLwg/3k3034YUNpqBPOErnQ7
74iTq9Zw3KtLlFVuXW8rO4L5QPUMK7hCkIlhtiE+59NzQvV6QnLYreESz2gIpEP7zDCKLPSXj7rh
GBgxVW0yY6SVR83XJZBdCJiFVrJIxqfeXA9ptCgGrt+NxkgL9E5HNMu6JYOYDGlFpYJzxeUQXIuS
cnt7cNLUQlK0P/EWzOTpmyMnpwWM6XBtIwpB/4M07VgoJe70BlzIKP9cX2Rh4l6CMInU/Y30oLGB
w1us0CQKjhW++YrTKwCjGNmYiqta9l0+gI75bwEiRY3RlfoV4R7gloZmmNN4cONh+q3gAArs7qMO
+/vigDQwcJHWhDPE1jNhQA3h8v/Rfw5nREQ4FpRiDpaAMH63xKJBiZCyXLp/aFGOU0289xCtbeRS
tYELYhcmXwiW4zJHMYMRk+05p8dhdFaVbDBS+kIBswipTi9yx/AqJnuJ6+hCYAbcyrSAgzobnMDh
oq0tivGe2hDgfWa4JISc7WxpP7Y4PEnj9T+yLpxklr1exCo71PrI0KquX0HWwuU/qoqI7V2JrUly
mr1bGRPYio78pH1Gh2HAuLSCo4UeDbtRIMkJphHPgM/DHF3clsTiio5flgwy/IuQ7q9DRWOGxQOk
ij52M9xa7ae8rl+awF4vSzWV8A35ny41Rfij6mAw2jG37P6kOBITBx99LHeYMPW0tYoXYU/NRTWC
qve8z9PM8DfryQ2oBcdp4YzpqU9bzc8y/KJU7h/DZlJObqfvFQ4dHOGhuoMj5Y8Tg7GxL012MsE7
7yqgdVAgBQiNCzv9hzXkjcW9xflNNVKa150UP2HvluFCu4BJ2qE/XpSAhtlK8E//z2h1knqpBCCU
12sdfLNx2rGXi1vKK78ueOmjWi4fzF7ucwlwjk23ZVQBImiajcgiMnroUGsvSBBr3qbu3sJ3ff2I
64NRTOgKOafRudI2fYZr5Rp6IAcd/T70Xs0FibteKqJILaJ+rxvYA7IaiXYwVCOiCRCo+YQw7+6K
5lgb7CFXGhP/TZG4/LVBIdNkifwMPLaYVk6Rd7TyEkjmSnvLpIYPxDYBaSwDAb0nepcCxK978O4s
ibRx6Ym1BDOmYikj/yuJdPm8Lop1rZeaxdKZlI01d3DmKa5tH3kSrDywMNPKXhZe5VE48qFVhHQU
hghDx0vHZEgMZFzJClkVxiy3R+VSfv5oSoUjwKz3UpMm1I83ndonTLuvYU+Pv4oq2umLaMRNlUtw
yBUwUedWjqXaiwV4rUYYyVuKBnU8/Mg4DWJettNcXne2bjDhrfQXyRbQMdPzjH9zm9MUD8jkTYY4
RQ/h2KW4uviTr54H1l8XcuPD5/VyyPfwtX3MIkJnRj6l05r/m9aXpIgywamk9l07YhS4eXWAsok1
ohOaXFHMWdEsELdBsP8mIO0zWTDVdnAeR93KNjlyLFacoEZyNt1Um//ArhZm+om8fOLQzywNg99D
DD5GtDkpqzde5Oilq0zPxZse7gq6KkmxKe5iE/TptUPQnB04BOAjKJThGo97u/l2xGB3QrHJmDKb
ZmeyDKZ90jTsxLbBFUYotaEnTUVTxa0Rt4Ct8ktt5tBPGnb909KYI7YFrcIXBlJvH0hsRz/d8wCS
VDD5xbZoFnekpAt0ATKEQar94GWS8i92Mg+le9oYLShF6iTjjIYCnuCtIwW4wOUvEHt1pcaErirw
Lpkzh7L4jBIRnxhhbYv4Xy8QTl/HCkBnT9q3iubsIMbMJk5MQ79PojJeXYZxL16UskcWBQ9iYaSi
/Yciz1SozUPyPGDfFPAdid5lVWmjaWW+hxBPwvq7EhP0d7fljrPpAEVqfsvK3yE+p5x87tj9GZ5+
mnDgNGQ2I4xmgVPZtX1winjwIqbdAUeO0wuWIvr6tmyMNZnF19MTia4PvCli7FHOT7eaNtXy1HML
Q+nc5UPkzrTUO5tVuq72d/cj47TRTr7DGxQAF3yyV2V8pLSdmwt04AGr0Mr3d3ttKceR7uhP1sBp
biVHH7EgzXEiigVwmV47NWynAD5rJOMM6Iw6I3A8aOX2I/mn3B2pE2MvcPt4bt4LZAGTpce85i8x
3OLXH1TOmydnCgyaGeYKvkQe1mWppCAqifJUBAr4tA40H7y0xxxKJuEvtPw/v+MjezoLMkvc5gKw
Nr7HI1XbmQDsGVxeeg9mUH43lYBfFjFKHJ1fAjn7yHuly+q/72hbgCMWYiW6tbIZeXQ9e9uvQU9C
p4eCLkPGKQkBjtpFEaoTG0Q+R0RFrDdcI03Xxpl52LOIA0/25xnVCIxJCATDZhrPNIeU9EPvAJAo
DIeZLSEJnFAQASRJJ2SncH9EP7KTyx+O4V0yeDXGMCca266MfIaaGrsax125phAO+rueK46/yvFF
AzTyCuS/GARcy61ii1scnmSVJnLdsctJ9/lvfHUAYPhy/gspyeGFZH1E7lYoUKUZ4noIreEopHYC
mFE3J09chRjnDMGOGUqGIzYo88TTcRD/3EcUwxolc7SpMzVN+o7DcmwFE0cAJlIJYIk+8+HZ1zcM
eo2nA2zuahOGWbOJM1ltxUpYaUC3F9FI1Ch33bJE1xNUNKhAY1tzCVqCu4sK3H7ZTPQT8BUMoZ4N
v4XN1wwdsVmWlXHUfRtXdNgtKg7UVHt0OdCSgc7e86ckwqODNAUxzLEhjflizEEP4mdpcGUWAVcz
fxXzpph6BptzOzKF8DgkrTKnBBzdlTO1sgpDB3CYZYz8s9cmW1Oz4Wguv+6iDgrdBnp5dFfuGnjn
4FPj2XH2q5P8pJmzpDUjHT+eV1zNjqz/hoDhETC5b20dKooZ1SwZHGkpXiA2CRpK/OUUIbV24eUI
/3DG2ou6m/tnxGhzqb3LiQ3iNFdU19u5wOJSxBtPoTM/+QZWXapdRyYqteySbAwEZmeH3YQiKnQo
5SdYIv9h9o769UC6u6Zv3niZpD0D8ZbzgXRIVsG4LSer/D5HpvHTc/S8pv1VbgFb7ObRyTbNzgCs
4fuC6RyTO+OEHx4tJmPqihJcKl95VwoUxyXVq8xgtucOTIRjsx70d6In1tZxLGzH+XpaR7ii5mxc
7ZdgP0VtMXHKstzoDjwP2SsM3YqIT/kjHbQltIveP3y27kv7x5h76ZruyzVcLoAvBNyRoeav5SU6
WSVhTfEc0HS++DP3BemU7lbfQqvIuyxCtRVzHtehLKc1qj30ua4P7+2sLRl6EU29n9per/srDfPE
FApjhoos/S7JcJn2uUtTES+wSrFPSKZ1Y/CTjS2/pGTEf/kyaUuv2utiQ0vdMBz86pbr2IMjkjvZ
yTswq2RjXzmONzS6BJomzl8cJMsA6Y3oIoJPFS6PFRDifAHDgNFU5r18Wflxmndie9s3a2pz0b+t
Shzj2qSqI2NoiRBKEXBFs60tliVFVhZOJOajRTdP7+f086K0JOb0nXQgZADv9MynFEjuJSvcJSs8
xMCDy7b5pkzP4gccyfMP5725asvYV1x+ZmCTZ61xjZQwtJjlRSI/iGv+L753rPZlroCaBbIYEBVt
1wWEXnrwpxr2pWN/67kWU1wpvs56GkObJ8fOAiQE/ecw4SFRxWtH2tvpoTOAjlBk2cT+R1cH7F97
atX3tB0Db9pdW/Eq+oJlfObgRQJNwAWq/ogUISCtJqWrSm4fzWgN39NNdzONOIliMpl94hOwx/1w
jrlu9uF6RLDc/npwxwAZ18aVNsGku1Qt6reSwtx2qNHSdTo88qJNrFvge/VGJM0Jvi/y7uuatXOf
51RXPG1YRJVxvmH5k5tYTHzdZ1UEIUguPnSiSTA1nEXshsJrkzgKYAX40euemeAtLkfGxLOi6frJ
4WGuv3yqnYzFIpmKk9uCmGdhxGwZth+VNXi7K3Xp/xUkz5qN4Gf9sR8A1M7FOm6iMBwuXVqc0nji
EEJSleB0KlSoKakr9pDcnMfwYRDSpFx94Kedscri+5ycYZjwB+V1P3EbWzn8bEJoG9lIRtAp9ac+
0ShxxibNYjS6zrPcNKxaGzr6ohSXtairXUISUTO92QLh2oe6kaEl92TeKS7JanD96AI2iNvQRbOF
0XvtD4yOQqvb/hTm9jdLAGifTc/hEoxIWuyPriJv9sAz0RGOGV06xLwD2rc8bogECW/NxjpUb2au
f2uFCW4+OJ5/do4QFdqVcSCZKNEwBVCxjVhpWsygpmVTugqNNEnmZCW7v3Nz4cNsbPClPAj1QlyV
/7LT9yFlkA2wQwbuJ6UYCFwwL05U62GvUxvxABnApbxLKmAruJNiCGnfnGzjuBLDL5hp3JjAMdt+
vRe5wwcSYRSfHaFmS4PkwhWnK+cmObjtFYDb7q2pplCo9Nowd+3Xb/OAgoULINs37KnVFhst4ln9
eEoImA1VbxwSlTMER0E24280tMNAmnA1NnkhijESu+ZtuSQPu7HxWaD3NybKtslAwWek40YhL5Bb
5a9xWfxaaNV4x6J7UoLpZfEJWtnFGPkTPCxcNziFAcjyTgBYMbXQYFWJFMLIHHP5Q9x6R6OaS/hT
zPq3Wr1MGZ6oLWqFo3xPZEWGoiK/Kfn+Cfcg0zPJexuYIvfpxeDRHRjJtdtb102AiT6OLe3SjW1B
IU1NOFkflFSUo78dD3Io55vwxytfpOHPS40eJ9EW4gQ2CYzgH9O9cxBAgOGoLGFA1Jjf91uFFJfP
CJuFyyW480k7RJWcI61DNjwW8yAuIeEgKywim9BrAHObK9ILHWkctnW7WROLA3YAXeZgKd8TdRP4
r21H68WQFWRzlNK6LXqrhea+Xylgosy0w4VAJUXkoKeteJUKG/HPOlL+k8IcfZ/w/X7zBWole7Ye
a2Fq/D5aBwhMwPU56jhc8qUekggpVEaQHdoLwBiQssiSLdkeKPXCFiWrQedpGs3NZtr13pFh9zj5
shEj3om+D1oh79w+SSRqqvZQSeYDLKEhNhEPBIXiPYhEBd1ugwLbANymmYOYqJciMV1EqWjBiu2d
lkYIsR0HpzdDTPDUkGejtqLuYmNFlOJDocbwxJ5UslktHDcrxrLkQZtwwXnQTDJLKWKbGiIhjvwQ
obmrszRNdeQEatkJSXNW34b1V1bpyDJSWAa+e9/mWVezbLqzCCI82N3LPG5fetxa+f0/X1Ygp7zI
QVVO1fa4Mx8hN39YI9Aot2zmKKH6qETTfg2Cf/2VVF/wrIi0zeFB6bffExWUzzAaBYBYarEZ5npt
JSTTpLgQli/NSjV94NcG7lkjODhWb7aLhsWnVWPYmd1Sa1zd8DT4IRntGaOJg9cqXIMIy20wIZUy
fqWwcrCZpNFrpL55nSa9qWx8O8xdV4o0tf52h0hWPMAZTf6hmszVWVYaREGSjOf0+QkfF28iM8ne
j93ODQuXyV18gjSbnfOXCJ65SFh5CVppRtiWiyMEJ3/tzYrm449IBsfDBAWqNkRnPy+qlRkfWRJZ
HHugBEy6KcjZMhRaHvpGGwB3LsQC9L+43p8BA1CNms/j5TZhejMiu2ty4nFHPHtWatsifUJcE12i
Vx60eSxeD55jXVCeXKkXwI8vJFtL5ptObtbNuhzBmbGpZWN5AVPrCK63o+DkjHxgdHefP8RKLQZH
ju5PiCIp51WZsTLK3qmnsui/TWw3/tyxDjErsBbo/hO1SOkCzs6KcqEOURTKQ/nCHLd5509rZ9M5
cb+furDORPqQvltD5Gh758dBaOsiF0Jf3gdSeI+C9GvRxapFLnqNIR6peobtN6IYkInSe3CjFbB/
eTH8DzLVbkOG/k0XenV61ui+1bR5LKf+gUzs8MRHqH19l+nLdHNlKpI3lx8gMylFMRSJJBE0RP5t
6/Qp9P+PuzNOsq//l6w6pYgi+dHoFOm8qLYCxZEW2UUeV0hplqhpHsMNB2rYGUMvbldKPFGIUih4
56xQtDNgezzaC8E4X8RpzXawjUVKApKU+Tv5u2yLWsLnxIrXJeiqXBSxFhBE5rwpBvUN56zYZTh2
qMiV57jdETkIWFlH9Yn0F/o2n9iE93MUjfS0YH0sb+poykooASBFZBZ2vyT/zijCDKw5rdajkCTE
VLA/kArkhxtR27m5BuFcwMEfltCjyzqlmUhgM+k97prt5zm5JLpeqGYD1Zva2XiwTBeYaRkVkq57
iAQTLSH/pdJF8kXHqU9nhGkLgs/xtIVDdwS8xQzCRkfZMJPEBL8lpubMR52jz6nwbpngD1Sf8OjZ
pgal4Rz7iR9MM1Xqy01XKQR0t5nDbcWekGIyr4OSnwZ8nl/Kz1C6w3Qj0qynVi6Nd0sHLioNQeV/
BSRkejLCc06EfW2IQ5E9Yb55naL66CKaE82rXlVoRI2uRboQ/SJlhyeOJ3yXX1ZLIDCCwNF6VtLW
uDu8Iok0I0Zk4dhpgbHfROiLPNR/DA2CbsiO40TnaG6ePejMXw7XGw01uq5UTa/uI09WSQEeKA5F
sSrgH6cN2Lo7bZ5/Pccx9aqvphe3S+HIRRao8w+u0c9hrzHNiS9CnIVsaoJ02oHpCrYlcsauBc96
zysX6THZWRn5ZDYLIbgfB3vfm6NrzgRPPzwHyveytncjB0+qsMpil1P8ZlTz7xeeutNyO73uFvyP
FbSYzZEFiJTeQY4b/uYZUYXLSD5ytU7SyOe7JLWS+sXlRsFUyyV51DzPcnUesP3FKtkDORMH+7FI
x4vVSU7C/sVoKl+TfLZu+g6INS1nF2nfp0QLBWjD3gnTI7fV9lZ1ifkWGbcELTIeLCsEh69yeJGK
8KptKRoqVqbvOj9ubOdse2axqSvu+1RldYNRNdad91O4dFNjlO7vq5g4fif0mCXh9XcRqlPE2WGD
6v+GZKq68gZw+sWVjLXuAcrMVDI2pW/P7+LxUu1PxVO+a9cp+i9YmbLEAjvoK/c6Jly3FijL+R8y
VcT3ZS6NHZFuO0L61HQlYln4xnAIiq5JcmvkDfo5+hq2HhhuGEDHellQq0yS06zKx3YqUDQxpqqN
apZWbhk00ddQIXMvYKDzlIlLsh6lBbPmLZWVKj4vWu6uBktxCSncZI4pOVcZIPTVzTlXSbWyHEHZ
/z1D+lWcnc1oUcuC2GOJua2fZw==
`pragma protect end_protected
