// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Dr2CzrSNFR56DdxWp8fm907uXOujQa+SkWrw0Uoqg3uRS2jol+DUa8+hez573tSqeFPKcAGYr3RM
w84ksM6n6mq4dDyCN0qszyglPhbYL2bi0N05u+2Gk4Xav9tKrS+/2TQgSNtTQY8/qJNsb3x3IlJO
Tkyy13W+m/b5ZPL9qrfIJKbM7XRTtdeTGutAoYFL11T/41SvsEsPgGLAWWyRxJqmrKbOK7l01Cu3
TBtJ3aiBgObtfhf4gwY3VssYNP2GO5Oy/g8FQjBzer/0n7p4nCVc+xcU3sBYmh2NFYTJJyRIex8R
5n4T2KG2OQEk7JriR1VjHIjl2jMxlp7c3PVcUQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
9zylwEn6zLGdZoT4v1KsZVK+tionfy9tNsDbDLXy90sa9UmUHboCR+fKroB/26Dp0yYERVtuDwf7
ezdXvXxS8ds3BAVr2bjH4f5+D50O/W63nxqsdOXpUHikHB/j4JxOxcclzh8xeqR0UQ0tCbY3hfFb
C04/9riLd7IxO9KjnV3m+wH+HEL+ztqa3XIcehgtTpqovxE0sZP8N/RMNJPTm/vLdEs4lHTLVZoS
pLpBqHhvHrDmoiG7VPohPJ9Wfh903UO0LV1eCcnZlP202t1RHwYMsCbpPOlQUo3ZlHqki4zrvJK2
H6GcUFBGZz/PbPxp/m0GjQCDyV8PRSpO8wyL/tqoRw7DJYXowcSuQy0EfiwffZqI3BvXbBQesfaZ
nWAHm87s0JPLBdrzrloLxqATAAoH17JLecQcXEtC6AV9fdlEE+Oshbopmr0P7CqwC1Z7VBCl+fil
h8tG+x9uMTctCX2Fr9hjrl6X2bDU1RaubmptG9QHyCmt7TpWIu6ilUcl27KVCld6IvSiiTfd7SA7
bJGlW5M0j4EjnJTAgRsTtXy1FmvhYEoqGQvANvlqNBHGYiop95ZlIz6pl7o2P4WM5NvqSTLv4Gxs
QB/PsMI1bDuNwqpS5BUjp50/bxZZSTG0X9t1fZ1jwPvUJttKR0KitETBi/qkgSGDSRK9Ll/Rs3Es
NdxoBZNvoc2eY90/UwgNSzfovSySaM9goEtcGsXkSBY+haylmQx7x+js3QzV8dINdcAWxWPD1Pz5
optzYqNTDzlXbptPGkFjZd6wnLfaeFdLFspXesKrfzQ+3GiMFj8Ol4wDEzLno3BteGyGsAHqpdaC
hLVgWvHKV+c3nTTKRBb3JnfLPTrudKI1wXi0c654m4OwB6x47YKGRHsWNnCncjDm93FBI0m8V/Vz
Vr1JBx4zFfoK7gxjw9nH11W3WmHNTWKu+xQCHi99axUwzgM2clHg7J7WBNHblHDOgimHa5rhVurK
Blg97xGoQEUylnBJ5mzTOEYczA1mptn176Cn5np7UFXcc34EXBHnd2JxNImR3yI7Bwv5tND7BclS
Yg7IjgKEL5C9Ld1hYZ+uBQ215bbQnHtZy9MRcuiXB3FHlELz1BzzuNQeE7NgL3FFRdWK4W3BtmKQ
I6/QsoP+VK1tDB3NezAPXso/KIwJtDTdYUYLEReKh4eiSzJH3krtTffPdJs1yUNHlUIgnKqSMI10
D6a206IFLgColGUKIREEt+AXdzXkrshR3+6YRV8qMV57UiOmoWP+wrirOLx3uGrMhvwtVdg6I7Vk
nvy9FXVEb1hb46kKzA1h0lqX/JJRl1pKDadtS8otM5L9zx5nKizrdlQaWWaOlznxG6KMJ8YMy+jJ
sspKF1JN+jsrK/0M7Pl6A4QRg0efb0TD2PErl2a3hwEIaWs74gDlIucqtE/b/287oNhRE9oE9Hnj
W9FJQCZ7a2/dFdFthfVB51O5AiHtPFpnkSncIKZD1qHUWOLsxgf5aFYXxAEISu79Qn/81fwrvcak
SEusUpyygUXO19LuIXLJObFUFPI0z8qMcaWcz2Nbdb/Mc/aAip1cMdIovmYFg+VxBePGrqA0/j42
VPERHAewW/YiV+bJ3/ee5rMLdmOud6lmmQ+tWyiAzlUpsVCdB4v9PryHYZK2vtheYzeqKvJv1VGo
mRpQcDmyxPDM/6asYOK6wB/AjXWe+W7Zo7BydYJvczlVSaG/H7iT9WLV5OR/VVckWTshY68dREzl
v629kvtjXPIBnYzzRfiIvshyeAetUg3RVEIAFtfYB4dEG+urzxQw6l+DjSM6aFULh2+9m+HRKam8
knLiXuxxShC80TUDFCYaxiUCMEFoh0tiGWPobtwLoiTWa+DwFnbHGWJiY945esy4JsBIDkNZRWMa
4cq1fADieeqadXMRSj3c8havbdtGTKfewNVO5SI4N5CyvYDrRKeKXQzYVRPRa2yKjdtVU/oH7qC9
T67atDmp4a3Un+H9SENIPuUybh+KTC/k+DQwRHFXuN8WJgzmM4P7NNvROiIGuMbBKPvrVOQ7ZjJ4
IOi+GqiZeXZTThMAzYDz9Xbtyjy37zTbOqvDSvwb5mhdii8CCmjQNm8k8wN3FLkTpNp3mTPElC8H
DX8+o4g4+q0XdV0E4nct5jUxh3zazQ8E1rDB3rFLdR/Fd6wwQhhQWo4exNQdSOoGi8K/V0Ym2R3h
KoxGBUUOa+8fRTFY0eQVz1QbF7S5xzQR3kOmEtpsrIWsnSODI+VagD507VK0HOJ0y1BOM/j4MZqw
uIvCAiyJkQqNVWHjVTtm65zuXj8wGa+eLiVPySlMr8RKNCarYP1pwTh+0hVH7WkTS6SFzHnp/Jcg
C3oKeV4ewOzBL4YJFh0im/sWLJL6MPhoF9phs2uDjGvsrRvQVQmqatgwMQe965j2SSPFT4QS2wQB
Wry8v6S5oGN8eoHkKD6ygWTIKNaTwwkM8ZjNFgE2xLmlCam5v21xWX3qh2WpO7uev+E7+26Yp2n3
aS0zd7XURVYiVEPypUaoOxAAAvJV9KpkAovVHL7nW0L3fi1jSgY2xuB6V00/iOKiyoZ9W7G9GsY7
dhUy5vJQvOT3qhy80GvhqPnI7K4mI7J0mmQYHVRAXI6gj5qGH29xovRsRClGPM45AWY4QeW2gNkg
yXAHbQSsNd2QCzDNIxDFFW04tGWyVf0Y8qjqsOormmD9aDgnMNhhkGfzcR+kHGB/Pb7Gc8CRsBXe
2dsd5OktSwmezwoUn1MX7bf40dbYx29uQdv0j88Qvg9w0F55MpoLeUAy7lVEGmcuFW+P+fK19Pj2
vKiId8pgf/RH8ylW52oJmFlOa5k0RA5PkvMqKlSp7w+jF6qVr+kFj3D4HLQNTrxu6BEvsy3Ao95F
BDoc9bO2taGOIwCYNHD5WmoH1w0Vp1lJAX0FnzvH+iJv8J3L/oOfdn8njQDg7MblFoqSwCGGVfyA
P9ntUNwiekkW2C8NmJ0cxgpXH6md9T5aHFodhV7WS6X6qEW7apjlC/2wFmQpnSbcmzBt7FaK8OSr
4Kk1Mw1+V6GTG9gOey4mHy2IqP9RQRGjd7kH+Tu8H0CvGhLIESmgatQOikNJh4rnLeaTxZ1p772O
yrRnLXyPaJjqpEykGD5Ptn/1+NM644lx8A9b7t94p3DRXUXGC4F6LvlOgWnAzyFTioxehtCxBeyN
IJZAccfMPElchcgE2tqpExK9Hh3yOY7FF36f5NA3tcNACz1tJi+jkzYjAxWb254ziWremVfqP1LJ
yeRZagynCp3bZxuYAmJo7sTXTgdC99QOXbjAffFFtOwglnHIPOlXK9hzynDV2RLOur3iCwW/Gmdb
owxgv0fBBKfPWg62jZgMpWa/pFelpgPR8tNVH/rlRK/PmW/7a7i14FFBQxdvKXPaS+FzOA+MiM0X
kWBuQ9MW8hpBlZu5n+1XSiMwIEThKLYGp0xgF+cb4BEhOXlyK0B1N+OJsgB1RLyM4Wtl81kOXfDL
zcPIbuQyPVPdFsWeVmToLeTK/tK+h3mkA9DV3wVlOqqkUIqx12znOQCta3NhhroDldmyoKXMAdSc
mTvqtPd9LcYy8/0cFQyUuVBE7P+8FVV0ySGkH17n5lbjBIUlUIFLOsxj8v17rVjcQ6hZTTR1+Ej/
xykyUO01TbHbttGtIR+DIwnachsw+AUu/3h/Sdzjb0vLzHD0lMby1gx9iU0NqMqXtj5P10dIhmVb
W86k1xPD6SbnkBjpzEQnX1uFNo96lsg157mtukR3ED1hZo3mhw7Pes9Zz3VfAV1hgohdKDdJ6UU4
jraA45VVL5Fe4lnyAmeP4En6Ty2F+obo1m1ffd6j5hzWb+1SV/aYEUmejTg+iUBzjjY04zHx0htn
Oh2yIxMDscBzjXYyy8JrwIACUQf04cAjXZS6k8eOayhnGxOGka/at7pkS11sSxMA88sSDE6vECvL
NQdxP9aGY1C6HNJ76OAyHAUUg9fEhWznPtg6tgO1xG2jGJ06vxu+/mozXlez1RDW+FWDpuMv0pz0
BwH4vrIGdYAOVLw53CWBLiqh/6lHDK3I7+cPgc1hh0ECyKPmsdybehNpcnd3SwTi3FpqGLAuGJ4/
Sl9J6z50CumEcqGi8iW/WsH2VJ0hgrj4Hx9JgOGszUhYZ59N0aOBPxWkZ6soJ5IXFGyjib74Ghaw
Qa/gDjods6NoevBmdPFSv8FDgS73eoQQh+dXkZnEHxxpaPEdb/uC5Ifv+lE30PcmsTlxSncG0G5p
Q3PcAzN2cCItWf2jLIliVpZYs563flszqN98qbL/8JZXoyH8+dOyIIuwEC5t0YG98IXcyHEDHpZo
VRynins76WSkStQU7H2d01pCQdXSuY/WtyJyrP1AiHVE6WMOrq/QXVIRDUKosI2AsCTVfWFdJRLc
5khKPdqjzGjxLYyGHXgg7BzJP7cy6X4m4okYjOj5STv5quo1ij4rdWzs4GsqCrvln93pgOQiKtKF
XCKQIPXx/RWBsFIy5QNFhrT+9WmY2yKikVLd7nDjo9Db9tGLmtm2pflqBFit02mFsW036xyfjP7D
YlqpjfFL0sazXnEQZ7fp84Z0Q4SGbw98RZKzVyXcGQNcXoldII53ZOtylSG1XgIMqp4bLKpP+o2/
OSlDJJ9Of7cQDuUCXYeBDi+a3czufp3uTkBxGg7bgOFRF6R2cIzm0YmqX2aTuPdAZDfgPWrxb+4C
38XVhXLYAJ2N3so6GwYXoJNkfO1f6Pybi5ZN9mxMYiEbfPsr38yRlDSj4SY2p1n71Su7U2W+/M6p
2CmrcXOslR4TbxyRMOePGLAXNCmBtGNpq46Xs/NJkDu7jDPILGGIk65mhU0Gren3CqaP3sOdq74j
ZPVrR+V/ykPQ2tEPL5SFhiojPQs6WuVK+xxke/kkrXPg8nhYMsxJG5jMDA1kDzPH3imPWWkRxyYr
TYRT1MzV/cTJOvuS1D1K/03B8gLdgtWMtEHUSLeA1dyfKOlDuMSmVM6X9fGnvSS1TcWiMAZWbM+7
ZpaH+0Q8VneeAaH35elGQdXyrfCSEV0CLZK/pkHTJNqvskHi3kMqRV3wDeOOE3dNUSasqUY/xtNk
oBbWdYZASUMBo6ZIDK+Xuswei5Hf0AHKHSuFJFCYwyIQpC3giEsxlEYqeeFSA1vYfrOVoniNAaWc
I8dvxwsGzBLyOhtBDJH9bPY51E1TGU8FtAr2T4/Isga9rFplanNa9jtOuJtGNIgkSWWJqqVfK27C
3Aityf2rXl72zQLnnumOBjwFa0VhAe4VPqYdOpc9+a8i/nOPUC9OF36UtrnDt8fPp5g8Mv23h0kT
W0zYZpZaXkdyT0WKppEYcZX3GOJMIbI1UONkuHB6BorafCirz1fYxsKPYMLB/tyJ0mAxJBUTn80Y
Qty3FLAhzkLfS4yMoD4Pe2WwoCd/u0jumjVtHE+sceKCJTWHgXFT7Qf/XTLJ69OrAthj9RnH+MQ1
9SpLU/Ztv6SRfu5OGNoRr1A91K4NgpzE6HvpsCJzCpYaZ9ylY/KGuvNk09oeSZ4dPgq9gtqz/NVV
bnJR4wLhfme6blrm9HWPANCuPw2l/sb47ULY+IYxY/u5Yio0QmCtjNzbrHLLKoo84UkJk3Vsyciv
fnOODnyMdPme0dEShgwq5e8LOfh4RT/tEI0oujXh1xa1TxyUWWD40qnaNPpA6KuHXysQ+m62C9Jt
5QhaFMeVzvtk4lDt6KMOWbzFPMk8nHv2RxLotJ+aRqQsaeiVROsYzATehy1e33hgW+D1WIlAbS+O
MRxfH8onsh1+/amvIPg5wizrh97wts/Sr0hrqok8YAHGqKW4ynC+0ht7oCeUtTlPqTsCaioiD5ua
zQbvX7TuYfV2Yvn+AMokrHm69zodp7RNqXCaKAjQRQeGwaFZIha1ykYeG4HZ6fttKVT4aMXySeob
LcNoxFiptW/oHejiWCUKDKPlH3bZz4yNHAthkm6AUDa9uJZBAhiWGJvMygSomm0EvOWOaIjWmN+2
1vOjVdkUwlKOrMrdIb1xRmLOOA6bVN5PWzrq0lRuBcwf7svvogRZTKNUpMoUfQoZWRTP8QlkI4MS
cy48KVAVDK0p5nu55ZfjWuTBLCFH8w+3rQpATWX5+9oU763cvKV6M8wVKAIEXk2bHkLpkAcbu0sN
5e49QobQHXcupsXHBFJV4ABV7UouDxOXJ/iXTWpokHjCDdfKOiCwsemh/7aMzd855HsFSG7kpDoO
wlgz0OymeKUW15F1NX6WStu81WXVg1wbnerg0x2QmnPQG9Y7Ha6igvzRViXw3AhTYUcf4vXQmxKx
0Gm3sVH1gborwS7ZQ+T0ipISgjKKXPh5hM8cAXdy5kCjrcZriZPIRXL9TF+078vH0nU6bCF8bVsA
ySVDkH+rqqOyNwNPGW4W8iKwyy9aZdyfWaLs+eAiFqTvqpQ7BVg1yOpqpg7F65v2NhVheq9JciFH
+mDA7wqHSjigC59d43DCb2Zg0KuXji7330JCwUOkWjbOEQdUL6GGFUOGgsu4I0vS/LaJc/lYDVWd
VOwPdeDgmrbqnNlaOm6k8eeFJDtNWEz34VVG7psW+Z+fs2OwXn5JrAPk4s5PCwUQlbx3iv5UuDAo
0uODGBXl/U5jtRDF9aWtyKBM06XzwMiRJiY0cTfAAHuCF7Cm/+CnKRdLikoZAUdvhbdp0JV28aK5
Xe2O3lctH3euRAYqLKK/orm2/Foo5zjcAoxx7390YeHH4RWjYiAFfbq7NkT/6UxQRfr7iKBR3GnA
6j6UQaXzE/ZnXwezyM5Npr8gC4XqjgQuIZqgj0YKhlML+2Qmqu9JwXaUDORScHMXvODG/N+5A9JQ
wSlgDJ6u/2aXju3QJ07inTgIeWpw/o/nFIK1Z2lMte86jCfW8fj+Q8fB2F9NuKSQVARwg1pskTmW
gTkvXbhKzZCDAqtOs/OlphDa/0sU0vsi3p1rg7St1tYW4xGH1JHyfh5VbQj6OSIOMubg6dhourf3
iZV/vIrvhuaFKfQm2ak9jH5bfyOle+NtmFwEeRaYg62T2oMFzZcdr5ugcWWlH55dHUuO09VZN58c
7m46U42AayjNl7NDZZNraasVH/sdHSOwgnUfYRyzYNVBkSHQU7978x/zhwkKtNk3tS5EmVKcYQl4
YMZQBvVMvsOUSdsozrf/PyOWtiEyXyXMoZbUnOUp4gvkrP+E2vlXzDazjIlBcQcbdEi6zgDW3/8D
vsMZPTPgcvIKiuYkTae+vy302I61hCppKy0Z8n+kgaDCWTEKez0WV6dMLTcvjbcePasSuWVa+/Oy
qWBQ/uzS8EsgC8KsWptVigGK+d5hBzUrfKoQ8A/yU2bccNf8bNK0pYPqAKaFPYFcntLdSTxDzgvj
S+BPvdFDUfcc9Uf9yyN2779wQi93+LC0PlLuiGdcTO2poBWOYSiH4GpKy1XE/zWtgBMNDKwfzX2k
4tEu5N7dJGfXgcov/kk6dgQUkV/3gwT4pkmvtZGuBeFSd0pHuPtfYOpArpJYLtfUzfDLbseLtUW3
MQmm7jMioFUgbWIfayRsr3e7fyG+viabWE1NTrCMWzgAxfbe3naMj9Tvp6RtxGL9pElqsNOlAcOa
hcZMPOgNOfDaXqjH9xyZdiQtTNJxRzCJxSZSMpGkSKXPQ96SW0PuRdEpwWHAu3BNjJbA3ddwHAFZ
3Q+dlAjOM9OR58ozmNe3t3jigUNWLeB6sV1ATMnN2F8npU2H/GsKwyM+sphyascAzkLdsfXfpmPw
07KMu1OOQ7/0MTRyYhGfWWNw3sjEQ8qc7MX+ysPhoGkjHEPham5q+dnfd/DE8mjYLHqyky6JcTPK
wzWdxxUwm1pBETOKzHuP3tUa+XYV0zhyWr37q2ZQb4qC49AUORwtuNU0JhBeY7j0rBtJ+UMWiqu2
wL/E0WmC66NMuB4O3mcmAcgZ3mGCneHLq7beVJaMo4jQW6dNeKFhrus3LmdCQy+BBNsyW1iKypMk
lpdcXgee0Ziv3UwIbkdaHQAQbsP0GjTg3GPw+XTjZ4jHDG5IOg7bnk4Pv10tBpCs7rPEc5SNJZji
yX3LthqnE00N2hZbA6v5VknOURIY86LjTH2+ah64mRxdupO/laGQVLWguxiMRzeq02iJeIlb6p/1
PLst7fClCFt8p70vUv1VtzS7yli04iv6ST8NMTB337i6980s8vhssudCQa6glLXSGzBSLlMenw2F
iIxNqKYLNy4VRlvU5PZXN6DkwyqCNaL7m/WxTTc45ZU2egh/LaGjJ9Mp6iD0vIGNA0aoAERqCm8Q
b1q/Y2l11tjaYPg+sqS+jtiBc6uL2Soq5L7P5bNCSGAi2NgPByynxQp/MxnX7JWhaMUldLg2Vtau
W1ALwtGb9wRDcNJhuteXurlXDOJXAP6NDNS8uAqk2HR9CMDYjg8L/vqj57YenQqoN4gE104yPF8o
OGe5jztPrb6IO4dHcVojFBV/AaATOWvQ3dCrqJzF4NclrnlAyPKRJKMsza51iScBotR1xs5jQZ+J
BNgHwiZpHjELadjYBv2a2r8gGYUhuWmEjjtJIjr5nL3PnaUJ44DUtL10qLSzz3hfClPo2Jc1fwgI
RxMdU2c9HOXLYa0OR0y8cTP8KkqT+8SjGTY9Y+f19FJnDwrow0cXJMr5w8q6ccI7n2Z+oiplAHuD
isPAF1WYnpK1oIeyZAavqjiUyuXBr3ULaCcP8qbDUmBydNZhyDSDx0gjFjLmwNBos3hWpqW7GL7I
xOYV1m38+1l9fPihqkNTml2+avngF64CjrxzYb+fPuW1sfILj8wvB3bPixwxLEs7tqV17EX5KUq8
OZKnpPFu2NWuRlTvBHyIsTonKT/lWZn2OAsFzaoNkQB2ClTU3jIuH2oZcRTD+bXgCcnkBg48HaLp
rWF+wSeQobA2IPrRLvEzjdGkRIqZVMCPU5Rawv80/8Rswfk0lrBmc0TUFEVSapql8AthCZQ0qD9g
NsxKsF1/+yfNSfWau8KNgIor9IGa+LZWV04zrYqRA1tRNQ/hapfThYmzgddKRco8Vj4g5hN4rK6h
Jz0uk5T/bLbJ98boAw5b+SniErhzwSq/K86B0qRCU++KoT1GK+CiLk4NolkASahl7U/mWZdy5Hy3
i553HBdIwWFUIZWLBFd0GEAO7z96hQlBo0v+3JAxY9mvJTwQI43F4p9ONgASMws7jwDhwNUsMz+1
StrjR/GSaxS2NWcytVihOmHC5IQkxjbj2a3BUqdugIpbneD2RFwkQS/99lIH7RJlvJRhYob9VVA3
sin4jv1xtC5aoqLPf2ckl9iD0L7jh2ogCAC5iS7BdtwcfCzqJiTBwwe5aLN19AoelybQj5ax9IHM
GSdIBcosVvuyrAWmT6wXrWLuG+ZDtwR5hYYcxfYzDJUTEvu1vpNzcNf6XIUcAhWWXd94/RpBhjhd
y6sqOt9iNO8mY3zKr2943FXDSPLfsS2WfXaCA5g8xVaGxpwsgFijymsiTjncAzh+K/FyUW21YwAU
gRj9r8lF0oD8Iv/ICVnqUyUIyzs+jNKPSuIxN48yVHwswPZsFB0B/jcj9cFxGG4weR/U8XGnslFU
Ryt+0c0+H3kWwQLwneSCgkLXE5x5kJmUY/FKSGP7t2eqCII4Yb0bnweCmOzsKdq5kpczVfHHz7et
TAflhcpLTczpI1im29kUiAu8NPSzyI/a9G8r2dWzCcN6HvI+EGr4GZ26h4RxtikinQJapTcOkfB8
L60VfwGuytYwbbDCNdL5tMRa8AKQjFz84RJphD+ao0qUO5PlFKnKmy7i0en0IIpWIXoISPIJhrO/
VJha55tWAk5EZLoetl0LV3R3+K7pkJ9LdWXyRORua34k+bO2+45ovCqmAuKgyq4+BizVaabwLl5z
1ZNy0h36ro3afDx0unTVu+2Uh7mJFjd4hkHfSte9I4DMqP9sE8AE6gPqQHVf+zgS/e2AQmwOSrLh
f5MstNRkHcO18N95ferff3JCwJ8CIP6OX4GLYTOlA52ryMB/CYSQQCkKfyp4306GiNbBmurrD/sh
sHJQLhjT68COpf2euckijk7OmzXtTVN4E2m9kZhHBHRf4k33uNVsbsCMnRRKy/bhe/MYBLC+v8TG
B5XMIg+F/43b6Uh/z6XaiSIR/F/cN4CdtuanS1DxSfyezAHHpjcmjxh+naIdJou8T6i2mVKOuTb2
VieHHjbJ6vtWJCn2yQnpPOrpThYGBdMvX4WKT36IPYr4jTmpsaGpOXcyt3Y4XqNjM6fXxaQzPNft
zWJBzRJPZIeZze3lA6nMcOYrxNHUvFbdMV7ML8rjzN3x1Z996SWCWYfQeJiEM54gD9m0vv4Bp/ZI
4wNeND37CuWh/bK/zS+GE+lbFq3909ydPM3xIQa/y/l1o1HQMmhorIZCmE3p140Diy70WofK5nxk
WnOI2jsKU8gxe7u/YD6M+NizuRj4VCVLQPfG+MO2Wh6dyMu4yPHCTYqVVb6EoeQamG03bjXHMYxK
ND/zPLdmGQItCeDt/4JpbVrQppQuDUBKnPYLXKnr96RlMDxGKAsNW/7Uxb8d2t8Uu+NIW2SxiFCk
1Kl8NFamyZqPczKy62coyPu9577XERyb2QcDdktDNQ/KtdFjI+nv7j75adhs4cYdZtHxWP31WAfQ
5v56TsVe3GLMF9SBZ92Hrl6EYJNwF0JFNPq+/vSAYtOd5LGz8YPiBpPzBl3rnJWZ5HQ23MEMFmRn
tvtqGidfDXmTf20TCcpUH05BygP8Fkyh8tKn6wSNBEB+rTfIwhlHZCGusFm6je3L591uTpqo3hmT
2lRacNxqsa54eSHpkwcc70LBfQktQMjZF/tOJiHHzVoPKkp2ZqCd2Fu4GTPiO1smkXQSybf0/1/O
SkdMRThPQkeqN+u4sXQrrSk5TJMr5JlKhOko1zyAbX5OKaHlHft64oPkO46+MVoDcmx2U5w/qtin
Ue59MiYdSfm6i6UbEwJL7rCPzFX/+NNODpZjNnCLs7GBjOPB/IS9xpVLMl0m1HZiap79s5DfTD9C
YdLeam9olCwXXQcQ/NUbzZTBthVveJAdIYhG5z/nuU+YbBlx12gI7zcA28uHR8pCJ0DJEkDuJPuI
UzuwEzUUnAbuxcxkmr6ocu4gPE744qLj+Y0l2GoX8voSzZUU6wxu2zkSW0Kbu4JVQSvqBpnWo86f
KjQ+jJklvEgTzPUN1BJ3/rJX3uGIweb35sw0k88IHJrv3XCs1hIO8ksRgO7GDj5Zv3JSo7uxj3ZD
lNN4Zaw8Ogmk1DTbukxb7Jw7XsAVQSaB3vyXuT34iilulhVTum8C9vs1T1stgjR9qxsDGdOyMJZz
L7NsSLZpdnsmY0FcYLKGKsc2DMkqwGbtdNimPkYFBzD2oO62Q8shj7x6YXv9+aFEt/Q6cLX3wv8e
GZiD7L3rJZmdXfz7BqzVgOqxmc7DwWZH74BMRz5Qazxjla+o7/6iaocwADkLOgNDLW/ITp+Orlz1
nUrW2s0ejkCWswEFereg6dTq080i48hVBFPwlGjAHa6VW7KTIAkpp/NEJ4CwSvoQX/R8N0kv/qCp
yr/GIT0pPpAruYbtsT1/ZL4EVJXRRIYXWQXNNWh0wdgt3OTZlvSYjY7prpxJxiQJGhqeNkOvn/58
jNoH6O1MphEaU5R3sOwkkqtwex05mkmUAGTmpAvfUlDRZljiG5NjJneonfmlBhSAsoWVvG7Ck/gR
QlOv53I2dyNGxMpWouMpJdzXG5MOLY+A8SDhNmdYSE2UqJETILdoSlmURCOD/L7vp7f6drlJiW8G
onsUZLfZ9rukcuNNoh0EdfpoinSQU6wrwpo74xiA5aPXd3uoA7BDka3LC/k1IvSjegATkoxZtpQX
N9QMTA3wWaonh1ZIFdXMBGhpbovJOCbFdrv54qgNwHWNd0RvJSXYrZjgKnWXZy+vuXKh/JqlvrCk
nCyDxpQN6cCux2EJ1Sa/ZKxOkeidhBNhb+EG+elEPYyRV5+FNPBwKg8uA7M16rT/jK029pQY4CJH
YEhVnozUUUjqTXWEDY4U3/ghIXNFCcV4lBrIzxhP71QYNb19kivGWpP9+snDHShhGZLR0kRqfybL
JRxHadARHku4eD5BWzlyDIhX/TbOwmXu5QKhM60LH9L6o87Fg/BndHOYBpBcG/mtZJAdYLwGIbAS
aKHwR1MchxQsNFpkQNJwwiXi8j21/xmUcgDXK2UKaxjbCsVMSOf1WdYux1KSNvj+1w+eKUA987N1
HAZs9LnZlaG1ySUnCRO/OmtL3nUZdyn/0qhePzNwqJVtiyRDPMjHc4fjJRqSXhfPOgMBankPW9AJ
McrH+rTwVk6EAB7XSPm6Y3xNKUdjbxdjJjEO9P6rW7XIgdRSprqTs0L2tidfbVtbFqYLX6b9L4tK
FyWpIBeESsDsgqMddKvjczJAUelvKipQH/WJp5BRe+4Fo3R1aCeAmsfpwM7Ypsazu5755q3R09vm
gAouLxg8GcUK/sdEqXaKaXGRxzpHAFH8s9BJ67X1ABmh24HlF/lMAgl1eFwR3X9snWsX+O1yoX+A
PDizGngzZbxDaShryDjTQKN+oLwV9p5weCfug8UKa1+yw021GzDA0oqz6Ggd/SVqSbZzT1hE6Co7
Lb9iYeHJTpVxW8oRAUm0hUDWOQkKo534Ref5hOqM3PWy8v8s8nf7eZQ2K6IXyKgybIZasLytkpR5
OFKe1HCuzx1ZteIz+a2smDiXzTBhS/UtDiYkCCVkNE7R4pflw1pRY14+2SvZiluYJ7HRusv5KTsW
W4D/wcnJW6QF4uFrSxCvRybZTzzs20fhSqGN2CtHDjv2VT8rRGQRyRrqase5x6WpTbKAshKowuZF
ONemqYQw1SuYPwgI/LDpJ/3MWfVTQjOxlX4Ouk78KEiz+91JjAUet0fWpNt2VpsLafejW9iqBxHF
olzLRjFTLncCN3RdvyEavVVp0FZhQyOhNdVKHmFzejD617c2d3mqanXaHc1bDcRANgfsAwgHEf/i
HWRJt6qXx969NJeP41wEOzqhuDNCZ41P3C1VWmnZCSSUIT/2p4eTJm6yk6LIGL6LZCE7llff2rXs
7Ep77cpWjH7EjOU8EImcqyUlE//EcYAcV5AYeu1Dyv+3yMSAkmeDB7Cy5oG5BABEy+/Jt4/wpHvE
d2oFuz1FMojDC6QuvLp/nKN/TqNgoqy8y3m+lkC9/BzFT7HXFefDWOmqBcIgllI9CBC/OJviOCFB
lWCPYXk7lsznSot4X1cYIQ10MaNR5Td35SwSbPpqyH0745XUdB3GXl2gQnsKd0Xcn/X0i1ZRSj6e
Lh+9NkEcgTwqn16qdBrs40tIeoTDimqXZPyPkZcVqzXmf2dGSb7KPZU/JJFMYtUD9gWv3fpm01SE
o/N3BZvTSq04IV2RwP9kZlk1/4oV8NFbztUaC+pp60szGIMebqFDaYIXPb872SYRFs7Y5AMpOYxb
qtb7s39hLz2H9yAfEP8yzzD/hOYbRnquOtnAazF9nYUZT6eK6tjNai5FapSw7weoTQu/GG5ZXRXR
kTjaN9Zre0/f3CGdDmhLKjMq2FmDse01i4RrROv2MgCtYHnpXmfbE/npDezwHfMGMLkwANJfvFuB
u4sXypk8K8aulvU3Z7PkRt622jm7oNF8jsfSXR2wCqxwh151QaJFSFtNeaPJ1fCB7bci5Ypcl4ek
1qsoUfH6g149m6m9yWEqz9av/XIyvOGbzKBqBKOnPsBru2dIvRVn9K2QXvm/qvlEJLGcQRtkcbKa
bhCqLOKXuwVXScq+c082GKkwVpWmanOZt632QBb6UxSQsBfDumQTLbh/0h/RmK6Rbldncv6rOJ8R
GPz1LathEQ+QbpRJ6JPnMwXv6IZOZ+WoBf+90XMCcWQOxINmMyO0vnUDehlLNEJAtBACIjUqDV19
5L/EL9qZDmVcgQ6jJYb1FH4k/5ih8TWtFnPtkyVUMPU6zjd+ASyYeQ0MloRX6kca0kFzRrVfpvhz
1DNjgbkccSAFrCud5/2mRfjalKsOAXgLVFV9AbBDPpU1ym2i8npDViz2uOVsETsHy8QFLBYNpKoy
EgdyyYwx7294XoLBgWO/IAhzgIHXfRAMlDArtVyBsb8ykwlAr1IRRTrWsoM1iEBLqzlPT0lpUa1Z
F+6xEFkMx+/G/NhclOLGNstCAWHNZOJapOj0dIARPdNQ3TGx/9fygrqF+cYabBN/fHh3nVg0gS97
gG0Ixcx7nEo098mdpWhHZywETVdkfDy/tzq32vBFTAbAaykvmugioSyTcwr61x2UKHmNGMQEV+G8
Fg8HnyjO/GkgNfxdtrl8qI40x91pWcPyhDlAaAnuy8fv3t98NeeV2wE06nkWLGJCFNOugA8+2gDB
LDAqiu3RJFOD89l1DmxHV/NCiWbrDKnKIitCPYWnPTArn/54zVXllpurnJ6KPfGAYy5+qxIVw8MQ
h7cgbUWwYnbwX9bs5CjeBLTtb0YkXe6evoIWZfwVQI0/ExD/xxxXL+QD2F1/WKk4xbocbIg2M7Ou
7EJMRaVYXd2dIaHRwyXO4oGFlI9N5ws8YiYm9nyxsh5asqhpfqwVIjLf1x2FHotYditwzfMdCD1J
C2ZAel58oKMR64rr0pYMkDrJHMt0OGFF2/jQI+bqWcoqp1//BC89fX8xge1O1TUQfteHGKQDuifF
OH06/mbuoH5lmtUKddx0ZSAtKYYcAm1Obch1rjs9YfB0fCmoIZsEyC8yQuU2leqrXY0cXx9H/z2G
mCv3ZGdP59J0eqqtfwxtpoLEcCl/ybUwfKR73bR3WER0MxIl/em0dIwUj2Rt3gdO+6lHnp194gEC
ydSwQTxQlGldUkhTX+ESyWbcMdLHNWcxPa+NQAaXgk+pm4ErYN+yrk7l46znETPSzV1swFYqIkf5
qBMxT/2O54bC14wchbTX+zHpNssimWSBf9eAIEnZQMy32i56XE95k0LvYbrTEmxVdCb6ynRDix0x
V+0rvR5ZiodZATuwWD7avP+cVgQ257/4nOGyu7866SEzjxEpH2CJs5QjQk2YVK8ytTOhc+6vAwmI
xeykG7LqjZ3B8HpVvo3QHXPZi1TtaeWgKVad7bpBJDVIQwFVfYXJfvTzry0oTb4NB7xpd9I0qvvC
hHgmfKPlgEvz8l+hR2kyh5eJbQI9iPihp0zqTl1yQsHCcvhNeiOIOk+/Vhr/J/UuHnP1c/Q/IuAo
2+Twl6rzKfcp+sKfA521dzdOgrBAv27k/pIhmwvpAk4JXELoCNJ8lyUNxsqa4dn1URrQFbJLVrmO
SF0VRDYNPZuedKg5B3g7L3zZ5FExqtJK2G3x9kGp8IB/l1f9vPCjBrG/xTzwzEFvL2/mGjh65AYf
M+u+WL1A7Nw+L5jfv5OE3P3jfKGr7jTnvU+ItNuyZ4eHeh8zzy0K/NmvxVnXbqc/c72vHetIbSwF
mZutEFTUF8TWkZUWCz2czGOqxgcCrGUJ/ZKPVG5v93ctxBRZf/irFgx3sWoEEYo+uVUXmXMb7ATx
UqNLeAiImWsqEtOeq3j6G78RW/JrDoZvZzVyQx2KH/4AzbCRoX+UOKw21tafclShnxqJ9QD3HHT/
yxJHM8SNB2soRMzngnVaw+KbLp1AJ+lzLPde2yWHCD2mNN/xIS1fMUdHB7MsaHlTP3C66QGf7wd5
9oBXn49yRADt7sKhwSWAuv20Am7ERk57WFvXTQ3JRjaJgelbKRXJPYWshzniDTSmdogqGsdNHK1d
LegYBjlyqNGgWtnIIcQzNagvHE2Ay1QztfmCiEQ9B33dStFyAVXjQVa7JtMrrr6RDUyfkgJ2aJcD
nscdPZAvPFYpGvYhi5FRO9slO1+gvkY81QTtrDod6BUdbwh35Ap4TY2K/gu7oJgJum2T5EdqRd3U
nxDlLn1cFhreYWVNxx06NTdlUSGBwJHS+HCvnF5PalHCJGBq6SkOJ0DeSY3wQgHcWYkdM2a5ZLPN
9QpofqOld6osE9e4Czadbdr/EJxdXLLDsWqRxd3ju9ZC5W1jkXe6ZTnnm2O1vE5xUep0gCCheNJr
MSoGl6rMT+HsQF1hODp5UmOYA1gdvDizvqkb1RXaSQGzhLgQcI716LwJgN4zwZdmGe2mO6FI4pAd
0WsYWTa/k1dw4QsEYIuVV7jMhaOP3nK8gQDZsLX+KevV1eghtVE9cIzlA1VylCNULeGpKXgxYvp1
Q55FWPr8aUGDdvSVrYMj8r/Pg6icUy+lsUmzR6shTDgjgdZys1SmG8a78z3dk4FBiIImKYB61pS0
fdrHrQQv8VV3Kq5yqYN2T+BOEMmT2AXIQKUhwMy0892atTBrfkp0mMtgxjN4ihujyORBmATIfi5S
9a9qeC88j+J9o1Wkh3sqqY3ZtlCc9bu2S8tjZaicnzJi8fEo23TBAS3NSCYii27BwzeVIXL3dPwb
lRGFNJww6xLOo1gE9MP3zRLWkxxY/zsMdNReih0iP02qtBEmEaETzHPAW6jBmT7WmUcMew+kde45
L6P8d7Smyu/3IQgPKEGPFG3arCnNlV77ALhdBYkmVDDDeAw2HDifupT/DFlsF2YpdhRpOCb3Z2U5
aALxf8IaUkNhXyRYWS6luY6iHLw/CHLkOkVAAneVJH0k6nWcvB3j68Kw7ympmqdg3RIg7YtNpGND
Z9Qmnzt7711QJEphzPJSCjLBgt1Y5pT/90ls7/LrOEVqx3H4xP6ItFdaPos/q2RX8R9ligOS8XoW
x2jludMGVyxtT9Z4SJD9m62jRs+hsflmmgaSO0xz42IEKxFrLl9hGTn02LTBNTblx8E/zsgs16si
0k9D0RToQywQre6TalUZ3eRorZfBt2+yrGJENnxsqx+rR7nucHSirnHptzUDzV40BdVanbVRvs4/
Yv6yIQGgR44OXk9DEdooTuec+lfhjaoUx4K1I46+QWZiuSL1TGGbUy4L+5Vb2Wx/8LbVMgyG/B2N
PCq2yGO5JA1UrAcg/xke7mGY53zRYUV88Iu9lPblg3kADZYTY1WBESULFsz6qVoOuwHcBqGKjr0w
pyX/maHUumQaYxLMfkSXwLAeDXVxZRUjbd5//m7ivG6LJdDZcXLo9Kjf6p89Ps4hH9nFUyujmSSt
ZnKrfC18N6VEVFr8AyHfJNgaMeXiLFIATsmJTUUafxhxX4EhLOUHGqgyNLbgp3QGa9bFyZtyuTqd
JE6pbUaN173KcMqugLbJAAcsHVXYSWLwaZJ+5bgOFQq1VRmq08qbmB9wEKRQ9ncgI1DAyarbVh0h
9aTDE1z185dLLk9HbCBE08dBygq64KgFWZq6BYuJTO57LOJ45LEA9hrTDQWfJQbud5GS/6qZrmVK
t751ty8FagnMLYEvAsO1ncV8ny0z3wemKvpykSQBGqexXnzn1bvgvf1UkZD4S+pFUnAFgY2rZWOK
gkdG0UcFu0rjkHenkaCSFwUZWTmHW8n0rD3Y6VP4bfnhqVp1gYkuaccdFemNP9OB8Y/WSZSczqnJ
tUmPkzqcAALyF04z5o5qQsmx/ksNg69ZF2JaZqnMSXhLUDHMAIVwKiWbeeQm2hEBgz+PDXINMYHW
hGOEKv03qiml/ugLfEeIWrth4rsEJWOM5rJl1JX30jeh62Yt8mZvPMWWaExPbQujJ32BKHy0z6R3
tC5XgcyyFPxZq2jEkdNF/sz/UfD0udJFzmZJkeg7bxdGHnTvTmzZIo7bXCGXzVsH4NLHnCYPVvZU
0dzu0XH/OlezvC9i0F4lxYbuPpzvby+tgyj8OxUTWWXogffWpiwSHC+ynJernQBwKYhz1n4H6gOB
EHSHrNg2iXAWrsowQvTUxdBuYGAi4lkIJX6MYy+r1bYZcGiudtLHUVvw8GCsvdk9o4GWWmJGcVJ7
7IbAO8X7wFqkRu0rY3WAwCz3ipE8T9nrPskMKhXm590LaAUydu4M1lfWvTniqnmR5aO+NAmCYTmT
bU6S5YffmvnsxoM1rm2TMqoXaL5qt+YliFcLHh1GfpS6hut0JX6o/P8+cubwYjP+FflnxZL6xoqv
K72FQYgH86QAYZf6aaXs6TF29xjLDf6co4K43hZgk12rjUujTzI0O4vf4zPcmwe+h7lchq7xqP8Y
lxxfk5bz668O262+Tuz2JVb5KADM/w4RJ6kvTe989uiio0R5pKWPOgT59zCg7uKBg1u2AGZnm71d
65gT0LVxXvkbfcmI5fDlphjxYsOg3ULzgIad0h1RL4yzgsaNP98hZxKk6nW78D5msGSzPICzbBAz
e40BEXCx0LhkBWQ053SGuXRw3XVGWIlRd5dnoFNYl1iEEBRkRWOwJzj1T7CQzf/rk9zpu7HQD+vB
xUIVR2eWw1f4WbbqokdxGklHjR+B3oNI80HU56eVUalDFwl1w0UKnd9QHmNn3xBJ5/vGCN4+c6Dy
Cgt94mO6EoFfRp8NbeK/fqKwc1Te4AmVUipwDGzNRONUOuSrvGwl2ez6c1RB4mMo8VJQwYvY90hV
u7XLzmLxm1ckv3EmFTN7QJUfnEKLnm07BFSoLd9pB8DFlDe3z5lCj6SmVSD7gCY3dfHkIkg18YSo
rqEsz2CvOKHghk+M1OmlLA80ItiCLmbbmykIqi6BkVo71LIdWlU+z3bxYaHeSCBMVuzzcyro1OGj
B24u8iZt6By4sO0f9RXQeoIH7pMtc/MS/LH0pOFzGfVrmIoAbHv7OYLhicQYrJSIVK7hZJVUutQP
hxduw0pyyurwQAugQ7yAJt5trWMxK6EL/yokL2NRuUyCyiQWNNcY2PnDzqMiVCPufbJwtTfvq5Ew
+ObBCTgD+Wwu0kViAOAc3y/iU/QbfX43IGJwYiXDjpsoVKsWeUiUawdvP+I1E7/33DPuZ4B7cpw9
aNWbpw8fUHVRzcoyy9qkzBtQDZ26QOQ6HJw97jcvGcJ1FUh8y8btRT9F8XgBEzd7lhQMO5PaBxUa
cDbha7JkX3NGBxNHW9htVzduPojyBMdPjebgp5GQBAcQQGFNqR86DrKrb1ifpzbnLewK2wejbtHq
HqPuKZSPxmyabJObXDhREWlUcbCzIBtTsENSmR73seIjRr8ocYl2c8j5BQlkrCzyhdaUYExK3rRr
74ggLanr/37jf4KM+XhM+t40WciJ5xRbgnJ3mFz8kQ1idhGvuHbkB0C9Lv4LEoX7xK2z3VaMDyME
hpgY96zUbME5mpqig8YQTwqX4JVCLxk8ABzE0bIo91HNjEZ5R0fnB4iz2KFn9zQwjzPnzFtRd5nL
f0MgfvDmcJGCPrgcOaqdrFKkYCEwYruCb14p+rtuPaXCPcks3Z26zoYEFxDTGgQlGoLbUiLSoO9Z
ctSfPMeT7ks7CfDXrw9kNlxPP589ZKKoJCMV61/I1O2CxXpyCApvTf3sDjoxTHY6/uFDeZn8UNNA
lv8eUA0REB0DjBLJ9t6H//j4Np6uhEfrdMMfIKeOeJstWX6RbMYnedIIo9VmgAZI0/S1cJei0RLE
Lo5RYlfoUgoGcKBJ/yOrbPdmwOkdUmrN9lXIGpZcCHnEGXmw1RCey/ACGKaUL2XOB+9+o27/5e6P
7PZ+Kp0daobnVEoO0rCaoEbWzXP+J0JQNbT4rKtcNMINZid2HXEdnNB6YJbrqGdPSTOWbySHoYoR
spA9epTO3kwVk4na7NYY5BTa8TvzKE7HeYeS91XDrqreDv4QJ00muYcfdbpsGkvp+kfAImsMQrnD
q2pWJk4TPHVztioGIcZ7ahwx2qb50Gl8eHlBpq+LkdD/wftzVVbjwClRg1uu6kmWaEq6rsXz5L1Y
+sxx/givlm/C47kcFHkDn5GB8CKciJYDBAvsuJ8owq1DbSIKx1LnUzq7e8YhdxiflaZ+NJU+iW7u
0t2cP5okSFJ6q3yG66JRIflZh82S3niPQGkP/F3CLVw14zBmbcKlQzITaUmxl7s+CBreraDW/A0/
w9JRZWPg0Fq0wFAT3drjvWsaQ4HC9P545HVgaAtOI3w4wnxbdlMpMm3C6ppFv9QbPOajZ+BFVYt/
owrYw8vNEs+pfDLIpWLo7yDeUggga0m5kaHQhULQs3ya1WSWIJI96i+PfMYaw5BNznS1RYDttlzD
buXn5PJ0cHNhKc0JmfMeZPc8h7tFyBWGxZGLiDJV7pJzki0KDygNI+8k0TiOyQ97eubJXCSGsaZZ
W32ZZQQiRgArUzU6LlSUNLFPhfejJkiiEbCpweLESn9UQNQuktasIS660Nj+GLcbdMEiIJqxtt35
jzxkhJAeQ2p/a+dz3ULqEwK26pSIfvX6bspoJddd7xEaRxitCoIXIdt06TCrKwAaZc0eGe8EMfp6
hYx3eQl8XCYEOn7a40VdnR9jQSPtjI5zA+omL+GHlpg7jJmPm+J7I5y+sF1l7JBheDZPkOazTNU3
hEd6f/K9PbTF/IzCNufyD8/hfldJTrfArXP1F8QWPtZ/WdLE1GwQyICbeW+OrfhwvgWiv6xCq0VF
EIlOQLkvj5VlahAMiZ0Gk77vlBovMqyDrqdFQ2elBoYZ9F1HVekBxIZiD7xmoYboemaS39LeS8OU
DhwcHWdHQlmZ3fh4HwemoA4zjlDkHpvjXs79L4Q/myWySlu+1kWcR63dHffKUgorrJNIXsfjqIrU
4JXub2gZJ/AlM5s7h7b4eQzQVy+xEjFo+Mkj1vg1JBk6Jtw4yGXIEtqjeF6Fv386siECBWkIy8ty
z+wmtpPORA+QN7ZfbbX8a+2xO+gTgIw5ILKKZ751fnPPHhk+XpuTuqrA74db59WalcuvZ8CsbV15
ZZAkT0fO/iQWpZcW7knuBzjxHS2RZoU0GSz5hfK8y1nSqw+QoUE72qq1Vubrck3F/mtwCCnVsqLu
K/eEI4J0Gm0aZdW0aM0geSla+vVqpC8MTJp1bLD80BhMEFaAKGM37Olp55vNBzlE0LgjWipCdeiq
mg2A2aJhYYwzXfyswWRnC8PwXbT/nGELVB2vlDp4pAThmEsbXZOcjdwbWbDIR6y1pyzqB5EdEpFN
sAarOOsB4HTn+O/Fk9KKqBUZJtvo4gv+tAfDhIcEVDY+PivIelQwEomymvOT/ZbNRMcsUj8EF0Ow
BSjyW2oHNRjYpNv7QOvHS+IN5agKQfwpXNJVvNv/zgnioASn9xEtcOtJBTMP4J0/RXzcOZjh897U
X+qUcznzwXjYsGhujLhN1hK4v3S/eHzBTeOffnFSvhlgwe5xjQWDgL9CwRUEwtoSJmbEfLxrH6h5
fhCDopLPpSm1nyCMRqMv5JJsQNLQehlqyPEKZrDgczcR/JzKgBATBr2bdG50CizAVQihu5DUO7ma
u7F1knHrSI6J5I3j1HiD/LiTzBIccgkpVY3ZP9OZMsmUS0eHAwAdKZqFPJ2cptXZcTVDgLE1etKt
ptZ+Q45jIy6umamlecXLhLGt0HmTSorRV3qOjpsIsMDuontNJjkWG13YvQwsguzXqul/2I4Yo76u
587f+CBOb6zM3FrcYsS0cbOCEY5QbBwkxpa/yOTW2XQai570EzmiFJ8nlL+Cj+MNPW9+nvGyl4jN
7QM+8cLYkkPP6CHVxkAK1m+WbWzg3wvpLIM6kb/bfJp4MWMWc9zjLj4+zYBZuWTIukmaqbzihqFa
WhzRlnfSjRgDf48L5r+2HYzyDj2517rbDX7jPqDa19SH7NqOIyFpYAeyb6qW+1lKWg+F4YngQykR
NLQ2NNREDGn8y8xRHryA7LutcSfT6G17aYwjB9isWHBWkIN9LlB288ry22Z3si++aU9JKZOYuBuh
qNiP0PSuSESlr8+6zB5Q+P4MtP9zy/mKAdyWCAu3TtCCZ1OQgigS0fsbgQjCdVSCUOYNmBnwBuFd
Ti3IiLYEQ7Mx/MBDtl0lpHzLcYsTO4m3ETtUwXFtwr6SbzgdwtL4/Y/mldDuhTAr47AeU/PPyxUz
A27u8onq7SQb5on1eu6r/ykixnXNzE/Ftwcvi4xbCaHu/amq7Ehsywl0EmqZ3rAmckgNMsNaHYVW
8y8QUZY5UWqaqHixgVhqI7m+43lO5vjTfXaAoB1x6J3mYzUzSuD3+osmc7DTXfZ+a8h9VaZLzqYT
fBNRCrPsjRplSE0npWpzg/HkSA3f52X0F3TGvf9t7rDz6xz+DmK3zBvVgbyTwP/NqeH+oTb9ox8l
r2DqeZcG7j2c1OL0ko1GA/GxmcRQ1BWet+zgyqx2HC6DPc8YqW2j7C/GGCVNJO1h7P5YR/hxACBj
GkVehjW8CDylYqNaa1Tl4pHCKVIRwsm0nZ+7s0ZbJ45xYy9cdXSFqY+lkj+W7La6Fu7bTeoXMgtC
UslfB89pV2G83acf54U9yfkyXMBYfTtBv1A8/zsh7kr0OT5Om5+aEwfuVqaZFpCB8764rP5jMGQ/
TmPEVHC5YJc8sjsqnWRoq8l79sEztmgdGputuJzjtAlqjsPDVHrKtLJl2hd565a8mv6ZBjgQk7b+
X0AtL2UHgWVEjRkA0DT+lsji7itbR2/ivdctCh3F+jzWUTSNNJXTQub7W9ATt2eqbF90eUT+KE3G
Q7P/MR4XgMFfqePzDAYCzmOep6kLJu3vsBakBS7ExC0wT0P/2QQTDmEXiHBrwdmA8tbM02fGDbNK
X32nvCGXbTg47usf3zVg1OSuO73zXWjZclzHCnckAxX9uL+fWnIhrpnbFPEjIsjfqN8P9KRkTw/q
N/CicbqTGBWiIumrj/9mDA3Qu33lzE1qKFUPedvc4nDDs1+rml8SA/yHcTBDwbqrHTvAfclYdoA2
QYKpG4uAR8+ms15oSvod3RQyoLtcguLpkXj3xC66XmAqv00gPmQf5X0dvbQG82yYXSJbTty+G2ZA
hdKVrfHhurOwBrECzo6EXNMzZugLSQnFF1EZzzXSPt0i/tzCe0zZyWC8X8H8+uxKGXwudgbaGTd8
GcRmQwJy40QbXP+NguXzQhFWhcXwUVoRtm3lOKO0OhHoIhsdhjapCAc/wPXrSKk9jYAhivCMlEqL
vXKqWUpGfdo9tRZbrSwY8bj3lvyC0XwBG1KVG5RWWSXbBHuiZYnAqfjMq8ZL2L5d6qaviNAaDK5A
cW+Mq7vyyP2BpsYPJ3sd44Ed29H0cbs7f8qPIbHeU7Q7XtBuG69/mv4+UixCscZYhLfItwOdzjd7
Na4iab+syfi4+UGBYviCHSOpz3onLWo7dUpig2AaFhZDj54DPhD7Zgi5rKgcZeW1EYek/pUXWfco
ePAb+d7CwGyxBmRVWqSnjz2vLIHtioHbDRXc6sCUw7TiHtxgCl+8TsN6gBDgQxrhMWOZrHq37pcK
Sh8ndhXBxzb/iDffRF03OcUKQ8GJzS9YSWX1zyj0uYWUqG3ip4JpU5bxZ/06Gg7wsxBHfoezdhRF
lpSNkNmyPFZvVbjOcV2L2u1hqRakmAfzW4zA2/UcCkPNLY6u7RxuRo6rZSr01ef/99d9gExzgBrD
TGTJ7vboBdkiwZhR34M+/q15lkGweOUFOGjKJaZe5Y4kH63Nem38nwPfzizqAb5UD3DrFk5Kfrxj
uGMXgPzZPXklQZsIprQ4RoGkrbjEsDy3ZUAJFdLSmy7j1hT7YW682Nm/aMZPWYl49G3pk6ES6nka
3hyDGhRTGCrnQSppXTTF0j/lyLoSG4+QTHWDQnbOe0fiWYuuKp7qgPihqphEtab0cUM2hy+XsnfN
3zm3IAB6LuF14lvjz/0dWFW7a7mYXYjCg1GH8+XsT/vDVGBgGwFgEPQn3U6XGnM+14EAEF3514df
SX1UQASmDjeMiV8g7gdpSp3W3B1ZYhASOkZd4IYBM7f/FEl1ZdbSWubrKkhmw5ZIxc26QLPdKYwL
/HgFcdYEUZUCGt2gkkIHbpNK1xRpaYimFUQSwtBGziv0qYr7GoESzjg7mIqXL5auydSFfoWqfRcD
fQyZMlmJG/Hb2Cw3T0zEX0vYteVfUnTFl63IW94ny9ScmHcdPJUMAV3SGQJky6k0Q1gAHKUxAgCK
LQVYAQ1vbWpqdulY+Nr+92Gstw5K3hlGwQn8P1r8rwxvoX9jbnOJW9g3C1ZsqZ93V/mbs8t2IGFl
7B95OYPZEPtN9aIDon2JfoD+N1FtW/llhceFgYYKla/ZhAKNV9sL2wOUyat6IQLVlfPpzZeJ8kTo
UrC/qAe/bvOvTTpawcUHjF9VrvGbdj9ZwfoHAyGY6oDAzFUbjHEqkcjrgvif0p//Pah+2vEzWvqd
UR7HQ6hmUh6MNSDDLNY0XytAbjrPNzQZy6jawh2Bp9AB5bzGNqAfhiEA0SISW396yKZIQK3vAFCP
D4o8Wg9I6heN3137t6JtkGVkn3pK1l5QjVP3MgQZS5k82Ne65gaWKHLzeMFK4KrunFN720mt0QOw
0wnZ8Gqev9TI4xxVRpgD5rWBrQga9v1Y5xHjdWt9wT6J0jO+CDxhLWLlfuEPuxz5KnPBfr+B4Mvw
PmC/4aYxf3bXuJ7l7vzjIzKL+k01HHGHnZWftGcTrL3VMJXI6yQSIU49ZsrDRNAFQvlO+3CYN56V
5IDu3O7X4BTPPFg79Q4oUQ7bMw4JWA5sZ3nch5Ekk/IYrb2HvfTVJX7j4I27q6X9ueGTRa+iZiYO
lUXIFkSwFWnuunsIb0PQ1Qv1WhyiF833SOuWeheyBlxG2wbLcBnoZe3Fq3Ej8dJLOAd34JYWhKbF
O9XbcU9E9vCaL9g3IuTo5iA42zeaUSjGlKvIYVpIzsReBHquXQqxmfjE4bjCIcqiZAlmoulnuK+p
Zs0oQKZh+4KYUWzlFXFBRvMl7qsP5XK2WKcwJJupgNSpxsZ6LdZeCbDf6ZLRlxH7iEax4PrKeTNT
YgswRECVVTt8fGRGNagGTkE0GdbM2XNeF89o8UFxf0wxRiMfRiP3hu4gJtdi8HRX9QDqhNi29xSG
AOeUJz3OV1UB/wLLyigQsULkBWOy8PcKTW3KNvwBLskJYVAwGz2TTKfe/ZXG17w7Dg3SVGxNgymm
bHdpdG3qnR9qrRWmqb69RZJhcVw+d8TJv/IaSnOJwvvNq2KfN70ivoPaz41lMCjGs2VMsJvOrxLo
ux45M2HllcvtDdGFiN6iIn6verSrIL4TxV2azLZVFI9DHF5tOrsK+rS73WSlCCOA2jvO+nw27Y6i
3b0F+ohm4mHD7Vq+6T4nZ0mQPiI+l+fJ5g7J+ldxnqe57hSjm/zCHg2WDExR7pe1mX1kbEowhCgU
aomJ/C90FjFreMVepC8tLuZ1dsMTpnas8/iYTddYkhoquma+GWkDCOTV/bDZwcRtxjv2q2Y+suz5
cm1iOVqkB+gJb0kVf6WVd+3dy1xHzN+k62xIX8fGlDfBslc8MtgxLhF0tpw9zklQiwjU5njQMfhb
b9bi/aVLtx0/z1N209qoN0Pdy6pCi5dfK9zwKioo11e84PDkzljIVOdjYAeGQUzhDp3AOKk9N75Q
v6HhNVSDjyxQpriB93ldbdvCM0KJD7z6cezts2QOsWQel8ttzWzJ6axX6ZPdtQioQYHqSZmctgtm
1Dyn1QxHlhd3cZkSMLRPMNrlgU3rVTcCdFmAUFhPsbCvUuuxu/Hm8APKl+g0Pwfh2TNat7crJgAW
r8fxB3DI+JTb1nq0W8qFoq3naxQ6Il9c597pv0yatcXkHG3Z3en6IuM0WY4t93DTeI84EOWP41kG
RCLjFBffal2bgp3piMKkSppeqc0mbTMIiRGEQDOElZmRlPe7wbFX5NqfQ8pNaT54vl9DnNFO+nyd
/iXy4xE7Jcr3ONOfa4/nd413MvS0JR6pfY5j4LHdaYq6/tRoPA/bPGJUkWdRfTblHmV0BQnh9Ucb
lcHS0XvGEtQD2A3CfELNAgk7FQN9O9y5Pjo+nL/W27G0K9tjVWWVtgfygMT6262LYx9jlSeedZ1j
z7Y5JNva4p8zT61FBUuFq5+8ZCluE9GV7E0oHHRMOj4v8Q90tYvCpNj+Tybn4y6DF9sT1pZGbSah
g7DJ49sZ00PqAHDwlVqnmeBBg8uHRAZX4T1bB3hZDPo38xo3vmOR6NWuqu9zI1eY/3fWVEa04B19
xs3E5lGom6qEld2XI7ZAz+Pq3kjP8xqqDkhGJHHngxpcCR0nviv+36P4+h5kpmR6FB6+yOt7Hlw0
/8/faX1sOZdV8hPUdoCWPe2V4UGRwzGY+VrMC7jDe7qBCK6VOJb9cUxiftDMcEKr4eBPzGq0jvLB
jeLIXXcwrYan6lABXGHRnvczeTPsvS30sJ/LeFdJuRvUuEzwTo0Jg+EEq4XBQQlFKqtdDtOBJkr8
CMqVyZiwgyIFFVeqyUCjpxjomV5C2vwCBtCQbw7ERNBoAA71UUe+2iGua1WBIJ5704N7b+1OBqZD
VOHahYGLXzY7clpY+k6WBuaQvoMVZ/ChePkCQBSzb7BXFdJVpCCJg8wH0WRBGjCdcHxu2yDCgTPC
kd6U1dlnEwkpZZt8uCIA48HFhhwZLiSt3dWmyc2h2nhFv8qu/9jqzjuvV68usoP9mwtXll2040VN
MxrvxI8aJ2wf1g/qHBuVYW3NKlcgpXtjreJW4l3xgSJCOkJCsbSzu/vZ9YSVmc4gdE2209Pbvmmo
TwqKChssc3RLE+DuzNomSc1xBOSFx5lnljDuQLLpqvVn3lEMdNnzeWjkKRwa7I0p6wHDOv10uTGq
gwsuNp57aVSWpmqD+DphLF1qzT4oSaqkds6g6YwDVH1TeOkYKL6eh71GAxFTeltEUoR1WyubgT7F
s4IGBf/v4On7N+pkScFDWbhjtr0GwcGkHFZi1ikK00wiIZYgF6xY1DRsiW3PuSVbHpJ7PT7CuBUZ
iFeu0wP4s2q2nyfEjnZKSH1a5blTEITQK1iVGEd56mWEtUROvWRtpVcB3asSmwDyzzh+5zf6q/Ro
PFLohmfTw7oKyklrc5YtlCAN34mBZNn0iLWYgps3c8tIs25PGOXQHpX+egZmLu6e1kSjnifTxY1L
GsSNOo9IAfRk0Svstk9Q+1YRwMu5z3KXbAZzQ3qu8H6H/v2DsdDlOEphGrPALqcPHAmyVtT44zOH
JHO5dSx9NVgjVspZIBIL0QK4BWOmG2STXgiufJEeHx3FDWHybQsbNjV4KVGtGsVORAxg6oU5OMae
M1d69cf61FWmqjVj0BEJs6wV/Df6VlRftiZ0J+TaOpoWCvRUjTxOhWvGs/YAQMHOyt+gx4r+z2yN
ZywvAEx0MrzCRolg6c36t5zbNR8UlRYA/i1HQ3Od8BCVS7kgS00LigTecwq2we49eF+86NY1QqiK
MRyHpY1OT+5rpgAl4iRK06x1hx4zuvgQAuKqJy5dv3OJ2KjgtbHcUqMxRoJ3wF3KthyoSB2CvjXW
0tClIQHbtX8Je55KKuok/uFzh7kmW4HwKvyxnOR+LXlsZ9TtjBXVOtOa2Xs4iawfMHigOFopHOTM
H4bkyN2BGHKpDdCTWWZ/XXPt9cqyWhK/hky506x/1YLtx/8Gxyv/ml9UoEFV2T6zBRK4tCOamGEq
ZgSX4zOlFMiHgHn9mN0YJxBsAcSm7iiyj0Lt+/3Ba+KfPwfIohA0HBhdmgSf0pvUmBOhfidIb6t+
b9FyXfvOLkOn6bLtF4tkT//BBZF90VAgg+iN/JuNC7CQy7xwbOO7r/RlcZlBThYJDUcLmqU/R6z7
32nJYcEhypsX27pOkf6bUL++a9AniwDiJ52j8GR/sRBMVm/2QBLpWr8olDgC05Pa76ULRrvH39hd
knaPPmSIb8+EGiKpfeqDaQakdGUrshj7gjv68iyZmjBwhtUH4SXxROcnKRTo6bpVZDG4WIze43wt
isaQgxFyXfBg4bNo4rsIXjg6Zgcw1akG6+Ss+QyNzFILx+irFo5wBjIBHC3nm7r7Ee3b9iakwrJC
Uf0RmYeJBmTMGfUKqCJjBekTxXpQKp0A0Eg6BiDaCdpYd22UgrVR+qK1sBVvJy6nohWCvnzsmQjT
JErgzgwNZdsOo6eFqmFFFMRaPNh1FtjxyS01i3naIdT6RiA1Y94SDXxlAub74QkPJAnrpvY2rgUG
FWb4K3U88KOc/nT6ecnyl/8W1hdnykDkgRd5o6BSiR0MHxrDzOgn3mGy1l+9PBWb0Q69k8if2eZY
vJjloJCU0Dg2+sFq6NJ2K8PW4OUp5XKN180ktvAJCB15dyDlqK68hG6bI8JFH3HVgpeQaJK+JkdU
m+b2NM+Ugz5Py/ryOgqST3eHim/4cSxWJlwY7bkb/f49lB7ru0PThUYC1RxZYdXqQrvK+u12+KJO
CJqtY7gfX8cbzoBy3MOl2Xt7SJ/Tep5L6NvOhzc8qLHcX50SVls5vNL43VS1WkkCGuYCOErZFfU8
L6GL3qRtyWHfIQaczgzVYue+Qd4383yPFBP9O9AnlaZCo7/dzUYJHa71yQM2e2kdzsGqrEZ/Xh2H
wMHE3KsqelRU90MoHab77L8Y/MuNxu25UAGsWsF/nv1WMtWrD4Patnzc8QHWxNPF/OhUpAbnhFAF
xFmHpaofNFqKN5UepC2I+L9TF+6H4bvM9TWGqkq09LaxH1jAAG3PnNmuVOBZVxZmJF4rceTIGhoS
JEeHP5i57JRMr6k/NcY22nZaJf1gENjCGSQpY5VvD4A5s2x0opeysMMiJbiKHt+J8VjsZWCTlXvz
PIi0cua46UCRuqq+NAPXOc3nvcVRxj6fdH9n0llN3TU7hAhZkGyyuKTTgOJuy5/qv1j2coFp1a+8
iNfJ+SX2Wueu7Z7TfXOOh49COLX7X+pY43Jo6B7iVlmDf/FLh/vicIEprS7GYT963Z7LXNj5nFS4
aPIw4aNJ29HiflUaDYxzWxpfA8br4Ar323qct7jjF6fsmHGapvqufEMTgN7GXp9uJFJD+hC2etyt
3MZBb6kKJ3J6W4Wlx9W5+Io37PPoyIlyS1dQ29fJXDghrg3H1Maf/WtSA4hiOchKIVWbzZHbx9SV
V7aEMGRnaD+MXtdsTDLigqRHrfnqSlpwJtDfy0nSOXCgbIduXIQar0BNkCEUOikcVjOOEm0MqJTa
JpJAQXCw4auZVcHBlZJPqg6LEieECBjI6GC3fKf7VMq9ZY+4kKy0RjypyT15JEgPcBF2zc8KVksq
SkpA4+DhDcXOxl0WpjnLcYNKnqzuT5SLwOrdQ4UZ8llSQeNNQ1xNwZuwsspvhNOHvB0Xzixgtqjo
YKtXWY63yP/STqK1Fk5MBGKnMKn9fkA+AD2/WeQ/g54HJHtXYio+zMucI65+7vFPjGe6HH9iC1aY
/NatFfzLncyA8QKfcpgneC9BBqMlmWhf4kdgoDV4uAK3v5r2qdcVayFdyeiuS0QgUpUkUwTZi5dR
NYQRhOUnMoBp8BfgS3v2JjHmy8yhICFaHCRqePfNLPqYci2oseIoojcqr/1z+LhMqsRL9kC0hTUJ
iXvHci+d4H33sZz9Qyif3UbHXP8AJ9hzVltTtrO+XDqkJi4idENRuSOuVFtdAtUmnOciP8VfPUiX
vUNQbnxO3TPJGNRpHAkz9M7cl11pq8zECgcw2Bl8Y+s+ePR9GC1XyV7DoYMDHkntOI56oEVurCw2
x/OHV816YGSxh2IIKBhvIlKwppBYchOZoSN8DTktI5eTrqSWvpe8pme2ndSIEY3ou8cMj66gavTd
0208OHqiN4spt0C7bPUwxFUkgD1ALnkc5RLjYOxBSep3cM4W9d2pmvdm9DWcR58wPgD21XACM3Oj
/EUTeu5D7RYZkUe0Z6iTyX2dI0xFOGY/CqCiizAzjFfzAMq1eKpzi0dBqGhiFlSlvm3shqRta4qz
bJ14PBnHT8IkjB7jmSLP1/unK64OwB+mEQuk7kZw331JhoBqaeg53r9nn83ySIoqeqQklrXAulXc
N+Aqkkju6jHZtQRIajlZT7q+76cMW5mCtQQPce2gbeRrKgnkB5JGSqimUp68MKGSVqcY/JoCHDvL
W0mIPUmRTFFG708DLG9wFDLGQDlxbVdssTQQL7GFcmKesmFYjtpDXxb0JC0p2tx0b6goBTrgnnhR
V7mDsweeOlcZnupbPuUoJAG0sqimFWofyniJ6Np+AjDY6RwPsM5oSrP+2sLw48qnkL/ixdkq3udz
cIO/jzNuXcLnTDZchl4qoBoPDb0q7XNC0IcUGs8HRH/ZSjb7qI5UvE2PwTbLqQtw78MOYcPVO3iE
jJBWfT5ZWpF10nWJfHSR4Dk5LsdS+pri4IbMbhvBIO9IAw00AiuA8Q4DY+JKOuE3FLDHqxpxYGUd
GwOsWRwiOPNqLNJUWDjvf/esYCwS78JCW3oX/IFaYcI3iMLp8oZ9xpSCpyI1G/JNJia/2iG8sb5G
riIQbcGRAjAkai0v/gpKyl/P1vkDfhLplRPs7ID6Jv0R+FOtPnZ4x5dkwumqas6aH13xm48Rwbb7
ZD/GjAVXrOH5lWFrCgE4m69+OT9QhsIWEkByIGTEA18jHOsWRFaoF9/0vsWvQYrUdf0ZFWFNfxK+
LnJNRgY8enjzlAUU60zniktis76aAHJoY2hdQu16GGsiioZWBiygWd3HfB/mw1BmyeJvY+2Qb+aB
/kRPeJI1cPnwmP0I3/H/+rtznidC2lZSfvsbGA+kcfiPFfhz+8v87SHcnk48DHjRpu5D8J2wuBrJ
uN/S6wEAIwmSirNmjvyiQIJxPZiwhrxMP3BvfhL8TI/pdZQkS3tdad6Jt9arqv3+v2Ljd3iaKiNz
jHgs3hzG5Mnl5h4qiGAnSYAKRmzFi3BVdUVq9Z0kQWJ+qpNcI6LEUmNiD9T30RNit/BYrY2lmmM1
lJwyqqo8p7/I8JFS2YENygAwYwNPcyPVE4LoLHBF7/INMap6HeVNIsNvbOnPqHker2YkEDaroUMS
JcotxI/31rsxT2JfwGPzmnxgDMp4RTeXFkrD9xgrTLK+69YAq+Zjfm8TA2hsCXvpiuy9LYzLXNHe
u+yucOYMOTMIClG/1ors/hW16/t9p7JBh2AN488xFDXvVkWZYenq1I5wNh3c8IozQZQxQGEEQkAL
8MQF87GrbXi2GyfRsneol4N+L2BKLm3T4uP44n/QhPSEpT2FT8p88c49gJK3TjhfHuWlMS7qQzj7
i9QP7p5ohYOdliednYzIt8S+bQGAz5+L0MUop/pEDi/eOt8UihLtQxgyFp2MvPOZxRtas5kBj/ZJ
G322tni5Ir+MGFPV5FaQ94SZXqXDNDJlIRKxfwpqoz6Z37cby/DYb+nVgG5HQBKkRAUYRcwJZCjp
B7I+kWRwDRqiCNi0a39bfmjlDjNcQWtZxSfAKmUxJqG3N3tQR45y7QSa+wCdNGoktSQt0tRcAvXp
R58LpchQ3RVvSpf3TWcv7noq5slwowBTm3Kj2ENlT3NA2z5oyV0SJa98oq3CBec3NhOrcHdQ+LBI
uZUJFkQk49H7iX9IGkfa1ldWRJdGq8owBQTio8XKZuxhds1/GFOzy7rAR2nVf0xHQo81A1TU3NBi
qNeoh0T5+LPy0KPs+mQTsKFEFdpmM8Cq27fmR9Ns681D/hDdISdSyHbaOjQkaL79PQwqE18+3Mff
crZLFFqNMBKtOvLHyvDq4Lj1IfQWbEfrZIcc0K4B8fHZTEHLx65RQuZh7CwCP/TgqwChaJuIUEZD
MGOqyIbmn6cnDWw/CfevI8djiamPVWkk8XhQbQ//xIF/OO4fPe4LnfWsnUxJmVB/2c8bsOZWkHh/
IjButqAl/kQB6/C/w24kFyRiHp0yaNUA4dAus+N5pR0jM6LzVVGB+ZGdjqdvsBfs++l4dZz1Uwrw
V38kTpC2g8hMkt3PdwaJzSTgkmgGt87BXxHxviubxTOr0yVqCexcrCqMVw+qu4ObFOoSsuFq2aTz
r144/baYjDOIVtrZt5ZEO/tLt6lVCYMoQI2AJZS5Q+xRAYbGwfqmDG50Qf4PBbSyRR6acpafYerJ
mHLA/5ao0wDNMeAZ/t+FBEF5Y5VVAmVyT2KqrbzNqeYtZuvOix9ClOJWYINAliwqLjbnPeGQh85t
CFEiRyMnAsWKM2FXBRWW0QO4FdzIULyoxVAh6WeWpSKFjQj2bZXnVhhUIOBgqnGmg60fwe557b08
vXwPlQJdhJpd4Oc+d08ngyGuQw==
`pragma protect end_protected
