// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
l7iaFCv7xTh3qvSYRtNxifqrCfp9QgyHWoVrpnW2qnaa9prxRCGet8wiKa1g9lh0
T7ZFbBiJn3p02A4JdUwhCGm00BWVoYefI+KwvwB0zRLE2r4vfa83V6yWgTJBBO6E
rqkJ7ztZ3eDHKoQR5u5cg3Pa5+Liq5K3HXaQum9ckf4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5840)
kHSXnuSxzrPty3p4WYWkbWmsk+JrmrF+8TnvnQOGoPTwMskcvcYq5kcElP7t3wI1
quLVnYVWWxZcOfpTDsGEQs+qdvwR6ULfZGEejVwzyOLsm33K5fYM35CBJpr9uiKg
SIIwjNxHEkAZ4MQFeuXUeMOMkRP7CP8otvx09s5uZZIjiFx743vwUJ0A+OHyAi6O
Cvx3c6C+BDO+M7thAGDlSCWA1wciYGwqiIR1S5tzww9MGmJxE0qjmybktC+vr+Yv
Ohf3fwea5umBn9hP+LI8P/S1eCmiQNxMAbW/UJHqgQ0IFIZyQIc9sHKIJgIkZscH
RRH5M2xH0ldwnS2A3A/oBOmq12k326ECfgT2v8FA/lvn7NEfIn54zIvtghhDlgsv
U1NcO/6O2GwRUjHlhn35ygNLxDPrsKin1zyJGGW1IL9mRCyL/is36EZG0dSFvurX
sUdJTzbhdsFeGnf2rvWSGZ/2NwywaXO9bwQuKh7eATH5OoOZgQvT+pftC7l3n5lb
IFSO4R8VPAFY8QxbTnQoJDaCVUzxnEITDl0G6kEfJCiQoGd75vH9j29jDTNz2l5M
VVrkVAesjZB909ue4OPjuhITa1mzgEJwtL6aBXJLzq4RrUNwSNp+5yu6I0QGcfjR
5BxvtwXe6THpgCBbkdg+rVwcfumlzwaEVzA1CaHIrMxSPd6V5dTq+WVVm4PXu9yF
qp/Y89Ztc5Y78t2K6BEKDYYKwQE/uRGbGYqoHZXts5JTdrwc9U7nRaMHBUzGYZbh
vJY27Xi8gvN36bcu37hHIFarV4a4xb9vGm0jKlXGeqUBEebNogNNhiqAukjAI0t7
LvmuQbrfUE05B1uKHvZJUVY72pqMlTZyeyddfVaFPAFKW3Sq7+HRErx/+BZIVV3f
0BIIZ3ALecTFLSqgaFHmilFAUxpVenGhFvk5irK5q/CVDBhPb9jmhThz4f9m83sz
wExPMpCtHcmQ3HWI3LLJZbnMLAuXh+xhbBVaF/c0AlKtK/8R0/AkdRgD9w+ICbAu
3CoFo9p2btb33cElqS1lljO1tKxFoMVs/A6b2SCBfnsKzCObTnX0XzbEITZJ0fbT
wXxfdm/DwojyiGF6Nli1G4p1VzAPhumsMTPns7rm2OYwSCnErskYRs7b8Smtl40F
CjWSh1/DpegbyophQPAehC92Alb6wucwlLUP0pkR6pk+olAVKytMqWakCf1dYgdd
v+htsuO4Ryd4g/kpH1lC2/yFxDWGpmxADwEvWZtQwirMAQXWul2g3yVgntOEoQCp
pTWe7lHeuyO1NFXfNY2yH1dYEY/TRrZZrgSmX8C5MBNp1a/B4lUBkO13QvIkYyhc
sFht+g9rW6CuYwuD4+5Q52kDZGhW+TIdYM1kYdVV3KNKGXLfNcF1bAfJwZ6si8NK
PDLqVVTSDMVuryCOGUyubYdiUpuQmAkLl/W3Y8GT0hbwcHSn8B8xoLdUE2sRoLuU
7pcMaeDL62oFT1XKDwsgLOrRKEJHhQRgxoMNnRWfDDw3UuWfNdZNYYgyOBllxAH2
f+D/9yf3+g7RTY5Ul67LbU+K6gIXRcA8A/SZkiBAQjMNI1FtU2si7IbBbHjdUVx3
6/3OMMvKHew2oR2CDSp5HU9EpnRIcmDpGOVQ6mECfU5mDindBeUT0/FFM1PtYKmT
gv5dK2ir4/Slk+px3QMg96da0cmWsK4oNl+njlLVk3XlbmcND0ZskXZAn9/4eNMM
iwEgx7zw84BH9KpkMkVYbijwyWULC3fF+6mOsoUMG07DQ95PQEikDtrhMidztiPp
sShBTA0+ABU3Ui9xKwsgnoiH0SrrJYb3gQicYZlmQoCvJdK0Srx+xLuy/ivDeTvj
kbSmyvb3MCUpvjpbIPEcwf8dOCNoA0szBJFQM76m9mPJien+yYPw3+JUrclXuQ+Y
IpY+lIKkNaiMvaZiwl4lB1Eq8VK6XP/e2KvPZbUdZWFaDxV2z6vN9WT8K2WbipOi
Y6nwkxtajiHsLoXXI6gtPuJFJ7jH6mJg9TsO1cDXydeFKTdMoY/Pplt7/ItiFWXn
7FMHt4byoo+2vFy1h6B0UqFQtxarj3ADn/3CmXTQ/EMXOtz4ppMSZMLgQzo0tRdT
fUoD+QCfHw4wPu4Fg4YO8neyhD96cUFY/o0jxj16+VTsEslFVGydPzNzEKtyGbwd
i5y5a1cOzRidiFvQE2O5XfBRqtBv3qaMQNA4GD6lWfFSf77JFF02rRXpFjnVy/BB
pFlBH/P9G/UB2CY/u66l/Id1AtikwmhO2BBt/pK0tm+tPnbChWTRnu5tmbxhyzr7
OangvJKnbEm9tC8cAzR7XZ0bQR6++fgbDf724MiK405LmDRzUDKBhnp612wHrCGl
Ehn/VR+baMkdnOuYwZAdPnes4bd/X+yU1biSMZqun01TDwpVcMsNxVQmvFXvHShI
5xSom9LVr3qv0mL/ZjqHWRyl/JLiitac9OYQYpWaP1EUmaJNB/aahqD5Pk4ZQwlq
w2nO080To8eSVvI02IyR/AWPPcFFON/POlWp3ooXBuKjIgfTyE0NPCCpdSo34hD3
1+3DbPggKUO28Re0v5eq2GC+gM74ZLHyPVE1j0JFciqXXlbiaixh0pVn+KmZhu+D
6TvdVsx7TnTRKOozB/WYdtQi9WDc7fwrV/VJs09J1Mkbb6I+pvAG6saMmReHhBFr
00+5C7HfixCx+r1/IWmeB8+nh3qZ1yfB0g/sIDBWiHy5OG8a1Ly+yA8CDKJtx0dH
dbhW8FoPwjypVdhXlZNIeLhh3u8CZSSckQPHil2iE1qGdmciKOaNq0o/B7eeRHN+
wwsI47U00/4/nNJvbtuomutrEqyl4h8se0cmhQUCvppRiktyAm4POhwIbTZCiLgP
pi5zh4rbbGZ3IlaLKN89iiSluTysTpoD9uvX7m04AmueqqLu6/odEXbJAnm/yFrx
wyLVrGW2HaH7RP316uYh28pFi4yVCADyBf1OerAAXB3lyQUOd4kBKNOW+EbMCUl9
mc/YJUqwl761C2b2STrmxh2hGSAs6QMNjg65Tf4OzRmohRJQJoZruQLa9HygfReN
wsZ8/zfJFRpBfduKzEutB7kBOy+ylD0kUvfpptXGlFZHsg711CXCmFtOvDlHiEls
eoxxoTSBxIsSPnFTKiZOzUt/hpXIOB3Su2goldy/3g9quWlKQNP81uaBEUQMylWO
xyBYBzBw7SYsHha3GkTqnFPMZ4O1LWhS0x3EBugxWRp6ZWbapmx/6AEHceuPBIHG
fDDGaQRCq18LLkG2GJUaK6ain4+6SnqHC5M44VA43j1EcJ9OdVQtEfYMrlioW3CE
BK+/aA1/xmfj6K22Sh+M7h9Zt7Ul1rKDSls8z0FsIeQDDTbMBRQotir/TKX7CLG+
KQV+SgXxU6+BKMZlgHbeT0hrdTDrSZEwDh4YET52t3RJmg/uOKkvAK1aTHaKIWAL
IqndOMfFrLQCEBHdFtY8MiUCB8VwVo+jlYSqhVptKQBrRuab8W+yfuoAZWDhm1YG
GL2c4KRHRWF/VO74CiKAhvlEGDl7Sr68M1jB1gwqQUXVJL+zfrlaX+75jpeDehfJ
mVBvcwNkgT8fvEy5m6p2flhSElmkvMRd3e0rWfEN7pEPvV4s7LHivsHsw7rpFoj2
jzAGJYi+dkOlCbjC7TrTb0V+YFaBCbyEK8NNDzvtoKRbd4+siOlv8LhEO760Nj8Z
DzJgeGiPOHtCG9PlykxR2uq4PXHObBDYO4plTEbHhgeamqAQTacunfFoHoCdSVLq
KnKc92gqyDoyvB2UGytEUFhVAtTo/TFPydXwpATFYtQBR8XeLYrFzZlbW8EQU4Iz
maXEQ1dk3mvwstqBkeu+XzigX8v/aBwoV4L008pM/IbcZ/y6sM68njI6+Eq8j8ZJ
H41IsXgXOJR+oi229bjL/JHSf5bALu3+xStWjAJIb2fKWR9LW7E4RYB5jvlAsAAR
b8W8gDdw6eNUyMuhj+rytQH9XthIQdIBLnE/DZyVbxEK6mb1Ivdzl90tiYBDNek3
mvorp9Jn2v1MVWRo0wPzfbDtTet/aT3y8Pkbg4CsXXMGJxIPHpqR0pFn0JlNMuHg
c76bqla0JCtlR+tdMPFHxXdWred3cymP9XYO2OLndkNThxjhbDf0g5RrowN4W/zf
h8azMkZswa6cKZ84oP2KNmdOtqdJLWwWxPLaAd+jPI3okEXSJCNsi12aaMT6aiW3
5AV9uLWorUCarKSTYAASa66EgU/Fo3DBKRhueycwiqF65iRZ9KOst4HPXm6NX8UH
JvhwWQ+Edeo2yfPDZQ7NQcG+x9TJSVmx8daDNSOk7DQ9bfXOSLqRJYUBK6N/EeAR
GmAH7FMBQGU1uifEVC4BmYlvxt6ec+emQnOMGZNtEJd5/01noqTWzGS3nHxzz1nE
VllbijEeGS2NTpYD8ue8JzX1cyxUc7u3ubGmwMnTXx3162XwPkqT6pbCmbWEOKeG
GIWKhDWY3QgsbQhJFGLKw/SKe2Q88hckf1V+jUbUB7GNm2Go0ws8ypm1ySVNJH8b
pLDdLl2lommtx7YX9CwsBY4m8cEBboQkEWvegQWLoYY9ydXBe6TW0K9JfBVbmZ0M
HcKVCEPPzaaBFw3lCfC/4UVBKado9m1UpqIRDhTBpBYtTQQpwJ/qdcUZBGaDq08o
xWNdp2zXenMBEiUbfamDPayHkBRJrRfbHOZxKKzM0skZGrgt0me6/r96K+4NMtQU
TqDxpAoxYiAHuJJ/on0AFmbJsPC+YIc7cZuAUMBP2dHWuX2zj1SDoTa4EKgB1ypj
RbeoCjjCLA6dFun9rUCDLlDkxzyF8MxQu1Jy7fwv/ckw7SoavkkBnzzMGeWaqekg
cYrNAkF/QYbmmCas06WQ7ydcyFst56gxj1KOCHWo9ufN8zl03ve5NVpGzdTsPNCd
NvbBBjhtZ9EipyluHt3lWNzgg2huQsW/HqzMJ3H5I0apBhzTMADeZMe22s4cv1Fc
X1nBY3wflaHgG70vneJXaT6KKOd9+BkDOMgnm0O+AhjlnUxwNL8Jfpp37q0aeIE7
RrN/YElEpq9wLi0O2FqHjpyRdDel2VOEveojEnhDTadyC2G9mQtC82TcU3X2y+HY
2DJbXUiRaOh7UMfD2vNe0BhL3OLoTwgTDkIFfKLWlblS3xgHvcsyvTT4myCiteZ9
BDWBtgaPHXPeU72zwP6k13Q1nFjKwrdLx5YFksoIMwahrc9ykW38OP3/4jAHYdib
VrnhtZbdptpOl0N2X43EJ8twPap+Wc+ijcRFM4CrHWD4pOW2XlSdsfIyhBUSbSaW
PNDrSG3AyV7DfjdZorXQ35aULTCPVhZUrlLY6wpGLdTcmsCFrQZdi8TeoUs35USH
ZY+5r1hYo4lXMn+tYfF7F+ptFQICwrKOF+dkiMwayOOQCTxMjAgwJQ/mON/keEou
LoPoGML15n429B2miZSOHp9GiF+C+LKxesQqLRA1lN86Mxg38wlNyyImwYmOaMhf
J/ARmgXEpNppYW9SGytGVJCgkaKkRRxBlXxaXu+59V2ysZUL6qNGUdTdWD0LOmiR
/TN3ngGU+r6qsFaLYLPnkom5gj74d+h8BwYwKl+d7dBJsE+Oa7xbvuXJxp11AuU1
YG/bE7vixQ4q4ASVs3DOI3h/BCuZOyTn1RY+SLDiXAixn+qhnmEU+fNPvPO1Ddv6
uaopm1RoSrXgLa+05qTBS8j417q3W6Im6VxHS7u2mA0SEd3lfZ1mOKq66+WPBbkh
qvc0kzQftUX4xxYMTGIdEN9dUK/72vG3JABm0rvF9OCKN0o2ZPpJ5IuB9e7XlFSq
xheVjAADiOu3Nf++/haEa/ildukcyGylJuQdOsDowiBPPi4SCEBt+RT/iVloFWUX
4rTfQkPLCaoFBXz04KCik2IUIL25fS6YrIBbMIfFlC8Hez08cdnRka7cr7Z8e1Vj
bedaLxs92Fmkpd7eqN3tUzXQ0xEFlHscK4xRG8xktxo1YZeGvTfu6CuOXUQ/z4IT
2G4eKreFQB8A9bgqUDpJnDDZ5gFmcM1XA4RsAcHV+rFj+gEamrIShiX3xFTiaNSA
UlCBJ3THd1EllxN3VNejMX5rC4L1vLAVJJlcxOZ2UYyTcA3L2ie86tLPE/o6CkY9
6vkf19IYt1yuUnIoHQTk72WlflTDbcdqPKc7N0L0f/pk9nKgxe2yUH/inTOhxjKD
hzwQu+mmCDoRpfxov8wiBd3acfodBLQjxHPOvKZwXH0kiGJIh5m/cxVfaY+fJv5h
kpFPNGeClVhlX6gZsgoKBwNd3RzA/2We740cplxnBWIAVH36Rz6V5hTuhIg3EaYa
7Y2xMxW+exdVLNZSfw1CT1dIek+0p+DKylDZQLb4XfRMs5JNJdZ5dZmj2l5bWYi7
tBpMD3OEISHZMMEVm++aizMy6v43YJZ7QU8BwAVe+PLyKjHMhah1FJn5r0dcp9n/
LDQrj7wK8+Cz9PduhgpFqLPJZzdSK9AN88LeUFjxqd3TvEeq7JCw8lcNCUT9Ig5r
bPHXZ7ryeT+2N29R9pJTz2uU0dvrbE6lJ4DD64hesBy1oXamXvAQ3hHzMYLuDv14
WFiZsmAPTAtsyd8hJ77BJJNKGK2kl4HcIjQZbtLecLvg2At5AE1hCH2oNVpatVIh
3wL4iW79NzmvmWB6wt6eLelzfE9eX6hGYxbi6EvfiaLh7gH+AfeSkbjrwo/gAmUh
mOT+k0w2W07D6qm/1/5r1+jl0TnkTInft5WuGKXSii4728OaceJDSa2/bSiarYlu
qNk+qr8IcmX+bGAP5zlvvPd9scjkOjtif0T1w+dJkJaM0gXXupex9woflB+NulD3
we08QQnNT8+XTY1LnrVDj6Izr4HfGy0wXpgziiaLLHNNqm+fMXUnITNevEWGJawM
QfiV/LZQaminNhuLUcG1lhr4/ziwYFpU9ALigABmeK4ha2kMa0D+F5e2V0MUOYZC
loBk89I3pqYgGXQ5fSBL5RxDHCISPePwBEVTVOAr1yeWMNVeeNyJsQC3Ze+fCr20
NS2t5XlWN/cSYP63R7k+XBPPERpSg39es6H7cESodsvuwHHKtM7dPlIf1Ul+rdMF
yYlxNbu4NE7PrslUUlqzey6nJWdOMTD/hSJ3I7CWMnacfwQzPvVU0EpH44xp+TRf
1G/8gZ4GdP+wHxZt0RnbRtFUIjby2F7nye4N4Um53Vh0a0ROF552EZKw1QlOwkuP
5IiV8H9ItLDISocNrBIqwZyau2VKX1Bg0i39xVaStjLsoqtUujdWB53jCw6n7f9A
ohf+hgaoSRFbHfajgctm+sfbtM//0LwJoA/htlljiR4yCFEKK4vrYzRAOAFQZ9Ci
fhpL0uvBH9QuGdU/RHyK4k1633vdghrft3K4gBzvHvq2KbRbQLWQZqRJBsBDu0Zg
Z5SupTnXSowoRc5QNq7kzi7GLXiHZTAmEQSK3KgJPF0sEFfhk3Xb1rdl8stoz0Cx
D1CEcJE+E9vYReDJX19N8GWwkllvFzWP/OPkSyd3QE20e3mVK8salWuU69Xm5kIg
Yakktr+gmwR3yWURtn6wNXVFdia2py3bPM5CKX7Mg8pPGFjLARfInL3skyi8SHJA
N/6QvG0XJD/ZZ6y1RaEORZkg+S9CaEBuFk80QVBikq2Q1DgmUJQNTOeveqxGSb9A
KXdwK1Fow6qgA1J3jEe6fCdzkRUA5uUvi95MB+FklUi3kuLjTydr3t/reYOETwq6
potsqZgtaJ89fGoij6+7CI9Zz+0FXJeI8vedZ5TKlB0=
`pragma protect end_protected
