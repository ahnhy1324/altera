��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���8*�"�Rϰ�NDSB�$�[�X�]�V?�y&V7翷V�e���$s8��5�IE�(}NU+i�O��҇^��<|@�AC;�%u��c�x݅���0>(���D�����EmX�(�����]�K���f����)l�P,
��d�"MX�� �=��	��n�ؾE�G,�c��%�w��9�v˹�r�6l[xs������Yrʶ��F�0�еk�x����;�~{���#���
pQ��Nmu��=
�;�`�K�_S�G�������T� ����^zRL�pˉ�D��c�t��T1yŖ|
�<.e�4U=�y�!!	{�A�@�Ҍ�,ET6S
al1m��sϽEDx�7�{���6n��4s��6�qş~,�t�4G�/��h��b��)G&�y�o�$���ݚ�� x�Ø"�V������+���@����}�=5n�t��h2���+�(�$�udsL팔�BBaLd��sv�o�Pz3#L���l :4)(��ګ�8��da)���I�UW���0�.�)��惌]+�#���ڴ-�s�%jկ�W�ŵ�7w��Jk!s�X�o�(Y�L��y�]��%e�%S(�"��O���V�1���<���5��0Q"��H`%��Q�~�Ʃ�Dw�)qP�V��ڧ�G��V�m�9y��]���9~���b}Ndz�����.qR�HX�܁P��EI���ݪ,w�9,Lw�C�P]���
�_D[�b����0��5������G��dϧ��Bv����]���$u��jO�1ЖV,ڢj*\�/��ݮ�R��HG�t6��2�6:�S��Z}e��#?�[�]�$��T/p	��i��#�at5_��kV�7�X�%.O�k}.Ż���"�����x�u!
�*�*����K�f��\ �<��nFɚ��f�.&V3�t�_z����RZ �UP'���I"���U�ϓЯK�݁/�G�5��#
/���R�|�1{���_����,$Gn���G�M�J]^e��Zd~;Rb��N>@���O:G��o�)��A�ڄN����z=$��TD|d�c")��8��|���T�k�Ҝ�u:�J� ��lHg��:2w���5I�5���R���cs���g�Xf����y ���@)����Y�GB�}��J���фQS�T+����;�}�ҧN���Q?�N�Y�[v��/&S�|,J?�x���=1~����@	�&�f�@6Tz1Z�p2����H�{��_�( �Ӏ�-�u	Y��ּ�.�;Erܔ��+�)$9����x���pǡQ�/T����)X�Z�{���W북_��w�@�,M�>�҉�>���y����J�n�uàU5X--��|�Ŀ�h|ݮ��N>��� ��F�S�"@9^��H��-D��h�Ep&j �X�U�����N	߃��N��0n ��Y�+J/���Q�4�P?�wV��QhU-g����+˲��Ry�i/IF�����%ɇ�gC��N�W��	��kZ Aa7�T}V"h����H}�L��2*ǲ]q���Y���,��btd��(��=cayLV񪼏C����#���4 ͅB����,؆)e�����|��A��m�C�(	�9R�����vܮ�h���r�(3����v�	�����5�j>t�I�&N��A8!"]��.K(��3�
�Eۚd'	��(�h�ݔmg�s����sۮ.@��`���Y��"��Y\��a8ZX}�����y))��2�'��E�g�w妀���PN�mfGB+ �5�8]欭n2~b�\h����e�Z+�{(����,<r���g�kہ\w�N@��S�3r�4d�z��D�-V� 2�K�z'��}�g�8����Jl����7��}��̆�^� ��t�<��3F�s�(v`��Y4{�S�9��|SM��; Rv��J�������/X>�`���p�f���W]I�f�ϋ�7[�9f�#ˎn��V�z�_�!��nwr�U�^���K8�習���.�-t�*�M�wai��Of�D��I��F�ȴk�5�/=~:!�ʒ���7���b�4�|��3��dqI D��7��Z@p,�Bl�}k5kˍR�_4Y��:q���`�@#�Îy�nf*VV�IϿ_p�h�ʳ{���;c�&~�']�ׂ�0g�|R0��}��tW�&�am-���˧XV �����9[�'/D�r�ݕl�?�t���Z�Q���z�^	�`k�Vn������^,8����`�Q�q�����b�\v#d��vM�M4���=���}�&^0�����4��pRp�ɁpR�g�pc�d�	sV[�,j��>1tO�Z/�=kF'JM��Oօ*gQ8J(��p�&�m';&���ɬ|���F�i�
Ǥ9�߹kCy��(��r���=B�Y*CT�
w�7�Gn�:~T<���'�*a5�aE0~,��V ���K�Yh; {4�D��Bouua}��R�қ3��"%w*���j��!�t�
3{B�!�
)�Mq��iEƍ��O���א�S�B��������p0�d?�bi4�0=:�'��p��j�"KFK��!+4��XH2ʏV��w*����z�!]E�z(�:��>D�UzsW��Q�"ܠ��c���ϖ1qUT� �4M��q=Uѿ i�����}�%��(^�����[�����E�փ�%3cnR9���1Q}���jNyR6U�*,�^��dd H�����4���1���sƎ�!�k!�\�A���]&��S�ء���@d�l<@�Z���Ԟ�@J�Vb b�%a��#�a�t���bUzࣕ��M ���mb1��5�<���JNq�� �T��SƧLV$3��Z��Sk9�'���]�ļ���s2����l�t#��wt�C�l�aqI��I�Axv��.�@=���#� �M����8���WF���u�Zou�opnP�y9�ū]���9,>Y��UZ��qY����K��XF7;�l��X�3T�OV������m����O�BwÞ���4c)ZLJ��8*y��:��歗��-��S 8BrR�<��A��h�VY[/$5�S�~�%�������R)���r�TC*�?�,�~�Yq�Jn����G�k
L�{֓�RG��;��;rྐv����dE5�ٓ�~�Q���k*�{�@��3�0�%������|;���}9&z��A&'�ـP"���`3�R-���׬�>�YG�ԨB�п���c���M��³O1���!�!�a�ܢ��.RuFRWr�na+v�`F �S�D�S\�1{�DI���	c����
d$2l�0��/�`x��p#j�p�[�9�x�Lf$���0H����~%!�*cC_���&��?ήL𛗾"�#o-�?U���ʊ�A�7��2����wq�3I�r���PG�S�V�S����`�)��آ�}��Yr����_^� \��Q&D��OfSf���[�V�� Sv��E���|%DR�.�HkKbb%�` �S΂3�Q��ܪ�:ꪦ.�7��>rG�=�����B�LF	ب����"� @��v|���Z��)�1 ��g���+ӓ�j!�̨� l�>(;[E���+{sn�qU�/#�5���R��&��iVRIW�StvYm�F/��+�n뱮�1�9�6����o�H0�J�s(���_���r8�0ҧ��X�4C���e���}m�7�_�#eU�(����K���"��ve�BGf�Դ0�ө>��R��%|����X.� ��8�]ZZihr�֎M���Qv�%8��2��_��{������c�b������Hw]�E���\sԯ���.e�X����o�ȝH�R�?n@J���ú��,��>��P�ArD�N�p��x���:���7õ/�����Я�bzu�j���k`�1\M�95	R��u�fb]��?��@��CL���m*��)!������ꗮ�(�9�OIa�{�!�iH��m2�)�-y3��O�O����Z���L�H�g�����ܩV}/YL�β7_���`EZե�J>�է�1��?�yo�1�]^�,8;6%�2�M��Oς�'b�[ɗ~�Y��� �
ԫ9�?��= ���:�����U������
�
����-�̴��L����؅۫D��k�����r3�6)���By:]r��T�H#������ʣ�g;����0�^���,�%o�g������&"�T�lFh9�B���E�t�����&�"���j���3N�!��p�Mq�9)��Z���9��o!����a8?��+�te�EF�;���65��/:֐{$q	�Nک<���2�:f��d�|P���|#�ݱ!5dG"��H�~�@mr��w��~?t�&�H��['�Y�b�!�ȓ�p��z��ZX��C�=�u͊�X����&����P�{���ض3W�0���	�2D�/Jq��M#�|ʛE&i*F�bQ��aԄo<q@��Z�,4��QFS5勇��Жw0��,V���yB;�Ĝ��_E�6�∃��ˣ�8j��8���K�¦���1(�����G��jH�����cC�oc�d�5��e����qfz�z��1������&E�*6&���kr������<����$]|��$���!4T���U����� 3�^y4f�tշW �zьtm�����ϝD���k.��y��9Y�O6�_���d�h�B�y����]��`�C�ƞ�r���Iv!�g&/�X~��:"�&� /$[������*�%�t(ou��$����@Ai�bW�<Bt�]~��i��v�B�G��o/�s���p�M�P�׎��o�Qz]��$�S�G��@����]��N�>���y����}t�R�9�{��k~������˕���Pl� s�n�{�	�	^1����mb:��2ɛHj��t>��o��ײ�=bǦx������HA�TPY�aְ��Y�D������:{��DA-�36p	$��AwΘ[Q�}�5Y�(�n�qAk���H��x��!��Ţj��bd�(}"�t�_�G�9��v�N�jpt0���g�����Xd&����G+��slgnkL��6r����)r�TV�E�V^ ��� ��4F����toZ>��݋��]��f�ko����4@L%���E���O-�Я��㏝7������%@pA-��w���LS����'"�&�H�
�EƚJCf��VF]0J��D����N����k��`K��o�)�oJN�7!�2H7��*
<w�֏)��j;7Z��ڞrqZ�`��^�KdѠA/+�Ld�*�4�(w=kB�c�?�љLN�3 PD���vx�Y%;�!X�d�7A<?P�����i�'I��"�����3�?Ӟ$�(�8imָ>w�jܤx�!l���7YP��TLE#�e���E�(6$p�J~{�bbvG�}06 � fŇ9��A�(���Z��4����ߴ�%%?!L�0J�ኳ�Ak�C����I�L�v�r�L�0�I��U�g�<�q_�����4����	���M�}�7P�y�;�1@��Hajp"<[\u�������m4�'�� vuںDӅ��� �ɓ���֎lv�)?��A^Q֠�!�ְّʭ��mŎ��i�䴵���zl�����rz���T�"�v����s�u������8!9�|@�o.�T�T��x������:��$��S��hTړu��ъS[�"���+��ly��!`jx��ʘ`�ז�pѿS')�h��ݼn�=;"eUu}�+t���|�Kz~�<
���-_��ų��3w�����X?��ƽ����ڷ0ƽ�U�3��$
�� c�o���P��"O2����k�(l�חpR|�?�$����]�ʩN�a�n�K��X*b�H;�]C�;�G�_�A髨���ǽ�����,�-'ay�:�H��;�����ޡ�B`�'�hU�|�4���oi���v�-�tϼZ�p����a-�3�yg���/U�W�Ic��&��J8���\�ʭ%�ĺ�<S$�$��Ԍg�!�^��Ml� (�w�]����M��J�,"���S�m���f�ɶmA�)b9 ��:��CҀۅ��g.",O��뀷��G�0n���i��er-8iL]=1���Tז���˖����e��J���`���we��i}�W�wʬ]��
���u�Dp��-��W�j�A�Q��������M����;���-���(�G3�UݎFr���[|�@A���v�zk�Ai�\fM�n�e�I�.��d���9ZX����[zz��B��v���*Py���2z�|꛸>'Z�4����֙!����g��z/
aCb��RJ��B���7�����a�����?�����t� ��Q
�C�0�;C���@��"h����FM���~0�Ӏ�~�;6�_mL�?>�}�����ƽ0��&�q�g��7�F�B[M���}t��AH-�"!1�[L)��q����	�:?��m��~AW�E4'<N�c6`�f6������ޯ��}�[��ށR���䊣��P^�YMJ���������碙_N�*�L�ȉ�r�cGRT��PMZ�_��EU�I�n���#t����� �mɺ�l|}$rṇ��5�V
�D�r��?gLl@=WY��7�sAW��IǴakئP�X��1���:�Gj� �,�GQ���p	:����:���C1�==�5+[Q������
�*�.�'̙�N�%%4���#b�����4э]�U8��À$0aV����nv�!�2R��ǩ���TU���w����I��)8�X�@��p��+ �F�~�-j��+S��uE {HȄ&b���R�|H����&��1��nݬߩI==��;����C��QD�<p�@���rQa��2��"/��n�|Ƥ�Yz����$�{*GA�E�xU�Γq�q�q1sN1���sr�E_r=�Е İfP:���e���T\��Q��>_�L?�דRr2_܁;n���U�D���8x�,)�b�v�cG����f�|�����I������.�|�,���yA�&fG��.���NO V���Z�j�藺f'���T0S�"j��M�T�F���3�p��<�d�t�x�@oGc���G~q�)\W��<H���RPW\�|WwP,
��dj�b��*���CP֍�H"��;�St|��]�R���K]^}9�.J��v�8ILAy}v)A~���(p(�TQy�܌�73ԏ)��,!E��}q��R�E���D�h?k�yYp�X8�i[���������A�Y�����,�;ƮJ  65�d�g�����#���0O�x�FX��=H����TNrhC,��ɱ��4���sz���_�_p��-��+4�/%9l�S7�KX���Px毂�����K	���
E�=�$�#}�q\�k5�� ���3�.a�m��P^I�1��w�=+Vcv#
��N<�o��E�o
�y�Ia�hmñQ(��_����Wk���h��r%�B�Hp[W2)��:o�!̢�fT�8��,��;`�ql�W����E��xI���s�K���֫�L���O'5�0�(����^�������+au���݀zw�L�S�-c����_��骦��*�t���,�>m{���`@�[�L-�i^$��~�^�l���z;�	�s�pͣaDG��G��da�ʨE�],��e��W�%�������M��N]������c|�)ouQ-B�Z��$~��3���'��U�S?qR�#��O�@ݗ�GSv�v$��=r,ب�uy��ӏ#��$� {���z�]A����힐K�
WN\}1�|�HSK��"��� �S�����z���1>%����t�(ge��IMJ�
)5��V�܀����yGM�b�2���ƶ�"-��<���9��:{��H�����Y�B�u�L�)�l�7d��u�M�j#'kYc@a�����F4�$���?yς����|,�i`�`�V��{%X��ִ�l�;�a�w��� F	VJV����:�F��\���2����؆�XE��S�=��ڲu��K�_c�Gd�:�sCҔ@Մ��F�=^��)���5����Ow�.��,o�s��n�ܖp�M��eir���9!r4>x�O.�)��C�����d��iG�v�]�/y��n�ЇU\:b��[�w��mj
��}���ۖ��`� ����= ������v_(�NNn���R~\z7����x>�!ǘ���盱�5�g�mj�6����{�뵪�ē�;=0���x��:�OLQqG��8��uc��Z.,>?:�à^0~��s���P�9�9��"k	�Q�3�LY����&�1��=���G3`6z��پ��z@�V��-��Vm����ckA}��N�n������������Hj<nZ3�\�����-rx�u�����b��m�AXg�h��i��g��S���i�)*��zo�r�Wǵ��,�Ny+Y n\C�9��4�ǐ��ҐT�
�Ԓ����(�\7�q��ʙv0o����K�c ���sl�&z�@�-�� �M�Ta2� l�_�)JW���Pu>�{�a����i�jsO���Ng۬n�����W'Y�'W�W�4�Z����~;@��#������M>�=���V�'�#k��NT�d�ɄG��yK&��.��Ͱ�_�?�Zyգ��lU�tW߫�p{��k�t�*]�bH(�����3:^W�~:��5�y�^�y
y���.�ُ���:�	�u7�E��G�����QK�#'-�պ��1�|���kl���������|������Q%2�)OEDh�����G�}�����gP��Z�=h�y�Ӂ�AJ�'=�c�X�n�+��������� ۽
��2�V8kNt��"j�Ҽw��7wP�Q+6VTq�9�
ç�%�[,@���=Q�p޴x!�KK�K?�8��V�}A�U8F3��ف0�M&�\	�/����2[����1/���X�u�d�����"�V��*���}Gв����wy�)��\:�ˀ��OH����0C���H�~#5.���,�| ����wFt�~��ב�hM��~:��4�!��xs���O-�c.�H�|!w�B�q��7M�T<N�ţ۱+hWZ3
�R���Qf��TL:�V���$�/�J0Ȥ��%��+-6��O���@�;-F�o�)�����`s�x?&Oֲ����B�(,�锘5y����}�+���-x��/l��	�Fw+�������.�Ї�y�`�Ç�n�[��?�Q����rt��y��AJ�;"���/�r���x�r��ֿy/�%�J�_<�H�\��Yx%{�=M��j)�G�aџ4�a��h����_��t�䅌^��_�3���|[[�C�U@UZG�����&Ϗ0"��0��v��{��똔ד�S��ښ1l��(��M~����/@ۼ�߬�I��M_Q��t�Q��`�$�S��%��V(��K�X(T�dm���5�$�O*Qw��Z��tө�1�F�>�����*.�������(YT;�J!d͎L�X.?�y
*Z��sN��j;qa��3��$�)/� ��y�/:F2�#�K��O0IEt�Ǻy��pl	�j"`Z�n���
�`�A"�b2K0uL�7(b�6������j��큲c�u�+T#���yr~�u]�Ki�EU���Xp���[���N���И"#�VEahi���Ǜ��j��0G���6sn�(�*ϲ���#���f݃7�cY�,Ջ����uE>�I�[�J���nv@L�ǐ��:���M�"�#s
��+Hܴe!J��G �G�7R�{��7���O.�IHMc���m/[I��,�`��������VW�c�S~�=={��Dr�/��ҧ�t_�|M�9(qpB߾^-+�v�\�nhN�=�v�cl�s ~�h����G#�^�2hvc79F�0ABM���=$o�FǦv��&���z~)��Q�����!�ٶ%�jSk��1����������V�#2�P���~T�A<G���6��{�d�#���11s�s)P��3�8?bJH�y��r쉰��nb���Da�F�G�7��A�mf����?��[��w{��c�y��^Y]m(C`��!����1���D��BR�y�����ۙ_hj���Q�6
�eU{	��S��H��U�b�=�-��	��q������ݙ�L�P4�ٶ+N�Ƚ�����dZ*�I�b-�@����ӝ_��Ԃ�Sk(�){��x3u�A�������`���xYF�%gi��q�B�U�OK尌e^���JA���#ЮU!�	����_��rc�[V6�c,�ݶ�"@��1�E��h&�-�]U��v����Vn@���{\cB���Q{�^�����2�%*�t�Zm�v�G�����#T���#�ho�3����"|f�0E;9<F��<�E��D��xRﺻ!l�O�0Z�K�s����&��>��� �M�ڻǟT� �oŢ@� ed;�����BM�_5��ݻТ����L�Ǡ�L�v�D��;l@��G�]�#�?+<�8Mᓎ�F��'!KL*������2�Яp::��E�:�N>�Bd2t������\���,�FVT�@;��Fl�<��~pLG&�j-U�62��,�����o��.�w��U�&��4C�g%�S-9�9+���r��%j�(��OV���R�/�k,,m�{Pm���� ��&�b������ي5�N,;��y��D�- ��l�S�_\a���H��
G=V�t������1���
�j��w�6^��++(�\O�'"\d��Khߚ04����ǻY�w�`�'�3��W�]���vH\��D�qXwd�^th��s�C��Z��*�T�����d�RA�-�c�ppI���3CoK3�|=,��Q��评59��������	�)����������Mۛ��'7�/��hW�n�!��E�

)��ˡG^q2�bƛ�P֨�g�^�v|�G=B�`?̤]�mZ7���fA��O&�{��VOcNc�c`�����x����v��8���ǥMM��!%P���ö
a$	�{ݸ������7���k3��A��pj�F��cՇ+\�Z�ܿ6�M��MS?��ĵ�>!�s�[K��P��UvOV\�W���[,��/��b�͋�9��K͙���wߖD����xT��T�,0W�\�F~���dF��-��T�[���RA�e����ʳ+�b k��E_�pKF�6c�`_�X��c����fV�[ז�㡫���0�|�^Щ*�_!jt�X�K�4��z�u~�_g{D\P�7R)��h��$�WMN��.�&SmT����n'B����%7Eh�ҵ$­�/��3��̆���`�T�K����8�l(.�,��xޏ�1z~.T���?���K6�q�4U �a��Ρ��Nj<��;$�Le�4H���~.A���AY[c҃FJ�?Q��sIQ
�<�؁���,6��Fu��;�Y#}C�Y�H\I3�at�G$����jHJͭ�f��wXs�y���.�����S�������(�;��'WsUB
�f"�!$�;�t���E� o����v��v�9r��s�U��A�^^+.>�n�d���!��,�ص�/�fv�A��ʳ���#+ˡ�����v!!���Sy���8��*�/��I����������0�J��om�l���5���e��+�^,(�'���$�Ӧ$4�����g�}k<���N��:B�n����H�S"*o�0�D��8��Lމ��e-��Eg�CT��+V��R`�T�C}dEvy=7\�8��oE��IY�X���n�f����u&�}���Z�pcL���5iR�d-���f�je$Wm�T@8�+�R�໹�'���4�#��#�
L��a���ŷ�������5�r��W�υj~��[$�b�`#��C8���8"[��tPY�	�􅔮����k�Hҕ�W*kk\��Cb�,)��p��BK\�$^�T�ܧ����B���v��A���B����Ȭ��a����"teu�(���\�(\��izz,|"0����z) �hƖ��p}Չ�U&5�?�;��H� �w�>v��/�AoV@=�f�\]��m�;�!�;U�4�ְ�5d�$򩨫Br�r��x��ApN�~8�?#WB�9���Q��>��(NLqBw�ڙ���m+�?;�/���~��f��S49�}�i4��m�/*��A(xEȤ6BQ���!r��
�b��o�u���cA�%��T"�w!~���,l�zZ���u6Y�1?��^��ơ�\٤x����a����[MFCa mMW'�����-A�Z��u���d~}guׇ�,�*W��!���;�Pr���~b�����z�_O:����g-�\ j� �95i����F��� �a0|N�|�J��j�]R��M�ĸ1����q��m�D N����]� �0��� qC&Y�<����_�#��"���i1<�2��/F��[�Dǲ�%�u�Gȭꃯ�Mm��:$"����v?�~�c�h��|�h<;�j�4B��S�b�itj���I�m�o�NX"���&��$�o\�(c]����,����� �����Y�߬��{�M.JZH6Z�@1`��ő��J^�l�0��h��ˆ��>���bX���d�,m K�,�D\ �Tr�]��b��f�����\���H���,�/%���#��n[1xr1~|��t��]֘)S���T�u*-Ov�}��!>��jd�%�d ��3�����6��Ũ,�FI�J����LJX���h�K�_	��;[�w{�<�D��Q�����-�Y��Ȭ�-�(����(n�\��p��=�W���A�Hԕ���r�\����N=�XL�<���%$	]z}�Z���@bzLd Ό?��Y��6����n 4L�I֯��.7��X�5J>"� 5%��;ڂ�{7��V�Z�%�?`xgv��Y��V[��@�P{��xRXb���I�O�19�+״��<��:kC���8eI�b2ϙ��'B7Xω��1�oN����\��Z �����U\G�5���j\�x�L�m� $�|I�J����h�#��1��\;�]���P���g~�)Q�ݚ�F#�@�'�����:����I�[Hyi�+�#������Jp�A����u��y.,eU�����J��Vb�����
�Л|(0�G���E�����>��
�Ȅa4����Q��XmQ�JB��;j��`�rr�ޘx�n�L���|J�L
sM�����Pp������j͸9M�;��V��w�oj lf�e:�kW�U�J{pp��>3�3���������n�Qs��^�wܱû���o�B�S�%l�ɨ�;@Ij:1������UáO�K��9�)wôt��������ǚ�Ϗ��v��Q���c���7�Xo�� �Цd��>%)a�y9��y�f�-��MRڂ��ٚ�ݖ�f��^	��N�=���Ia���L�?�]�㼬��i�e�F�����>Wb9�|}a~��ME#ύؖ� ��q�?��YV�=�U�L5��u�C�V�S)<��(�YN� K�hG?!,�zT>��霅F��S��p45�,��� G���H�g~�jgN��0@.�<�g��7���L�
I�M�`�n�u�6X�l���2
� }�"���欦���W���hڏA�!��*����y"�@���;I�-=��3زu�BQ�����D��E6�f\�dq;νC�^��1����h��r�Ւ��/%��O
��}� Py�Y<-M_�P1��\w)��� '`)2KJ�<���?��c5�^��ۚ�
TE�\�Āa-�r��1��u%)�.x�O��t�3܀����KY��~;l����^m�7�9�,���S�*�J׏�3��@լ����� ���h�����ˋ*>G�]0la6Ha�o
y�(.��-���9bzO�Xi��$�j�$�k�'3w����u�Uo�@42�`.�m���,kM�i���L@�|ߪM)�W0cD���J��֡���	I�c� ۤ�-2M���5$�n��rl,�0[YK!��jj�Fym+"re;
�GV�x�8�5��ڼR���H,V�QyF7X��d�K)�����8V�� �g�
��	��,��*U#�����@}]|���Ws�2�b+T���m���u�Ү�>\��zGQ����
V�����t8��2`N*wij���\�U؝�Kb�G���_��T�ߔz��5���6P͒o�t��2� ��D���).G�,�bP�0Ҟb��.x�>��C�����e������p�	��Nk��L��	�L��z�MN:�XWɴr��2jn�C9C��_7�_ݣ��R�wW)�vhc��~"w`a�VDUh�HS�]�&�8s%~gs�����5�V��f��}I�2SyW^��{�
a���z "�X&�n0�T 4|����jyD ���������"Eo����6*td�LS�S=+��{o,;�^��½J[��ߛmU�8$���ޞQʤa�-=cd�jRHJ����c�N4M=���e��ȍt}���uk���p�J�tN���,���	L��H���|_����l�k8�Wby�
;0#3e<+��UH�埞S�y;#'��s��G���L-�76��*Ĉ�W=�X��`n�}��3D�ZC�~՜>�������4��q!3��V��A:�EgȣE�{ay6o	�\*&�7uV��SC��&7I��U�|�h�ԕ�極o!w������I��䱠��:��$�$$Z����|`��˝vY��A����A&=o��2��LV��kn�2�"�{||m�����`nfq̍7̧kB��p����ew
\�{F!����������ep[��H���y�I�im�	&�N�Q��9F��+�&��X�eA`EI������bQ�ܻ��`��m�%x�����1YD�ǘ~+�.���R���N�������/��n��ƺ���n.Ap�b��:TM��Y�X�Z[��~�/� ,g�9�^o(a��=�;�U���9qk��Ӣ�i7s$�^"^���h ��	.���}᮸����7"��y��l.����*���Ò8Qn-��׸q$O����.�2�5�Lle	,�b�'�7���qc*�`��HV&m�m}�\1�����M&A��B�8���X��[%��$f�ؙأ�F�)���T8���Q.X�=C�.��FF.�~���L lhEy���ċ��]};�w��bM��(+�WE�z*\D�P�	d�Fs�$�4jn��h^FP̋���~�S�9�9�����wv:HK�G�'0��/ ���ԛ�!qNM����qX�Io*�g�uE�+��t�o/~�v|�$��R�#�����|Ŷ4^F�7l5Χ%��I�=l6`<"�{�k�$�
�4�i�b�i��(Y��赈��]`"��T�q~Um�+]C�������&J��	M��h�_��$p�xgK��/|�J�{��%��-��YJ���*��Iޮj����K��y�/�ȉ��P~L�;��*�TOr��Pۅ�Rm��ǖx~��Z!%E�G+���Nv�"��;�o,Px����_�a��۬�������WִoJ?oK�oH t͍�ҽi�ۥ$e�H�ܒv���&ʒ��O������ak���"�/kl�-�4��I鎌�D9v`S��޻�5�{���(@����-�np��%��?�a�I�������e$�px�M�	��&����̽d�i!����@����b�T_�ڪ��pH��+Jl<P�#��la[�+̩Ql�l�T=��P�m�g��ay�1M}͠�܌qB�B�uڻ�wen���Azi�;�lp:�".����I�=y�u��w̎�dOη��me��_���+�`�<}�]���L�\`)
y@�bi&����NN.++�cl-y����{"l����:��� P���&��=��Y�v���@�Ѡ�QY����p�䏚 ��<H9n*�$Q=��Z|�@��8@2�)������n���|=�$-�(i�g��ֵ\�w<d��Qq�
�^��ǧǾ��/Z*'�*�H�3�^����Y����p\d�[G������Ӥ�����3pl��{eԬ��c7���J#���W�5�lG�'�kw�%c�m���$� C�z2_��r�ɬh���O�v���/P�.[\�6����D�70t����sa�T���^��q^t�u�TJX��d`��("��`x/��*��Eazu[�t��萤�˨�K%�:p&w��8�/J�1\h���� �z�2��*4k���_���;��k�:*�d��Q>%��h�A�����:iN�!�3�%��J����d?*-��o�~!��F�țB�F�༃����v�3��-Cm7EBw�m��#���Ƒ��O��m��p�@�����㒯d0�Σ�m�"m�䅠����Cx�3��לѷ�O.&�ӊV2�-�w\�N�L���rŲ ��Um%���Esdr��DK�~���%���=�?��{�����cOCWR�ڬ��V3��wŐI+E̾
��w�\�~٬��̻CYc���JP��#�*h׋e�Iȫ�zS1�w��=��	�2RO�0��zR��J:�9�b���9d�
�Բ
(0��ǃ'�]Y�y�똏���s*�j*���oP��TQ��V#)�O�������G� �`a�s{���tƝ6R$�.P�Ri�*VV�ݪ�8A���Վz�΃ `zS�������Tl�֝�@��v���!���2-z4A ���9�p��/B��ë��i��4 �����(<�V1��RP��i��Ͼ����C�۶l�|-�@�"�i���8��Z2�)�V�.̜��lJ	i�x���t�sF��5�� �|ģCC�Y��`.S
�(�������4:,�&L˕s��dT�w�#Q��,���f ,>\4o�Z�[D������%@,Xg�Z-�P$}		����/Z�p�sL�(���#e�.O��`��O*Fz�;�@j��j�Z�ŕ��a���cמ���DÿŊ��r�ZU�?�ڄ�GQJ1EedWp��p�Vkq]~��h��,�ce�A��!�q�E	����וqA�r��@ �l)�I�D��c*R@�%�)&�~X�1��5��1i^�u ώ��Z���pb�c��j����Ȥ�:�hT����ř�"�u�&S0x�����8�Z+vB����["�$�9~�,�GB�*5p���B�6���PR�� ��o�g�e!?��E1L����x_S�z�*KǍ�J��DN�͝�1|�/�^�y�+:>r;��4��^l� �	R��,�ڥ]LsY�����j!�h�zF�L��/h�.z��I��q�(�B�ԉ�c#s>��E���߹qB��jL���0`����,xv���x�
<���ܿ�ϠMw�G���Y�ݧ���_ѭ�Ts(ty�P���s�z\½��:F�o�L�z���/�vNu�R#y�"� �a���!`A �� ���|�6S�!_=��A^Q�eS�Nk@�2K���I44��r��Y4�(r�b�����w�a�����xA���_w�z�
S2�*���~�`�ꫨ����d_g��F����z(��4�i3��$�z�k�w��%��3��x�	0-����1�� �/x�j��]ΎF�U������J}�|F�d��t�e��N~
��!��7�	�9����;��q�� ���Y��!i����"oڝ@Ͷ�J!O��9�$��E�q��fʂGdf6|絼p����t"�t���	���i�.Z�����a,#�j7�B�Z�YmU(�a3.$�
����6u���a&V����u&ӄ
�iCʵ���JBƇBg�<0�Rf��@ά�}2��M��؛��]��1�(���rF������D��D���E�>����x,��`�0º73r����5h,� \`{g֟*��}���ِ���KN)��"����� :,��i-g*�ۍ�ބ4��$qƎ� �J~�O�f��x'��oؓ�Ԛ2��}��)�s[d��$����x�G�p�"U�1v��O��M4�Lf��7m���ˀ�UV�F�C4b �� /�� 	��L�6�Zk$.i�^���J˹ASh@A��>q:����r8�z����v�wѣ�8�{(m�ݨ�=���u�k&�M���Et�?�z�Q~��֜r8��d�.d�g�.gģ�:K����{��j_r|��.W�M?�B����,��S]�>P���'k�Ɋ�����M"+ �(ڥ����/�K���o|��O�I	:e��a��(�yDzh]5�~��2���F�C����F�� ���C��.����J)�s���
k)`L��|ڄBe
���4{rjj�d�`��Sć��cb9�:��I��%�+I4�����B��ﶗw��
�S�q��,l��c�^/��ff�|�+q�z��=��R9H�;"-m���Nx��������LR�c�����`UW9�ʲ;��L���L�LLP � :At��4�N��DTU��w��q����wd�>�`�i�F�f��#���Y'�Mda�)Z�BS$� �G�����P�q�\�.�;�̒=V�nu�c�>��,��ZZ`E��5�}b�[_v�Vh�dy�O���5����q �K�+u����"��F�(5 7R9db$"��?mP��b�i!�m�]t�F.�*�/ϛ����i�y�L=#���Uo��v�$U�a������{+V8�����k��
΁�����_h��������e�r�/"��j��]T�Im���	�&K��j���"j��h>V��ZK�$8��B�O�$"�	��=�[ɪ$H8H��_�.㢸������x�	Ϋ�]1"�Ϣ-`����[��?x��ś�EO���9x�^��ccn/h��Ғ&%C�\��KL@r~���<=4�bꥭ�d�{�Z����2+�L�tsk�Tx��=�EQ,a�-���L��Qs�{u�n�ir+#�EK�9$_E�}�Ԃ#�ǜ��˱�٪��a��	���`,Zֻ�"uNj��D�׿f� �s� ��
^�ח���Qk��0�&��5�L�8�&��ޒG`)�C�����x$KN겢 _ߩZ�4�Qr������h���a$s�^R�Q�x��'��~%�$��YO{��r�� �9mb����Le��d@�P�Vw<��+��Uw���C҉u��|g����.V���QO�pM����Ų��-+����K�X>�w+�M.s�@�{��e\<��L�"�.0Q��L�2�C�6��&�ѓw6�%N�QS##kmM����<�]qDoۑ��=,�iSr�L��겇��m)�/
���']���	��r���a�|R둴�@Y��^���t;�]��{��Ay\��n_�����9+G�A|�����(ׁ�
^�:������(øA�(�v=Fr��ªVk��4[8<E��ԑّP��������C����z]-=?��~A�y �l0�P�3W*�YɌ�'���/fR!�!�Е����/a ZI�n����S���L��6}:a�T��9M]y��ȦP=��Q}�Y��&�h�g���DE/i�H��@R���ۦ~.]��r�weh	�Q���Ym�F{F�$ź^�A�v�q,�F���g���FӋL�$�C��Q,HK�MD�5�q�9VY[w<8[o��:F�6��J�����(0�@ �v�.�z�>GL)睅\��7�wg�Hb���GKRM	������(��|��E:��m�rl�µ����������q�0�M!+[^�e�#�c.�NV*� ���g$i��o=A�7&6��ξzG'�0r�s\Q�anS�q��L]ٓ�N<�G�
���uY�#�P 	�dr	�_�G�XG����58���ŵԶo�Loƫe�S���6�X'j ���f�T��p�X���	�ɐ�^�%F�A^�Օ݀a$���O8�6�����r�����$������p�ŷ��9/�'pIB��� K6 d'�f��u��\Mz�:�+O�ա�P@�uT��Zж��}���V�to�Hv�L����{�Yl�Q�1H�i>P���d3Mz��NµC���)
ݿ�#����$Ju��E-�^�R�2����ݟ��߁pT�������I��ש���c����gE��� �k�lҪ�Z����_ҔDf~�(�^��׳��g�����4�%�$z�s_��0��@-��i��=���(I�p����0[ƥ�����A�щ�ʣlC�H)�g���IϺ|�1y���r� �~�)+��J��[Z�el
�Y�����`|:uf2�,pȂW���T�zN��{}��M����X��r;u$�P���"�g�اs��&��JO)a�㱋�J���Oh����J(�Ⱦ�:��ηà�L�8��3H�ﵶ��Dw��~nk,c*!��Κ�����0Hޱ���[/��:�ɲ8�h�D������S�\��ѿ�lX��$ϊx�u��1X�ц̍"�V��
�[�UX�2!�*G�}H��)�Y��Hbu`�a��8�6ݮOSבk`W�X�-���(l�Gxl{�~���ԧ��F��X� JS[�N�"��S�k�M֎�g|�rnN�D�L�7o���BC�U�qȎ}��h���}�#�q4���]�x�9se�7t��Ƌ����3�� �����N���8�B��&,W�Lg����V�&�t�髺�l�o��o�tȎ[����i���)]�d��k�R�<H}F�`[�_Q�JP�|MG4:�-��P�{�
��<q��Yg�I�s��l��Sdsz^�m���h�.t�����䗆bC���|���Z�w��$M4P��$�����^�f��Y
v|h[�����V��jvP>�$�B3͜ȳ��.
����]]���l<䤒`M�F�W�b8��䇾p��ߒ��f����j]��8�?yc�;aIJ͔�Lj9��<J�'���E÷�S8s:�D@����p��3�&驂��������>s��Ќ]���0leW��D�55�C R_�q̿��~��\]��7���+�+�X,<�a+�+��V��k`�0	�>)��bqN'�f0 ~�e�|��i*p�I\�ڡN��0=��4=q������q'��jM��d!0��ϔ�u��"����$�ڐ�:3+�!��	29ݵ���D�y�y�M�ڃ�'B,�e�^�S�7��A+H�$
��2������������#N;��WHF^��<���_�q��MO/�=���#��������x�-�������a�\��M)�K4>��L/��]";ޘ}���V�ύ0V
u?�t�B2�N�_:˨m����X����_�D����C^������r�k�Ŧc���we��N#�-�o����t�i��D�5�ȥ ��_��RHԐ��A �r��6hO:��d�z���\����s��g!�V;�{.�	��>j��G¨���N�Q|R�,�0���}K��,�k�ud��T������QR��k��ٽΧ��ԉ_��
��mNy�����Sf��w@^	�c�E&�=�>Ӻ��\�.�|��q�%�hߝH�(�Q��>�)U��Fm�ۗ*��.�aI�j;rff���{>%?�+D�2h����fT�v&��9���}
X��g����D�X�2�LhI{����dX|���&�(������T
��.5І|�'`�o-�Y}k�9�3WL���0�Eݰi��>.;l����dV�$�|/l4q_�?���n���v�7��yQ�}�i�����-�D�V��#l�zWh����a~S�a�B�� �N Gqr��M�����h�1yfw¡]��mp�C��/Hn�Q�PE�Cl8-ib�S\B$4_�8�l���2ݺ�t_�?WEKr���d�I�iKA˝��}�4f��2�����zy�� �X���_]���^�,3o)p�����9��)��l��H�Y����+c�%��~�l�1C׎긶6�ng��3mMjG�Q��V�A/�b���>��J��� a��q��'�*@�/��-���S���s!���ڹ�pύ2��fdS��de<��(5����7QU��:>��p��W�[��B��-��xy]Ç8:E�GR���[�Rښ�/����6d��]e�����Ɍn�}O�$ӝYUw)�ج����έ�\�>�u��F���f�	��U��
��߄]N��m�]�o�r`p�mGYVl2gkj�ʚ�ۓ0tI�$[��T�!"�&"�v�E�L遉,?��J��'V;.Ĉgq��ﵑF��X�寉q���)_�h-6q�]P�v��O��Z����.���hNhE�ʄ�t@� Oj+��
G�;�)@�sm����u:R���W�{((*���z^��T	644l��$jw��Uo��%��h�8�.��M&��j4g�{�߭�k�]z�c���n�}��&/,/%QW�[!���ʎΆ�8\}i�xƤ
V�NM����~Eu4�t��pߴ��2�R���IQ02^��i�7(�MK�HSk��R������N� �)t?��"�ULM�e6ҭɇ`ɦ��&�����k� ��>�偱�tfqw �}]�}'WB? ��E���5>ӟ��N����UHG�+�h����xv	)>�>�'v�����B�~�������Z�T#(�:��XAݻA�:���7���['�g�5�z�:,��G˥��(�Ds]=�V˂�W�S�g=*�i��鱃�s(Zt��:�8� [֜D�N�'�!���	u�3 34k.��cu��]ìZ����h�6L=��;86��-�X��N�3ԥX��c�z�ƾ�oA��\dx�b��Is�C3X��V4ި�u>�`�۫�C4�Vr���^�F��|	p��� 1%�EM6�*N$����
�@�c�����@�����㍝���tR�rN/s�f
y2�ר�de�'�( #w�/W��oW�U��+����U����ݑ<��؆6d��hJ�1���4M���6���ߟ��&���F����Cq��Ȋsv �Q��"��HZN��i�L��2;]��z{�670�K�o���S,H�A�\:rs��;����O�l�w&AW�H����*u��
b;�n�ۗ�	%�:�)�֖��o,r�xM>,|7��c�ᮭ�Sfnm�>�� �B�(���y.�L^}jF������N����{m�tR�\TB��4͡y3�x&3�l�D%3�!�S^B�J|�KR�Tt�W��$~u