// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NmwQxthNz120JNiFXVFwiT46aW2tlZWsnGSgq13cnADN2EK+kxXfXKfe8aoIKziN
ejWpFfpFbl5VOxvneEIgp5CvF24aJMMpYAwzhpFxvlRj6HVNEfbN4vPgvB8GSRzL
5Hg7gdsh7mBsw0SLYXx23LWAeVFDtMwhf8rNoct6RpE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18576)
WtcsdEEGhRFYXpTNxgFfxUWYkcYQ40JGK5JhOU2KBZl16Ma1fw3oFnaE651/BWbD
TEorz8sitDDQaQ5T9PIlZzTfwSfM2Y5CcSiw1EYv0JY8AoOOxglwyGlBXOzgSdjM
Eht8NOXd5AMwHOULWyL5mP+RI7JQjefLIELFyDdJcK2M5HAjLSZAokQ2+FkXvfPx
ewegtnqz14mCC+7yEfdMkO6YLmyoHJL7QIQ7AGJMmTfdGXQRpbplKMG3725hknXs
egi1WL4GW9NkF2Zoc3rahGJf+jJltK+2urAhUe06T5tKH082+CC+4qp/vzI3agbe
5RfJLrrcAsYMGCGh16m5XsH77/5r2EuOnrI036lZe/5PrY2PsZ7LCovihIJ1QRpm
JVypi+5miLK6JnzwDhb+1I6J0QCRJoK+TRQ2G9Ae/fiN6iMpxNXgEtvZ3Tun0Skq
fupAn8uPA2hix/pef9LWtXjAhZCJdw+QfLRtPc2uDzbY2QN9F1CYsvtIxjV6GoSc
o1ryI4BsfMkpfxqitH69MWaVlQJrRq1gWleNc8QTDRCJuqeAl6SzyEolfhaqUrUs
Bye4TqL9YJU40UPMtzCmKrq1FxNIOsYysXAd3iTarspO5NqzZDtqJRuO+vOhA95A
52j4wJLwI3DqBeLevZApUuaTTl4JgIaktLE6j4jPt8xrI5Y41IxSO8FMhBW0/weo
I6Kf77v/w9vS12l4Ma+jzEsXYDMs6T0yPnR/0BNbWODBSck8gZnQ1A3pkpJ7aC+z
zW7gDHqkO2GUlf1VLhb5LF4N4BNXxdHpylefy0hEbCUjZ4Nc1RuV7LcRggXs8eTa
ZF5HXVjCtEZXau/1/+EGCKJyWYzZiuGhPoH6hL41uX/5zvgsh0JNfKzVWEcuH/SJ
P7q+gtqU7a6Ch4zlS1Ip9XJ25E+g2QcRi8FNJHhrYQ2Q9KY2xyeJH/ORKaC+kQon
4n+SifiqVNxXIOMWzWIdUmvzoO7LcXETW8Trtwpmn79yEWaEl0o1CsjKdYLPI4Ib
uQPrKRjN8H20/zNt8YngiceIFbMcU32KCJiRKyjKgAMSofvQh6Bp0UHu0C9mHdPd
tMPy3aCx8EcR40ai6+8yShSc/+WxdIAF+w9ehRvcLzLlLtEqji5gOkpOKqu4yYk2
ugMoywKy0aBZFrm5doNtljTVc+u26W8AaHaaJypKB1pJViucT/+uF5WKE1ZBWn6T
Kj5xX6/11EtK05TEhM+t14NCCyMbKqfroOx8GeM8fWZuRpGCrOeVDj+B2ULo0Trw
qQAvAOZEUPyR+NleNcrpE+YyXijyBW9iCXvfSYdzNs6tlIew3gUnnpeIQEIvh0Pv
8o5kNu2XueYxyZeg7VZratYaYpVHdd2NllRMQXA9t2Xya17SUj+XeKtn91bdBkSP
akf5tlqSPpUjv7OK8BW8pta0K2G3XXpBynUK7+IRVgiYSCRItD9yovAOLgpEv8kd
RGnDPxtH/wb7as8R8KJRlwepS/B5sSrZupXUPmL4NX3OtMMxXFCb+mdXCuPjoceM
RyNwzaS+gDovMcgGm1buYLPiSws/y0HdS6ZSXW+9G1grXpxjAPiXTkh0BFb8+Zsn
r/m6f9UwpJ5dMdb46KZNztgYwX8S2NtSjQt/1pErO3oTMUOenpUknZVYXcCkDk5Y
YymEhQ2isidsJvLaICuT34VJj6bHac1m33OL4eB2MGLxwgSBC+6YUUMHIcM9pZvu
LE2Jz/fR4XMLaMTcDwFsKPEWhjKNAVJc7y4Tzl7QcxalDc1JHDbbk12Bqifch4jt
GomNYd4xmgztTIDlCtf78+rAUafgaPCGeqKA+0+KWY36QzvqSFWEmxBC4/K7fyYi
fdzRC0YS/LG3zlSuN1mteShKi++tkJQIIhi5soVztKPSSnK+HoNvR0b0EhvJbz0c
1LUFmNw40XBncuztkM1aBwRgeHmFnFpfH5bNNGBAOfZSAGk6t2fUJXkbw4zgOi1U
WA4HNFd2Wp77dubOPcQvNdT3kUdyrpsvEfwjU81W1mVbshVYh9UyUJj2J027Xwn9
rJKuPH2eyLQWS+CyyNXBt8j2EtFTL+4k4mNkrcGWGzO43Q6RC+So1K0U+hYKVlok
FYz/FDvKkWbHarOZwau6TbFHp0IDolTi39Z3ZRoPtmvINMGUoq/O816o/Dr8EEQV
mvtJepa2VhDGO2uJevjtl0QMcZulRJi/C89hF64+zztkPMwU0nLCNR26ARKSFDcx
D1CHa1J4r536faytSxGpB8rxq4TolSNalCFAhmVaWfBJZ5Oq1DEph4BnthCZ0yaP
u52U0qe8C+LsKvbrv/7drS2PB9oZYoBqtCIYX7bxDGdS9ChcQJNH+F+fwmhD76f1
4AgRUI7IP9cjvPlsXc/ZHCQ1mMzyLMw44AdHxQk+rHkkmy1lmt3hsMVBQx71MerP
73hkxf6QVn+J2FT75+haN2W7AdIfhLNTsPgR5R8unNRl33jXj95V1MabDhn5Fm4n
faNge31uRmAinDgwcSmtaepM6IOQfSmHu3uGPDM5zPXbEIYqC8WwytP2EzQmW7W3
FNGUFBBqhsgx6O4fjXu7+LDQB2K9y8SKmgOrvB0ut6urbu5iF3A88E9sZwBaXtzv
09XgWraHPadvuSKtXlkDtClLbhw0Oe9AwtlwklwipcEr0So11Z7nfdolouKu447w
rtNZb7z7RWwhcsF2ICZxSR93fKfJtOhEOQKjJsHV/q4dWSbPmPVTXR56rNOPM971
ve/yG3xu7ZL/Mwmt/nrJxTYKL5c+hQ+2wZvJ3qaHJ/yXW9lICrhYCCASSSOxy8Sr
b63wTIQZLZKUhs9v5ab7dnjlOt+XgVuPBjjYJ1taUJq39rIcgiaG1rWBcWmgOdvB
3RHkNx43IbhXfwbldv02un5LkoNjiYiUxbaVZaC09lTKSy7n5SlJP1LzNtUAfvOx
+Nr3orz2kURDRJDAH0yc0L2mGA/GVndxSy9dshMml8QV8+emwXf5cNVaGYnG0Wgx
DgvULib/fKS8tv2/cIYC2dwis+YkxiTjz6GF4pYfG1rRD5KqrqQhXetI2x+KT/9F
IBenfikalSEoKwU7zHN9edfPc84/4JZjMqSM31xyOzUQnxzAwxa1bkIPFrMOv4EQ
LezNvstNMo47YiQpm0L7kL0YKe95JdRRlHrF4l7A5TcfWmrDc/UpKbxqm2znBUwd
wcxmGVPcdjCDaj/J17MVtBYcxvjYnN3dAGVswaS0Ja2R+1SO6SuCTpx2GfZ55ADp
6lEKuZxoRTBIvHzBYXbo2idZK327IYiWBPLBXY3DSpMk49a4AOIUftnVPMTyLQEo
QEuB9oaZZZKXAdvDmST+RvsEsrcuK+SFR3i08hW+Rp8PP5XwOIgxnzevi2AIhT87
lCefpzRjNvt4l6LuwlqReSnuNX5e4gQXKDtvRXxgk+ohA+9c1WfxVcboVOY13Oyq
n2VZasq89tRqZmAH6vdsZETzmYr4/eSNKIR/HpGFgod8TSXXi/nM9Wb3wO6Rsrfb
9Ih+ZTDQGkEkLH6TJeEPIj4IxnlJFtPQ5/FEUpZ/8PM0+TyGY3T35ceRGCgxMFSq
dwULAMwNJUSyY7y4q7DbV4BA6X/VwVfoyfyUOUZ1qCbs6PCIP6A/QoUdbw7eKNUc
obiumiVD/3uSAxvtQbpMH4+ZZ+C8szHHrGyPeWuAlnS+r7S/L057iuEF3hcjvLR5
fVp2LhrlfO0AwBWaOe3pZzYJJs7UceoWzv0RNtF4svplGRr4NsKxFkiSb3wjW26M
shIak3tgSrnDShMF9QsNDNHP5bP6YRvuF6Yhvzu32M2fiiRvWfUbG+uTQt5wEdna
u9SXEeKfYMIxiyfSeGjSVyPhSsYESKX2vcWdW5ROMvXbEq0056CUpAtqLfRlFDRa
B+mfqaTfyPBQTNllSn0h9UWPWl5WRfaqDSD9xvGcvr3r4GtAo6GdCe3dlhCelaPG
PfxxWQMPFMaibSmW+hVDE3N1sbhq00XQYlXUvH65+dJfuZzkOnEJgaavMovcdef4
wIzPrVxDOXPEhfgry0fGueRDYJ9BtWM/vIsy6dQS+ghr4uJAtm3LG0zcd2KnNISO
Zm8J+WgQEqmcMx9xA7zbXgRKV2RLhYzVshq+DiRrk+mx0KnvNlLGg0azmFIfthts
LIMteLF3puIcRWGR18Py2wTV3jJk0bQQjOnBxm7aYN89RISicC7H4QTY6V3mkPCA
U3INvmBwAsywnfavpovASOmyk7E4TxcPU7BzbeKrziFE9hAg114zo0dfEZRzrJ0W
XgLX7lykSwJSInVGB+NekBthfuMCwDqAvQwvCkZX6GS3lrEND+W4SbKH5/4r0Do2
eFNOROJs8xIPCT1umyvkd9O1q9BIQOipNjGNMhfVIZiMxvJJTTjYLt4SiUYiEeXk
PUZfUocP7C8caEifjOP/2pCPJ9sEy3thHo6N48k3X9mS+b/KDD1CXuSzMg6AYmxa
A4ewjBWbESXbFPlck5GBL0TAlHMEGFvFuz6ux6n1AUavzCvwtmx5RkGvqXrLeWOz
FPNCJgnffaF0xVc803/eCGp4a5PKa9URNtiitnESdqGaLcS0Lp4+1uFUhYIX+7W3
stP8s94pwGGGD+SUZNBvbJ8vCOfjPzuBUNpB7fTYlUbHsQI4SBpEGW8OOH5TFJDf
z5wX/cAYRlho8KGvZQaWQY5+/avB4I5oG6tzRfpXTxVgM/N7q4vf+cUun892ccpo
VPEHX3JWrbp9SreAHH2G+udIEDO91wGPNoYyKpg9pYu5Z5ihNkeVRYiGNCo4yS5s
Fsii+UmJMacx9wvO8dms/Hv4AyABm8pG4xhppr7MKVKEqVKiSknADpQESS0U2IhS
Y11/UTqks4SS3un/wOye6jEn2Tv+cBF+ZK70T950iZ31kz/+eHR54oXSYlP30dsm
5vm/bTm5RIyc8LQLix8Nh5EjCBPguxRrgPySuoLGVASmZ4L8JnuHRx2m9PyFcfaN
NiKq7WRZJa2mspRe11ZXBI48rc4sNifSROSQUKf3yDBnT95tOMMC0DcRVp7t6ZAb
rlInCCRLE1kN2iX4qbUGcc6X6aexXSafeP50ENMEm1/sXP0fVzLTaL3o7F6l5Bxy
iaB3KqvFE+szFa7qZ6IhT6tUjfb5YcU34pyxNqDHyOSgEv3UAI6R43fr8ZfSFJWo
O8km8ZmvDiQXYcHCHLIsdP1HKRA54z8VzERdBwWAI5buNXjRTQ+c4uof4f8pGQeJ
KpZ00j5HZY8pfIrCfKw0dO0aClmF+neC3+d4SlA3yV0PLvzllCY2LV51H3j4GipL
5OoTpsK9hr8lcqhqJeTGLCpjtGUju7xLH4rQjGVSKk3DT1nOSSq3JcNK5sIUmmw8
07peoUysfE59btutdMpbk5/dsnEuaHIBtYnSO5zbHA7WHJZ38Yqce0oqVcOyGr/d
KZb1M4ZSqdM4t8T79p0FkCTM8gxXtNsVLD1iLXu+7+nuzKHGLWTqcMOGb4jahctZ
RWgIhKrFJRXNQpQlgTKyA5LEUcbPgcfTht/bJwI5ydWNhlefHVXaowL3iIVIJNZU
P3+H/BuDCOMdlC2tI5juGBbDpVeV00YHF/nxvYncscn8mKpC4U6CTGdLL8flk8cS
kYCSDlkRkkEkk39zbP2iifKzhLbjNq5HZM2xfZoOwmya557WLrPeAer4GWS/jD04
X16LKQm82o1bYeLtW1PeLZqHTgoeAw1INk/3XLAr53Ecmh9j3mtRzS/T8VF9aK31
7LeQ0AY6REj1U/w//NjJNZv/0SRzQfNpiV90OAiCZ3hja5cuClx17Js0LGCA2vUE
zSa1P8pTt7b5RXLpdt/e4L/WzecGiFIqyT6xE4LJF3Z0m5QUaUrEjOEIt1gillHI
1bvBWta82HyvuP+g3Bj4lW5+w4nT7EJpCsHjgMzZeQwArZjHTRPwAQV5HK8KCR0V
0odyoKuSZtqwRjojuN3JvQfIiJamrP09DpE1qfH1mbWqmjWscfgTBP0qcv1FMc3+
eTf1wrjadeW9FU+PBK31GX3vRURVAXwzeuypQNtQO65h+auWyuPUdyCwwRtgkHq/
boP28ipr4qwrDPzJN65VcNMNu5f4OHQHiwnoUysar4TW87tH1LjFnbDiNjjvl/ub
br6op1S6a65ET+AZgdnoiDsJsdygghDB36WUdpHMuMKl9QAGjva9Xv8bQNLK4DkM
AFpTyzCOUx1yJ4km11mQ3HuaaMgAa1Q5k74DTFGfWR3JHUDulCOXQFVraxemngjt
0zP4nWtvsqvnyFNkwBMRlyP0VX1OPR7NAaLCsh6fn38Ara9CWK+HqS6yNePF+BNU
qMGOOe15/27q5PrmthGt5LRhr5L6gYd9YlQwEVCfoe4EectYVvySvOxkPTk7G9RR
nKoznm1vEt/tzXXv0BC4LjDgF3TSZtTESxYSknvnlRatfvZGLFSS6m32dyp1a2su
rqKOMZP2YhVH/nMXO+g9CVfAT603KyAW6u/4crD3hkFg6qfYK7hy3G5gDQZRdApD
LU7yn92PW2RdMZywOsV8OHVJxF6UUhbps79/NMyqdM75/j8OzfLqzNvb/cwd6N88
7lEnXPj1TGOmlgK1C/j/2901RsBvf/nU1SEvBvCRoYrOwG1wxdK9fn3TiHwaP3+B
PymuW9odkDjUDyxswRTN+y+8iQYgkuLvIucyC7IqdDHT5usZ/AOoE/iffybVFHnb
xprz4cH8Mp8MR7dExHq2bs9TYzjVKH9KDl6KwuRWHXiqA/6tf2c+o0vgN9A8omFy
n6eERnx6z1TMEnzntI3DCjbSHKBh2goIJCMr7+Z2XVeudsZncJYyKlQ4YB+DPXuj
iCUnTR6ZLXGxULbZS0hJ5H7qvRo5TnRykfB4OSTcSYjnFLP5Y3ZfgFq7XxUROIjS
FJWqenGrAA7rmTfLP0ynKFJtfY/8GaeGTIkmPd0FHKyLgXWstNbHhuoDNZ+hpGF3
lxvoObd1BdSeacnA4sXgW0lWay8kSV46nYwjWRBTFptfBd8gmpBXbTXna3xVfFzH
h12I+YzehhPtnue24vjD5zpUQE9ZK56WA2WyfjI35VmpSPoRx8/1fj0Ysh1RFK4P
ZytRUA5wAyw0lrTz6ymJ3iQoLEh19fPy7tZRH2HxLtyH+IhW65sFXBhU+ZtudYz+
EQZL0DUNpsQ0eEt3A1kqaT9LYs+6tlFRULYEsKM0VnHKXDkpIMvYbFNawIk6qUd9
paAx4XeRC/q6s+WaDuLqdGQRUCuubmKAI4XvnDU2JQ4QkYmLTT8uKUGZAP5+XfM2
EToDuivVnN1fIMDCaSIH7QjRC++djz2sqRIiXp4801YUoC/POMdrIMfy4+jh7Lrx
dCLXWNgS18D7j9yeXon/E0JsPKuSgFZDDNYSu+iHQq2zzP8Mywz1tlLttMb5Cey1
GRq/1C98o0gF3UzOpO95MKLfWWJsZezTRXPU/Rp4wFApGYL+d34Oy9bsfgHnIApf
EQLz6DtZv/CrqWBEUG9YlIQKIAPOdEW7c2gnWH6LdEEDaXmNNEcf+E5oYMcc981S
zcu3q1y5sKloqNvjODhRz3eQ+CEjwURWLKCKqWaZmjGJNokAynupmI1gVDe81H5U
ybjT9sb7d5VzUpDbHD4DQA8JhpWfcER1oUdYVGAeWf0ANc/yzlkmxKfXmcdBsYvL
k7MjwiQMtG4hX/qiO036OwpTBQOwKDQsMQDKY0dy5Nf03ol+Yseivwr4BHNl8Emg
Hj4wt4GmrGz9J5FUV0Im2zTFapYMi1IQ5etkD+p9TCgsdCCOfN+0S7HHRwpgdCwB
lnKV+KVdLOxAYJf2zjLZRpiF0t11AR/piiGfbbf1Q/asXT9wruo8KE9q/3C1uHxa
laWZFmpPxtLjimmqDTyQcz6rUolN9OmD66Po78sGeS0TAAz6u6R7h5ydQH+0QO5X
tmll1QgHitGkx/jkxIwDExsAzCKfBIeM+BotBdSkpiP2FoJXOTP97oJgqdKsJP8s
s1aMEtckEh+jbawsbLfLjRDDUuV3I3T/gkiiVzFSPMhwEHMQ9WqP7PebZC1SsZwk
xCceP59UH0bSVUypRJKg0cp0vTQpXUINnNTl4mIfJHwwwhDTgiyDCgW57QMbmStH
uEmAT2yga2TiFtZBlUaDxlJbQKKYLr1u5WEr9i8cFiYER8APACCpveItjOUYzik0
KXdEjWIGzVkFlbFjzKIekkZQnTbAbKEwmbuGU8rqYfbCrBbOZI6CHRBi1mng2Ad7
uMnC8y3qmLrfzCMvgPkqoCxxoScM86SOnClcyX0SdL8KGOWO/kEcSKk64vbABxIs
gdoLBSitNVH3UxQs3WXvETyxrnOd5j0i/QyQ5xg5y9VzM2NjDCMEKNKU5+XGbV0w
hqgHwXAX5pl7DSfV0NGguXAxFv6gWLvfc5uuXFMVpVzpSGa9VCXBcc2XzQqX/oYp
5uQzkqNnoAp9igkh+vC6B6XVCZpkNrjbjqFMY+Yueuw70VNLSx6elVhocS2K5D2z
b15ZjvTjdXvdV2c5WxBLIi47meEv9Yj0kMzhD4xZTfVowS9PpAU0163oXg6V/3eS
xafpJ+jkTIwC+OE/7H7VQayeOA6b8dTIPL82ZUH6m3ADqELp0/8jfBlVckHg2nXl
dlrWRyXVYHHBnDM/m2UKg2Zp+kifmWddWNRP5Iwu3vo4kcehLwnrwSvVZgE1wBpp
slhZ6dc/wisZT0G9JL6tqwJ5ySwj58cznk5I9L4DuzR1Q7IpRCj2IvWiRgPLwMgM
NqIyJI1nrw9O1ClhOdiw89kdO4mPhgwf7hsQgz6TLFCEZ+KTxb4xXS8GhrQ3fjPt
3Yo0Y9+oeXz05CHM5HnjUI1g4yxW83Wq1K92A/8DsMqwok4m80xoxkPyTQ5QjU4t
97jdivUnAx6kBpF2I5+Ca56XBlduwnLQQiHcKMazTCOQ0yOMVCag3GYt0+W8K5jD
I5KSDGbgwsjqW7zYzy96pQ/naR2e/3iOxAhlwDqU2tu2qWywi/Rih5rckYB3SQQM
SKsu89+IqZsF6ho8RBkWBv04UamJ5ZjRmXl/l2YLminKRKLXRl4t6f8XYnfQSFj9
S4eUBqCj5silQCwco+P/StY+ZF/qXdIbUSVS8eCGhWWzcAObdz/E5fugysnIMc3W
7vzgAy/M0MVcCxq/VG9/kMoyNCaIRdmYIGy0J71uLpx9AYmCm7prPlRgjsWQd66W
auUGGMoLsQEt8k2ZFmiCHJC8IrHI6j/5XbWWFPnpKj1+ph+PxrogQGXzMTJsb5c1
3TZyW8lAy08MT5lMhA3dFBe6opi1kBsVlkYnmqoGQPa4t0MYfbGXEQyb2TJatDSW
akoYz1jpycSLpY04tIom3xzBycN7GErMmQGBhqzTygXcotuVsh7WQETAumXVA0Tn
aIMnDttI7qBpSdUXuV/9upPHjb4VVqR7Fj9dJ/CK4Prr6aGKW/ZvuZI2Mc7K1jrP
FmY0RB5S9wPIRhp6cabtJHMMI9DCeG2s5Eo1wZqTX42QlPd07nxtdLnjlFlK0/GY
0dhQDJeVJZJoQSMtcGXD9qghu34xEJgYHdpC1Er8dPqN4ZSrXrgaJEv/WZEeOgkR
SeybWGTHHH1e+RlVlwkBB0Aaccuc20WJAvq03lH4cYazbJv2pwjPm31Tl7E8OIM7
mJ8ogpC4aDPjxrb0q7rB/VMe7IQmSYvuWtMsBuiFZafFhxZaS+WEWPVmvCAWYLcK
MZVAxe2AuALPZA37xI0FY0w9YUqY3Q1rFRdE/4ctEWLf2uQJ6zjAJCWy5+HRF7Y/
HU23V/pvCAnhzM3+SSCwUSkvuLH4bWfN3sfo6P5I2WDk3xDbBApJcjswG883ubN/
eJWi4l9kJea25lNRJTa9EAtuNMdUg7H+afLiPxTjZN7+u/zTXDnYcyU3J3hQ+syF
SrDYixhJbJhORFM/yjPLx+akZS7aKA0n4MePRii4Vl5wojrz7Q4wOpMljbIhkiti
5alRypcv8IzS4uYCq3KvlkfidMk8rvotJLZHKxQg4t3H5b/KZEcrLjk3Tekwp5+t
UUSM1HP1ufPxQMA8NCx1zkyecLVmzy4DQDaIuOlrcTt0z2mfPQE6jcdBgejcWAb6
3mlj9szV+k2Lo74dnin/S9Pi43z6Twl2pzeqlU+FsTuPpCOpiPSyCK5Zf/ezXQzS
hjIPf8DHmVOKVIiglFEq43eQ44gpVwHA8txJvqw+E+4fZPz/ub07pMpmg8dgCqob
p2o+U3lOhPhtRgVlOyuEQYMveYtQLbZpOP2Z0SEgnEWLr7K5HEf4ZWY9NaXNiZEE
djjKEkOSesoft/43xSYHc8y9ubg02fH/ifVZBtY6OEYfzR2fpF/ngnICGydxqHjx
u9idCo4EUoLHOYphgvjbBDLnPmDqPV6u8ciJ4UKEUHjsNqsxJCtlfKdQTwz9Qr3f
eMTTSasczHgxCkTiXNqCJJE7aTH8ZNXMqlCIh1ebXjIyu7Cj/dRHdDtdclMBhmXv
bqICCSLCXOtSiFGPnQdb7ozu/C+mbJJGZmTK8jesNsJg2ZO7haZwXanssRPspzfv
4bhxw6UZGRp/YgSqlbiBBk8G0I0vMOP2eQYMIzm3GSfOXDZDF9430lU2wMopSbPz
EpEUVlstH9O81xG7DE3kAa6yNURu0+eBCzi3GTNSC/CAF3NgMDzdjKtFl2pz7nyu
1q1hlkQPH0BAtLP2DFgsWZHKsjR7PfDaxu615PfA0NKqBtrG76vJnDKDWDdI+mSx
EhetALuKdNxv/93q/iRVuGUMekHOtdCLRScUmIhOWtBWY0OzrZU1VwQ1uaCe49Qe
MdwiIg1WOssbcQN2C9Ct+6NQncin/Q11h87udLSx7uNDqpWTRaRGC/J38Hzepv97
D+BrhBV8+CAPyI/Jn8yoaqCnH9y3qY4vISiKjOxPKs1zlEkqvxBy9b8g1ybIopLh
dq5oen6LK1CYvRdAe3K/WxAnW8fC5Vps0ZtM7+Hx5HcSq5WmqulLkd3pcC10sVSc
0NFAtjXGYSqBgU17EY37sq6zJqIDr89dZxnYdAW8diEQ4klgR8tAFUVhQqwF5Vqk
w4snzVeMdK7581CNIBlIA6bhc9ZekZBSGejL3mfk5n+Jld6xwSruibvFbrMqOK2x
JYza8vdcEthoOlmXdZVS4rMaPArl4hibSZN6+RkfnVGbBNIXoFy8o7nL9FHB+Tzo
Kc7aWEIbr8U69Mnq2dZOo2WWCZyAoNiGzcVYerC6bs+ovwEC+ZJXichIyED+oelv
BLu8TKUYKucgNupVQl3m/4+5B5ZZjA29+JcOc6xvks4DjOhWLMmiLQsX4k4H4maO
7/a+fxzO3/sV3JH2TMyHtK4NYUHw4NueF1ElQnmSz+4daXRugFMH8kTuYoPRDpR0
ZUmxKWFttxg46Eld5XY0kDRrcG5WczlfLZSBluoFfjh3TJsPWXlwon7kugHEEqvg
2+4mvekLFvXXbkPpErfCZ+Uo1O82ply45x4F363FVPbD1bmJJuJYbTnZZjwM4p9Z
pxS4HiK3qN+XdKMg1sXEzdP7DpadDctEKpglbBHd8ysl1sBTXgZr2IgFP3nYNv6Q
Q9EHIhNjac1zTUM6wmom58+qSEdirwlsr/O07QnNkT5s40P2+Eq9FjrWDZOGPxEq
aYMbbsS1VDJqIGbUyYvNg+ytem8cuJJpM6R246bprfpwYtq2/nye5zXs60wNIrYc
RomKF8gbyuP8qeQKdGdQt+8+28OMShZlQMOG9NiOv/aXLaAfApXwGXBYU6BSzjwh
UprjG54SvYQzg4wZquJ0EI2sbCFVwvUeZaq7HMUrjKKJlyixrN1g8olKUY5Xq9G8
BmBMgyKT9ekkFs+iIpJsD9s5tgCZRHlKmMVaDjoIdTvFnrkBAoJVAh1Eo/akWpC6
JBRiKUqPY27nGai/0QqNDxG3G3vujPEU08VSxTuEQEV6/sh0oPuOXi74fsGuZbH+
6iaCpW7rEtq01fehKreWgZh0ka7/lTpsh1Hdk4DKeaTRACSG4lqDmnoxSzBYKodk
vFO/kESTorz0xnIesk9isRAyL0ULwPccdc5+Nt3RXTDHpxmlkFAv+lWQgb0GoTc+
QCbQ6RIwVK3FRUsRvaHrjUAIDrz4BmNNS9zD2GyyFphnNAhxDG6cHP+5sVVkvAMa
OJiUca9Hp7wn5zSZlP9xzbsqwrr8F0Ta9Gwaps/vvoNNsRGS0n+SklWBLqg8F/9+
fVUS74iZCsUCFzPYLXMI5ZQtGLmpuz6rmzO+2DAUrakfdfAwqWeUzOzFCfARW66w
aKfuBieWffjmT44pG8mnrbPtH4QHevztsFm2URYOkXDEFuuDnrHmjrBof4ErAYtV
I1DeIsrDacUxtyzQmvXdXbYXyIsFjGXmbhk6ivoassDnmGrzCCbvlExFVHjof1LB
gl46K7ITmcPvzMx2O6ewKWErrL7sVaXPAHle+LcjtPJu5PCw/AIOyGeGs9xJ4EWF
JWPZcke/d0scC9/SZaY5eMw/Ye9QXat2gBzJWv19rdZcmJ9pjTdef3H0EfleCqWA
cJP9mXXwcqjDgKzyOLo3G73eZa9OhbW5lA3VycwgPzhQoQA8Dncw2yCGC0jL1gtZ
7LPi7uRsEMXiD6XDyYtDvJCFodq3iZPou3RUlkGF4EGuODwCwJd6PlE/0MkjJ2G3
jW42R84FuGhNuQC+O+fWrVuorYlRFW1jlE7Djq1edrSOwmJHtulPBBrMif9gpNfc
wwTxw0W1SQfR2Bx1OYpoIp8Fm+kYp9oIzP2e8POe7DFisOZ/XKeWO1I3DkrjJwP4
5D3loK9fNMWnd/6lErZU6t3gTiBs1ADSKMW5XX4lXv8HtZpUihN6xZcDh+f/PipQ
CeY4o/Yuqc4OwGDVmtcEgOVU0V5hhEM0I1/T5LaytL/ZS+LqQjJZfs4GP9OmOIhm
akpixy2CnE/GIqzYArROyBZg2iolNUq+KwsDxDPyVeE6fsb4wYvi7hUytB86RN9+
5AmSGP0m4boMG1tX1DmVIObw7hrP3kjj83ngbPBnMX8lRXMc8AIkNYMwBAwsd7B1
SKe+vSv/j0Qpk0lIUPj9nBDy+cuWa0r9R3D6iCQwJZtrSqzwgouFZQryXjb08TZO
NfZ/15gArNd2YASxcGMgj1/Nat+qKJj6vBb5cnEEV3NoAlzDqlb91VNHw08vpykg
0s9YNi4JLx2xiVqic+Ppp242PWxBUydVVJ6N92/WfOd6n5s3rGeaCPr0KYPZeTx3
n29DbS3i5YUajnEvw6CqvNxwDUqzZfMKmVBsUS2OFzqCkSBqUdFwujEUqBNvn02I
/fEnLKMzbH39GlG9zSevxdC+RTRpauUnNXb14aq77xq5rp8UcebbN6lXvQys7HfN
goqau+AaedFOfyHvPHFio0HDdR1MzDCtwDFQMxeDEeXCM1x7ZGKFUpCqvoIp2/p/
rS0rUGOCcExtw1TH1v3EYsHvEcZorH1B/kTxOr78Cj1WvQx2iv3tc2J2TXGrwg8E
McCj7ARVYCZlC/RNPF/ZqeaGEL6ZdcEt4vhATVE2cVE//r+j7pgG/dNaU64I2zzf
JHXhBhWpXLr6XdbM4xIxv2N6wX2grgLkBEANhwCyGuJUiARk9/0qRIkffyjRFeJp
Zwxxaxi/HPKmQ9dcAV0yjsSIds03JFEDvB7kKlMdyfrwONhCT6n/yNAhubOF1N1E
qHgDU86vAae+xKqmD+OzNw1USGkWjw1nQYOUdIbEAP0N5C3v7s0hX0TkUaRSOyhB
VhDKVQJ1zXxMM0pueZ/hlbCWTSfXf1My64EmrBVz2lJRCU28JpukZjPMs3v/4uI/
kwmOU9LP0aT4qxNAC2oef/NxL4l92Rj0tNIGSrE4L2SSu+gaQ6yoL/FDiNySQRxL
1omLely1BIeVhyWeZas8Ka3iciPU+FdgZWCh/yS2QmKXXAyoyhm++BsH+dOakXhQ
lUrKumMe7X9GEPD6lknRMn9qfbjoljVQWcTWjg92RjIjNt/TVyzbhxrS6J1yrxId
IbRHJ/aRhWDLNTB8jzizX6t972uhzc1TTaxs8VLLB0VnhCGlSS08y8g4KIdmG8RX
XI33QJ7fz91mnG52JmfgfwDUnAGmOINpM1a3KmOhHjKNYIAUaRyzf83BEaL4/8Ju
2FA3i6hwWNjpO9OKuh93hhunFNYaSXkFrvE0Va0xxBU/+YYFid4u2PkwryG4boMg
W3LpBp+GYffkZa0eyGyz+PL7aJMpT2qizvoEtuoPSIPyqCsuZkmKao+zZmmndIo4
OVcyjewH9fwsUKcci2uUWtzNeFvPdQzEbY0kIQwk4jExfTpXuyTntcavt/6Rooi0
8Y7f+5iRkZz5GrNhGhkggo+2sesncSdFDVzG2GfqXww73MHCxvsV+Prcidrb1xvn
qhpFXw7RW6hXYNlBg1Bju6FSUc93F1zbW6Q8xTCwGxINV/vEX0m4Au5cvG6NvBzw
wg30K5K9I8Fn/RBg78kRZtvdvJWwn/E19bHxikFUV+9Vawgk9MgBe+UUCK78BgfA
cb1BGBJ2ULKR902Eufzp6zGDybvYBStwpDb6HTk0qJbEli4SAOQWlk1z6sTdLO/m
0I16DkCzodmAUS29b1gurg5THx869I1lw6wTDYupnDvTWpcb2hcouo+uyENVjT51
pQCNb8cx3gJxh4BBIH6vf8S8h1kRMJz9DI91pp1FtrswfPP+jBQSpkCuctCSuWWb
bTp/jJ/2DxbU0skzNNQlg3pTcvuHpR1MqUsbZ/k11h6UbmjDw+MVrGK1vdMX+E4k
btMa1qo2ZPqNMjQRX0jj0DJD5WbBoc+6UKl4eBWtZUIXKs9ii7/xBoQsHAM4fRAY
K3EY8WkWBweuQv/JU+YR2EB76XMiYo4pBZU+ravXPpeQYrbfnaCw22Z9fW2mMm8k
AwymYYCN5AlUlrUJgQvNMv1wHo7/TYQK9rUmiPW6jdMl4L+8CfFrhcQHoEz9nNSl
aRETgzFY3Z0P9JFZ3IOTW39Fd0y6yNobasi+885ZK3CMZVd5C9RV0VE9/DQY9jWA
+x5Hi8ZBOQsRmemowYZye9x6fruUvpffL3MUlC5SZF9nD2Uctx1RVrF2t2ULywGR
w+L8fQYNCvyi5lAmWJHeTeRcSbo3W0y15C2myVV0MvvQI19Wq/hT+4p7LHvN7Zb3
FcTpHoMUTiim9q9KYlfhYa99F5shUK1JWIRF+WtFiPeZyjebsH5itwD7meEWxrkc
D9zYlwf9ebmekkIlKXeA8sCftluBOxNY3LP6hrTr6GDOmiUtBZedpdLIfi06r8o1
/6TAXeh223rM6nSfkDBdrADBy0+mk/PfjwSOKmFlu49hvpZyUXKam7hr+/QtQxC9
9gp7SdQZZV/XQujWIq2F/6insDlyoyDxUXzvqEvSYomP0oMChREubiJ8btZIW3UA
NjGQi78+j4sns+GgQKVMfo/vE3/TEHMkbFyaeueo1s1zbT8hJN37DYUa9SLr1vQK
RysPrxGsU20Wn/2y2zpn5Xuh5WcQvTJ4iL0Q6YJVsF4OlnYhLx5NgmGv6qnfmRCv
rKqTjAchfsNnnJVwPAeC82XGnacNzOVu4Cwjof7wEmB3c6UtfNkq4NTu2SiM5p8O
T2FuxKOo2EsmbcKgN4ZaNT/FOYk3bGpe0+ipli5rF2bv8l+cLjQuZ8PvtVvAtoux
i8DmuWgoDPz4eZT4gPPHQa1x/ESMQlINR9vEBDusRtWMjGFsxti5Imb/mk5bePWQ
gpOJ3xdT62/kUeh3nDZuhJ/psPRyqaqE89nKwbO5dnRaCt7KQTNsToC09VXXenCz
ieF3JKH5FrOtk9RPlcMUxEPl8ltjuXQTWLpOKItjk6KFirNgKXRrQpnGOB3GlsUB
AXfHU0GdwbOcD+rzh1kzMZS8PSVMclRcOE3rj/4+nRFXPSj2nJkylqkF2iRp/NXe
keYFcefPpMqjzRn/7T/9n2Ql+1jdVa7n9ivtS8G7j9GpOgIq3VJB1SQB89DQHit3
KE4+fGUEzCYOO31Y1qVHJ30sKx1NpzKU3wV82GPK6qBZygEpBO6UeiIAjVVrEocQ
Su9yVBnWVd4Y2y5svWJEaYcBDjIaJezyrU4BcNSuclYl602GAtXfzD5HE5jNRj04
G8ly9piEa64DNWwonkg+VNIjnTdiT6Ys4WUs0g58cD03EX6VEyflEm3TpXppxtBy
iUD/izmYCj8DrHy2fez3X64MNguQVHaItPzZL3AhNyEUpn1m+FFhFCQfC79QiprY
qFg/HVpbZDusl+g6/TtNRuddZ0Exi6A0o0Gi2BFrjxPrT17EgbUmI5j7LnUFnPyI
P7CtJfuNL3dYsow31Gfr20LBHheCtQrml8WXSzMN5Gg6cKt/KVp7jbuW7VcZcBIS
h0pZzxYRQrCzJKDnZNfkNLtajcQlMIKK7eTe8dzFbQshcoLxLUGZEACtWVIKcBGF
b0f0anA/rNHdc/cgsIms3gR5LgsHDIFJvOcfPRvSfCeneQ+8NkDciUwpkkWjvzid
zPPpqyDyws8fP4p3Buc8spIAiRSVlOggg9yIpJ0joN8/oAVcdJZfUWqVYgJ01SkB
ymZgC/QPIZBs+bPzl0Mmvi8atYRThQMkSCuoPVxRQQnmOQ5DyTwIBpWBCw++vY0K
ujxoq3nKFta39kzIHF/ZeKe531qb1x5Bjo9yEh8b+XW7ForkmYoHqpUNL02e7ksU
UqL4icBBZ7Vg+rDjlvCCWqHz7V/xa1jdgSF7xz5hBT7FLL3hB5ahzIN7bEHnTFIj
ugCj/XbAVILYpPSFOGBpXHRf1soW48vVLzmv2m4lw+265LVqOz5w0yJa3w2wCL2r
v3XeL1GSye9IIOgAGU9VUt+xsKdk9mzw2F6cB7w1cVQvh+YTVYUuYtwXm3wX2zp1
e1HxoehIHZzFN4TLCOOA3e7lCEqZ3qHSBRP5M+4Cqo47cGxsH/FXed3MvT0YK6gB
zxKQIaQGCWB7WBzYC+L2Td/6VlLpnEA1tBC+QD1sS2xBYLnP+hFpnpa03EOgebqU
0AQst0HvMvdGkKCc+X2iAwnZnipEvRYI4UK9tnai1uCVyw9Wns7D28faNvp/J2LP
/f7DQHNJzj151SvLQO8F0C/H33YoBbc8njKwiduXSrQ1IxFJgBYjYMe4sEW80GlC
8VcSsVyKq9joBwE1zq23Wkh2NubvXkpwy7CytD7JNNTYP1/A8zSlueBOuM6rQ3Ny
T9NjkFMEO54q8tDeN4UGqsLlZQu5GVK7Rm8BhJ3GdydlpzGk9wQdxwYaTHky07g+
/zX9gD7Yew5im7ehGLPvFIKb7mSAjqeQziV2HP2GtyIqj0bSr03ZZL+ndDNOsrVt
uNHH4ZESG/6dekh9ivugyz0lK+kCRgCYLOycIHYmpr7UuXek+h/akm0rOXwlnz2L
kUD/3EHhGrpSW8Uw9/U2aWGVigmv8AarWgE8yNcB4j/WMVmzuwgg4LRqywF+buOz
S9w0TIhucQ9B6ffYuzod6ECPpGX4zDnielf/9NRx0kFEuXeLqZt1X/G3N7lLZFuz
EVqZu4E+o78RmBhFsiJrpDBOoyhtSj58FFVpqsAXJC/QtGYitNPZbOROQINaKh3i
cqBgQMRGingsJv0pF+2vMS3IFdLmkJw+Dd3qw/2ZVCYcjM3XxzzXntIVi30Tkhiq
lf8hXS36PXa7NYuC0hj3WcNy6Oh7ZpbZMuX6QB+QFHq2ZhUuc0n35+VbXmqxDvLh
oDqRlDLV3s62dRo3duDnqGqxyMl2zujlu8iColp2yvITDqfDx6g7RT5NeFqAol/Z
1IyA8QpJJOV7LPtMNRdo9aecP8RuquMHLEv3sLhsHFpRY6Vy0b3lcjV/HVpSHVrc
o1NIznRxLQg/Zz9mFhOKDZ6dRWm1W/Li/s6mEjUYIwGlERjLmMDxSVZmfDqhutW7
JJ/aJrmlMRZtRysQ3YhonDcU/nEczwiFpXwdQk2yHY+LcIaiS6vjwn0+iHglmFZ8
qjdsF/SVKHDu+BMJurMXhLMZ1F281KyY7z9a904kFKSUH7qE9fEC94tMOkNVEjBz
ejUW+6xJYX5w4NUYqtx+O2DjKov3ctqAzKkJ8v5BhfOPegbI66+8QGJdySOqjrHd
az8lZ41bs/fyouIkkszwTZeh08kBLH3eQLad0pwgaiiAJI3pmQ5bvwI9OUl8QDrE
fUhxo7+9YjxzF6AD9kjnvNxOu6Pt0wYcn5/b3SBRXJVz4eSX8vJvhqxZPoQhnI+K
G2+eRpxDjQuvCYU5byzk6nIzhT1pLIrJkeH8DQ/Jgxtp+eyAFnxWNXCBSlITk/8g
dENugKBa9Et0Y40kuDSWIzZZlZ2mAXUhw+t3uu6LXS572RjHaY6WKcDQ3+N4qamw
Jfv9S+BCHzxL+yqCkHa+Vmt8SthoLaxvEF2k2DiLSdD447Kf9ZZjNoXU9g7E9j3I
YhJx76Q/Mpv94elYPM/MJCEjFNf3CM62F7UdF6SCaubUEoAXxwMMm60+g4eTmDSe
kY7AOHd99PFE3cuC4f0FlPWcRAIRzPvn3Uk4HMP/9q2YS0gT1BEsp6GKlan3HOgx
+H739NsUP/F7QUxrRdeqyc8tceLlhF38mchDG/fVYPkbzZ0WS+14juPhx7hb/gdE
J2G1zG+lLe0KuhEgadxSULtu1trcaOMaoU2HRcxALOAvG3445plE3/Nmk9fM/E2j
+FPnCZxRcp7yqpjDlIo7f+/kWgPaRd74K5ODcl1gkdJbrxU8aIaPnBCvbj8smqRP
W8K+dd1GKQEDHfsERjJeeqcHgRaL+K1hIGMmZpPMxO0GN3osbFDHtlRY9IgweCou
bsbDzJdx06xz9M20VZU29EtSN9FqPw0Wq1jkk6CeNIv2iKye2Exfa+Etfuhf6Rsq
5B/bWAvvwnc+n1g/PPQsajcOJNOdDbkw9pMTRRE+exHfSMUHyZXfn3fXmqOzMS66
OJlq8O+8slyVxLdxQuWzK27Q/3dL9T0ZtoxanWBy3bHhjnLFyU0vpcemBcJnMW/k
Dpy4Ruz4fVmWcxNDkB8PDSvqVVPC1eBUd0omXGsmSGHuq0xekAhXcx0MCaYYZRBt
9n9TQvyyCH9Ua4BofDU3p1ApGZ/jcvNpu0e8qVLmXs8lO2l5ZBmxE4PizTYt893N
XWyCGJ+U8KGCDKf0UA6tDB7Aqeb4MaTWrM0BGWDiA30NG1MPWC2IdHejeRULnFKI
VAZ0kUDs2PJqVxpXKp1BgelN0nc31VcGjYzFzWR1Li5pTdtalfExro7CFivLvlAz
yUBeFIl+rKhB5uxq+Nvq5/GSyjcWpgrHwCDPLIRtV+A5d7Lbb+yQmAdJopt3q2Sw
sAjE3eM9Sr6doHl6e7d2qUxjO0SAWfEl48vmXt36NgLxoVJENtXlt3uIXdGpTiFd
/oq2aAiiLSORv3WD4kuAOiYcwI4lZGkEpL5Mu3HhCJVyyWtOdiXXc3Gqnf2PsTyW
fRGMvSbQmgpJrMs5C3XpK9uTO6h3O58zvtqhUdS1DGzXsUsOK02QGwOTkS0cHvar
aZIJV9gU4HbAhhJaSvnfClzJYBMEs9AT2Ecte/H6v+0WUkiKX6gH/heFeczMGuqR
UEBmSqi+DAlx6UbRbpsxREBRqs8u6E+NqJ1Jubl0aVOb7A1mCpCw6ZSSlQVU71uJ
MB+V9tJoJJEdxfM3INjFRKuWgDpvMp6Bs8NEiPH27IHuv/F0YHFjfdBZN3Ee/GoM
37qcrJ6jj6Mhtx4yXjbeX5lK6ssko8nIoVSG6f93MtehPla+qOn+eDfC6AtlwhSR
DmDjRWU54Lftb9FxxdsPXCIPNOTwOTAxpgwWD8dT/QuqUREfRq+6Xt4SNmAg/j56
opXibXwNP/I616S+xaguO1pTxagOmotqzLvzCDWlvuVmGpEz/WIC0OM50g6Uav4Z
13aQSA/tB5l1+nVdK3QyitB4CFixmmAdSMwjpnKtALdxpvN98IFTKTozEHNm+4UJ
4JmAcD7w7TI+Pz70P/08dUAp7waxtbAXp2EmpAqhzxSEfW11JdnIXOpfBNYlVrIq
AEzq7li9eal3G3sDeOnEe0/u50LX4++HC1v3YzkAHWj/X2DtCusQU9YZ+RwMspz/
8n1TNlQxBCFYIKroOd1hl3ZmtX4xOiu8stX5Ws2JEyvtwvt6aKhOoeEFpdh7o0J7
3owtFfudAup8AZxE2T8325kH80NjG+zz+t6Mxg5PXZ37KFtB69yW/MeXIPVcJLRD
y9lZnuTVolFKLzbtReMWrKLHUk827gsaeg5tdyDAwIpQ0q7xMtUz5jhv4OVgkldU
PXdCOGfxiJe8wZOctg/FZw/fSqn1PWsz7R+UGld9zBMGc3GnUpDW5VwEEX9bbfgL
x0dXlhtGNKgXKAgFtekdfXZefMT2oBtwh5fw8jAVwkINGzSwIrEDCt2uQQtJtBEV
dBVYnMH8LXXuXEALbxiqDk3lS7ouxf54JFXBIWbqFgGSV7JFUxBtdDESrV824jqV
YQlIeNcSevLyiLS/QOOOizN7GBkpxtU8vCnvfUw3RS6DxXWBJm8uTXkGYdpr+I1e
y6jmgsgXBPbOX02D2ko91XWQ2UeliGSkNDGeps+pGYSsh+a6nlMkIhXqk2fs/0JD
gqlnxKEbcdbHEpxSRFzef7lxREVbnvxoDGmtZS3CTz3/BL8ZKohU3+anjYCvlWLj
ZXZmxK65+rsbn97vk070pVjugBJoGUqNnsxTqXbt9DlsDAvCHfKIfDgrVA0wND+t
Rb9cBXJ93Z8hXBI6+qeSiRE0IrLZeOWcRPUvpBAl9qdOvtwRN6TQIQOIfKIjXaNr
KkC1g+MB1iWCBIJKzLiwgYgTJLScWAnJFSayvpEL0zm8I6V9g8BYh3+d9OJun/qX
Fxwel5DFGyBzVv8ukACvdAOVIUFaNNU3664wRu7fq/0BOe8NWgxLoVelwcN8b2PC
NNEiMZclq0UKZhSzqCDXJy1l7BuGBMLwHlwQ0VM1hhEcGjp12GE2Evq/SsKLjHYD
SVPP5XcS0nPjRSS1gPa1BnSs6kRU6qcNmXiDjmNjhY8ShYWm2FbsYiDj9+5jTgSI
B0IBpA8mwZ/wy4cOp2v4HMJS+qI+bDcAfamdYCKMnxGEjQpQ6pV0HVDRSJ1TueRH
hbWaMuz6+6SzymAAyDQkgdi4J75MEPvddm3OZ+xMnlinbb9oS5p9Ntwlpt2MzKwT
/7lGV7kECZ06cMkS60e6KMz7sJ4b1SdiY1ZlWm/hoCjoY1BOoKdhCf09U7wDqvTq
d+MgRxkuxsZHq4JF4tZz2dptx6G45SpizOCwdpOF69sf7/LcbDgFMVlTGBeNccUk
c8SFkDZGg82ChS63omQMqRDIb96DEO78uuAEsF62QU2L18SvoxOYk/rwifbfs66F
utbcLZ5uAwZ+8AV1tAGTWFeKgluH0hgNFfryNBxBsuPNaNpnAHnnnmEl9Zs+ea39
ftFLwcDZncwP19FjZ/hke1Re1kIiCve2UrDofOcMzhdA+6iVGir5Aenbiz8vZuKK
C+nhAUo9u0VWDUBcsAD5lpZLN7Q7dou7KgflsNFTpmctrZLVqJUT06nepOinuAxt
Zo1EvpG3i5zApPX1562orONOUky9AGnNupGz5LpNZLbYF3X2NCacYJsnd+VgIVQK
HvjWGx3u233eAGUqib4da9QRBVaHz3xs7KZWqdK4UDANM6cJyb/caTuRxNSYGyCp
moZ3zlzpx4EZ+dUP++NKhfai0SrlD+l5iJF/3C2mCMOUe7LE0gAINs3XdMBQRKYC
p2lHR07X2cQxH91jErGhAKvu2ZlBMl93nI8lOCJdyh6Sp3umqfnWeryEMiVKFCNX
hmmoCcUphEApPiv3U+/bWy43RV99lez4kW5/4nTO8dt4OQNs4oD24rH6TDvXdGAi
Zcfypph1QFysF8HlEGWkR3eIvifOhOtEsCL/gsxNmOM5c7oTkVeCr6fkaPoeRffI
cyuxo5ivDjTHgK9xRT+0LSgFRHY7vXDZKoAebhzyg5msRQtN0WDnzaD9Dvip6XsC
9Gic0eMs85yUwSSgTiGI9oGG0y9yBJa7QMQ6z/35yn3vazF5ZQsMXmusDKH1UpDC
U1RkfUFern364KYPx1OiHAbXmSQCX0IiAmE16vl9BLyOiPDAunLc4Z0l2nc98Dv1
25ri7v/RS+jlpXFG7jGYZnCbH1QByCnXYtEoHTWrWuuryboZ4/nyfiiB+f7+0RqG
8ComXYLgFqkKPz1KjqZMF5yvKoVX7zoY/axaF53rG3pKY5+Lf46Stp/XVMVk5WOs
6xnp2TawEa03iMqH2Svw+oOOKpb1d7SCUs2CiRdLbyE9CWRJpON9KqyYu/O4WXlC
kDDEm868G5vCxEar59rgxe8HN68N5VoXwCziGQp3WAGXLXGe1x8R66XxYx20QFds
CSyvacb70ztEl/5BWaaWWdcZLTazK6QoQ4d9jhMIMawxf2uqls8WjLmdsBGr8GJ3
ZZdj62Xz4S3E4uTVWmXoZLl29n9edtItpIbm/dlHaWJ7h3OxSBqKF6G4+fhBX5Es
tVnWt9pw8b7UKXFxntSlWWHT2817Codt/P8rKEGANM/EWbquAJicvcbfYB78QmMp
xtSEAyQbiPZdjI55AhhAN6Tpfy4KGj6p+5CyknboC41ged5XuJR6yfOzeZB3QeGU
YH35TlFbI49MOfjkorCvYaH8xyaPjcSqtji8l9yiS2zU2o/1V+r4MEk4UB7Z2Ipd
skJxiEDzxSpVBLwjnK2rRO6fX2X2PHZcSjGLyLU5jKMFWxSBy1X93JxJ+cUtP3re
sJxvDaHofbP6Mr93KIrbg6/79EeJmIYE5WWgRZWCu3FkmwYqXuprhIMcbwUVS9Vi
vRJzWLP5hC8PSWXUid/TB3GYMmMB1NoXX+tWgQJJv2Qf5r/8/9IZZQOztSOhTOPZ
s0QOa3EHUIbTn+1DfWao69haCTAb7VtJWu4bWBR17bP9M42E9kiqniUoxx6X0tP8
SrtrRd7xt9PfxTWvBOiIFVxq7cu8POc8THWxqyYwxRm05hnZhYdQQHIz1nV4+Qf7
cpq7b0XeeyW/U0mZoHOAmG8hNun5rQ5pVnDey8pKB1lbfGGmJ5vL647tfRgZ6RYj
sLAdHFF68bTzJVoR8sPrByTqsTky/HBNXVQSzDR8ymFyGr3PRwfaejaeI+kseuQh
vHkccAUSDHN2nVe3puULGMErNc2ZFIWRIIWaIr4/IBf+8N1x2+ByPFytorZqBakd
uXgDLGNvGyGrl9gOrvI5U92g3MgU0oFUlYQybJTt9WmUCo9ya22zW3xxQB8c6lbK
BOxbF9cTEO6YA35cdgltBjoYXeGw6VRUUeHzbQfOxp5lHRVm6fH9gcV2XdEdxJXt
lHThMtp2ZIh9KHBXRtfXcBymIukyhzRhvVpeMa6gsJnqPVvkCeh2uyFye6kb2wS8
F0aTLbOJFU3bYCeC9nz2HkW8yoVsU1Lo+jwNlYLYSAv7RtuZdtuc8fX4Jz12DZ0x
P64o2tMnyyuYllqFOiTo/Ker3w31K+7EAJ6A+3LgjV9cqqbXuNS+4Zj1l1TACryd
JmZNMrPdG7a5FYptOaYpBzrw/8Ia9C+7kb9TfkqD9FpnfOatXFFI2+UO45WVgceR
t23sg0EJ589BhUVZr5iQDy/W/lBoaO+KToTJe0Szk41XqMexySDo+D3xRgunEGGN
Xyem50LJBhjl/ZOS/rPfKDe0YOmDDmlVBk2vuate0V1e1fN8v8ppze0MWLt9PWKw
xsEYg69RmUJNJ1+I1ZaUKmaPVeMIvjkuTn4MApWLNET/z/QBNmQbHljZkXkMuSPL
FQcNn+bxwt7nXUBUZYxUbhHHFHsF2qioq6ZrU2EB13a0ocUyU9i1MbodGDWQK2da
ei1/T1WqWSxu1pAUY4UxFAUw8lG8Po3PQBpgoNhq8xqLNpN/Tj8D29xR3BOwSLur
9kcMzZAoREk7uljXQd2TcNrZN9JbmMr5X3idlj+dPbKbeFQrD8VKInTn2lL5SynV
sHeCyJWuBX1GgLk8+YzixOVi2KTXpaxW+upTMaUvUccAZOvuR8PnRHm1xqRHMm3h
I1uw27oFw+WHf5cV5mVyT7y4aOupqYTagsYhW++NbZFQLmfdIZiRp4mrDKYqjAXu
KO201yUbjVeaySpT+eJ1skAf3tbJZptma+9uV40bnG5kkNirUfV7id/VLYhlCoHr
AMzYtsqPP7cehXSPDO0LVMDytPKUfeiN2sNA+gR0a6uw3dYxvKrg+Lt1tEvwWOFz
U8oLMh/IurcHFcBhrxxN6JeBBWg67ZgLKUqPM6C3o6p5yc/BBI7K9wc3oOY4BSb9
plmu6d4QNfah92yPOa8B8sg2WZXX9dnR9L7d+5xu4BQSGYH0G8jC6Hpo7nUIq18h
7V7JxQHkUTkEPJNHXNqn2pKjJQDrv2qQFDJT/bmbfb3XRrh/TYXNOqYxSSRUfhgC
eUV/OoMQA8HvVbsMIyFBsqT0iv0lvBCnFXXVXgRHAg4uI3k5CvTrodtdtsWHl1pi
D2PZlIGGIkE+n4BU+NuO2tyO8XQc9QXKIfHc1Rc+nwYTCGMyjzmQaRHBTuCGcDMM
EaRPhHdKj0rd899LMzJSViA8+trOXCGMkzgPV/dwCKb8RYaW7X3E74UWtWve3uHa
PCh1rZ5asihP94SbzGTK3W5bykMDwQJamdPUvhzNYeLYCV4f4MlkbRcBS5CKxlhi
pRl8FSQ+FfsTIGpKmCVe0t5DQzkON+/msmVe1DGaqreDIorsM1Ds4mLwa9Xhtb3k
`pragma protect end_protected
