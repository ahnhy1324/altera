// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
kwEq4h7q9lQ9Sqz7MKqy9LSvGHJWd75fcg8cBpZTyKWhjQL+YFcB+JKbHjSIldeU6iawuXawAN+4
/668UJ0lQMGWUzT6wRBn6qdXjpSS3GfCoQsz8WWuIx/MUXmqiHYgxDwVX6dKlFY/qdkHFf3BfjiH
NzZDwkuXIDK/myk5am5HiMCHzMIieBbcrqTNSL6eJcHCtZ48pnp7UKBKudgYlKhC6Q70jBdTeyCm
YaRFxCUUm8zXYZ+eZAk9tduHe87F3yO75pQ8lAfAuaGXKMLOMNmLlnluJUweDUCbcyitb1E2sPXZ
EWbBqTcp/+AJ6oRQU411DUYW9hUVtiDen8X4MQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
3mZuNW56p8H81xgB760gjJxuvehwjxzDjlNEZod9XTncOp1UsPbKzyvvxpfPcvamoQ/NMjpvd36y
wrczmInQHegv/Vq3KGAaw+/lsi9+xVU0FL1MHIq17dYRz/5CzIdMHNOKaPkXfaJC8F7bd//5ELIc
uCSuafVMr0mLCAU7yj7CnJO8ZvBQrWnveba2lBxmijAUFEistfzMX2X4uiPxWXTTx91bvpjS0BIG
K+PEfH+eGvm1CAdfE/ay79bI2pGEJ80lhkARUOSrbCOmAO+5z/NFraRMTrkNgR9NkJuHW3yxs9Jn
33L0+vreINHuxJ7up0Aid38/MerP8UrZP+zXLuFdbmL9JTHlSCJFGRq6ngThSO6a7cSbd9jfL4be
A2RRbC1BRGU8r7yQqbkdl0lZjwAuJA0MHe9OS7TATZuaFhN7NpBRBkvZzJmEVMEs5HXxvadDSw9V
jFvdm+CdtOR/K2VVLPdM/oSUGfzIGAO9DNCsOF4UoWIGmuc1IL9iafNnhxL9vMkDBbnXOjBwrtoW
sNBXOzEuSH2WNA+vArlOmsutdd8+PSe96dIqhyaX2pab3SPBJwnTEA7HT8Ctxj1bvyONnj39uXmv
1T2pa0bxupf11zsJBMuAuDp4BszkoMTzb8whWgrg7uO7hIwpnb91a7lzJ9qAxNBMiqoH3aysbcwj
I4bcUtE1kDsk8iUAWdhUHt3OyVhIbfSyDf1jlmtabTugAG6CvB+N7Jg0LCqU44l/7OAtPd/yL6Xf
RNbucrwF8LTklWLFee3ginyrDi0pVak6qTASefSiWskRf2/aIPuaDyv0ImzDQv7lbk77p1uq4hh+
ylPBuz5DU3XjE0w3OdjfzXrjdz1q9FJfX+nC3t1z7ePpcMQrkwBHhN4KT5LpwNX+nmu+OguPQ5XN
rH7+BbuYl+/2p8pwIfNAwtaJ6t8H+DVbzrin7ycf3jUtMzMKJm/JfGRjLgT2tm5hKhYen3C6ENHL
Tai0RJIFuJDJQ/G7pP5t+aqe7GkpPte1wEWFxISvdnu5LtoUsxIUVzW8cN+DLJyowMecVJPFwPuG
gYnEA4iiqhEJHe80D/7IzAAKx/miBQ10l4z1JfRsW7Pmp4m8NgKN3HoLOhsvvuO86V48GwWPLpYG
KsNBpEozKHB80tX884i1LzVJTCoTK1zQQVV2IXDBgtK7jmcCtDUxJpPR+TEMv5/1y6fE+pkunr+k
M+ROhPbqxiGA57aI+c2CvIF+zgJX1CwkXNr5Kg/lvsFc7RsVE66ZgbKr9VoUB8MjwQxJXt9QOIf8
w0Zfocl8Qx9cZLxYN1yqmmNlcWqKFHw1p2s8gVFxW2EOI14tm4kh3bEfnyjfmtg7+JbTYtDw+AKw
VJDo5A7RCBv22Hlubr3ZQx+DsqL5ycBjNNt1aAzvgkIovLd86M4T8bopfrw1b0LZAEIUysXKnXQs
5XQqehewmLN9AoZxm50PZTqLuMKFHuqttdrUcZz/oR//6Dl4amzgVVUzwt8QVv+hebico2NHD/6x
ix8h+Jz1+1LXMZW9LpjENwE+d7KWD7TOq5kISdGOkH2iROAPFVUqGFngzVvkjqpHxAQfaeiR5E3d
d5smpQ89yxkqi5YtUaG8B5NaJS0Pj4zaL28xd+0X/+kqD20f4kiKtvgfWs4LN59fmfUelL1NEuLX
Z22F2wzjGHzjIci7/6PcusCVu2M7kAtz9Rhf4f3487bSG6wRO9Lm2Z9tN7+I/wLRiHrO1r0GlQ1f
VozefgBKIgGAzsvMf285rCOfLfghXo2DFXUebKxPAMUt3a4DjiIy6EALsDptulDmUBGQK5LN1S0P
+0efnM/0MKqqi6NZbb+5igZDbermDyU8jVdAq5FjQgE+PWeRmpWDjqLtHAtXIoH/QWt44Mly0b8f
G1O+U9KtcRusNK8AetZ4eLs7x0AYrTCVxuyUVJ1P/KIWd6wRO4v5jjdz9QmXwsXwVX5WIaj8Cg2v
y2uhHDsLs5A9iTFRs/13ph+avxIw7ideWVQd7gDriWh7x0+b8oc/d8NIVMfEQyFpgmZzSjfjujjl
hzRQELSrw4wYai2NJ2jZsd0FSRp7SJrqJQQVbrL02cP3OnmwxKmwYLIMiVkucwN3TkHwkK4XxxHa
d9C2GgJ7/TUqcJlTF52Ch9WKCJi3c3NABPfI1GDhj88GQiVE1f2JqQ7e727QVUBsfpkqAhKZYcbq
CcinKf+yPCUzxCS0WPU+GXtViGj7o323i6sQyD9CSMrpJCnKivYznYYfiovqhPJMtIfwM3ZfGgTo
z94CuPw00zodbp2YIl6N3nOgie5oGTLrf9uQHhQeST67akkIj3lo8b7ZUBY2w+6UnfbOGdC1TO2Y
HSBWxVCDRJo7cesSrQuvTZC01WGfm24PH7dCl6bhm1cOe2Q5OoVYXRKUCUiubRCQfyyUi6RX93Gy
j7cVfZ369TAxKtHAoA1E2ZAStQtG7gqoxYuVbe6B13nOFwSA02jdy5P2BOUOtnN6n7uVjyOYrTpZ
jU2mWO5YbP4InlKSCgC1z/+DHa5hKeLikCTMmTD8Ru4zeNEUdztIAI6IRsW+bpwg2lpV9lhZBW7A
deDA0gB/lVhYvjRNogWoUPEBX/G+l5lZnIbkW9KkQJ8RidXEhDGjOd3xsGPj+zxcJ2CQ3IGygHVJ
iscIonfkPmQ3jnr+NTg0oFAJ4INWWu0wiaZwekhd7iS2WGUyKO2NFdKJW3GrPMm7HVos2Ufesp0q
UE1JT0DCXiD5FtLG7mYS6veTa8+8Qfviqhwj1dj2T9IzkDrvG1kxzdWm4GQlUkxPlagbqsWkAD37
v8FsHBUcYbg+4G2n1ZM7XN/rGKoiuyN8qPa1wTYf8c4LhGohCAZgy4NnxAWJV6Gw6DyWM9JYHomw
IMi+j/LqUd+8NPQOIug80eaWQrBRl1lBDtACaXxI/F/FIFEHOf9CDlDaS81pg2ccKdEGLuIxKS9m
oo5lDUuw/ntrHRwnzUPi7JUwhQeEVvYUS755hN73mpGl/8sqPVr4RXRQ8K1A7RDkb3/saOGwnF/T
LjkLU8XfTKHvHueg073bhXJ15DMmt58O0NEpSFGf3vjA5WkRL6HMv335qK+SuWMy668/2Bw5UJWT
VrRgJtOGoQi1DP57CBxix+ZfpoXmFYXItdHYZNhOUBkHackhQ67V5fq33hMJ9DFaHTB6IFDCjr2N
pJePUcX9zZwVQluPDrh6f57xZdro3ZND1k9iLydO1VK4Kc9snPFhlAbgHgXAs5gp6wATAFGwMwz/
rwNPXxqMdfrijLmwvFXxtfNtbt3garm6l3tFbZXhhAmSxsBVW+fy9jnk0lndwDfWQ7nb2N84oHcY
jeu0CZATsZueiRx8Lk+AsbtlpWtQuprU0YzRMmgwGLX5qpKTw0hR6to69+aTdXspxM4HTfC9Dxmk
/A+B4PT8tJCvMi4aVEtqu+a8m2CzNC7OFVnfanWan6UPSChy/iB0gwc9WZy7t0PyRnP7aOBCsxJ/
IqcGKJdtjcyLASXtxRYDyNf6i097h9ykFKfOurtSOsnWpObYdW75TJ1kpdXv88+tb1eCmOyX4wwD
NRvRifbKb1e6bmOOV140oES4FJcNR5ywCodtKuVqzGe4QNKG0oSALRHR4b5Ao+gMtasAfLN/KIiS
hEAFZTuqOnk0PHgqD8zdiHQil59Iv7qiTKMX3jqK2PAurfTSndRU4ETrH50Dt7uS0IgAuWsIngCp
PznR2+ZpLK/n2OLzxuLkZco+jd6wV7IYumc625+oWE/uld6D+T+/vKL2ZnSAEPvE2E0Tzmdr1QqJ
dWLD8F1IN+B+xTzF0jwSe7lhPjxLKetZhDQmagHU3Ju6qf1dtlkbrT8RXcfEoH+8rOsYIVxgQwgM
AR9choMupil90MXuHrn9tiWmTpN3MpJuRQNAWlOHjXHJJewIZJcM2GDVwh7xRe3F2a2uGY5nbTSd
Nn0YxHotezQITh5dY/QgJlvzSLY6KoSZn73mnGbcyi8CKXLSMC5qr6dVhMNQs0P1MkRKVciT7Z29
uiRtjYGBUJVxe8GgL5s7CWk6RLnSOr4i9YJuh2Jcwyfu4fv2EPysLOsnaN08judKhaIvL6qyRcIQ
xVXYzx4klZ6+p2XtOaqeuF3o7QGek8xq5JVW06HnCtxg/XlKYTC3bCUZBne1dypr3eHXwvXkyb+f
8ZaxRNnaI2yolHVhNUlun3Nxap/zie8C4Lpcb0clhFWRrFLW2rKYV3+5TVQEbJmGJcD/LUkOBDdl
GEW+N/QdMv7vZqXBbTLAR0YUObg+rP2bB6tb1dVzMW/so8pBRZ6onwv8L4QJey6Uqc74lUApdLUK
l5nVdpjaDQofDhQ0QPc0PU5u24fB/6XYs3o4Wb6pw+ExNXSPdIFJLOoozt9g7UlYCwCWJZg5McRH
OQThaCPpoFkW/93WoGXOnM9hAeAMPItnWIASCqBdiE3SzXJlJ0araEex4c5uBkin+Sj2zd9iS5U6
T4sIT/s7swTNXBGGp7+v4HKsV/kT+nALF2i6hf2m9R1Ys5HDGRwQITVhf0gP8LhOIKmFVh+gUwbv
jQ+BKF37ymBOHogSKErE8ooucDU/gcAiCEud07U6XAdUZm6GkplrXv8P+sK69JymntSOomz+/MXJ
a6QR8TrD82WcHYmkZwWdedVolzv0p83eVigse4NGuL7loJ6yziP/1U/ErzgH1u4rv9uwCJoxajSO
sZnfZFzemofQmLjF3BmcpLofpzmXcK7OMTrRmeOgkzdd0hQ5C7Z8XN/TUSE5h5EybayNyq8tgnV8
iyhwg7qqWCRinaVyaciQjfAoY3Oa0NuU5EjJYeCvCiJ0dkKZiwGqT1cqh9pI31aJeO8pWdPDftWc
7iD6pcOw6+6hige6/ZBnhW4zJdJ0iOdR864ntJeV284+vrhX8fYi5GgVg9zsMWlVOg+uHJfoi3Rd
fWr2xtWR4BCWPX9OQi7FTixTtZe6S0yzO+5jH3hvmiBrzaPlhF+4v44v6Skf8C365u+FU/lC4svK
Q0BCJYzWdg24FMuW0qLtwyhCAoyvXXt82TW6LBbEEYwHlppJpzpmyn1kpesjFMFwk0KzFhRl1S/j
4l3l3SRP6hMavkJmpDPmGRzGdXSb5mSBkJdSpgt0klKpJLdysRw+YuVpsgsrUs8U72vER+guaN4u
bg63jl/5yDpIGUyZoPyROxC+InVU+LFAIjnbrOEHPNqzvCrY/JPxfwVSV/u31S3w/wr3yRCo+qW3
Ms0ka8yBNcL1aYRPESGA0juMbykiMFycFxOcp9wTjrJ8pF/NgtpADNei2FpTgu5U7uRLzKYm+NBC
Rwk+Iz59BnGVCKBbZ/pIk4Pyh1oFpQ0l4mJQlFVU5J6hwnBhTiVvLpucw/u5aUcqMC8ioKfpTrTg
SxG5pLzDThMGtpNRyse6QAkfei58yTs3pJWGl1U76/zmTPNqhYm9QUgXo2tEDNsL/rdxa4ttxHdk
B3pIP31CLqq/eoBAzGv+bjUFNbi99d8pBiZsHv/GlZ6e57Am2dWnjnfPi4cjjTcfuevOXw4Y6i+S
/9/YyPonFHKYDWg1CfZVoMte7kO4uLOGbFelTnlXW7UN5pfSXfLVCNeOGlqQhETzF43bM+8SY0G5
ZlFWhEjPeH4GcxrZEiBg9cI99V1H3at5JTHr6AbrpJ3GUrPAnp+0FS3jUN9jTXZ4xMSkY1AtpUT5
f5+wlqLemYwdQGrFUCeAZYfZcwuTUyC8xCZyT/htUnLUEDcTG4wANmifxiWi4XdTtwZrl5hWoHS2
aHOgPZhGsVmJVQJ61yT1vEIZH5oNnrUgBKZH3LY05JANNeSQ4I07eop2iZXslmGldq9WLnd4/Sau
IeBFeeKi8Fa55E61vi/ShGGDg/xItgseiZPDek/mUYv2H96bOvOLxkws6fsd7Ow3vE5Q7DG8VKQf
Ym/Zdhbvja1BXFbIfQnVle7inWtnh3fj4mkwlHYTJPw77e2DhydXA22THl5eW9cJH8lBIGhJLlR3
RaXFU74PSn6I+qiAn+O+KEM/ZpdiuICq4d/UzoeogEJj5Nky7rpkElNsJFPuyqV4k/6g6n6j4z16
SuH8pyX3X/U2aUMzwY7lFZJvrs6ZtEcMxUCJsKg//gpb+6NODPgRs/y2l0L2ObW8t4PWFbyG6Aty
7TSvERVixkZjg5TvPEW6RQdZfvg7cUedSNS8bKIPZza34t4mgYFSd7fzgRYryQkB0u+MfSZImrnk
6ya8RWypWPcInkEQvPZshQgfRKblicj8nnIfYJy12n0tXWuGE1brSe+0solCvsUNxHZIv2K0kskt
FrZu96agl7qHQcvDZHE1u0KgzRmjDj2+cztM4G1kXYxLNPBC1vReIIzG8SmN9XciMGwRAnGFBm72
w5eprUZ3rnhG5/Ufl3f7eTpN2WgF0Mk8GQqyGOms3vKXPTZsEQBcr3w/XhRjhZRryqvcn67uClgm
JPH9ieIcRArjU9Xh1Xvz8yZGd67DScRnuEa7fJ6A+B9py98QQwOgvXP+5owuFQ2POEFFuIvluPw7
KBtijodw8jdrtUOKORhr0o4t0b/pNZNppPFzgvJt4z6u0xSLVZ1DWS6NuTQdXyUnriTi+J9mINb4
mu9cZeI2y1el2bgy+aycUja/xS9PITljHq01F2g1pdHi3s9xoL/YjA8KWGjdxDFn5sf649nU0uNV
B9a0WJ7s/I156Q41kU6F30y77kDT8UBmzQAoWqqV7R2XJAnu86HgHBFaSzT2WBoYWXy15DQ5lmIR
Zg9jteighzF9H+NFdXUrrXQBKgqKlabaGBqcv+k3Mwf26FDZsehD+2iRA2zoc5C2vN1Rq0Hav4Ri
0P4NoKEvcCxSC6Fkl0LBaR9XGltsQG2SHCA1E6xUzGN+P6T9aVDHJF5og7PFsi7N9P8LswAY+wh3
h4HvN61IsUcZS/UmlH/923i9T8N47KRpbOXXx3CjYp6+4pH0AlYetqsIW6Figwv+AKZe2YmeoVyS
wrZDt9aEP3JVMD5n6i79A+myoG4KOhdXTgVNpf8zGytW4Feo3EKiB40tqmC3p8GUBH2nR3SeWDw2
EX4WVtTRkyiyYKK4WuPqMXW5ooNEHOlWfzTB8wYKJRIzTWbLs5QxuSFbFWcIQbuQHLFCrnpIRjgq
IrQhUFuyGeLVKbENeamegIkkq7OpdvujVbMC3gTrtnvlGKSNdW6Cqh3Un9/oCmo3l/LVHw8W2ZtA
7i2XeyGCNcgk0+Z+G6H9bnYvPdXqkv2XoSnIeQjK5og4HghhFx/w+Yjz00BD+uXv28UfRWG0sP7z
cckGbq5WYfl2TBlv7iqnyQYBGIGI7Rx8AOlGIrgi7/vbXy93Lvkmr/QshGaS4Nkq5w/OhwskIp/8
NXrTIQOiOrlYirjD7m7C/lQ4gf0X9thHIsRWHFX2M0cxJljqurIJMi3cvHnQBUmLGQ3qFzNWYVZp
l/HdYxPniBoKsZxb24lSNq1hgoJ84a4b4hnKk0l1STjANP6rHY/T9braKXZKgBHSD22fymNd7i0S
HxT2JkfYScGwjmPU8IWvb8TGy2ek28B66JIIttMpkfw8NhZR1wirAe7l092KLMP4sAeg7XgI9cKf
qbizxpX+JAeRm5j52Vlg+2UcIN/O6GVLTy6w6Wmyaq2CULpyPrWSerSTwnh2gIWxws5FPJjR1e4K
CaprMmzKtPAM3rHispnP7v4U0/poaq/zTtJBL52ox8GAPiMHpQx4oKCS6pMkmFS4e1SqvE1KzxJ+
zGcioShPgqXkxzyQgH7jtZtFlDc2fz7rWfpDghrxGgJp8gkNO2f0AyM661TcizJzJ662rH4BpCXd
B0eT3Igy/mHgxWgv+xeixye1LkpNfqunm4nfZNp+yX26lwQDhw6LeDBlNBuGPx9qOJB2ihADXTd2
ZxxR3zN0C87qu/NmZg+ITZXk4iLRp19tvOVvFWJp7m2AkVgHeVyw+NdL2+u9IPO0P3nBQOKi/jW0
tOormC4Ogylt+TPDgrqnO/2FDKF9pXJOHGHD+GQkwB8BZt8hpbLTy16R+1s1TQH4T5L2zOw9xSOx
y+c7abkMlQC4EA8uZWi0XMjNzaaQOdnpy+GQQJX+1u9VFhpi1IsrJVsi7HY2b1+8shh+iUw+jqW+
pvWI4uQx6874in2YOJXz+KRqJD5DPPHZ4ZL5/CVFTY7D650K5qnrEG+yvt5LP2ur+/3hStNwkjgj
TFRcBvoUbwYuYzK5cz3QMVIABDNb3iO/6wdArqm1ofq9v4UALux1qAZjCq3U1OKlRKykJ08k3588
UX/Lmdb20avCqX/oeJKxUNBseBbtvlef8lGysz/TXQ5hDBS0uzVs8+t8M4lR1VctN1U19C0ZXhSp
3hM9WGy17t7sNp2MhnEKt4s19gZfvYF+3C4gEcq6ZEzU+kdeAqT+pzjyEY6zv3SU6UGSquAdF7vo
XTKjHxwi19sUpq48LHoNdVEYVhY4J+44DTwaBAtEXsIH6vRkWFiKwYbdYdRRV0NpUQkOY1wspPKO
eT3dzbuikabO93bbn8pQZmVa14NWwkcAIjJPAxs8582v2r6AwD2kY3H5Pxzxi3Q1QrJaq+BM/Ie+
/gcy4UpVc/0Sk/LDopj7GBZtrVQGBSzaQxazczWW/KSFeLCS0l7Cio2CFuvCxLSwgLiW1m9LqGks
Aq+0aC1eAojFkCoOjtmrd0N0B5XYJ0NvWm9avXCk5y6LajCBMVWvYO2TsshkM8a0LZ7IyVEctSAv
+NRt+dYFYow/kp0Z1EjVCCAGtOC/DwviEPcEMMGr7Bgyn9OGG3h0eD8C133ayz5ime5jXnvlU1JY
/2MbfxlzXNi+lAL96R50w49fTDQF9/zjI8vK8hk4NoByaIqYDGGVdHfLZozDZN2w9pDwTiuyAY7e
PvdBAedmTfQk/zPVZux+obiYI1qju1if+BbFB/FrrjcBUjJnf9HJkLCwGtGLJbMwXnqsseqKfX5C
hjTOtLrj2DFut0FvIJAqJI3q0HeXDp0pDgt3iT1G1u4tImIXf1i4NV5iP5hYyqKUF5QEixmKsUlf
taqUgChyUfkXpcV6p40zzn+IFVslE26HhMh7qkReHOBT7lzyPusByyR/8uTN2plVFvLOLde4My8J
3FC2GPyBmpaizS7G0Vx9E8CmtpTYZQNq0hULyig6bIL3inDC+TC/M0kz7nMWVFso6pduN9VG2fcx
GFdwZ8goyedlwgLFjIkSzR/WDLbL8PcCMJgrXlH1ARhRLtqOShtpNHyxVrO1wEZZkiVN5PDvwN0/
udEa7Plz66FRFZrT7kPAZJrlDI9PJlvvTeH28IAQMl77tq6T7DjLf5UcWpDRfCyPOnDkkR8aQFUs
mjpwEoejkh5Rsq02hw9i8VeUAcXiYTHQqV6cBASkW4bKYyM/pk0LmRG+9Uf5FLL3z1ZT38mOLjjo
a9GTCAZtC98VtAHo1lo7yoqgV6KtbHiq4jv9oJXJjfC5pEW1S2WNEmNIVTofznL5UAzMpf/pSRYs
2pcBFJ1jeUlw2dLfzK81KBi7o+q5odegwEz0QCLS71a2fzpH5ENoVBi2E1wdEgUPAcd2ehZayvXy
oTljOQN7XHptT1ZLkmmG5Bvzf4dfxzlwJNIMw+1ttdVMf3qBpucxj1tlbsr+8dUCIZTiAWurioXr
X8YpIgxzOLeTrim8fEdEB2dno15+dP3qtycKxlLiYlHyF2CDO197HQlKoBxq80Avm0iHnDthRVgf
gtAZ9BRTvrpGeT0TWjhC27itrcG+SdX0R8c5UuB+K+3TepmA+y2A5vDuv8fHIRnShmiWQp4+9MFX
rrsdHxTL2FEvaL4wdCwhoGJySmPolDTZ1T+p4w85wrLYbfLxAmW0KsyjADXeC5vr8ru2ANizJ2D4
sNShCXls7Fe5bMn4YZc2nYpAfIhpoD23wYdKNldJIj1w1/owT8nCy7dPme0fwfuf+OX1LO/EjXtv
GTJ3jQ7YKjijQx8u3S4q1z1YDUlg4zqGBkg2WrjVLSLUCnFZJGBdbo8gEbhGxRIqUXA5oKwJG+B4
6thmm10chtB5yLEIP9GLKd+M+Gq0hPSIHlpMH2QkhnqV0pV/zLGxBcNQhEWcK0rsuYGqyBPcyEBZ
Bd1SL5cZCTLf8O+5YhIT5J396Ew70AxviDGTg+Js1R1eGOcF7BQI8nKYFobfJlr1rQts1W9wSHOg
RsUx2hhudG2zqr9UXX7uz5/VB/coFocVTK6Xk/6pxONtXeqQ4fr3RhOW69UMV1NV/+Zu5tmEnS7f
zkqwniDtc+5DqRMfr+DH+LdqK45+FHVovg792TFHVnRnRB0N+M8gdEySSRM9L58HysFB4Lpw8NYv
aM1zct+g4Pw1SYoigt5yNqewCr1YnB+sn3QCAxwxC87bEA3zw70TDAggbz1x6xVuBihrB3TrUbli
SAOZ/nOrlxLKMWQ4Q0awZpP45pg0kTXGpmMzBVm8+7hdFqxatY93o+u+573v2Ud9czeFzAzeBPrI
kzWvLniqFwNIqvgOFKZnYGl8p/BBeTE4lJB1cU1aTu8dXlHQsKhL61yzAku50I1L7vJFxuabEGYH
gnX5qOJgOqOTaAIGCA==
`pragma protect end_protected
