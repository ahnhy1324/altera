// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MlLZiwpBKX/WBrjP2Fnh08QWZ5mVQMtmg3VXhYMwAi5TezZPNtI9jIxdrxAXQEUb
R1sgb2jApZ4csCFHien2c5i4L6vfZYvU5NohdAKhcqwdNu22u2gIWqUxAO3S0y2z
ggq/GAHLaHwVCOg4O7Por2/jRqbosoOs5jKiWqc0N/I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9424)
pTrdpb3/f4YIt7AedNvJXzZfCPEKfTVQPIl5Z1b8jqHyG8rIxkg0XxTZedG3tQAI
GJNFSJ0S5R4+Ys7o2ikakTMis5v60MYRbK7WVuxLz7CXF0/nhh9deZAlcifwSNkO
HpYcU2UE6LnrOGNKHsAjNgP1unUI02uFNAUnV2fc5zwZ2N1IgDHmzsLGSXpuFrlX
B0ds7lzxxezCLWkpok67MUOX6mec12+OYuZNkn9B89HePD23X05HSm9/r+/jrWwN
s9Ugxz8AZ1o9xLsLMk2dEpaJYIWLiMlx5XR/Neskzl9uTYex4z9yRztagW/DqLNj
x4TnOSpqAvE1uiv1afYYx+5gDjmq4PRRD31jOgMhCWZoJP1I995IfyFvUxhTm3cf
mEiY8XWTCT1Ltg4mJqaR0iP2KJHAAXQS8aCWZB7q+kxcnQSp1lqXJOtPalRhG247
pN3CVV0HZNHBekHxwGIwPvu6MDN7CVYPuTm3LHfaX22kQ7de54eEnd7J8KmpoTSK
7EuCOoUOLw1wwSokqUH4lZURgdFhadReE83ci8CeoYbMIze3GfHIvuA4Lq1jsh1X
q+OW/DKngIu3hxyJBQUOeLNnWPV3PS3JtoUCXw+YLFQab/lpSeteh46J7ZJzqU8n
eleWBC+yWK4f8XCVs04Ex8R24VNJraSW15QLq+L2UsZX8eLjSOsCH0BDNn5I4oGq
Fz31HrNpBIo9zyUIGp1fpJJWmP/764KaEROrtkllJD7aBePRFBjMqg/Vvo97l8nA
DrJLP6camHETaSUYEi3yVepYloUwm+gfcI/MOI5hWgxj9qTpwgO2h6/y79yASKl3
KpasFvBA0B044aBqsW+sK30+TNIIVdZlArfLk6LuM2gn32J2/pJgZ2jZEmEGOJZj
hwg0F2AnTpMXh3upb0BIRedFeyqtG5D0N+m/+xaPeTnalBjXBm2/ga4H1Dl6qF23
5K7nTEu1Rnp5ahOXcy6gAnIaZeo5WhMHnkth+ReKwAV/A9NCPg6gFfn2Xv4QNWi0
8AYR/nddD+VAIQ2mNPZp1hhoedkQy31y2LZTAxu61ejprQM/28w7wbDsJrgjj6sV
DfJG5CWqjaQ9D+MOfS2auNGyb3SPKZBPrcDxIh4cgSxVnONZ9ywbEbmSdjufNwX3
BWOJ0c5CqtCLJOcx7qjasARu3YeuVpUZpU+qXIstutwV+m884esEjcS0Zn66qVpt
MqnEEqb6WrJy4L6Y7YxfISMdXdo7u2QJTwh9w7uGqYmzxXIUwIdzSZKFdtDVE4eL
DwANusEPVavk3hzyJpZN9w9dvs/lizZndlTphYCtiaqOfHOWS78xsXH3nIVahAY4
uAq3yxTTmuZbuGx31lmi0gZVdZIXhAHUuJPz5Rk3AOQC5Twk4Lq/l9aWs9VQVVqL
FHhII63b/jJynu7gqTUijZZWlVLr92G36YdPv7VR+qqQ/U0xWX+mt0kPUjopbIke
2Y26IQgwfTdVA+Aoz0OvPaQ28XWbBIThB0AQPtKG1KUrzHnuA608QqJ52Iw3E9Qq
DGdK4JEUvgsEuy8mThJu5XHXPdCSZW/tbmHpYg35CEMVS8iHKJYbH1dnQaHYotL8
wSUHAj9ddTJFJhNn6vYCqVlCU+NBQ0nPgVmPlanaLTFkjUwc6VgWY6dsH9A/NTWm
G5QZVoMqFGYeF1vMVrxQYetbl2nFCdtnPyLwfqwPDGdkYXUWgJnCJpziKowT+D7O
ZSMiA0tM1g5vP02Sj+s3rPR6aB47GN08Q2sanHIdx8/F6b0ZqvhrdU7KBdUmkuFK
hmdBxN65zkFr1OrgZhHygcDCCb+XZ8zbZmSiGNas54WTlHbKKgutmkacgaXv/hXj
OKvKpBwMASM18wZaee861VclB/sx4bvuTdI9v0jDSWumSBWSRBpT5W/OYaesHJ+U
YUJdjh8Z3uno1NlHIphY7gxkByiPJnCq1QUVqbQhJm5ISbaKJ03/Trd2CwSw06/C
SBzysEfA8XB3p2C7/D1OYfJ+jYku4A++IZZD0DNInzmoH+0vZ7Eth3FZTMD0GeuD
DysagWqJBq3g0MnAFdrnfJyETBiP2AapJKK+Z9+JZdJ3YUAymehArmRvpkeHg5NR
dsFrLPJxOMkdV07QR8GgaGz2PogfEZzUXRARSvABRNtLhrYHJDWwyUKADYJ5ojqs
ZygiRo0WxVXg5itKogpIqymhUsA9A6kVLlkgyetziBhcaZYzY2NUZZK5Kx8S2Yoz
C88GSr3GkGcjUbyVmfxay+hUobfYEWJuu+nVHXrFRn7+VMX/JC0U0pIolbb1hz+i
j1di+SVan79451fM7cdIQBzGG/pdW2mySGrFenZ+StRI/yxJcIQP7OWnt6hbCsQ4
75CKLlAoO8euHYZPgYS8t0oz3dlI7OuZt4kiopusYZwl8Z0wCjPKkz/U9cBp3iz4
Pa3MlNNeAtSjsiypC3FHPNuLXVqGHQeKmgBIPABXrE45waKCSZECJEsbak2osmP9
DBb+WxFVoj3CbZ67tf6+po8NjYk5kFUAsYtuKUNkmpDN/VfeBlXvXwW6jjZ3+PvW
CBbFvibRQ8qEYn0/ePTohgqPumafbA+s/W9xZpFF2M6aEY5juqFAvdyuOo/8AhFM
18OeqI3vDjTIlEgkj9tPK2NYfNdZW4VlXalnhEIDtZ6GDUJL7G1tSadFGG+iOeMz
HLE73k9mBOKiu6l0aEe8hM7QlcHsy8r6RGhuML9R05Cjt/PJFhbx65oVKQydZ9h0
yW16M+KiGM1AHnjNBklv8EQNlx0ynTsV5k/FcCbqbLJVR28Laifjc8UvgMgB5lKv
xxQsWXNh/CS5wuc8A+Wu89dUqTD+508O7b3ZMHUeIe4kSKln4YxvdWDs7UCMThWy
k1OQ4CpsYTOTpZQUqTuTN99PLoKU9fr88m+ZuWcoofk4S1HFKhBd5APbg+aekOzA
2TD/VaAuMYLh9VBdRg0l+qoBNYw7n3kIIICgmNOa3jyWmvb/Cjf3D0C9EODnpirH
E8l2uO9X7omnD+5G+yWJ7oST50ygtI3T41wRq+DfAphhwm5+GysHuH+Ynl6MOsDc
j6qRL/iaYSQEQdwu8jbcH2XN69ePY2030+waQDuFNo9fI8dhpZS/NUDMB3Prq8uQ
4NRIxzJDKBOytxFbFwpimldi5Mp3325qJKNgEbaZJ/33BP5oQ4VEzrW8w1ML2VzC
dTF21sM8qDA+V3Ro+6f3LNtCKhomPH2c7hOJc4jCoCRbo9O0krk26DflwEPuPNLd
a6X+VPYmh8LXFPMuDI+zErKiqTIWJGXI0nuegCyvrOb3GKsaAxamWhAPcZ86COK/
RiA3YSk/ehxiLMWIdyl2a1mhJatYN0crnkR/q/7Uj7aDu2n6F0nFpgeaJvrmKK2s
VeWA93NmO7Ow0IcYEdsBCYMm+MWd92sDhUWvYZcg+vkyDcPLx3jjMkdYtMqs7QjU
e/Uxfzkv9RjhPDERKUHxS8Vz2mmFh6+UuJr4pKTfhJGdraOh4pXSxISaY+PFF5/H
x9DNYvzw6ZJn1AXHYt7EU0/uKNmtulog2fnjKY4TtgEB/u9T8X8HXPXmHUR/QtK1
+o6LvoOkuPM3eQ78WrRziqrhk5eS1QH9SPoWLbNu0wsW68ICT0JVr8ve+0nz1PRg
ifFFFf48owgUBYas8aJlwLf8vZ7J0lzQcFWoFoor7S14FuTe8KRSMp+oHuBP32Fk
nGXLSB+OCjzG7YdznKU/5spOv/v0x9weHEo+9RtLo27/w6EyPkp2zVJf6iiGsOTm
nuwNnL5OBUIp5YTRXEvMUkf6Wf050BvdI5x6PZiJAFFtnVLV5AVEeiS2rEIC63Xs
y8js3Duh1msfKYEPpFz/6PT1v8fm24iWXohpZ6M+9SGeNEfInHGfdv0WaRleajvY
fFac1psdkKd0a+GY/LhWHl0xG9XAAIRpH+wUu6fexhhLhLosCYcC4Hr92Hjjhnyw
as9Id9KQbHtQc+5xlpcD/kK27Ul2Wbg+YHePVA8StexdezjGInvIgD0nEFanj7ts
ss1tyuyy965ke6w5IbYtXq36MfsfFKGXHSatIW/kXQfHXX42JGRMScHT/MZXrfQd
vsl5JSQyESonGYhnn1akPIu82l2A3hD0cc0trBIJCwp0HEIifAx4T8V7doZt2aU2
4X8cuXqIX4Yva516UbwsFXxxyITQxKsvEwgMgnTwLelpJWAjsI1TgYw3DQh9nmLg
RWuS6xLZ2JX3E0BWrbwCufl5HFmXqXPSCUGThXm0kRzFRHDihOjSZspn8q2xmk7q
ELwuFV1hC0tDoJayg7rLjx6QnrIWAm+lnbq8G1QPT18fR4i0MHsVoQV2GrFHoeU0
k+nqkMl9XBvru5WJKeJOar2g/yetECE3cjrjVlZA4On6RB/pfq51nsHEiWyDnP3Z
MtmZoFq7FZkgigiOcTQDtYGlXV7lqMnaBVC+ls64et4rFvq/K4BR7gJlYDU2drmX
9XoXGe2q4u9tt+Lj+u6bMCzb+1W2nLuUtqflCZMD7WA0nF9WtajDkljsqkqVk1Iq
YgEFwyuKGYURiTCTwIwzBImaVW6rWuYu6cLivrhpjkeKtSleq9ez3ysuJuvmI//X
U0CPw+O3IuB4aUNRE4DdrDOWCJ+OnBufRdS7eUZtHfWikX5vD/W5E2j7YoI5/CK7
2+z6FVMrxHue98QOzRa2QrRGoc5MAjpP/l1DsBuUHtvdmB62bis1oWsROB/IEj+v
hOApHnBZEI5XEBdTtdM/VtRPuGqRi7yqp0woM+Ub1sVhhh3DfFSn5/x27/vvu+By
AeGwzDwekW4AVQM39TMsDXtr/4V0A0+niVBzzU2C50FvhzojvlMzHBF/rdIcMzgO
N5Yxo71kegYj66I9Aj4z/be74f3RHoDVKqMF7BK3RxoLevhOBWz6+yM688FFZwzJ
XyaNAj/ZIuxlR5LwXVSeQM5yrGYIHEpB0MDHZeZ7rIbV/UrDVaQI9QxjUbQhIULS
pp4Yg5omucAGKgIxjb43zS/dCLs0VsOhC55Kqs7ktDU+RL8cm/+LRVgSsFP7ziu+
ojrvPdT/LTCbrcygLYUV3SKKeT9GiDYLnGiME0f+rvUyhHdsMqg2T946EZLZE8MZ
OXddk+8Q0GjToP/4p0nE9ffRnRLWqGYhXyvql0EsS2Pxg2SIFD+2DvYi+B1gPJwD
OSGoMs154nbXOdkkf8HiRpyS3Fdbk6E1qGwVqvrjHYVIHEScCb1Wq/Q1SthudXlo
vq0q06SCFNu2DtR8hnVA6Mu3A7qwnfCv5X3nbEwt/Bo60WN0mH+1UOpXtKz4pSxO
PeNS/CLhNoKA+sfQQ6sRbQl1mTn32rOQGOz7dU+R8+r5yS2eIyqyKZtbhD0QUPiB
WEVe+OwgoUJ4mMWEFM1qC23/evkKxsqlbdDKbh53DY7sFzVFREjJhhvz/QSGzddk
llUz3U85tcCSt68SSj1OxmDymkrzeD4U69exdry/y2yZsgH2wHjf7IG3sG1q8rJB
8N/1rx4sYBzDKrnuwDsDM3ycT5fmdttNSXzRkwrU2Xy52L1aUgm5gPlT3uBzwz/S
5FAOw1PUVh7Q4iGT4vPpIUr4use8VzSaDhii2fTf/z9qru5SpjWotzDGYwRtvKb3
rkJVQkd/SFnSCNwRAvpvpSno6p07AfbElVOrcGhc7IbXnLYhdSkxsc2j1iDpCFgn
b5qwUZCn7/2oR2sLVqLZ66KO6wnmqrdOK0LJpdHHcaEsi4b5gyP2Zz6ILTkHonep
gctJz1n1+3GryR4MFmCSbYHN9zCFHiAgDGtyn3TYQ2JOM4s+v03QbxMx3yClCV/m
U9Dh0HDaLZcrUVyR/CVvgU5nHGg+q5BrTu+j3Ua62fgcCSx0sYu+hIC2G82sxLzM
D4zl6Q1vHLsbadu4k1czNhTJesfVicdKN6zqmbhQl/wXJ0KZ4xCI12gXCQmMv1Ab
/48kPnMFAgwRIo0fQBbO6cWz+RyFb2TClVuWgShCbjW8aYpg39OcuGiynOozJgIn
8fLfvbu088yBMWWQciOcLqdba5vbmNGxze5c1b5JyYanQbotcvl+09spkxUqacU/
pWUbe9+k7oXWE19jz4sH4zGpg2EQGcbqg4DjH/str7TaT76SfTse2UxAOwitquQR
Zh5kUK5844O/tLHeDtarjdnyXkhmpWfL/tHgQLji34RT2fZNhMYGQHJvEHY5k+qU
8PNzymB3J3SFwrUCIfgvMVCqrQPrg3ECJUm/30OvU5q8y72NOLryw2VJJAEHn6mP
0qRWQTh22/TdRM6gM2a5IGBCR2jtpppA9jlIDDkmjXxZANMOnD+8190qHO18QdEu
4xlYttDKOFQ6NYipX4ETQVYnuWl1AdFxgXr7RK0ceZKEeV6uG5xWPpnQK2CSKfCn
sKXkn3W+8wZmcwe5vI9yOrplIbojt/O5i3xLTaRGUaNFP3eyyYEWj7/r2IBXkRbV
b1eXVSxbYQtVXkFx9NWNBUrQWBtLfePTe9dIEno2a3LTyhdu1MajzXXk06lUwgrc
fdGDZtp2uc455UJ1ACUn9BLJqGSmSYCYVpTlkdkEuT4sE7BlRHPlhVm/Y4HPxbZm
XjGdecprdkcfP2lDPgG4D0i2W3v4ARFPvw2kAGnBz9QhREPoOB5f5ipoXjWJP8HU
qLSQc2Or6ita1LCpQQeJURcanM7cGiGzlrIID/MMRUSBsZQC+eKmcqsxs7Vqf4kH
L281Hvg/SgNb7ny5wVo4wpq/yfyZim2YR0r89v8xZkFlIzxeCwZ83aWLlmWjYVro
Tz4WkD9lo+14H/5PnxU6CwZJeEKex0DQSKJcEy39Ne9LC4/iKTKvDyUd83MHanMX
xLUfpHnfa4r7gst5BtEEMu2I/fI2g1PMb5u5gMUv3Kz9F6BVwmaaP/6oRg4afj7X
TzSqvXMHsVq2JuRRXpJyg6mh8Vkkh43STpJPdEYlcGMVmhrXCCY7v/NIcUYQIDJz
HKYzpl7EZzIywK+54zndSCXgW9IsHZvCO3aR010WWiRjN5JbbjFW5ANRzCXmncW1
6dwbKlNPTYvVaNQ143ko8NnYyVxKkxEcdCWusAJ37fa9DwcF+EvvRQL/Nphuxu4l
g/1S9bbLWd+vPY4Sw5TL4amEp0pHr/fKvluJRNlDGlQYGE8xsZs2tj2kWCDmqUVe
EZcL2VmUNxbyyMxu6FVe8vZoQ96f5RACnH16S+kNwRAAadeuclHUrXjOV47CxVh8
AiKIr3mmbZZoTDLtHFhp84VKt2abyPZ6x6WXX8kgE4263IWscmRrRShozbE1DHYy
YoQEqJGGG8x3D2cRdxenKA06quqKg54y18bwBadUP9/kNrpOtPdfGRUbczYmgIwY
SVOqRWDsitaBb6AlIuHWa6lFNFL4RgAfK+GsznpchxeeU+tyx+yqDIDio8AW+756
DMrTNpfokPZSlhM9eCp6ZN11lFA3Q/xIcnCXZkn43gm1zLsYGODf7rabnvhxuexT
H09U65tB1Li+Aw5UXdzaGBjteAWXnKAfr8507SozK8bgBYmq4GfEVU2imAG7GLT0
MS1J/Sjikz/bMKyxfSizJbJ+1p6Imvk37ftHNfpvvrEicsshdb0dttGXsB+oeG2Z
3ax5RmiILzTL6iGGR9qevUvCBhRPqL8c2NO+hJSGBhQo1bVQTWp3fI2Ishl9vHgz
MlD3ylFTlHp9YT9uh7fGpMit+HJOy4pkyqnJ7DqheoLFnM0iFNFmGOxkAJ+jnsPL
Sryqs3FMu95x1IorAzziJbQ1Y+DRKrKqAeHPvu+HvgVWdUx5gNLX1qvKyn41Rlii
9CLEo1CGJLMx757cv71txfSxbtl21GSPJI5aHTentc2l1Rnxrv6DYDNEfvpCuvsp
BXO/vSbPDgEyR0hDRKKn1mE9C9sNtYRsqXgQuhF+RAeaB4SBxAkpsbtLW+g+TVSz
2PO77A1aE2I09+tnk91MPGgC7Fdezp2EZ/mQUm6A4RGXEym/6EDBFmgLhEJEsMTe
sMVJ6Tpu9Jjji2FSKggErcsgU68LTvGvhU4ySUKBxdALCjWt1LVPITQk4S8yzyu7
SsZQ2I3rMHHOIHn7WwLG0ocRsElDNTOPZsLEjcKiUHkYQFbF5htiTuhQ4hta4yrn
0df9QIV9PysOpNUjqxWeGmO5HSIX/I3o8fe7NsE57U6/kUKSFZ2Lyg6PKCZB4I9O
oP9Ul6Arn6FJ62/5eBeqkcDx892LFBtix7GynkQtZM3RZTFv4qM2aJtBiy/9nOJ+
ClbU5r7VE4/RxXY37hqAOiS061v+8BOdYYEfTUruwznjevI5ORe8PBr3mccES/WG
hDAQQUzM4ffVlTTF9M3NQfbeCyyM/WGlhIlNVpckipsdngBo1F8lXQA89lOIDl5i
aQYZ+aaAu9wA1tLnOisrgP9y5zDJgzw+geF7dSt4adpRSsATiWm28xaF/KqU/jUA
y2D1oZvphUhLngbLn1a/VZA+RVnenrZ8FtRdQsP4P9QVigAErwTPcJgeteJl8vyx
F/jzMbIR7p5+zEKTLch/u0Oeg/aF+nt52yuvm09JB8Glb8CwWYVglcYQ0CdaAS4G
NLyvAlKltGEnwHXrEzrqoahLLhjmkKbaogQ+hdOce0FFbc5uxRup+lAjwObbldaY
UwE4QWruqLYFXomiEIgNy0U6sSrM2K3atL549WwecGXc70qbEsslvNSDm4/1BVB3
ed8H6xmEHdWqDpBMXwM5TfqRKeU41gTb7FjDJ0IgnRbGMytC5M1FTkg8D955nll2
5fvrAuB/ARRzcIbGWFGu+mgenMV1Is1HuSRqmpduVwVaxieeRujMhJL06dKeXgx3
8nH4s307UpjbxScHhpljteVkOdszykIBmvBzrfhdOjPsu1T1mJCnFZkE+QpLFsoz
wCftAS6fw3Tw0FVMuw1DOY8vFfrLjl6nvWUlZ150VDKpJC20Yd1XSbepDbWEH43Q
sQAvniQYB90/m5NjMg4yI3e4Y5h9k6AB8RtnB47t49VsWzt/h2vQSfLfVaxe6ne+
4vfBus4QCf+XretXi15gB7lMgwZjLpdp4xQDQISHcJ+/sf7YTn1MRuHm0SaUC/3l
t3Yv18Tejab8yO2PJSUfdfyi10sKfREhwO9YbRP05mjFPV4wU6dqOo1+K0AL8S0Z
unISt3raJE4LQlHsakhnQIN/XPF44gY/hkbUMrL+QjNHrgZA7pdVyeDXIfIuYdki
VSD4uHibbzg5BDXH9bi0yHW5PkE1D8KnaTwGdNo27ewYR386c0/+k7LXC1743Gqo
fThihMRA1EwY/iu+G+/8nFn05RNquAAjrTGF08Wftijp+NDjZt1h+TedLjkr6v5n
P3zn5AbY+9NRrTDDRWH9/xpPbJXrwueA4Z7SqhaXdlffzzDigMErVI+xgJJkC7B/
S5QX03o4N3QSedP7NjHI1yPRsFVjbxfJf6TR8WdZSbjU0E5WPYP0LeCNrJ4GPqh2
UNeR7Beo+KPRKT1L/FZZINLqXN9TrewVjZgdxw2G0d0WI/tsK7I4a7XzIPvXJZIw
K+txExyItFquE8Rvg21QDVLG7MsxHBPSQxt38BNHeiWwYnCq1BawyLGmLIVV6tRp
6SgbCVYTBguA6ogCNuPEVxdW5q54rsuV/RqDI/dUdpEeyylUhEBcURKIKSzWYc/Q
DtyhPmSSn/3oynw2t6cfkcHcA4BH0KYuJ4KDqp5c+H/gWN881mx2bK2R2yMur8SS
Bdd04lCBoRY18BRzXTAMuY62ZOw/kAs9jZxfkoDiVw99/L9O6K4acABAUVJzCRPy
LfPCfft0iiX+SgHic/LcQeVjR0wSIdk3i0KYZu2CXIMW9jgBc1rawMOtHuc+6Fmo
E+p+C2lICC7Y9d2FUO/nc2Y95L/1jSb0W3uY9hUuSS1Jiv8SI8qwRykSybnI3win
tedvkrxLSG75xfKrg4ORf5E7etoOHZhhrSdjL3gCitmAVZ+i+hi/LyEOURtj1NBC
Rumer1tAD9tNfjsQ50zgVuwJcPAZrq3NpiJDZJhFwH1sewwnTeRHeiO38HIDL4As
UUlaFabw2uzuBCJJ5aPx2ksNy+YYICK0Ip3UjstZZMY9HknJnPkeJZ6sKlk50c+W
YbnFcuXAivH1Qk9XZh237S9Qvd/bhSqtbGy/wkjF0PfydJdwe8zJwEmadWzI+pEL
3Ek9eC/QWtWGfcN/ptYDQdgWpJ104+uWyL0Rr75dewawiyI3CusE72mOpaHsiuG2
kqnw178KUTwuQzueafgfD+qHOce8EKCErX+bKLItv64GV+nYgs7N5o4PFhIa09SQ
09EQR7fch/W/EWdAiP1DuyBZgBovBI0lIetHuM81k1QXgpTv2NWuY74ewJbupNzo
zs2NiD6QFA1LL/zWlgyhQdC1QC0mHfhn2NcNxEeU4cnYM41wu/y9rfBrtmN2PMMC
JEZuV1BWobyaL8RbyGriPwidN0tJhQQbrGzy5yZxrSmFoWRtIBnUYlAaozDcGq3X
i1q2rRdkYCbRuzrGdpMrTSAOlYIVL4vWppLTphHOUcdlH1T1AaDmAQws3uffn1ns
TD5Pl/FTLgMGV5gDUrfNPJmxY116+H2UO27IC5GenWv1uAfLu1IwpIwDxnyCnyq9
P1WYtZRfLk5ako1hgvH/ptb2sRdSj/gojWg3CU4x3NG4Y0V94JrMdQke+S7tS6vC
CNxmQWFPIN3CJuxAtOk9UsZq4RHpVWqfThH6pL+nsr+ppAvHiWu47e38ZSv07hWl
jrUI7ZuJTuMJIdWbWEpXsm36Wh2pAwZNi25nmi5xnc9iyTA1lMl9hHmiOLWYXKkZ
EJhwxVaQCEM1YJkfMwyOjkhDB1BOEwaLaE6dO/lQoz/cZ3iQE1edo/JrOJMUVBTK
xwTtB2iJEvkAYayExB4HBAr3gOtDLLjRzHHoEdHotluFnkSvgVOsOiudheTgdzyg
Sy5pCpoXpCk7jiTxmRWvLgzZMoWcWfAuqhbh0Ey0zw12kqlghKbCLlvJfiLyvjGP
I0UZ3D0U5QYoFYQpl6ZXmH63wLX6YiymEXHY9JR++CP6LJScWZrPYHwIqJx398L8
ct7bgimiSG92LQryVDRO4G6vX3DkeOKq7GkA3m4nkSBs0KOyX+BgsDzSTGP4DJj4
fQ2yraMhz//P7L/KEDqtnYaqpLTt2YhQKZYBvw7/i6wIoKr5ijkYgmjc7XZSLHDy
FW1t/mrezCijfjKop/S0ktVFCFUE1lVwdv7X6Qxj1ZQqUoHpaDg7WMyZG063C9/Y
KDvebG+wRz6Gfm2Mjl2fI+by/baKRtz+3ui1zRxPUxEIEQNnVsciuQwgMHL15Fki
FW3LA9s0kvWUpS1H/s2qgrgVLam8YeP7QKSgpQ4v3bh4p47Mq9k9lLdjA3+TRRYc
e67PeFrqtNldd3yQ91JbcYX9/ymYbMv0YIMH9eUnwnZeMpdPZWeWIgBov5kLr0qL
Mci1sLwWMyx29FGIFemQA8Jk1cMOIyrEyzeiGPXS866PfQRiU57fRcCi8UNMHPos
bJ809sjmTp5Zqc3VqLb+Y0xXj206kkd5xQ9QwvnS2QA1cvX5F7f+OFHGjI+QhPOB
0UmGBdFXAFA+nrT95RpYJXnZ4hNmGlaarTfawHDt2t0+2XhvmZBQjSqpvOWu8Jn7
Eq2OiNloWzj9LusWdZaHDGZduPQFY2N6R+Di9Ivf6wIJWhdxo4Cw434jrDeZBUcl
eE49jsU//1xRz7S0Z7WF7ijCQeraUZ+rENxxxknR3tO8388kcJKU+49Ni6GEOhxc
PJpBqKL90CgqqLNtdHKFxNYE6n25cAWyzT7bM7Qmj+Hm/47JDOekJo3iu+dP1JCa
ehhPzBN5gp2GS7YZ5K/OiubBqzyWAK7wCFCrv1CoZ976rS+gGBP4085ZMHVFQ5gO
OvT0HtDs54n2DoK6tYTQ+rtwUcRzYPnot+lBAfvksIX8jFHQXWgmYUJQivF9LLC4
rNM3birGJ7g6QQqfFZYQyNYZ1X1n9DDD9X8/S+vNblQlG0phqw3a5/WbW3GzES3I
eNaAQw6dyWAKfmrkp75YmJlR0ZoOZME0rTJ7J3+JUDoovx6CIAMAgcmeqjtglTGA
Ut2SdXJvJnefiGwI30cyEOqdlkSkeAJdg7qvjWKZ47b6iLNMeawf7ZUFO+BqRLBh
9QmR70mRmVyQHKXUa4s3/4AmtpZ38WA0J/lFBeZvEqug6QgeKFLmyNDmcuSA1PfL
IIblqH7OtYEP6BJbff85nJoWERp/mK8d5uaI1gN4sAwV69KgQD55nbCeluhtQYUG
lEXZqirFOgIIlbErkk31T5u2ElGhC5O0ajMqyILq+Gv6a627bSIClrzpSdL+N3US
+2vA8ngihxZwOvrq+JLqzXR4PfzGrbiNu3vODEJhPN2KepKsugkYFuWShm/ts22u
e53t5pZ5mZZAtqfv0vJPRmoMxeCMHT7H5DToT8S6Wh1/ouHWtWiXbDLLEHz5Yriv
s4J05XSnAeZdcor2yqbGBYoyB+4RQbAl2UG7XNA3fBkn0PYuH0TJnv5163oS0itn
M8FXnFJBqDNxPceTcQzXtw==
`pragma protect end_protected
