// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gjlWzbmZevZlWtnzWO5PsZk0VjSVzSodIvKklAJlzDq/YOc8ghvIiGC/eWSzMAQ6
WTk4l7oMUohJoWw6jHQKQt0SG2s+peHFCKAvYO06IFUxWCt4dPuBb9R01gFGT2pX
ZWRGxzirY4ZtowwxEYQlqptcUpw6jJwe1C8/Ti9vKD8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9008)
+lfYcB+N8dHeKpwEoum5k2zsvuBZkkKxI5QOyTv9MtZn2fjl0ethOLP5RGii/apu
L04av8H+1fCrwSnrRBSBFKTOgfW7EB6otWwI3Jj4gWQB750yrPwWkfacCx2Z0QCY
mdRIATo/imXNrzi0FxZ5NmkobK1sfxEXVykzGWv+FI/hkoH3M3VeHZ4PhAccK1fD
0GnSlPcZFSizyxvycAfnjn5zXl8eOrR9CM0DapcyxtILFf+F7knE0m5PRLB6ElPV
/HpG/oPDj/eRckuki/6aWEkpb04CjMDe5yh/+qMLsf+bQxBBPvMt145ZB/Zh5A/T
pXDzrzP/TnAlDnUDOARXdsNM/BOZf0swepc3XVuCb4U4BUc4m4Jy3V4R8+4JFBzm
+FKoymK9y1iMG7k2zuejLYKoW5CE++1jYYDC7tvIwIN7ihrIRC5CsCSCDEau/bzU
cvODsPSXwnKO9MIuy4AezqA6CRvHAkIbpDO+DQdZNuXpKlnMiazv56TsorFc/4ra
5Cfmn2yerb2Kv2I+MV9+WU7dbzZJSQux490odnPs3UeB/wm6LRv5dUkn/WIIPPjx
WM7gIMg71cDGObgu5SXu7qeEA74h8u0bLwvM2pNo2lym/Q5U8SCnL4ZYit41nOEZ
mA7Ye2+YTJoyMasoqGTWXsUNR/sTtudrA7wQq61lfRf4HNQ0hN/7gtNjOmiQS0WJ
qtzQ6mu2hIHSREVcYZricqHtD+xws8I6HunKpTFsuIi112WjPcJZP4pq7CcsSpQL
7NzBDiwhhGLmFUzYkj8sl76JHHeaD/UPrUcpR7fc0gFImagqBjuQRDlUo9GaqGxe
2N1Nv5yKJ9PKO1zqTTc6OklyeqdbxjAvpUpHzOzVfoiBOjd3FOrjpsypt4ocyD+S
fAE5Ql3cKSkcF0BrDza1jbrUkYVPAjrpFkpzRQsqCbVdyNNx1nsekhZPchxy+7jb
PeOLcQ6lEwXy4lUhtETwmkn3bE8Sbmgbi0vUY7Zh5ZyuxOYiTNYDcUMe0B9aw9eM
a2Ot+QgDYNI+gRuoBt/u5SG+NVBLK7E+eGOHjsZJqjg+Zl/JU06W7J70ydxweH/F
qNS90cyFZxGyCTT3BqnUzat1Mbu1f+FxN5czmaNOmLXn/w4Pqb41PRSmDferqpWC
L78h9a+wuVRXTK6sGNkzsWsEDZiAu0ARJ2Ckvnwxf6XDUVXoD+PZwI4xuCdAMaH+
IE5E+4/scXHtTfmzTzTX4rrj1LO6sbbWgVLsvWLIUsSv3cV+evXDavFblKgufX47
KOY/kxGhYLS5Sr4IKQd0+TINsStLHF5CdULZ5xwum64KgNCMuzHejKqkpgPg0ofD
Y7SksBUtv3nwk5b09HNwAGP8DxcRLFFJCjDX/B9vNSG5R2t4QgJ2EkrUzm/dZdSI
HDPBp4Qvs/tpU3L6smxOBo5ZLkohLtzCdsW5qoboZSRd0dzgfzu8SdrwpSW9Si4q
IrdJj2KL7oAEKEIscYhb9Q6UWM70n53buG+EF4+caDE9a0VCFDymtNjWj9jDBD9y
M7RXrgBxpmZ2wvlvWdth53G7nTPv/PeliJO9hmYlLKlh8tHxt+pjqvih2xPObEOb
i39oyj3x05TDCe2XQUfvHxBur+fFSWNp7toN+12zz85n1B91K7dqGuokkGRRGX4q
Up7C4TCua/+9dMDEzmqVG8g9CWmv9cbAe1L48Dd0L1E3Xab1BQZedOOlzBgG+3pT
1KPJaf40M10u0yqD2sSb+gGbbLhiAYQ1N9LbHGPNx8333dGI0hhAsEvaQ3RCYteo
kLf4x/RHX9liUK6x6Vl5oxirav47vCIL+j4lFu4zhEp0nJ2mFzc6tVNWxWhzcm+N
9JN72luRD7YCQMr4t8tGkbdP6XF3zI9gdB8BogdrWDUrMeNYw/K+8sconIIadbJv
wDXFhx+4pRC13nhcia3RLJGaDDfM0n6+qVneHIsr0pgA6278xf2sq7ye+ThUfuQE
RgSBTfeuUMj7K4hnnk6FWfNKcW0Bz6B6rVriBdFwUrru8ImgK2bvryAoUHK2yPO2
4bT+T9fhoD1o5oKrrnJfzoJHuOm8TCH5z+QJVukKauOgvDNlulxjkQc+8Mqog+vU
QhY+nDdw9mJdNBRnoFSL96hG/8OEzFDRTEPY89aULmLE+5KAAGxWrn44eYBrs1DI
oYaI44xqhzzlTCqW5xHSYXA17GqgOytCdKw81PtoLdx1jUhDxaepPcZe76+GFJfe
3uR7+jT3kQukEuKRTM+9Q/K2mz+e/4WuqweRvM2Uq7Vl0+TX7ew+QvbKb89ZphrZ
/V15xzGbw8brenyfrqqPOcz7E5P5qu7U5wWO/aDS0qKn3gZWV3WXrO+/T5k+6euW
6XQJzG8RQLzKRFlv5R9jwRhYeb91gSkDTmaa/nI9T62bxFwCFsNK3zCSOfieTTUU
FWkuSNH+ZEbZ2w/WofbLygQLDGcXXpOAIa3WWC/AOtWRrrzgZLb8SWVUy0GasXdi
jd+GDD9DMoLP1cOCMpIWaNufglicIL0lt2zy0QWh1rmCv4vFwTm39k9Re29V0JQr
n2LoO4QbaZx7xCG1qd2pr0bGaCEPFjSE822oV8M14BGyDXUfUIDOPG3uKJ72wuBX
9Xofn6/BY+2cGe9Pt1iRAloZAcVhVKhS2u/j0RCCfgkapL8XFnmpOqZ3Bw7S0obD
E5GZNv1B2IHToGOsnWH1nWfLPGMfejpr/E589ZCmSD3XsZgtcX0U2j33J6LlqfBI
yVpzN6d3SR01b0xa3DAeKvAIv003g/8bVbASzlt7sdS5xpiBEfvxauk1qguEgs+F
lTbeOl8YrS8uZwzrHxXfb2K7CQjk01X7WyQtdlQq8BBT8TXiYW0oOJ+bX2N7xvZu
c6dvrjCb60kXUywT5V/Zm1zPKxhskZhaVFO3nWuoR8JQ71EQKhugxmpgO6ai5I+S
SpBHsBxWaZxU5uzI2QOI7RcyWEcl0IC2KiSfK33IuuDwV7tj5c1bIKcQ/Z/VuigT
Cn1CGbQWcnGURmdiXFAe9hERk6sVykLTUG226WZ1Ht2k4yCE9mJVz0g/Xu27ug4O
UIytI2EN6C0VgjQWuTDSc+Z+oIVKRw2TVPloEYaL2emZkGsUDsTncuZidPLltvvA
OEJZ7hdzwHqd9iPpShcMGgKavnb4rfIwrjqPA+8dhDUS0w9W9Mai/YLUQF+9xtFt
4Sp9KXFGDc5Z37KxH8A6e82Yd5KMEOo9NYIxkXsSRsbUosO7rZzUkjT6gmvx3MVL
ApGlcCGCUohDAmaxH+kOONP7a/lGUPX4fsXM3KHM6jj1iT0lc1NBQzWuPjnVexnu
Na/dzzgS7BKZY4i/B3rIuQ2sdcpsjKiJm0aueJ0rTYtkuibcSxqf2NBc+37aLCMg
p1z1wdJkrAaqOkQ0f25POoMixQjXJ7/Ci2oVVtd69rcBIIjRgcOlHPgeMl4IUUfy
jYRc2ToeiGyyoe4NA5TIA4XI5Ejeqhf59+j5BsR3vkc2ontiONbfO2SX0W2Jiw1Q
ahLrTMIcLbGXbJv0XxcEtzt2BQzAJBC7GlZsNS0jV8JoGvxuc5SCR1IGq/PZ+s+w
M6Rg3izx79KfncK3wnWsfolFSzI4AY2VbPDtrUpBClbljfWwnckM77MlC6Li3T4/
NAROT6FOr4bcYGEnkpe7lGZpBoJUCp5vv22hmwf260xJbAyfro0uRk5uIZ1dNOLX
FbDlXEo/Lwz4oVZneIqqknY+Icm4yjkB4i91czGGqRfGS5a9GymcqYuHtPGy5KsE
Hz4xtr3PcQXBqperwogdcIRA0h1m/OBN5MQ0L0jKai7nN8rsuOi2QZiwDtV0w7hQ
lxtDLGemeKpnAu72ZJALf8ijE3louvUkVlaGrgfuKHWYmiBHlgLLvZYdYSip6fr7
neGIBFkL02bBQ9gOvjH0RMEXieI3Zd5ghIgfMyy/KCK5lPmlAIXAyjPwH3F5wJA1
htZsWGGRB+X8MWGrJW6vN1qlkxn4yrD4hn2Mx6crnAGhMhmFgBFrYoAVnDgmrsXd
oB2VpIDeYX39/1s/wolK3Oxda5kvLSaLqj3EvEn+ro6xs0WqqNRMI5UhRydGsi1e
qdg96kZsfk063aErvxlbwyNcFfdHQEsZX5HMOkzqqMFmvftxCvoJD8swFgPED2ej
l+rBWdSxsO9zIucfQkJI9c3vhxqVe5C4uojjH9wpnrRztHMQiw4n2cZkqsfD6zor
KcWbuZx25yhGG3v0s+C/zaLxBuU/TozohZWU/YlCbqtILwFtT9h2qCxn5eF3Iivy
CpznIyJRMrhxfEJmMOKFm1kwz6urMlXMskWVIVkirrThD+xj6iY5vD6jXX+q0OEy
Khp718LGXdteEHt2LP71oik9O0GcEdHuxa495tfgbteQ2UYMpJfgiKVJ8oDf75he
Dz2avvGrvKLOJ9O2gMPqm7xOrQntNbcH7ppI/bZDEiNmUR9Ey9xOrtcARCHo3NyW
CsvVn5EtnBYz2807k+qxPfdar5zbVf2WW5KrZFQrhmGHkZvOsGH3Qjg1Bdptmbd6
bgypb2YA6YwC/GhhlBvHwxzDGdonTLnzwyNGWv/niN+gwmS0mHTDPv+s7WdkLACh
LMoC5cJbprGVayWTuvSFBhP5zfx2mkzC6MfX/jP0hkPMeW76kFhoBLos4gIJjc7h
4BW6LOlqOOJrhtMHvMS+umnBSSZ6cfFOzLzCn1p0vFTtRuJ201Jt7y4nBc3eIkTv
HhXviNK902VtIc4tbpaBQVsO6kf+8+tQRb6KYkkz0uLP7wZwMQYXP4Amt7ra+iFj
S+V+vHvyp2eNqhara/LinsMXVrC1yROpCQoP1CTCc6OymwgjvJ7amjM0XonUH1CM
VwSlT2yf+YfLege+8TjUlueVRFneW6yl7jlXKGZ2QCx9JCAd50902UwuPBP4Xh1W
AhoPl9Z1UtmsrjOwF/Zq29uaBAFx1rIliUyHdjFaIZgC/4aunnsGoPdYOpPjyJgj
OaAvMz8qo7J62dXE6pxfHrVaIlxnZC+Q1eA7GuvoLIsoKS+gWhOSh9w/tbYc+9RX
5LHiVIcF2j/WRdTnFk2OJFTW5KJF1nN2p37HxJcJh2tTwvZM7mfE+XAxDT06c6gd
wMueMfi4/RjlW+BddDxruW/vuFpjKEdffxf9Enw3GPV13QAuum2QyzluRoyG4dvw
xRiJxNT412TjNTqs7ZJLon4en5jVFnRrsc9jD1boaBMH/xFleSjjZsUwbYuLVbBe
nyfG3kuufh2RJGY7/LskfFs7I/7F+tLvKjWjNP9HNBFhE6EG0HbiYK1T1LjyvGDG
tMo5pOB+xnqu9XyWbGVkcRqI5YgmoDpx0l3TTOMBi1wgle31xDShzE2auz5d2ozo
XNCgFhpXm4VQWZua7AAHY+RFX2uPUxl28ZCpvIncUkoYOhLouIF1ao3GySn6jprX
OCAgP03aKMiwvfG0eCpCx0VcaPq8TiYDZ94EzO7bYvyT7OxeId9YREKEiImD+qcN
I5e7cappihF/TQT2EK5MZ4/lG8+FGAFnIrPQsqtTPspyelsUuD6tK+88a//ZpHDa
tneJToiMRse6hlr6+T5ze1Z4G0abDINoHzz80aaM0KLyCPOrrU6TQuQi6iv1BmfM
HzlDR0u9v62yWT8YJdOxMmB5NGUtsuT5F8D/9YknX8If+9Gmpo2XMlvfW3GAli/v
7ktGu/PVZ58Y80sqme5ANNWX4TBFLlXezMFR8K7dpGTq9HdgkNTK/sRRKsndUbDK
xaJqJnLdmclHMV65Gw5yVY4wYL2eul4KPKOZ7VkzbYbCzLhglIDFF4zfA5+TVIQd
Pr8xJ2aTgi2tC14lZp3fH4nrpr7mAxBsZMGCpKRQ2CTG2mFAhiyVrGiR5lRi2XCI
sTpURSIS3u5hF8Jpc06KtQ7Em6KAu36/R5FtdVOECBpk4usyMHOsj2Ml87gYMREP
WP56MhwcLCUFJmKtyrmA1Bi7kXt4FczPzXnH037lP0UYQbz3uH/a/HT3L1Xirno8
/PoGe2fpGbOsbnzuL38cgZEGTNiIZS7Hi3gx3fM+eahYt8SgEEZwQTU2geUujJQs
bQiMNNjdz3s7Y37RgJPqkyharElNcqWyNMxGK/b8o8mCYSI3ovqNyKYFSMt0S2xS
k/trcpo833gFHaWpnIYW+d0fGtUVlLkgFer4y0sZcMrzWyg8BoA6hV2+0gMCCJil
9GCU6HVkQlME+w9h1CgCNwQUmlMWjxev/YnYhR6tizjKpQ995cSP/lVt0b/jUl/u
ujsNpy9iq3CUK3UL4Mg+0te9XGbT0lLmo39yXyuWRVLBfbYC7TO4ohlFAWavZ5e/
uadr5tngC/WzNAqnlDOvbQMk1e9sUM5PUiuYnctizw1yGY2qeH+iBcym0j+dnfK/
x0rH6PAH0d1n4UDkJfCp9wQwvWCiVdFivrPztGIBhwYOmyUMhA6EbLorMtxJ7zBN
M+Re8sdHuEf6O1zECzm4qfRYiA2h3DyxYHej55QSiGueMDCBMw+DlJMWTrOfWn6x
lluxvaz3ChsNtISHgTHM+nErKuRZcr6LPfGNVA/hgwVNX9URwidt7YrwojLjKBTT
2NRXSLy3hFBJPXXmpitBr9PnmGz5hz0+8aZRAd+GTQfejrLDrONZAXhpygq2Sz1H
SgyDOkth5nrpihW8/7GF7ti5mNJ3F0uEtwBUP1s5Ex4Ly6WxzTFriIouQxlMrrkJ
RbasfU8pZRE1QuI+5dn63gDQY631ETVSnBJm/j+DruuWucL+DIZZ41SGDcArF6KQ
A6cx8Zgi7llmewWU8LopFH1eQ6JBV+/XO5H7e8dIjNIIYTr+Ll/WGmW+aIYkLEnk
EU2k7oKsmWEm0CKPl/XaUBSH8XNI8meHbnhq5TRCjSVJqzgy0XSWhuBUg13rZVnP
0Atm/LJha1fSwxta5E5fDHqB3zt9W1i9DX22SiQ0QsSF6l3PVhvTTeiIkT+VPNER
XNyHrGkYW8OWEhOpOKlt5TQGQ+dcbrcP60He13fkA7EJMi3BBBKKN6qwlvJRGLh+
BIzypcsUyNJ77tgdW9V5zulWfwkqPuOGdZcrUl92YHDnIpF6/zU3bfsbBfWpVIJn
nhW95+xoNcp/N9VRDwf8yocPorgb77m5vrwbpkkMBaJL7wFMA7DhxGA3l/qG8Xjr
uEcf8JgvHER3G0QOFziIpS/ScUY0+PqBoLmIq0nNq8nLFigLeruXya2gm1TH5xcr
bSwKaUIjXY7EwtyBiluv4KNAZZp59QMNB6QS/tG4zDotzYET9qapLMFxCbeBZFWR
dZUR5dd2YZPTphIfF26z61bcJT+UmlI0WTM0g6FZ1fQXPPpmUyE344up55dM8Fza
H5HRlXBEbNh03Owdm01igJHom3/ZuIHolWJivyd1XQd7P2Mh49YUY4KIrvQLRzzt
9IO5p2DX087vrOW+32btqaCqXWLv3C3Zb8lSIxs7julOODV8ZQ6BFTLmGEL8owOt
cMwo433q959m6Iod/25azix9nQLNPh9mJwO643T2sKeGEYDTsCDFDo+laLL7UgeG
zAe0Hzhl66MvBt7fSDjUJ+5lh1w/+ZponFfTAlcYQhMArpfXfb5KwhZa0VWFXVgI
9XqDO1W+uYcTC0B1nJSPqYHkjwb9CTcplf/6s2gNr3bhreoF7FKHHSYVVhb0SQXW
SXGF+biSVW7mbuSxrCaqECO9XX6Y97x+PTQy1jXKBXiMl8absV9oQj3RnD3QXdF6
18JZ2h+4ANZrjQDxjgWbE7LCqg9lufge681gFjrYQjMaqF07R1tsk6gXDnZwGnG/
8gYx600xnrQ+1KDMwA0jjt3myVzJ9fKKyv1QrLq9p4d0NiYbCZ/8x1lhtdWphTEN
4TCMYjApF5jgTgnhbKN6+tZV9B2gDOPhfO1QBqsNnryGtY8F1a9aqxQqguaPbmeG
I2HtvpwBY+Y0uHwMsnFilJEcOxjRRECqU/1snJRA8vh3X8TNuPGet5cN0L7zFNPw
ES6MZSBJHAi67pflgS+qDjGJNn2/bWeuZ0IlYyMpJfEOG+BTko4i9EIqSqh0RHJr
RRQddol+o1KNYZ+/yA7TPfyNS4k0U2r2/d1rWACso6dUN2RvLl3IqKGd6qBnf2hx
IJvOq9T/Kzo3Ds4foRNC9cxIywagOrnFRanW48ykzXS/8FEczAF4yrkrrAiyy3VV
3IvangDYaaCev4t3peMSrc6axri0EtpBr5Tu7zz8vD+p9zoIbiTbo1cIpmNHVajO
P/hS3ZcmdFmylixEo0nqFNeK2Hj5V3HrV1OKiGJJ69+Zd4oilCWU48TArcZMvoPb
gmjXooZvoChN7SsL5RIMbp1HXp6cLhnkMe2LgEoIVHelcHX5Y5vpwz1bevdMkh1n
MHxKLS9QE+cOmkis1LsNOcX6UtgcZRGpbqcOZmYek9Q3zhhssqYY/6cffgZyKLzE
To0fqLKwgE0+CBGgCKbNOdocRkY842mEHjL6skeVDtpdjZCC+b4Usu549TglgqFk
tRH2tjuAPEMYqrYG8WYEEgFretq8wUpslFlrg9VfClSbN6uiF5kAQ8Fx9HdfKMaQ
oBwJnYwV3uM4RaBmE9i03Fm/qYhXw3zQ4ExzCRc2bel5DhWWicP5Kefjvppu1kab
HQcpaxKwtGPCga+LxB163LzXQczxJ1K1vvFEAo66L7vybyLdutuOMzk/cHe8qahR
NCS0S1PBtRoc0fpkjQm71P3tFXePcAAy1o63hSdHtzB4kRR53wEdL3mWx6vtsJ5F
ahcmd2ya16i90O8Waob0gpTFSfut4SolcZ3ma0tR7I+zlbcGTFVmvQsQu40LQblk
XRriAhILio4zTCntDt+BmODl5Ynf6B92qh/orWx9POLsQ6MGmma5gOTQzcSPRiM2
nGWh2tIOKLQNyVh6XLfDwlobHDwGu38jfmZIxvXkxNo8wWpGr9QTJkTek7epGi9+
6ptOlyvquLiC0RqpQp9I2v8DjXYTgSA86oXHPjdyO5+n91QAHs9IkanXGUafY85V
178BCmQTN7SJEARbGNturKOePzv79RRAB0R3V3r7y8TnmP+inves0YYCl1nxx09k
HUdMHskRyzwFY8BQ1j2vdnEuJxt4MGgJJnchPwSbVm7VBkibsugLgSuKY2ND1F5m
DIjY7/Bsbhgl1m8bNVLPSnr8s1z6uio54ezPr4D7mUin/7PxVxjKmBIGsCSgZiy4
VIFS+z9H1z63utq3TY+PSFVT99dxiYmjtzUf/GyytXiycEvuye0hjsMwCs2ab2uV
ry1cuGysK+tszBblF81A+tA5Txqs4kXiT3KbhYiBR2IX4D8XjeYaGawTHMkIL2Qd
3ILVjVD2BTDs3Aa5CeolUtCUnkMIPghB0PncpqgVbcXbOT14SUvdVXuLmpJMTn0u
8YIJz89nF24+88i2c7o4/mrtvdPsvO+aXRFe4cDApciS97WWSQI+yZFNrnKfkUec
373sRE9171FttTc8Bulrml4fK15JfGqSotqeVjmCRYz5sOf6t+T8lvw75kPpo0AG
VwgTHJ9mGMkwebZTBmPXqlyCVl/97wrouf60KTCNeQyAKIzD8gop9WSlpjcW2SXr
16BHctH25tt7KqylStkkuXzXt6E3JSpdwpEumOGFjt5suAebhJFtfejvrZNZuRr/
Pa9YL6P4TylI0KQnzf2NakEUnRlIWUpAofrFv5Tub+SXGpExm2ZwyicE6dEWle4l
UncwD0DAJkrZJIlCkvnhNQQdVLPSeTDoNMFYBGGC5/5rdXd581mSEIR+dixI3bPg
3McXaVHeIiwwOk5mbbWRK0xlARIUY+sEAHHm9yRhblJ/3dhxzoXYNHQFCqXamfOT
MYv/Sc53f5e86grVmua6eGJsI4YNCfDCZQ4B+9IAScvHzhITmfwmXd26B/6lhVF1
SMrR41xzxgrFYNR5OLAEawpfeAHbU3JZ0no44o8bCKeFLNoGAJRtvNvePZwbbdA6
J+Ph4Retmnlw1xsOGZWEiNZ9wyluQ4wapQLGgLMJdlvta3gfOSM7ZdBCuafyXJER
UZfXblwgMsJzokyPllc5jodKg9VDbug16Jfk0Yw4CJkgQljtffp6eBGUnZHmlWwP
Xt1N91RXbyqurGt/iRvCSVVHdbgqGfErn6cCz5WhWenz0n/IIv7rMTBEyPphhBEB
BCbIGiQYS5AlyQ/IfUxhI0QfGb9ebRkF9rc34yMfiikzakQXKewWCEODIhiqfKi+
pqzBcHd2YVe4fh7QPvIs2Kp2/hbgCH0o5Lw6yqdL4eG0fq2siImJB/dCGz6fXZPo
10TokW1yMmIX5UeY3tDtDsLLhhoOkDPvNWt/JDcm91Xu6ZCnI6+FOZev8sBGLV3Q
hK1/AHo/6Jpomh65+N4B1qwi6x3MkmslDh3+7uSHaMR9gNtmOaGbBANwyie/aFwh
wXFYhSeMavk/B7Sj3J+2iVr0KhiOgjIIkmgqiY45vOTfKY3D5oDawgqC1eAcSIQG
Wj/f/5/qJpVR31ZqJX3eEAVku20l+gjDQIXeQbuzTIt/5T0Qc2XurPPADjnsOfDN
1Kc1AhkdaVuFx6kML2euLRwsWvAVvxMaKHcz1puCsY3GjyICi9hnL6G9lopi2XIZ
t/HKTR5QxA2HguKc3jiE4v3wWL7qCCbYfQLr4bagvkL3Zpguay9uUPpFXJHH5rbA
lNBeOqhb6UsEHBQYgOIUbYz/QMSZZ0LKFcUy7gEHz4OMYJmJVcJ2o3vye3zQoAqg
JHiEpsI0SaYgSQ+hzjgcEZhqDE2TdrpXr5R4xPTaSmY1lQ/ukdE9w8AC6+UgYMKE
DradeDHQgXAw6JM4GHU8ckC8KjKqhEARpB8ynHlLvnFkGC63u2MwGllA8JpEgoN+
NogZXTO8MTKl+ShyQSmiKwXguHbYCE26qrIZxy2ocoCzWMbH2jb0NgOxGm2tqvj5
BLTQqHInxccQ71l0u6a0NROAyVYOkAGYBYDTVfX7azopvZ7c26ap0NK2LA0jwc/d
pjOoLDjHIpuPUNJyxAEPe8KYpHTTyvIYx4soI1+kJ3Q1dMtE9LWat7+cG8H7zpuT
GU7xiV+jo+S+ezdDS3nNjRKtAmlw+bixY3UXcwjVSp0jMRrtIfXkwJiSGuiCZz6S
8+5+EQbYKHAAqJXWMLKT06YeyliP48fKIIh/gpn1tg7MUwEOihhOJGQC26Xaspdk
ON79rLHYJwt6Ml0WwegH+N873eTkPvja9dzgKcDxlB4hoB6MUQWMnEXCYRqLCVCr
UBOtkUAApx8X3U7DYW0F12I5/gGjCtdRotp9vzw0qPqfVQgJ1awLXti4RYlQJLsb
kWuCp11F1gb9Jjkj/kZsA40IA/yWK2X1QsclMCtBuupS6fzrNXW/qwaPmqzmpNk9
D5SRJnUmfSBwzNxOaj6U1fx6z5os3wMpor0zfVLYxVBsTgjq5WYymWk47WpHNCtO
AJZYWlFgJWG6c8zE6m6jgSbfIk6sYiGQdmrmWbQS9krL86hPAEMdqpkePag1Y8nv
jLbsewHQZhCjgxtVj8QqaXXX9dIuXDHZNGc5l0EeJWhR6SkRzg6opPOw4Saa+wux
uVZKq+6Zm+qZLGjGCLt77OLsvIT2pfPbCKdpZgHElmcvfxW7eoE0MmfdjW1BcQng
ppLkAw4+p8WxVJSBUxAYnbipyEQZyHhyykACFJH2Mwi4mtbTudmNSsnp+onFMgVi
jfRbRY7sqdmM3sEpfXraYKs+ZxNss0+ltH2EgQzz704w8PWDCZjYP0GKn1oM3l4m
TdilB4Y/J+c1cQaoHWewvAmwqGSHaXZTNu/S1UhZlUoKKXdzjzT+tuzYs8mb7Zcg
+3b5a9FJfGMdo9/EhMoS/AMQNsfGgs1rNbp/DiMhNDtc4ithM1Iyx0GEouQ9YjuH
iMlakXpL89F3k3ob66jCoYQjWWH8xmKr96WDFHa4dD4PG/2xg+xFvz2jTRp+CR0O
DItlkrx/fVepzEFulBfQTeKfJd3koQnetpoy257q6SY=
`pragma protect end_protected
