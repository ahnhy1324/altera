library verilog;
use verilog.vl_types.all;
entity lcd_controller_vlg_vec_tst is
end lcd_controller_vlg_vec_tst;
