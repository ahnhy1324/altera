// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SUgouXW2TAMno8yS/B6L9A0xvC6gqfsaFa5We8ESs0lNERpm7JlUXXPzmGuIr0C6
Exkzv3+3yMoxe01o/edtLDBfm//l+BeqYV9Y8xuJJ+y7c4vwE4W2ZBhmTvu9bAJF
Jqdcr7yVszkxj6JaVYEwwQ5H24CfJ+8Ijb7dA023XjQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25056)
+FexWSiVrCVFRxI5BTIu+YKNsd5RvwnNxePbju7+/tkIm0ML+M4VKIOv47uSHeE7
8XlekMtd3HwDY7nLbdDXOJuzR8naVAgFLPtQ6dTqakwjCPDly+6ki8hJERXmfewG
x4Cnyami8ErxXaF+rtuF/FPghLwpPZiBm6nPvzk7zhd1Sf3Gc/i4p8j5Uxet333x
O1pYYkOuRPG1HISnRaI+o9fAbYYRSjc3SR6AAIdafWkEMh5Q8G0NbcdPCvREyEnD
gp/oyt6FlQeYgyQ+EB4xVuX1Je7JpluCjsTJ9sudD9IR3aDWD+9WMKbIRm+GkyzE
hN9LfGYPevU5utCA1D8w2TxYHWo0MFNsNW1KSNaFz+mQvTvo3U7b/V/GigldU0SB
U2pTvd0u8HFvn1AbXxEGBG228/p8Y8k5II3/5NRNC4r0K5fRmT8gyMIeM/ZpD5O4
rZKAUtN7N6TEb6D/8+todl8EaSkO9jqJhk7CPdp/HVJXcYEd1txJ8fBLMNJA8oQ2
6KmMQPkrpLZ4AATh6OB/BDo/FY9L5TiUDSIViP/QE3ON5eH7oio6lXmfNpWwxZFP
ljyUqcjSk1TQFhFlYGTq8QCaVOD0iiE3QaX5LtAI2BMw0jdp5FNTuY1KNzvjjqMy
6OA4qVvaHgY6CQ7Jj6BczR9wyeUei8ZKCh4MgKL/0k4IA1Ks+G7qTnUkdAWGvs2s
dpmBKl1WoQz8VWWVlyakJfpz/2dTxVOp5NlhDEe5sKJF52Q34w0+E9xuZFQ8Xg8E
g505iL2xpZNYYIGtpUF31iCvoTcrNZVLHMgEpWQeSJi9V7WHtT5aLH4D1unMLMwl
VD8CVIZMCqWx+97SJpxNG2FNXzOza5rMz15PRp+iC3Igqd9oEF42IdaHkjHayNbq
Ia/kHQd1SiuZnmobAVmqDYcMz3a62Gx7HDKduOiGo8fpQPKRQeCMdFWDMXKZ4TZa
vDSPgSgZu0K4Iyz3YXlPFA5pxJ4ofAEmBs0arCCKx0cfh6KqM8uFNXNw6y6dO5BD
WwY0efjPFK6uQMyJryutcK0C8Tu0C5c6jFXYqQqCiUHU9MClyQA8/Z7Ji4rv2063
SWuWpXEhhNyShqWQhNKlxjsI7ShV69CF2qkJdVCxPq5F2ZHbmj0+T+LBLFqAKk9R
7ghb8INXAi4uaFHOZ/qaqcLEDqoT9agPsYk1McH0Q5Rmuj7lag8wSsMJP93h65SG
bkll39nbJDjzZqxVFV5uV8deLawARe3ny/sqI8Ibhb2gN/nPh4gkpF4XKSJLiSvl
WxhzXHGPvW6U5hhCqAHycc08T4g+sN2q9JCqLHqtXW+xzi2euKTsxsxBPBrrlNUS
nnZEqt8Ynm8EAV8PCedVzG4feHXvVEgkstIX92NCvHQsoQnNuYktdqxJdTXzo9y6
3830jEx3JHLB/lFLb7U9tqOi1JT2GlmnEzZnWCYaUIcAfnPG1Oz9Hcnebe3+WMYk
vFJdf3p5bdJAguSA68ovlfsjxs2bTNF7H3GS1zOzj9dkgm5HDgrvY0TR5/F3ji5l
GkRM3KmM+3a3xrHunfJbp4DkQQ3uDhS17nKWmo1BrwvTA3kDtr3zcMT0n5Xs9zcr
zxRMhBfDVvWcPcT52A91tPN8r3g7zrcnknJkNNLwBTHptjzQ5Or0bfBortmMomNy
7MHSJYwF1Ymb/raiOYYZvuI8kx7SxCpC97SmBNWPNgxQUTOdzdbiOh5mFSBejPEf
v18trnGnjKyM5BvhRoJ9rDr80Xh41ffGx+/A6HHNcfUwfKmgPa6gs95jHkHJX+qr
2BLIsNmKVtLYUJsHtC2QejyjKEX9TqJ5703PhMy+A8zTTVEDGKeq1+iNmodcsEVU
dz2qnZ/IBKncucBr1Wpqw5XGtdoYU7Q4Ux4JiXfdaUxU21eF4j80TTmhlAeAZ3lb
CFf9JlhJjqEs1nguON8Uq+P/eOe3IM701YvFE7f6trKZAHtwu90y6pkfgX0qFeuW
OO+tE8xzTb7tUtbyUeWqiaqUV3jsCE0Sy9Apa4GqfDFoMqD5xDy6d0RLYvzi5K7e
/wpJhMBoCNck3nlHTnUfvr/87YcxJ9AtjuvbzzFf34+x5/3d1D6/ygt0um9bjZxp
+YOJ76ilinU0ZOdE1nT3m+cgxweXkrfKrmh0iD+x9FjJwCIXw6aLVz2HwC7+ATOT
V6FomNykSFs26aITy/3ePZ3OFzsR4IgCMb3OoqCwE308gv5/ysEMPg6qSiie8tXJ
qkcXmOenVikJLu2QDjiSdc8Yg6v/oFLo4TF+RER+hfs2KKj89qgvXhDbGaePr+uP
wauvKshg52i28nN9Ayb414H9slqzmk6mp7nw2SGzqSqbpr6b/5AjGqm6UcRO9TMb
6E2oALpSYFd7wUcy4sg23jx/ozRumCeJgZdlsKDl3XXDpTxTTGoWOC7VuVbCzoJN
INxy7yCl2NQ6UJNGc8+P9IFA1nSTwKGwwV6Od1bwM0HtkRYqmjtCWYNWdHi5sLgG
nM7VZkyPYa9ah3rJBfmFR6kSXARqdAE8qYFt55qxmhfUHrbO2gdVO2LP5CTZYFdL
eXKSGGR38jvaQhvYZ9oD0t38ZMwvTQjBsP1f8PzNtwDksTVf9+jzyayhHh+zp6K4
N4HzIsTZUAthuMzSUdPL7lD6T8lfcLzIYQz747Mfuv0CuhxuF4qlBdQdXM+WCYr6
4W/YIpWlp3soeynZODHAmex7ywzLTwDZK9GhWsmf+8e0W5yKH90jc27/AO0BS1fX
NmvsqgtEgeQeo6jefVgrzpCpZ2BkDBVgbvKdCdZ97QTn2vDVlkKY4mBryf6/Whse
iTe3BinPd529IBVlAWkNAkA3R6S9njrxh5OX6ZkZo+KPksuqCVL7xeH6RTNdT/hE
frV65ukus/1dnhoPORwaRmQp4fkUfgrtsWpoeT/f5S6lMcYvl1sT1eJSpMVuhu3P
gqZECP+7jDa+S9KCt+LC0Zh9CIRjdnKfBBU1fAUKHnTi3c6bWR50bplpEp0pvYiC
SBUBu95a+eR4XCzL++VMGHoiSvGIo2T2V86k8qc2v5UIbxEfddml+Pdc/aFjeDmo
vfNMP/Akl4my/oMs3ZwtkvadAYnJGYiibVrJf+U/fYTsrVUI52le9Qn46AHEik70
9fOCtLwEntPk8Fi5kKkV6dsy+gjvvD30tdPjy2FjscOH4/VBR7e36atVMFb2C9Do
A0l04Y6Bh674coRuuXar9LBil5BPvv0suIUU2v6cRpn7+Ikjmoo9PCJU3SneIGli
SIqh3Pb6ieh+3sQd8iO+51DXESHQRyyedbcCXFsjHIl30ZurWNH/ZZkmkdzNr0Yi
HUR/JHnPdC58xcrBxZp2Wfww83Z7r4jC2MVNTXXJ8Am48Oa5hyayo8hWqg/gbcDo
2kTcRVxlIXsMyS5iDOqLuyJRtX9ryj1TTr+mgUoIG+1ByfG/eqac48oTkG+GAtcy
FUzpz9YYyFTJE0fyG0lhuXyCGID4p2RAXtL0cSLd+NkOzOXMUVWx+XftvG6K+oia
WYDVIyolh7qQEnvRtBtWHa0bUYvFGr97PGedTJ0mJklPZJsVBqawPL1R+cMayLia
SlbDN4GU7/A2yT8H+KzZYbjfoJLlEyuvCFpLB1z++EH8dmyzm2HkohujVLt2loh6
MCFeiIy2wQKTw1jwvfEj/nKJGLMXI/2AoSDS167T/wWmG+PQfsCzLUUxVu4OzsUb
g6pDpLHBVaDQxI5K0vneMwM3zj9oqmAV5bJ01KgegnZFZ5RkEM3aKt9XWOOOX1Ef
0ivtcEJYGjzt8c1vTX5Wy0+RZwUiI/9Zqklodj9xI0e9holXr4HOP1Kvq/lb4Zdz
lJdy3l7+xWnIC3rv3vXOgLuZ4pKO9kB9MhzwAQfRCxvcFZqhfkFcTrKJIb3qnx2v
koVCPM0XM1MJC3rzrpzHbG0VGj5qbGk3OeLPKL1SyLotYzRmkNTbmXkLYVJ0oIcb
adeDoTkZ+h12AeWDaaLjoi1QoOO+WMRH5BusmcTpkbUMIqo673kFULFMEBgodk7f
6WhnaAtksC5tEcVqK0XHwERgEVSl1MsS1OEce087E4W0gyuQ9Vg7sLF0MlV4CUuV
7OE997UdZoYym4ZLWAZ48XIqoAFH9jzA/Gx22ZkitkArHmLLXAa2lOAdewiCZy32
tzhBP+pgEsLmdd2ms9KadVddrHhknhu+ZmcvfEZZGY8n9qVZ929DU+ZqZafIFFxV
k7JD0hkC+1tcv925hnQfBZnbjxOS+SUfNd7Kic/XnFpAyW7SgyUASU2NNnp+SOJy
w6H7uwOUgpdeURW+cyXoDBx5dUyUNaU2nCIXD7G7x3xySeh3Q5Io7KgUPmHx6K26
ids++E+CfeFaxIhXbTw0Kn1ziGjKAkwZnlKSaVyxQNT3CEs7D46DnJn2zzG/tndb
hsm9ZuSMtXkIyidHx1uPXnmpGN3csAHdCHYGlkMhVAmKU6J6vMshgf3n6/lGyYKh
1FnRaqwGZPXcP5y8gHXLhw6HN/vrEbJ2QiRbr4BomGgwSPyHu1EpL0PLnwjDTdLw
K0oLYnYb1cQ0H05D2ncBEa31K8+nAK3UfWU57aqS8fr3UlXB42+OxXMWmoEcj3ot
9AzccCFDjPuThzuPBF3oIMyYzoS8+VshSBxpvr11zvaIHpaiucUdNCS1rP2vYXoA
TdYDrY5yDhl3LGIScGJQSIiR/0J/Jj9iVFiS1RP0Y9l0g26pcTcVp7U4Qf+ORyqo
DZMrWS/Afc0eHKmBrDsHTywcvpm5JgCePM6Lmk2xJJw//xeviiKPBlQA70FNGIj4
75xUB/AChNcDFHquruudpiQQ4hRAPmm6OfN0ulQy792FyCeYZNIi4V0XesUJ4xEi
XOXAlO2CsAFZaO6ZSBRz35GByxHQqGA1qE7ZlNd5OSENg1VepJJOqzLARDlyJ/Vq
QJ4ZmT6R186nlvBD/4YkAsDqFZVQoZpl6KL1d+EFVelz7G+MRIHslQ0vgHJT+OUR
pE4wU9mKW7K2hD9RSSKNivJMSUvS0rsbnUKPSOzjDxnF8QKLdKocBn23KBE+HO9J
CjUG3hAivTFyV3w/FCnTFlzBVbynVUm1/OBP5GjgqsRnA3MU0PvnHP5LyTcE4DrJ
hSDMfdbLMJccuHSApbIp0iu5xxFwc+FQCxUUFvy5xInYQ3rV4cfDpxZAfjx3tUDy
9O07slkDm3tScJpMklVLNlrEaKDKnLtyq20stCYBGvcOMqBu9h45kgk3x5Y0lWWg
W/lAPmAMJi8Pt2ghdQZcX27QIL1tsRP2sPCBnezVi6BmmGV+uJ4SYXgFavhObG2Y
xwHmkPfSoYAYXcHAU8BOkEqbh7/OvvmmGMBVsRobxExQn8hrvx0TAnC7Ya8I+vjI
dQsHbp9YO0Z+YIZa5wbhpqRwbcFygXjmB/8H7MwudTorD3qhdMHjcEL40GTWDfCu
J2kL7lldVpSz54TuR1qkRDjyfLst4B0nwJ/dJsZPE6o7q6j/crUqCOBsKpnm6//5
3Hs3Vyt+QsLg64gy0IfrKFzoQTdUHJTdp5UwDMkPA0BUn01WMZ0jK3E1QEf/LL1T
Nbuhkcy4TifTtDOEXo3syaQ7TeNSbx8pHy03V6tposXW8WOxR8TA7/b0VvpiYsEv
SemOyMjsinYEWCAVEQksIGyZwy5Mfy87ZxbKSq+pR5EyjfR1oAfrqTKY83YmgIm9
1Z8OSM0/rNQUVdIHLhr9/evok+3YrUS14m4ZGc8WtvzCYpRP1LVxFup2Z40w8ww4
U65C3cSW2TklpqRpM/VCIa3kXSMkLZ09OUIWSvAkHrGnU6864Bsyqu+3hZsYoybQ
zY7Qev/n4lDpph85SLgNqw7FDt4f+nsDJtpMqzrOZKCtA6Gwy/u+uxNMW9x2OaaY
/NiLytoHUQ9GDDYUph+nR0xmP008OTcasENV+0SAZgLC/gQvBWoA5qQzLpbMCXNw
Jqnp1SGYcoPbv5irSr+LBjtwJNNmHEj+ZbsxOTAdUvwjp4V6cvtkw8xkf4AfbjVq
/xFXDbM4XeWQa/5w8Bvy/meA/OhBAMuiCLAMlhsBGre5LH+DpQtYHwopnUbd6LE0
mGUH7HYiSCXHuXIN3FBRVtcm3D6nOQyGVd4kuJBtQcLvwl8jrLuczHS3nqi77sYQ
/hzna7Py9NQbNMP3Drp1jp+F38SMYaDFEm6g39EnWYBwkr+krcczaJ4kZh57K1rK
kAGS0LMApIQ0R7fWnkDDRoU6v/JDPXgJDH+EP04pCpZdRDfpwOKbn0BHHZjTuzzB
63mVd1TY4B95CuokORLGoV3bUVtRNBHS7DSR/z2QiSq1CxQOzuu7sGXuqBNK0IZy
nzmI2r/Nswwk/JoWT9z/h7sbpxXIHltVexTG0f/wqcdu8JPavEsEQcWNfmHqbntQ
r7SnZtuPiyBYL5ldoFT5UgM5pHp1xOuc/7h9FjcBuZBemPx8nKHhQXDoeSMlHVZz
vJjbR4L1crLtdkX+Tjn7LiyKiz76TS3zocP+hfqbKlCK2141mMboj6j9EBH1wlXQ
VATsttnDsGldyJ+HMu66GvuXGKYpOUu/sfsY4F4TKnWYLg71nA0PbxGIkER9A5Uu
km5DyDyedUnTyc1PuAzLHbfJbi77gnDPAkZCyRN7bHUDnLictWSN8dpcrya/zeto
V7VlTC+Gg5C6Y7cpKEprMofc+tVNwT+10HscjcbqPudoIT2RmT320sBUNbKhwuCS
AhLUH8++Tc4nm5KPsQGaNbhBHzuK9qpXd8qJkN9orv6U21sw/IP28ocbd8VZTl4y
QQ1SoDqEW/njFKcXMhGd0FIl8MFRE/9eHdFnGQplOyrPZjoSz8+3BdSCKs1sc+eU
1AqVouZPgXkTLsvMqj9upkEe8q+KvEoaQpxlP2j2gXZXnLQkkvC4EaUELoVlAYxS
Gl0fKcsPrVQ1HKhktS11B2EHrkKGwKBclJwNQQr9V9aTuAZ1SOfnQ30iZFJ/kXPo
ntMcQQwlfBl52ZDPxKRvtLF67JAnYktHvhd6OuiMv+GltBssFMELXEohG7AUkaaC
S7/QjKmfQKbAP4QuBGNOKfdEIeSALTsTMcdeNxYhInsXX8QDul0HZl6IygDpd28t
1Ai8deSMCDInTiErmxUgUebWG0PGskUYRGCajuAHfDeTzwkcWQG01lrGRIF0hhaC
jqPYhuFWjF6twhGwqD8QIS5TBItwfRcC2zb7d4v5uW8Nq73JGJb3RCjrcurScHj8
8ep3zIYTQW/5ZGJcTtyoOuxymdRxrVnD3jXtAOqVP2dLhAGPDO80zJgPXt38x6yR
vm1pXvWwlljZPXL0B5jdU2Zl3ZkrdQg1WGCqu2Pbj+qlyNl/Muwm9lORDNWqkY83
tT2LVn6fQlLXEbeIDb1oM1IV2yCVKkbczjeRMc2u0euHwyEs0ka5lUYON9dkdZOJ
U/ZN/bjoNIKIVnocq4eOsTDQKPIfkxgd+DEE7jTxbmVSUKMiTA64rQWzTxlOz3QY
ROm3HiUiE9veCZo2sHvq3FTBWhWxDw9PAR93N0O+b2MxQuxHVrPwz3BBcjgGbb6S
mN0JcJBNpQDQxiSIzXM2FfddUzR3XcIgHSSjIZxoW3rXEstsyT1h/eO2Ct2TF7Nq
8ab/Qyka+I8VBRTKvFzvR42w+jqNh2Glb7febisbA2Zyix2/s27GU0bFPA739hoP
evbffsOFSxer0IALKDdqNYTHS73eN4YGXrxTY9XT2b1zMUMpSVHJmeFfOZodnSTw
pMoh+vqL6gm/IYWvBmrlvOc8+MmXMBbPzTB71yFkJf5ZePekTWVUbYXDTice2tVv
OG3N1fSX2owp6qOHinhzWln6c14mLwAXuIxGmujsSEVDSQiCcT0d42OLAgAC8B0d
IpO8wqE0x/OG0gdFryK9BTubRYyJDjLtcksNarimkFuZIicDsyos6jtG/zN64qfG
jcfTlFvdt269sRVM5s39Srf7p4bEFmVW1tDMEQU6bfN8QIu5kYaGdvn+rzAymGE/
o9Ou8VE74H2HIOi0mdtbKB03Pwy+UrTHxTH4F1XB86bXPSWa6bP2x1wD5M2RdKV1
sUx5Yi2wmS89BXf/8ntuVWBTZ2z/KKAKnW52H7Up9GkwTc6rdBPAXNcoo1JJFPvP
uMhSjDog5GX5NSgNKjEIVsoefXCCXuXziHedAkRrUb2oJATjKvzevCaHHH2AT9GK
OWqOUnIt0eTnIbaFE2AfpIcQm1+oHdBkiQLiHPxlGy4vqKD1LS/hnGrC2XUHF/hj
H6I4FDeU1HFnZhhw8m391BW20/Pd+r+r3JRbR0fpdfwtOrapM5UNsvwKXIdLgPbH
64MAJHhitCmkSE7fOiTuIpo+fv3L9CtMCIPneg4vnijiUmrLjVAUUN/RnbEHm79S
66rEc/gQ55aPVlF33zedDDyi9r4BLZj7iHqwC4aCkJEqTUnFeXMD1ksOlqGKmWQY
pl1/GsjNUguaXJBVKna4uGZxC1Y6RcBh7Hwz/QR20A3c7/+fc8G6WncX3lTjfelD
HMQ++Ox8ZIKnEwvsKzZuSh3P52jDBM5OOzhJ3K1kCCa6beXkzYYd1ehXcQjD+sva
TpxGQEqnU9VHBdOH+UezPXRL+ZOU5g7T4sGTSpLLcOA471nrSlFVDB1pnHvnl+V9
dxWvHPR1ybwIRLkKI6YjGnjMgnpaDMPLJ+bdICAKG35PmgPi5r7wqMy5bngpgpFj
xlOe45Mrb2ZP81vEvEdIT2XK0F1ashkTc07Gg2tDcDc6VypE6YUzMqQIbxLG31RK
2rXiBHn+XXX+vW9Y588VAQVNaGRLFyvpqY3i4QNzmUb4tPIwNw0PFzh3DqfnWJAG
f1ZNrUqi6Sy1NTJxoMJDxg8iw/9uXtin7YaH8bdzoC+gJRagG71EMfqbRlUSrK9G
dRjP8jKol3sq5Eh1fbhhhe1Rq8tZCG0CUFnbcNwN43YC6KtEIs8B7xskNRGSAyfI
Vzr+Fc8VmZmmE++87uAGfVE4lJq0l3zXNQr5rAnHY6RMR1nNWGOhYT+5eQk266fj
/uwlN/LLSR842irjjJCTSsiQ1x/3wRN/MKC3zkfQSqMBCiG9lf7gh4AKDQT+SYl0
t7gDiweGPtCsI5xjKkq/N479LAZmOUN0nLK5+PsK1Z2fzOHA4KQtPooDeDrkFdQa
m1UtcLm3PfY1BH7LQMyTAFRtNIchlMCOpO+2iqjINFEPBm5W08tUu0eog1hbbCVG
J+s36FayDosN2rCUxqfbNqNZfI4I91SsOnCsNb8FASVCc6fREHWx7RcKa09JK5fX
MQyfqxYtJBsxUzKWe0F3oCFCjbeuST7DtQBszxub0nY/hrKc8FCdTaLhtkJFQr5u
W3or+ERn152Z5e5N89eXKMqB9ZbjuB2QTVs2kOGURupN81H2eaLOH1CoRfRhkCIL
79axgvksqjAw3K9BvMW0r2R+zkjBFBbN6c3Mt4RBmf3hoaQarUZYKiHTvTuSF3b/
ITPYa9Ka+R3foWotOqsP1msfEA1fKr4CldxMOhPzQ5V4Je6/k3MkgOwP5caVPpe1
FqhWTWqeY42SPQLZN4U7H+a+VCy87ngDlXgZtZt+M5yS4xJBBsyeU95YJlcUIQAD
s2QaMHZv5XVK1srgL5gUKaiaseegJHwwyEwpNEmMm8f0HNb7Nx0IYgccr+nq/sJy
HBOCK2R7tRsKnlaOy33clGaNBJs8/qiCmIoyFIlh7rGZp5Y1jkQCnpVHDPivUfmt
ZgBf3dl/HPss5TP+qfNA3A4rcIn/HQR0A3jKg7UOenNwUCTzt6j1d1cyjorjlOQh
IwOcIpuv2tFf1U/cXgx03sbXKQyjDfvbret9umXJ04YFvFrcUZ8p7ykup+2xLGNU
uVto6ImHXr5FvQJPNwhdA6F4kXkYshsJxFelKF4nJeI9F8Y3ESP/n0+aBzLG6TMG
aGxHwchSy9muMTu8fBR7GPKg8DvsVqHSrsd8dmZXm8ENp+3hH4mvm+R3VVG5bIW0
YMFP6dAbLq3byUWvJjIIObNz4TWWJ+2R/Z21chx++jqc32J4og/htTge90w/pk38
/FMwL1FZN+fOa90CmxGwV7E8bIudaJvhdwAXUmUFVAJwPn2jWoXQcyZelMdVQM3p
AiqQ9pz1h1q77pQGnhaj5+e2llBiqppMlelS6paLQgWhGRVyJnEjC4DLMVxRT/eu
cXxU+21tNNSvUNSHm/lVCw2W07Ap6AK/t7hhQYlrNT5gbWpsaAv+97OE4dgRDl5d
xD1nR09vq/QpZefjC2zMDqyRpc8Vu+2t1ZNvKoh9dLjXtbitRIiWz8+n4jODKKZW
7M+z8xVLpYVb4StmQFPytTkinXB/Z1FvPBtT1mhyZnAGKdlmoz3ku2dpvdN++l4E
x033SQvPCwytVSTGoer7Hd4Ldkf+3oCdz2D0A/Si/zLn6xN0Wngor4KizaeGvZdq
YYljeP1CnNYdapc3+MKIpsb//6Gx2fJKAsRPYL/LYxh/XFTgEessfEGyvq7xZJk2
ao0vCt0lqNPmYZbv8xCL2YYMx462K/IVM83OVVviw8yyyrRt3f+VGS/apcOCLE7d
ewc21sOxXzrV0R037r1FpJKKAmYONEjXZHtpiwdEhc8yu4mdCQJze+NLkx9sDVP9
1tzXO5HwRAi8XJQeIn/heBsgxvg9QloJlnrw8LRgBifjBO300vGZY3s62O7KMfMo
Q8AvrT3XGv8HDBJYjVjiZFeMExtFLaD8oYvutLbcEu8yG7cozu6adBB3jmmL+6wP
Q3yxnshuFVjgfZmz6j6Sqxh7zWfBArB39M0BBRiPamUvKm3erYiopohiX2vbmCPs
hKmMx3E+zPRwMy3En3Bd8IM6n0ZRxD0mQ4DTrlgYE5YOkVr/zu2HsSonQCbtbtUW
EPUNWEbOVavak6U1V8nmOYuVAAFkfiP+Ud7GFG/6a4siSNL6PtBGFNZC8iyDekLL
kC3KXH/cQosk6b9YP85qQU3aZPMnyceeHHbZhzTo8dP2EcHY8ko2cS9MhsSYaZts
8MrG1HgzU+hX42JqTmHDzzvcxVJKMj2xOMiZ1qRXfex/U9BG9rh4AD4HsWJ6geWz
x5qko5DV0xGkqMTM8QzO4QX+9SeSiU+LI+pegkGMSFYBwzqvF61gX6pFdBTjGnU0
DY8zHQSwV10jGdXLSjorCLV7MGuU81bHXJB+LbFbyaacxi819+yBLYLQFkkvukNv
YyDeRREDtTNpErFYeVyAqyBXmjWI9JMSvpG8hOxyKq9ewy3sdnfz4ueSBJhLjeyt
XNnHh4OmysAjB4XgIlseeUmzh8z5p54/cRe91YXSXNuDkAuTdPS4yzvoXd77FroO
8qs2R28ODcNbPgI0qxeM25MbFJXT2bXWDhzAx7NnQBgvsJe29nKvot62t4ofLkp7
qw+sNUHdZEAtEAYuQb3tTNq4aHeh58z/tgcXTLQ6N51aLPiUov2NaI5fJsD+KHJY
Th/cibv2uSLJKyU60ZUQelimx0aah8UPDA9t47sSuFHG3I8Lr33xingatbFvSroO
iH1n+rPqaqBXEcDv/2WhZELDYOo2fli77uCGrXai89rMqEV50LRikK5N5cn/Zop6
PsgOhtJLqM3fCMGBnL0NYnI7FuvPtQpkF4sFFi0PoBLSjjde63qnpftXWdIbavqf
OAuS4YlmhBBwnnwUmVUrVl5IP2/GH2Uawuhd0HodGRY68noFQxUIzzIwK8GGAKmT
FdZk13ok/NHwQZKpybyvOsn7Fh52Wstnd2Knu6sQgWGbV9DvxzhmRKac0y9AinbB
weU6eu+AwwWtqPHrd2MxpSmhyK5NP3x2GnXNUYolRfUeZIGKku26ik3exontSBwv
BXnFcF9YeCPF6y9iqJfI9ZaGnyol+IN9n/nxn2jWy2ZdL3LzDfMsey/WwNvxgyOg
USrFuumpkSa42pcxjxIfe+1CfDmr8IlxLF5vu/JBrtvBkiWJO5OySM/BDnmho5Td
mAlLuZxTHLB5zg8HebO3lc/DoVBFDd++g+0l2AW990Bc0NgwT5/H3YDueJLSk/JX
n15bDUUTUtdTEfflWGXCyPz4HFpeLg6sXIvtxlH12N0EII8hVTg1TazPAfjiySU7
HMdVGOcW8O0LYMjWYWSeX9rS1sO0J0KA7RwBPdelJEVazr4EwmPrYu3a/jw2Ctfl
/5TxbLKr6pXR6G4KL+1tO9TYhoKwLlf9mit6t9i3njE9TV1Jr/EdtOq8esNwJYZg
V4JXbaVS8fi3q8jocbA+l8N8KCN5Qe/y5awZ08lgLhLvLWQP375W4DG4fg9CBhII
BC9lpNy39DfMRBcHKaxIIVjohaYaL9QG8JvBbLVOxpvHfy8C0se+dve1PutND7VL
l5Zv334BYR4IrspRxEZHEEaGAepMHB9z7ZtfyDJfTeG6yLwTKRy46Eg1i94j76U0
eyDcqWkKYRE/ZnRPVsSr5PgCSS6Dul9u1b4ODhi3oWoAkeNFzFvuuQ2zAqhSIeJn
/BHXWpp1jKJH9XX1IyWicKk8SZRey2R/qFNyKw8mYlIXuzjqKb+7hSy+vInDR6Gt
D4Vvw9+UUug8OPL4KnQUDyjQ+KbmqCBA8WPp1kla3zAn2I4lRmxi307P3PUEEDyT
NqIKLOhreJPFtMHHiytsHvwLFElaNk3T5MZJ/Z7r9Zzxk7fsMrDF5nT2qFMBDWzp
ev0aI5IOZq+YeD9pWwLK7XsfRo0doiETijx104/QLk7hfSWNjoR0LkO1ndTnRe2H
964vnHx64PpSU3ENvcdb7trl2R9Fma7uEv0PkNYe3paz0mJyoPrFcEhRFon/9but
wnJ4mYbLx1tRV6yOwTufYfxhHGg24mNVCBbPwY41+u3d5no4LP1J6xuQrNZKgaXC
Y9kRmkhJIRbFA1J4zDcsBTYob9VM1yvsPib60rdsflHHRl+hylcwWVjrxF90v0vU
mCmPtJTJVYFOVh2DUQZQk+TcmfkyWz6cdrcbuWpo2UCIhwIYzT4K9/yuZC0L6xP1
VdF2efWwAKDTazJ/rRbUNZ74LfyFGq082XJ9v6kQQwTWgpJuCzs3waB9RN+ZcbFv
uIQiN49yj/D12VKmt9ujteCKut7iEe3DUxmLzwRfv1gyHOIT24FKdzL/fLiafLxt
lL37ElcM2jorzSrmMOGwDbAhEGCYjJ1qwuhwBaBja07EyxghJr2/i42evr8Gqayy
TGGa5R3o3RLt/+eCTuJ2m84Ep5FoCQ/LFOpRefoRT7LVeqQXZV4Yjc+TiipcaNrn
XM6NYLKf7A/mElRDEnlw3ksiMqwHtNsTLLW0p3RzbFL/HOM+5uu9M6z97fs9BNBm
rur7Jmh0+mKTQHiOn8IJrEP4xeN9n2WN87o2s4hTAJp2NfXSusjqmkXoExoyu6pQ
wp2i1kuMbWvSyyMOdjwxBB6amwi2ymJ5LjlRY3ZzCG1+wfEodrsugO1thG8yrQ+Q
DE+yfvAINljfWiMeC+JHrldXJ0iYZt7lCASMZHG7tMFvA5uarHnoTfbxe5FssC/3
LuFJ0EzEXRZyqO7iHFo2IHFD3Bq4tnJY2qnB8J0/d79O400h6iwk+mdmp+9TZkzv
/3Cnglrg6rLjDxFYj58mTJeNynJ7VIIrDcSdeJhYHJTtcrI6avW7vMmyQags8E16
l/abidmg/gOOmxQHftHwM2W77Rs9R3f5Xx3C6b+Zbmy+xlg7JVmVy8ekNAzcNGeQ
b85sUqF8wkEolx3dAffZJ/55qjoRuWgdIJbTw1E0dHqvKknrt45xvrj5PuDeokJc
bkX+zkpd5I9Xpva1OOwy8oF+woGoxC+dtfWZRnZ21r/5kYlEIHjo6od6WtqynnIp
YMmfPeOB7sEqA64bo+qkIL7elOZRMbPgfm824amsxQHjvjTYfItmXmgc1Gzd5wa8
JwMalX788JY4J0Ay9QY3jbUSliSs9h/r2s9UzXCLqJURyflQBKU6olYb+1jwAe4H
ncny/fXcUnWRfw10+EM1wI2gqgUWWSld8MIwp5MZphTjGb4V2LMxX2Nz2lsTZ13G
c09MY4DrAF419s9HtRgc1qPGHFcCga0yUWrI8PMENlhJKosNoXqXo89JdVhwceI8
yAGZJ79yik/U1XejJUDNmo/oWLQc4dwpKs+d+EFRMuJfHKCPDUJrW2pjYnCRfuzV
nhU/ZOYH0ihYsCDWBBLmjxOIQ9jzRjutcJL3v33+R9estcxs7KIwS4Ta/WyizO/5
XanSB3Mpvdp4NUGxGSVcBWGxVBq6FEPFQPkBCxyE9/B7J+UXBQKVD5Q2okjx18UZ
VuGmprUH9Ac8fb5gosbLoEvP88rhdtIDrTEZrZVYvqlBkE/s8jezDCrkt6X3Kge2
mvpUyD6cZQ7mp9AcmSvUJtQzSghioPSw5Lvz5+WFFkjZwKOwD+cqM5F0UnOjpwje
CgbvB1bDCnueMdb9/c4+N6onUAD09ZZeUa6ZObMIwpjCut9UaLTMkdP9mK2ih6IM
q82H1B3REjTkogF2FPxe77T8+yC9ysmtwOeWRxFljOq3v24ltLxmfuV+FC/hb1ge
kiznYXbKn6DLv/FRTKb5e7rodXEZEPyZ7L63jlhPbpYnqQeLssHz72CZcuuNMcJu
+xzCMkfa7RWRSy9qp/DrVxrXEBVxrLpBacpDZmYHJh4DXBiN5Bv/bj/oflgYoAAn
DEk8ZgWHBC67yXRfnYG3GuzRlE3UMvNg7COXzix5f3I3KLhtTLBw+kW5bVtlHi2t
7UxsnG2O5CgCH6j4twUoo7f9eCKeAbkK7SZMCuS55khuDPD2XRmKapV5OZYcmdzY
nzh5wpmKwH3bwR/X5A//fMr7ZcE8xoUZEbtAZm0IKxMx3HRmVSAV98I+z8+ACfgW
HfTiTR9mIU/raI9KfWQ4t1Xok7H6qIq8E+6U1KTIhiZTXHBnLyO1SwzJs22TPGng
R3MVZZI9txEumYGrDJXSnSeoP148D1NodykQoe+NJc8KHlRa4W4rctNMEIwK93b8
K1NxBGDNxpayO9ma6DgdCkWfmHiDFLOg9wqnwtjHPEcl1MLNtof1CnXXEFZ366hM
ZKp2J8b2WmBhYXzG+S9zZ46RLcE+OC+2FMSVSjeCKbznhv8jg1bM7aQ3nD6hkXaR
SF0cXZPz+7ptEjgQdONyluertbR1c3M2NMlnnFWS+qCnTvV5P1vnSgcK/itL+36q
TYGtne3Ldj7J6gUHeQFRiuvf6VqiwRATNv0KrMaxshFh/xsKBn55vGlxAqW41j9F
kg9g3oujSZgCq3vVL6KOQtJlhl8GOi25pWJsmN6hLLbjpBq91DQWY+COC5R7RevZ
VYhu8xxYAHDfvpc+9+ZLJY/6iyO60OBfm5JDYD3NslKaFbIycOLISZ7fqp8BoxfV
3YxX39VR6iWVnAZcn2XhuUtPDKtW3sy+PvRLXrFXi+OuVR+oMUoZ5Mics7mRllen
yeb7jc0CM0OwpjXtmMG5GFYfqDRPH/bRjcL9ENYPGI6FpiLoUPLrAozzXHun3yjV
srIOsawM88gOmntHDgTGggnsKilFPABob1QZlR81BLTwj2juQ7vaXreEh+PaHkc8
RcfRVASjN64OUL1mkBzCdl4ArqKBydVpTyJR0nLKYh8/rozO9vMe5z6NZJ2wwSak
Z3mhirFxX9DfDmdkyVEpBdPVx3ljDhz1+vnKpZ8WieUlZt5AVFCQTylCPRHDoqaD
VTeMpnBnQv9ua6xkqD/52q5NTsFoXJAd8vJm76e9URM932o1xS0JZXdEjHxoFNho
iQXLU+t5X/ZDB/tHydC4NBsTaKhK5L1LB0kstYxDS3DyqPjtSK4Xeuv+fjLFE5IG
5pzr/7KbU8DoZjNXzyqOljdR0j5vJy9ILDB6sxdJD4cBxHyWGZbiyOyHh+oRJ8Gd
TXj6tJMpUBzdIMUaK8jltRgA6Rl3Fpy4WgQRCZ8rDBHyK+UAKlwIwwaVsqvnFODK
lPEMxgGRgibf+Fay1bzMbL9kxoDvTKTBQLL4/Bb7bZihCloUZq3lKIbY1OYTe6zF
WOyveKGPddcD7G+r5HtWXfNnOOGDXR0knx7KrzmC4n+bv8Q2u3X+EWE6+r9Yehbc
AHlNESTLvMCsyw0SmHyn1FVczrFz4taNxGS0DZTqMjQuHGt9LN2XzZtffXKS7ayV
JwUv9/Bvm3LQhLLbQ0pivMlA11VRG++GedxC1jgTMsaSRLC6+qScOaYiQR6EMQAU
Bcc00FbUGItYPBxfdgQqUAGiDv2+puIzr/jiRJbm0GRvaVPNCKiJZ+KBnbaAVCiK
q47XY3R1V1yzCf/Jj+4ETOU/nHF82Lpk/gpXXIehPaOLyldaK/rfGCIi65UEeYpJ
IPUyqPGUiGSahVxhKa8qmiLGJYQNev5Ssa2Oix5E9Mm53DVRevDQuwxWGvFtsHDc
3EVTRjcQHTs0iloxrHWl++DrWRX0MCD6j3aqj5XSH59lLLKo0MA5RKr3rdhcMKNW
Q2I80z7k01sddB276qN+72eQZseWdBSrnJkOH/YCB3ZlW3IofmVl/ISY4tTGM5I+
BkH1PyeswrwfbedInqvqPLAUaJ42BaAWDVxhNsV+sv7p3WuRA52Msp/MzTQgwMHQ
hgLtCHU+cuMx8e4t6cwpFcYNi1IhFpylHY/lg0XP+TbfVe1gqzaKnBKZvcSJlOq3
vph+dAYnNCDUzV1F+kQOSs4lnKTkFIk8ckccNJixkNe0l41GS527M7H/4HcLQx8L
1TolmKLRu9PleNX1lq35+vuV1+ZXC3yBc+t7Z+/lvyLv9tFt4Qd92X66lsZew4Px
m4rKBxSb+A5RWi1HM85a2ls8qFO2PHRtqb3k7B9Yl+Io8kD562CH+BY3gIRSfPHN
fOyB/MMi3PyB7E7hLI0Pejl87ZA3jAMavVp2nsrrW6cI8g9rMeXDwQ1RrLiOkNax
Tysq+Q5WW7BgCi1XrYSQzuxTzWx1/lj2VYUp4reB51h0V6iIvQIm2iG9gnBYEt0l
Wba14Si0nn1hs1NTny8WzegCE8mZR5cCO55L8Naa+Yj+ADQ3LxxaL9IanhlwHQXm
lDXnYtefBJ6LxpH15bpyGw+w67Nx+WmtOXnCvqcS63Yc3e9s+OpYTCTAKRIVcDrW
U9F/9GdHxY9UDdHcahpYaKge01m2SXzjCWuJkagnC6gTL431fiSvyS6hYzBmQcU+
rgpSkSyCGbLQemY4C0T1JBcaVMKrhKwhzcGEnsBTut3AEEAYQQ6WQ4xX/05PIGyB
YYTFfdhPoyThSWctg4TE8MJPpjgDni/0t8HJsxHLXNaBzGnTjSWj7eSF6ioG6yKr
Ub8lEA4yO2pBeFNHL8C3tbyWoCq5IwYLbHRwAVAof6QwtX0b6Qniuac7scrAfyT+
2Dlpji51D7HK2QGpSMgvadh91rcHJd//5Vxo0NBTrIfHvxwMgC58320SCdNVZMQG
P5UaIf1V6ue2vAqcFeM11Iab4S5/RBbFYLlPcCQpZvko9hSz+hvuCUU3Jp9Xf6kI
LHL9LinaWwc10921H2j0WB7uGj3udjXyiV92IhqoL+zq8aSC2rSmxe9nxp0J+jPQ
bZ6q30VmXDyfdBDe+s4XtTVbZ7tqzlgW8pT7dEa7uWzTHY0aZTYkKNWfNRINWxJP
QE05qzwuKq/UlwqQSdz07LUfe0H6H8EQURCeD70gMDu4sJTwuCXREeP94236Hfor
wcVh00iQ9UBdS3KowjSO+cJRcJOP4xr+zW1nS2AjUW+tldmrVwPiAUXpC4gQl2xd
7thxgSXMSkdoAobxDMxZGDWaICsGMXlkNLpgS5JMya2MVb6/r+L+Mi8ZzXUwyURo
Od7MZbfyocRvCn5A/zNhA/y9MXbHrOb0o74W1BYIHI0Zo0cVQWks5WiLaHLV6A30
In8kbAav04+1a90eFNDZYu9bMlBJcgkShqHuJGqJUjXVX2YxKetQn2xXItmH1+db
ENzdF8R/6op9Aiq+FJIQOjDGFBMcUo20/bSWelOJHq4kVgxyKaQBe2FU1vnGXo0e
LX139Yn8j7zEAjD64t9dKUTG4JVQC0EPkU8cDxwbjYPDl/BA7WqXOP2M8kplZYrq
gXfvRMxWX5mr/GQ/fyPbF7qVu86EKe/Ft8TrokYkd49HCtCvngds1se63Bss1mH7
uBwuQgi81p1o5QLXQJansMHh4/fggyUoJ/wmHrMI4pepd5kRa1y/mkP24ku0N1Oq
GWw89QqZVKigLTmTueO67zuZIhympDTNnVqwNKBC9LwaBiy76G+0oOmM5p1iaXsH
UVewP7g6iqY/J7s9enDdTxWiaW+Xs6IYuXOyZOo9PZeOflRUHYSFtppVmwdkHf86
W5UmUuXLVYGnhsN/ZRLfXZ6Yl1q0slqtyGqlG/te7X9T75iXT9FYIiMSODbWo81s
aPJqmksUU+TQA334vkiYCVWkaCoq1AkxSnnUD7sG3p4FiHjZcD4Rtvsv3kJlZnGQ
MTspz0nhBKqH/Q/ZTSZzwE7HDuyZNPmi+OJzWwPx5zI7GAXogtH8B+F8LqZ7CI3S
MyQ5Km0yiJSffRq4EiI24wIDp30NlJQI6Yf0wGHxnDbDWkL8rtCIWj4GBA+GWVHh
DyNB3Jp0uCbkCLJe83tIRbhwEZyf8MG7j5Dh07HTiqQpzgIOo+JhH2Wj4M12oPi+
kdVfuTi8/mgaJwWC5wVVPOhyZ4advqVhu/arxOhhzuD7njDNafbSvgAn7f79Yf32
1xJLjAZzPMBqXg0zuHh3MfDbuL105q9g2DOAlNiiAzYPdw9elQ/yklAiR/h9HR2a
ovTYBqTHr7pdUh3toL4OJ7Tb04z+YyKq55Ke8/DmEzw9QaoC0uXFNujB6EZVmCOq
CbWdhiBF7f4j77J0BneOwQIngPvoX+0rIue504KI+2KQqbLAaJeMTIRAq5CLxPUk
sXE3pEqb1Xuu+ovHvfAK0DYn/vBAXnr5tLgwxEEHP60+uwFJL8tiFv3jQlPmKj51
IMqE8TFzzW/dzG4/vu7WnGFYYgz/qlS6hfLy9DzY6vO69gTE8Z6dogZa0U5MvVmc
gSN4QLuTOXc3kmQvZD2eQlqZCHEmB3fjcnT9Uc59klgen4SqXvi3eMvoQakhYI6C
Q/mX0QIB98k56VJMhb2rBp9QFyo2VXLQqdJPAvEiVvTvALWymveXQzPTup6WYdSi
vFiUmHEyABrYEwtuHp/zcejHU0MqMhbSB0bvtT5Qwq62V5bCC0pJLd64vTTDajZ2
xqChz5j1RhhFP5UwoOHH/iJw3aW3Pjw7mfhSUypjPIRBqS6EZWv4Z4+qPFrOD/YH
8EnCpRnlwykeVWMS/8T4JYuVcXtAKbAY4DpfIkBkTa/AeHJU3b5EuWdbwz5kgrg4
KT/RU1Uq8DEN4Ox/zMF1Y7OQ/dr8yU+y4SmRieFyKjDU4wHj2dJ1pe02OacrSBBx
Hof13vvR2WtcFPSyltwxKn5kKCCxAja0CCqBpOhEgHhms7e/pGJlHkRQ2u+iBi4b
KpJjyNOz+R4gxxtQnyowyxQ2sfBTuPgos+4PXHKf83kY89+YIU8LONZgXkw5Ar6X
Fmv393QHwbXqy/+Ef9Wl+kDyQAoRzZsASi72lmlqRNhKcx7YDw7jkQi9Ztjm9IWA
kwsSheRFyBDWvwyTCdVQIYmVaJF+YbT+XDe+56iGQ28iuttoLDJTlrXdn1v1opOJ
enBUs6ZS3MyHKJaPBxpD+D4R2hUKkUJlSDF8v90Q3I0wnk+QJ0FbO3yLv+NVfrch
I/6MJyDUR7HOehKSngx8xLEGr2BJH+bEam+6xXErLUs4pCo0HCVVrm6Glv/MYyoA
wgj4QDKWYLciheCmRhuPW911lzDQ6eWHFVyBs/F+phUibbXY0AEpSjyPXzvEVtPy
WjiKlpiQOWz6Nsfv7+CvvLd0OVIiT+w8An3l4IocF3XF4FbMcc6m/wx0rcNfTfzB
9WSrjhNvdsGfXBIvr3Xdbrg7ojDrhB3VcsDfYvAcFOqLTWpnsfWZdHjU4iKV4M1o
wdDfVztXtCtqi1OzTDB0N39nulzzSMgRzopxS5uvkiiTVsHPyKjzGFgk9K1KbNBm
cngrgTOxekWBPgp6ZxOXVYNNiG0BjU5PbmetfxMjJ6YTObtNBzjv321GV9+06SZh
wGnuYjGPgu3UK4sFCqHbgulXiWlh21yoDbTnGOupNyH8ayD4Yyi2pY2ZFO6075Zn
bFkiH6LerPcQaU3V4NZmu5LG0Fff48RaqXXu+0P9zCNLpVK7d4IJkhayajwhXFhD
Syo6W67640B0gmxGiPhjKpudyRZ4qc/1HW7U2NkzoIAjt883cl09XoGWpZYkdweX
SMww51z+eKL7huEcjGgTPzPI0XOTR+/OMU+aGqz+FYxI9lpxKZnsNRFPK5100+fl
/Q2fsiXqI6SH1EuuKS0Hjexf69XrAKnJ7Qxo71tX1No34tsybbSVW1y5zRmHvmBC
aMAT4p13fb8HA+cTJqavVWqg6qn4ejv9eq3LLKeKRQcxOjxcOkhYcDUm5LKm71G5
E3v6Bo2KhpjqxiypixoWYd0FleMcux/Qh/I9ByUHmn9iyhnII0JdNVBEpwpaTukV
AZ44bqykTs+4VmgJF1VeER4qo7Yc9RMkl6i75x/Bb4J/UKrZ640p+pAk3CmCoRZs
9OtmUiCPUnotg1d/QmeL3UrepSvKrRQQVVJMeuqvbvZbFOqe405rWDZSo7Xj+43I
rCP8ZFC8gYWV0U7zfXWyI13+r4Y4dvSDvP2eq0yTq+1gJgy6vxZMiLtnGvJex5i5
xi+GjXIq3Nz70ms1R2aEYnzSVLpeBu9QFEC2Y07+jwfxvM8beUQ9Q04to3MbRYmW
T1f0RpU/neqQa8F5/lzp06ZYLycFvhLeIidsGK2Tw0jTsircfhe2GqRB3Q/MDVc0
0mDAyDpulT/ct50sFd7jAm6TGPrJsah3j01h8FNIt9poQpIA6zom5z2PxoiqkRCP
+DNYGKxqG+uHY6Ni5/XeelhWVDRGEuPnIKrDqWtt3Stj24a5yQDOxAlsqmJ+QyQQ
BbrZW7Q+avJF244bbmwBLujFZKTDdrWCaxTScrpNhHMvzO75mPt35uMXvZkeVkFW
ZnpWSHxXX2/EmXHK6zO80g5q6PCDUHG3xoQYi8jJQO5w8VgxetXf7lFiM2f4aD5u
P1T7kBo3Tl4QxjDGzQLw599qy2Bna4F42QiReSdw4T71YsPu7f+DWIt+i1NGCwPa
vrQbVrf4c3wIf+n+2t/ueQisOK70vaflX077lxb7t2NfsGMo/rdQXZUp4GNRRZT7
nIIroWE86DeT2TuCS92PvwAsezD8oS2yyK0xAY827RyalJ9WSbuBAMpdjqzHKuhN
EnUff+Bl1Dfgl6ljzP89of3SJ5l9Q5lTQGMusMY+2jExIF0uzC9VSH7FS/eJKhGO
ITSBr43miNpnm3n4n4xHr+hs3vP5D13EoQsmIX64e/3L83Oysng7jhXBRbz7zifu
3CElu8SYyAegksqziEShgT5Mheyo82VLQuacbOAbY3DVsaYuQhw5fHJUd9vFsz+c
KBFjumZUzMc0llP1iSVro7tO3FPgm2ovrSbr9tpGnCk6Ru/k8foYaz5I2KBnogap
NyvPumPg39JKD7koLbErj+p2KAFpdCkpV1FNWvxvKKQMiM4vYQ4ii5088lZZMM7s
2UJ1mvHj0+kjyVkB4FVA8yJvS8/gdLYvIplohNiQlaSWAu3vg/KsE0rw2/Qzui5i
TdjON5Oq7tyG88zs1f8pUcosXtSZQU9xhFbvcnQuMlDd7K8v1aHf14vTcuWamV7W
7HvU3qBqK9Fj6nwzwKXaY3UCBXauYZH7es1i7IBWTeC5Dgs8PYOZ9vxZGKp3blsG
jMPFAzXlEYkfByghN6sRCrpl+UKQCZ/Ou10QZhkFD2Gj1eE+SaeU7NEWdTvqNRHH
iG3b4frdHu0FFm0QvBuNho0SLOnzLr9xsfY57ZcXcWSLpwu5ZGxpUOpz6t+6uujn
feXsdtqcStgBcOi7V0q2lzJchJkTFvVtiFLtWJasSkXg4/lnzT11hl5efejM4mK8
4nAf7OVeN+P/dsAy1gCZvN7GZ9F0afWEV8sBgxj6HqXf70wvPzpZU4xIA8aH2/8u
uQAaCnZ5SZuN1F4e06gI3eP0M7CA78fSeQofTxQJCdrCoUCr8Fw82KfxMT8rs0Qd
RbJw6CcPlS3sGeZN1t7tEETkc14y5tleQ20Qa8KSAMPehZpRee4Eubs6bO9WUVzY
clNebJKn9ukqaDnZnq1YjVxLzwHCPxR05U3bnxlhHugeQ5XidkY6OiH1vfZuP2TB
MT0zG8X875GGQDRib6iYjJTyMdRN5vKySsT/jfzT3+PVrhVQ661je1K22nhJ2a3M
Yg5SiOMZ/2ihLieBb0HIT6ewV9tpXGAHGJxioiBMlvdJZ/d2wSs5OZjAE9/28o+n
ZwXtMr3OygWtNvJe6dGk+/C58shEGBh5eStqtSpQYZlGh+V95T9OGQ9aog9THMN5
qr/P6e5XFqvIYfgIOEDsiiDP51aHHkgCEzvYs70ZVDyiO8YfpDQMYm7Qz9MNVvUd
WWE2S1nwVy1GPR+g1bZOfi1+6qsKn9DGxzMlBKJMrkGgbKjX/gGZ1zzmlL8Nv6Di
KITJYVasKCzCKshy7sgBg5i+F7iVjXwHmCVjFqLO9mJz1ovoDndZUSBAaE3KPeyr
anSs9JQN7+82jqNvThO+eEcU7lfajSEyi/mtHXMWCR3qEpr9cO/qL1Ux63qmzF7u
tIXWGStiAQeBs+CZH6xH3NrOziTQLiVUcgagDw0m1xGiQgNOsjQBpIt2vT2v4oJd
npPxEt7jJPuf4a/wzaydbByFgeV3cKa9glwGoqMXcIFHESYMo8RQy0zOlKNFVw8R
QNBQvlWTAwtGAoyub7vFl5PtEWQ64zNo8GPt2x1Xh6gZvYPE2lNBI+Yyo8nGevJ9
XZrIBhwOecKmR7Z0ncRnzE/608wnpA7TN/5hw5qXOLdjVyZPtudlMOVdWntoSY5z
qa8M/sQ5aGAbCo7+iGaPvmbPjxkKgRWPfG/tn06ZnMYj4B7WtTzFedauoo1/c1nG
vn22vTHzZ60/pNwBTRV2hKLW/nDuuXXRxF90Ny+lE7PCelVBXmMOajyCywfxmbcv
cK6Xtf8czayAeQxN/faz2QRGZJFMYZm74Jfot4jF9qCABaGttyFjRmDEfcWvhMug
0pKyr/rB5VmamMo/rZRaQQr5OkUZ/RLDSOKXTVxSopPF4ozIZLffOPBcgMHxV/7e
FZkdp+sJryzNFP/SyBBmOhSnMoI1M+uv4J+AsTcjK69kC0NkkVxxklegWOtLt/RB
3pZfYDCbLL0YbxoM3xsqmMQeq424n386RatXnuO/GUXtyWw+LeDVY9/IxKeXtgsD
IfNnatNZqcbf/Elg5FvDqmv3MvFGlwTvJ9pJQswlxaWD2Dd2O0T4pVuVftqtVEwd
MnZoWU081hwOhWb10IakT4jNkD5l9AaAokmHmYxCbvZBtu9U1xQZh6M9sHumpjX+
znas03OhyiQ7rqThWVp9yOJ85nygm5YJaAy9VwxK2MD6Es1FLhVYJ2kEIwG3Feeo
PlkSI+iNyeBx2yTfiOVfP/6uFFHCzEvqWjErm4nN+d0/kvTr6WfKaFs2GlhSxl/m
U7XLYFKJoLiVnfKEfkqdwHz6/1/qrYD4GMSVRZkxsUPSqCUolpgVtmWkCmk9sKNE
NudJJqW011ePF6I/vkffOAqgjqOc1Fi3IHWKW0+NcljAwNz2T3vuBYm1AvXscsI9
1LNgQkirdzXMLWLGbwOtfcKRbAgZHYXNaoVUonOjk91MjNMmft7QclUOpO8MZ5Ma
fQFrnXOwzARE6K2V1tIVpqEOZOKYzt7nq+nP1UgiHfI5jy+gAJAgrjJ3ARxq+/Nc
6XtwBWN0/7Hs13lajSsr1rTYs8Oc3S/IM87JuaUvjXGNnITdIryqldGHZTPWu2ZT
B6KGPab2LaKWzimBMgjX8Z74deJmb7ZTB7xKYVPHma/Kj5/SlNUBIbEO33lJbEuH
0q7bfCDyNWS9ELZa5IoTfHcgYowhaB0IyC7kkDi+RIAZzu+mqYlqVb+13fRNLe7C
zsvY5K3qQc03z0IwjE2hl6FmUm02arTrN9bcXrD4ttggpmaIh6KacNxcbT/txiow
JmrabR+1z2A32U0k/KKWeJ4GcGTl7xQ8V/1Pw99I3osfPq1OkNomArwRD8CAXQtb
5oJiTK/p1DanFDqfi5mVu+WcwOGSM8hf+sHoEuF0mo8ZMmDQTAsqk1S5amWEVNw+
YlDKDsN0zmH54nd+Pf0htmIErzsI8lQ+NWmrcQ6Wgp36kf5Ej5j/+5V3I/qO5yMZ
UPPQ9biquiWiygKHK4FPjhfYOEvBB/FJ8TYbjLQRYx1xs+h4XypFSMUk41Npt2sF
GfG8J5QIDYZ3Asr8yf3cu8FFRiRxBf/N46h/TuHa3UPM7W9StfMlo3ilCr7FTRyd
Lizld9fshxzSh6p3x+DdNy3E9oTR9RqLMj+AhcKk5lFGJpf7XVotMOA+vaeNGGTu
6hZNGB6rPd5l4TDwDKCwtPAh1t4IncXVjFtTIMvx6SW/c3Ugu1DHYxYjVofG5TQQ
+ccnZBu1avLQvNxN6JTJzxzldv87JLk5YTExoJ9P+kfbWfxB/OtaOopfUxO4TRMM
YBhvWnhZBmETbOGpbbqDSMIdIzF8RMkrIdRlQ0zij3n1K4ohPX+v0V2xXMM9FT4k
jQ3dbMQKU5uoWg3CEyChFzBE1OqLjde/RGsl5wWLmTt5Tud3e/Fs7JAzj5C7aCF1
KkwCz/ssvLvM776M67C3bWxP3rAq6AhVDVCnIvUPCMaGP5mYrI6HW4wnSuaIKWB1
w9TD9pCUEivviTwvzlKZBqdOa6+qGt4WyyS+7I733YA3NIQzHrNpHXscaSvxUAJW
hWgVBOJrEPElQ3I8o1kLeAiOnY7TXAiwrak/zND9zL8hcmL75/3K3iGXbFNPjZ2w
hEVBPpApokmgwvNrzahrJZiwY+fghh7n15ayYgXd3ym4DXHINmHJ011lAhp2wuSG
YlYy3uN2dAenLr/4eIYEC7Ofm5FoDiPQ0NYB1vbXGSpJcyBoiOBYs4/TFDq5nspM
/0J15wtkWxR+8i4VlciLddNoFkhzIT4f0e6uzEJLvz8Rs+WB83sGgWaMueUFWBJs
u8XaLvL26al3wYO3cNhDCV0EJZdOsoHMJEYL6a/5kh/NwAxVcaVXA4HLqmKtXQ42
p3tWskrr4SkgraVvlpD4b9W2NWtywHOtfQIw1uefpmLB2EEmuQd/tRwfaqgajnzk
OC2T4H2j5urRGmYpom5BozcSJo0VGFGAABtcRE2o2+ge+bBdFh+hvxI8mPbDK4w/
VRErU9oFhWBtCLAM4c6RwTaJUtUh3AZeD3kMlNGxBHnFgfwE8y4tCVg8hjD4D2ct
3vjeE7nFw0VthwO8Qm37VgyYLKklDaS2LyfDI3ioXEturWed2OggLIvJeNuQcXhT
FPvBp+3sQOaSlUqVbdct8SGWTRTB54ddBR79b/xaYDGqfprJIwgXB6/dTb1eL/4r
fwwlPS1jnqYd8MO7XnIN6eGizdxrQ5u77dd8Ga2YTTOMCVxyes3DFjd2kbGFnHTA
uSwM5x4t7HqGzmXftJJ8bEds67E8LqjrFRBJuot5TWWZQ/THrbaucv5cnlRj0gZ0
BdfzSvOW/S5D9lByLCRQL4qlkCrlU3164IlKaoWUlClC3KROfB3NdliXR/UPJPES
Q44/5pNBS2esNT0Fl9ROl7KT4d54u66GhOIyz6lKmS8+UEVaH0yxrTnHnMQ6DIkV
V7a6B61AkTSGj+fFf2/7h2WxMbuHmdVLF/c8Ukl9wNO4nKu9lbRIXNVBLqBDa+2A
ls7e+/F4EUnxQEunzqynsaqMw9JQP0UxuHNuOb4JCKx3AdRubJiOnFq8SLMnVO+Q
FIMf61zoghKW2iP6nnjHEJp8rudeLoDO3Yx20x9hfdPcvAdB94wtabDh5bT36GHD
i/okkoi87Yxmbo5/mora4+tXMQRtGiYy7Va/m5koSIc287BWwRToDTMuv6ZixCVA
2kTMtDFFuH8xL1LCer9KA5rBslGntdKNuwdrhHpNAfP32WwmQ9kBXxZ0JRROdxEZ
FNlzG1Ew6gbyv75B30RbrjU8fuVL0ugG9zbyB2ow/TmBZVaK5zOJ8q627Kx4hlsL
BRKgjDbuTam8u3hiuHoBIdxbUeRDN0Kf1GdzkPG8WRg4JyUTM08uSVL5mHkioG58
rLTNHuATS1ZVRZBjCuQfPZv+aTezzJOQ/YF2+qJ9h2J3RxtxjcgKn7/7d1pcvG5Z
7vdj/Hy2CYUoENe1nypQCcfi9Ys45DvcAOhZob1VRaih/373r7/4eHdg67ywi5uM
0rresAr0Cie8ypWCO0Asp8IUOI/DMo/ujMYpKRLDMMFTowTiuj/xAnWuZQdL2Ro+
0uvM2qYZvl5wgr8xlqv01fofliNDK34gCAxZKoj8Ha+AjXl1lIAyYHHWsgXIAOr2
E2rOCabvP+uOp1m5WTNRI2L4k27QYK+9DMyrlggxoQSxSk9/3GCrmCqwPOlMB1aL
gyHBEuZml7v1dig9z6K1tuP8jShTMkr02rDbBBbLi5PKyd6HlrwzJ5oYZwtUSNzF
JgIfni8m23IqwEUAaI3U4a3kP5O55YYGYxtuHv9+X6kZTTjjQBoY52y3baBhgd3X
uIMlvtTjrto1IkIxiMO7gXDC57MbTzg3gsOsita/gZJDGs+l4uV6f8SodP3y1/Fg
DbxrdG+pdxWc2yU0M7oZXoza7paC4+2GYtElRkV9onq2qjaq9wdt/iqqahz1t27w
EACxAKi1VtkUP5jXWLK8cOCir5UoNt3epCJqXYfcentnh8ZKxkthziPT8cIFM8Y1
qvD9UgaRei9FpGgTWBZYpkx7USVxQDM9tvLTLOR1mfa8SKFMIBETCvLX1nB0dxSM
w1TWnhHskg9u3h/A7sx2u42+fCv3pgf1a0QMziJ22WeQrNpMKKeYIGde+MWLOWbU
y6Bz9KAAouDzZy44zy/LyH27Cd/JXXw84YVbOBM1B0HYkbcR2ep/LZjDchnEiaWN
PA9Q2PrWUyg0vYH6xHvJcbm3PXKWGoWxLs5Q0uBH1wtivFZ3LFM/bRP9GFFho63/
A+wuzDRA9WTq/gb9ksQenGmIffFozHMGRYHxMKUG4meKihDDkkUWNUp1VVKSLQiB
sbpO5HS3CLDgtYduUxINHWq4vS/xNJJWiNp4mOoNEapx2+RC7V+wdaI3Ug51+ohI
kSLCNIkRCLYoOvl9zGbF70X5P+ZEnzYmwYJDzJOg5kHLcrfjPx/5KsazjwYoHw2y
+y2vUGffD3cOxtvpC1NzfdrNWNx09c2uhPhDs+R6pgHqxSkD6gmQwV6IoXol55+7
zZnmr4Hbjk+X45PffArDJa/hyj0ec1DNccztSPiWM56Emc/7Nqye1hP88ycZ5Bj7
PGGZH+yXPfpY5gwtd8YOU219ywdsm/wvICkNflq81a6pN/DgLWf03v8+A2PAX5gn
goXMCQDDXwi/yppMdwbD9hg9Gr+7svvkULiLUf4O8f23RVE9xj0ZXk1DwRA+2QKW
71mluKBu4F/sEpfEXHkrm1lhiNsT5JqWB4Sm+mYVtUTPzKsjdlL2m2Fb/bypqmYr
ISzsZ2NbeHrldIgTQHoF9bmjIHx5LhPXYDc5ap08TBwj6e3E35EoEOMteeLp+MU/
832taNdlJO29kDfsiXN9212TU6G3R1MWNBdmMEN7PmAf5ah4fi8VszlKPfg99mqh
KbZsv+/nhw/n873U3h5rIgw9CWL8k8NepUSJVoLLuoq+OfW+yFaONpOXZ1j4GoIq
gD4fmRv1FwhovnO2SvMydVrDn14tIBSI+2sBZ2o7fpmJn+PlkCJL69f2PMUU8Jl3
qpoOQM2EoYbFwF5cBt3x9B49tAPEAd46lNyVS+mOlTuCS+6fdXl9LiYqRcveAzLk
4tbPVrioOu3Jp/w6CI9ogzVv3tXdiLMR5dt4gZcR6o5FkpZnQr7tQwgLZYyEvSIo
MdFB/jmomXhpvM24ptT0+OalP5oXEHRIrZ7wXnGVlFfiKWNLC6y+d5PoHv1a0jTj
gdsAsn2ApkpfBt287NBWU4zGDPxY6BcisIN2ha0BXsNzAEvhfqXWSWxtbLdQrW/N
4DzfjNuZPq0jYzIw/5v4nVFXWudQiXxwdV7ItLzAX2sybLB7TP43X9R9rhHos+dC
N4FaZqQgJ7odcg6mQEkzvdDa9qoyqg9udmw/oPA+pT1uuvg+ePYZTeuedaq8jtxT
cZ+0PPVX4rQNr8vxIOyqSgavz9TXxt7gldWSMe8NQ0N/HklkzGxIzUIx7xl6sQBw
w5pLCL0+s6LT7h8Q+PsGFcX0cTopLdCxFrY0wep8vUHyrl/+ykoILuzP1S1fDHwz
NtO8y92T1SOZebrlFsCI92DLzyWq8IkrLWoaCsyFUuIYKzxh045yURqT6dUcYDey
zZ9YGfYVgc/N6+xPG/3c+pXY87b8vPg7Fpos4t235x0F0vMGv0/eRqHvQOYBpqPL
5R2mPVb1iHClBu1e8uThPe1oLRmACxo4tme++h+fVjAPpmy50k3uXlFtrcTjpdGV
w0et8EJK90O1nNCE7NX4rmrnGBuMr0+erTozzquwM7mVC7gkdWYm7fd6rhxS5cCY
ZQ4Kvo5jf5ReyxICcRJ8+U6FHeAbIN18+pile88/Jvjercb0o5/DnyHb965WExhu
SJi+vmUK/PP8+v1XjbtkdTkd0jceVv68VhCx0bLfv1Z9ik8syo7qCsuwXZA8LXWV
FimhbccB1h+W1QADH1qOZuVhzxGonqDR7frwF1x4IGlOjmAAeO7Y2GIMm5NWtTGI
D57zNViAj+LO3yFqHHn4QXonsS8khl8nQaLwJzkGjVPUjxkvzX8Z7JLSTRWWeLOH
PcWkFow+G3k3DbJP/eX9IPiyW/vKbrKBR7G5ICDVeuQ9d87E8v7WuqaZCxoU8kyh
cfq067rq8q7joAkznbZxQS09VGzVLExhd8PtgeuKE4NU9iVHzNR3o94kjUUJz4f1
b0WuOpMgp/dYv862SARESk4MCjDSxgEZ8MNqwI2NeOW62xTB3EEaYHY38rp7Tewx
HgbC+gGXQNOY6pu1hRFd1DapIL4NKrZq5pjvTY2XLFf9GxLKORmP7RTt1WCpScHz
NhuovwdRFCCpq7rWLElMbrrmtPu6XcJ15nLzIeIYW5AGia3CxLgSDdcNw43nyBMb
WRAjEt5Zsh80CYIub77xoKEx6XOfYP3fG2eYBDpGMaQ/KfTGjh6gYJcGWemscs4o
PzxFeql2EGMVfVasLSSIEE0rDygXfC6x3TKacReql2ZRUe2D5VdgNC9UwIKg9OLs
93R/0ZPDKpmZHG0U5+gZG9wEna4o49u8+wOxx2eUGYsT3iRAO4cMecrmMySgLVam
yG3qkfCz6c2zvV2YnbuEAsV6UYATpYwZbY1wgrzpA+2gDER9FbhwrYgubASF/9Qb
6zYfC6YJxobQ6TkXqs4pjWgRPBP4ux49BXhD75DXFF+EPinmo01JeIA4qWEmOspy
IA6KR0jtvJ1zA20oK1xsz4u4p4qGlIc28UXPGDSuUleL+FGPpWgFSRjcVFgGzOA3
cB5gQJkoR6Rq0nO80XE8ojFQIC1AudVJIu5Zl4EHsUUQPbDTQ+6etAZu1CVuH6CM
M5Z25NbQLGNtWA3HJUciGeNqUpXVgoV+f2KZ1vlST66NTQq1NXPCWNK3f0HWjnGy
OVGLHHOppCQhIPB/CJA2vP/+l2kaomdZkTJOPGmpFkl2t/7ym9cVt+8k/HHAMars
5x8J/wYkIkZilxh+LRU2WH0OnNjF6Qi9N2zD3QsSwCzfU+esFBTCrZtzVMzFdSKn
1aKRKqNniZwXMp+gLbIMgKulX9Suaj6S0Lr9yAnvt0YFWhV+e/iC08xni/SYtOh0
n6JoUsCQt1rAzbim7j90cg1J1RnTaOHI0zzSAt0f800UTcHtY0w4CKmK7VEJM9Fd
QSJkmNP0zbFrZs0v/aZXWnEgLOJN2P1PxF33C37NB5RVJhdnkyIbJAmYx8WnvXdp
DahMNefsHgyfrpx9QZS2jT+J6Dfnw+QBEFzVBb/VQowABu7uoJbkmZe6I4QpB0hA
CfBR4RV2fEPxqQ6gWxTtDgxQaKKWDZG+KPNC7UZjy/o7bRTmU0NAIp1M0C82IALe
fJZBXJUby5e0N7zgjWhjhzD/YU9dArZX8NXYXPZx7YCaHOAsY+AHClxp0xS5TN6I
S/hJJoiJ19CbocrWMu0KzvMuc/T8ys45ThI/2I3lAY70zHKi9+JyHiGNUJ75ghMe
lcurScuR284tDjdBIdnd7ljMn6lZOoLcrDOVzCQLAxFdPkVBBQbydCu8hzpk2TXI
BoxXAusF/s0q49SUOfnKI88Q7S53h84sE3ZczCGskl6zuvbAWec4k3nQGGwflcuA
DeJMd8T/gNehvrdU7Bay/bpXynE6eGb0/rLDJ/sPSVe079jz4MyxpyaiDV6h8g1a
mH7npP/gFzGhQcvXvqNmU4mgMDHi+2BSPv5z8eFugBnxnMjMsmmoig2XgGfuOmm1
QtkA36B8DbHTCi1CRKFzprua6RV+4vVBYFRBdP19UqUKQbPezS7csFSW40fLVnmY
XJ/sHlyKqUj3k3gqEnsLNFluUNXnMtwJqdNO2za9m2U0R7hAZi9VjBYHtGkyqUix
mZQCRMzrjc3d8vTSeahPy4rBOMZWnrf8zHrjgQmJDFxTrLsccGI3GP2xyprys5bj
E1sd0XTS7kddpNzs0Q6IQEAc8YStn+tRO0qQPaxdQ00jCRc3qgqVzv6aOaAbEPv4
6qNMuo3E983uq2uysLJZtqAKW93jd6O+kzqt3affgqQAnT1raTB8T5/sjpE1YZ4q
HnSOkxWgtp3yrSuDtqxmbZzNqFBrcLt1F/wmUCucFQV6ZFQIGPjcofP0RRpvcUhT
/Lrr0RekUAbA5eZHsYjW5rn9k8Tig+K7ILOio/bwswTPInthgrbusWeEuJqGzqK2
8PUhVobVQnZhhfYvJ7zVmc6dsGKqPJHJvAYslDe0wUxhk3MCz2Z9gh1A9aizapMK
5kbAFuURTfA0u83g0YVtKMIih/oY072hTtmG170DdRbHewhJ8vsCxPmCVaPsD+ea
ZtjRylHrYL08WhaJlqfCRpVAdtD4RcxW8zAGm2bM5wYdZynqLCUoenyIpAKw8Ib4
VKybLDxn/1LVlDBAaSXtfMP9BlZu7aZUIALUEx8PTfv6z/tjpRSdOHhxHwhR1/NZ
npO0goO8sEFFgJiacnWg7Nmem4Rpp9nmaWsYOMEw3T2bANuoR64jD07dIW28PUNs
sMwwmKhAbQuKfGLQcElohXFXjig7KwNu0EqZ+ORwd3zNwOCq1clQOkje6RDz3dG8
GTEc5Zn6xLbpQa+POepJeDBa1b9T2PCBVRRUj1M077v2QkOVPijdJ5t+j16nfxPt
NwZpfC5pPPNBXj7+BU6o6pueF5HuxXtA9FRbhSGWr5KRbusT8wL49bSGVvzUr2GB
adiNevVJHZrhB1S9q7YHErl1KTYmfWjTGmc/ReHoKM2PHQGTGoJaugywaPHQ8jpv
RmtYttiMktrQzL8LlyLi3g2Z6JWcKlYvMM3EOmtFpDc3P/txpNDqZBbOr9Z1vzZj
QaAi7acegjV0Vl/MzsVkKmkaRq+aPscHqhpxr8XPrRrTyb0PkvOyo8bMm1jKmFvc
S/Y0iU2i5L0F5Qv2bVmvFe7SRXR1loqEccz0Y1z5pfoqB0bK+ZRZ8PCD12awcZw4
OoLIxMJtARptq4iokQlH4MNx9oFnwrpL/9Ji0yAj6IPRUOT7xDYsLDNEsVJt6/RH
OkHkOSd3mQBljeeARyhIcpTBFCMbFYxb1cQV1zRjP9zv8Kb+e+EG+VFUBcS1Vu2H
KJrMYYsaUeftDlxKz44sN0Xqb8+BrWptWKMeU5ywwJJzfmSo5WPlx2uILHpiTCh9
7jAhkpYC+37sdrc3r6mPmayBdX1SKMQFfkneFDAUfxgtoR9oHcIRW+MtRw8rEizb
M+LoBvO1ESTR90jN/aSm1HYZ7YA9WQorWth5rkGJjS5vzcAPNODbCRAvtO6yO+pR
jrBuddR+Z2w9DGYwj0NDRm/MyNHjxP2qLwzhO40RdhkdK6zCRk54/+8Km6VE5mYO
KtZlvwPGikuBC4m1oWuVN2ZsOAXe5S9IA7OOOHKIq32IiJY6VYlgt/gUyPpkMV05
qexMLGU0j1gC2NdEEzpSj90fC7LanJvSKmz4TxNSEog8ntbgXTXAF3cWYCBKIe/i
nOxg6dLVNcRrtymfg/KUibF85U3u0QEcOPa7BFnTzVKeSsCc/jMx5+XFd/g5redF
YpG7DyLk4iLWSIYlU9aHzAk1okGSKUZPGBdTKsObspU7MumS90rHSR66PFuquRFF
Im52/QgJnEoW0xRFbw5/sh0Y/6E09653bF6+oryegDpQeNv0zqVfnZvxwPJXUO4C
bsUh/Wp78UX0tRc7A28Nz2JDe9Qy5b2AxETEdbtfFEliX0cD1okfYf1C9s1ynU9i
liYidD9o8DBtXr2ab02XiDaIRVkwhP6FFQqsJ2VfKt+e33auvsxRFdavjuZsFMqj
DyolkmfgtVVJ4NCAOoUOwuZqr/VOuQaZDz29rF8OmIm6e1oA6frY3GzocV/fxYOH
Z4plD/KNXSmaBxxlygJ5P989rvOIgRFPTky+QTualaIBIAUdvTP6ih09YwpORwRr
39zP4iF13YRQz+Bo12+pP8fEq6XBPDUjRLfXA98Akkw+P1pGADbSa0IJHa5cbhWF
gXmypXiW4C1zle+fznXOq83CPGHFmHZ6RmWKUhvtstbmOzU6E4bUsWnnG00I5Y+B
w9wzIxRf+5e7QxJhhDLjMNraKO+t4E9uZK9BkTq7qEICa8SFwT9CFtopV/SneluI
mcX3L/RGBehDZGC8wglR+rSMHotxd+irHmPsVeRGsPL3CBxNFW+JWiA+q4dDjRXB
+JWfqgXLnIkxSPNnOy5n7i6jVaDn/iqTq7w7hUtIWa5LIKSgjdtbnetF+aVDY11B
0VfG+hIuWysrup46r1XOXvdNhkBMrMuZXZYuq9VzXhOLtwj8L5H1mAuR3MQEJvMA
YFDVkIwB8eJx554PtDRd240ThM5g9luy/Y8XLgYnenDBMROEOilLS9HHjyhdBJtf
9IQvBvIrUJTbeyIwHq0HyYmVWyNuKmmwSzOqpLLfNm2jePz84mEXyV20xpqgZ3OY
pfH/UI9cJxRzFRQqNwNrNq1YaNl/RNy0X8JKFBiI8s4W3zc2Zic8mL3lX7UokJsO
X6vxu9ctUuNxqPSbEMFzRphtFUkNojxYuZ5EVnHKBgYHFB2ktmxok3Y4DtBmZdkQ
`pragma protect end_protected
