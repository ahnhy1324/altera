// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GHo5+RmLiMIaGJXgTSwye+RP8Ku06ZQ07aeSekxP3MaCriEL54jis+kGM9Bnsuj3
0emXDWfP5C6V0rb0//OIk3zUt46Njb8HuCjF0GHsMAgH1++sk/s74pi8PT8aVR22
iDYQoaZpn1lO8wEQ0J7ckZBggGU56nt6kT2kbPM6k90=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 63840)
BCR45BG/RhfQRWqSIc0FRTC0GyICZxGnkjJ61kF1Qy2HoZXAL7TBqpUIERn9v4Tu
HM3xaJzI2ubsvIdhjwovEM9b8dZz1xrMaNRDQNQD94Y8cV8xUvo8gWvOohcjPPCI
tYmR9rR8fe3O4ASIsUouajJe6qKQ2hWDkjv86G8LMpv/fw8/7jmupxbbgYRVKka9
VxpG77i3Jx88A34GRjxKf0yTMuPJfpMa6UWzXAKFsLZyeybPIOj4mthrhZubTvpB
2CN3rbEQMm/Hco0bKC+B2rJd3hHKjcGbtSo2bKK0MpG9puM8mvOmmP44uYCisRcf
lkrMFgXmt5pFF3myqjhxn9uJckpRnwpGoVolgF4XmNFPU/eDZHuHyiTVNoJnw5Yz
bQL2nUCyKPd7VZKM4SzygemVm4AWg2J9MQm3kbjoCvvUJbtP170DboctMhJdEBNj
Vu+bEzQpLP1cHM1b2WUE3GZnN4UsBcmjXHSxk3+Lv2Bqcka0ZE2gkh/GMNWa725u
opbYcrhse1qKE0vAVegIz3Jo/RNrw9wDP/o/SxB/yd/VSQgoMUSJh3JYp62Roqw6
Chfo4DtZCUorv+ZpRSwLh0Nq17C2eeWei7KInPAMoXYATHHmAGaq73N8EgycW5lv
hTyNK21RFBDzYUzW79RA3TauHooQlX8CrHtxJqbv+KPzes/UoJ+F7j3iPrT7r6yP
EnMUy+mJKFcby+cbiLMSpPo6cwVKPWo1miemQw2SHoj7d6iAPtbRZXw9V+1kBV51
p7lYIczGMgkS4IATM9hrOFX7rHNwN9CwK+1Z6KXU6SSeKiYICNl5OwcogvDmqyiv
aMbJgpGGHhc5PbjyEz/2tcwq/Yb0hRxDgZBMeLzean+4R6AoSaXCis2EtLWbxf+X
rGK/PaIcdGhqU6VN9/A0Njq4vfFNJ/O3ZJCYtCGfZL8unX3iw8fCUmxrSRwusmdB
ryQ+rBnpJZYCZJq+r8RYANyxuARq9oR/ET7k1yGZHV4iqWiamwsB0AqdD8rJePLf
aZ/iripohngTPvaFRrcl5yNZDrQhosJJX+l+jKsR7KkVO/zh/DPhEWEtD9NoO53k
1a532ZY9vt+X/3iur8eJKAKCgrK8Iw9QLWkP2pl8+ZazlJJgC9tDt9ZBV0XqvAae
GQQBUhj7WQwcLbZTKjwtgFaaPwUDGlu6rci+2ZlnqOiSoyl+EnaHg3bWL7OOruoC
dQoKXb9BmNY+W9/pDoTo1+aTeIObWvUUgtH7dy5yqOFRqAAteWSbTB5UErzlimEy
1qZgEui2pe0/264CKACZkcLGAEAx2a9bieCoujrkfJGZW3wz8YKGp+zS5GhJSjPG
B2tIBIaTINVQicEh/++BhCQElicXjmwgW5Z5QsYD+tYerqaKt20i4xCNWlvE/p3q
N8ada9bSryiTJDaOEgcPEow+Dcvr3VbN/j4tctEpDGCgr3VwjQhawJv75IiRGfnG
YGvf2vK5LUWbXMphPwu1ZB0/d1kNPOcBegyeWmCgCUZPmxxcFAdr1EiBzu6ePbP1
d0rDT0hcO4ilT4wbPamXc4F2LX+EE+EjeZH3t7etEOD1iqQngMZ87b4B5niwgBjN
YdD3yBWQ0wIMexn3CFJ0vwy1KGrhPNDtX9080TB58U1eTqO2sgcOMx0nIgGIlaJq
u50oCPrLSOIJ5QBDg3OmV6vbCrSzBG74RM5aaaDi+m49uN94bpYT2aAMxSl9cNiZ
hnXLtG9L91A1Fqnh/Qe0aJdABHoRvCvu9bbDWRTOwQ/c0jL3JssfUXUJ52PKDKC4
j6UhkPnYrOUFZhZ+FLhVVyY7uYoGOFXyB1xprsywyfnPgDOrTzQWGWZ0fy+4oLlY
21ZRs0qxv6dxhoSsoXxrMHKAL2pUfAfBZJIqnL4+Ia2l0RTLjEbaa8M7nSONOd8B
kLHUuqzzchkqM8blfqchRh02QqD0N+0kpU1+PvfcumpVufjqkJiRsYao7xHArT/K
MSzz+SDxmQdj9qO/R4bjfWFJ9OBgHEj/SRXQFpFVJ7mfHP6nvmVEBdTB7GWiyqyd
/I23PIyDY1XjSaoZtjsEiW1WLCOlguJPYZZx1/Qo9DCzHMtTswmn+hlc8esez828
h4P6TdnodQ2u+4OB/L9+4s9kM27hMfU3VRpnb+AlOmmvQssbU9KbnmlA4iIPY0yK
b1OKtiOsHrytv/EkhTKesY6y94zUTJSJAeamgwXRr3j6+NVYnZSanICb2CBVo3pY
lJpjL1X7fiPcEIiv8qxvGfIwr6bCiu+OX3g6S3X8Wiz1xEpOS+r0B7foGdxdeiyU
+rxD8yWEYC4SCwdd6E159IdpCT//D9RIyIwquvJ9TCIMOkkgfgMxGBrSBNoRa4dZ
tVRdOtj/SuCWz6XwhxaRhQTg1uZFUXWOWUysndYuk03ynDYXhUrl52WwSnPWEytJ
B3HlcWcXmhhFxR7buQZGfoEnv9bj6K2fq3InL5lghwvYehAKOZSIbdP1TI8oiPgD
BWgisghBLBT5a38RFlyOfIvIsTkNzqswFBzhPBV5UpR6Sy7mF7Bq/Up0s2hH7WwP
RCEhVGTEJ62tWC0HuffrsmE3B81axLKrYVRr+j1DRejC0gmdPZrnpthWQbn59W1T
rHpbU2mJYaQqTit0OAzCv24bQox9pd+YSVocIfT7Ts9hEtCF6F6Pva0bbLan/ulm
5ZXrG6/0TuIEYW4gGMBQS28y0Yc0R2op0N8dD0SLXq7ebMaSRSIRiaSC6RM4Y8C3
LdNmq6lMGvSuDdm5Leu5cS6BKUuMZLd2LsqSVBOk6HPbjgOs62/MQtt8/zTYgrQF
b7gEPtLWDqmA3I0OBnIJOhZ3wWg+Nql4H9Syw9meaU2hktVRwOF1f7CnCTLv2BiF
pueW4EuVg90h/njEYxIBVoH6bEmBfE3SkpfnUmmttBFWrBIKkMb4xORRg1ULuCjn
y8WXJVHSlUfrz88iHj2j/FlX/AWzw+x8zpZ2q5PAUeSY9e/MkbfrXINgo8vonPde
9K5Pn9fp3bZqh4N9DQ/Ym58Sm934Hqu4gcfyLto4eX1rIzaY08GcYpZbEZyE2rnm
FhzBT5tm8QEddmPCmWjJgLiNiKYBl9jHCsF/PPhXzY5YChcbr3SuAUTP8WZbuMky
GW9B1wveSvdHVijqLGeutTTgm5sQcOca96Ns/5zt9kYavnjlH49hx5bX/TIJG4B9
2LlBnNZgOOEZ2vUk3xB7/i6+YFeaubzqLKtGsP/70n6uEKc+fVHhGcw71Qdd+B4B
oxLJXfqhB9z50EA85Ydco4XysdW9xOF4DmNgfFJbq4FKudydufLTgbg59aFvinKw
6NIFh6McmoBJUAEk0EouUsKJSnBN7G1hRkIHvZEfriRBtahN8/vuHDgt0lyR97vw
x+ujqD45VHeF71b4KGsDY4NShfortxFInCJuzY3Y6eDA4OryDdvlpB81XBBwoP14
jWX4fsTXFvLH/j1MOS8DbOfGoyLpRW+Dqtyl+OMtCJ2xS3t7rleLPAC1JE4NsQET
KIiaRXh/guxZal/wvDoSR/Nl5MRhZgfB8TvS3JkWpbIlJ61x35/DkZhfe7c1Oywk
OHqmn/l2UX7/X0H//FciAbm7p6Mj9awfG9FNmErrsRow/eiXmBYshtsm/U84yifH
/Ugxe5iPxlnwfVrU6FN4g0GXcuicnJHoykzO72Q1EoTkMq5lMuGWRxK2d0Lsl7rL
Nxqjcpjfhb72YlvI8DeKYUwYQ6e2o1U7VdZkvSkGMuSo8zZ47LywsMahRhSnvLK/
kNyWhGDPwPNx6487/BIkcImjD3NewKeMRZxBmk3nz95d2EeB7SS5MdARS56MuKJW
IjzAiJ6GAr05qvAjxo5tMgrKdn6OxTZXeBYEoWMaXnT9QjZnEcxWPCe6Twp+xprF
ogSECjQMyOYdE/K/uYyDQf4XocVmAe3fkBMui0eqXBV4/tkOFxKWx6qjdGB/HoH+
xCVGLhjg5gl7D5z/4TeIxD0cCdQG+yFTxonYXdzXSomsUiYw70zd+T6wdZJAtBYG
KfusF7duaI6UVSsc3SOtv3elbQ+Brh1yOnGNlkUnBWbl2rbq0z0cju6s3+rzYxiE
P753F+fNLDma1izgBFM8LMb95E81froWWHfDUhHlNdcb5cxvwCNuWxrR/6HHtpOt
C5348DjIYKTuUnVYG8xPXFeEPuShyaTsRA4UxuNaUYUWaq2mY1y5coo8MuQPf+JL
knSOu2trodtHN3oUkhHDIIbKXDR0ToxHs+0pRVvY5FCvx2P11nfyLV/k8t1+GK78
CzW64dnAzTnCr9C87jjU6bMMEv48Sn352rg/+89HNtKhWYtrOhFVr35PLUvlRUet
uPbUFGeOa/vzkGalX/+rmt4bMiObDmEVdWhyEJz5H89aTapCnX7ZaxtmgAZ53X9c
mOpQSIIPVcNPc95Azcbr0FTUjcucCjkKwexEmRqMBxK8A+VHKGeVxUnTplcWH3AO
tgEi7Q8r/zYWRxCkmjanVM/IArgJBjLEqLQVsnKTCS5s/7ThinzE74lmlkEREVqg
AwOqFpgAtw2nZl4kUmytH4z9+Rg47+1bzey7KQyNicmwYla6bwNGzsEQuOXZA981
Jg2r5hVgY47dadybZfDg1YS0N7fpcUBicPTwjI/Hb0NftDvBnK4+RlTsRPC+AC/z
cD673k7uXShrc6wXoYL5BpXH0kMBYFrsW9lGngtcp5fFtRS+grNH1S0Z3blT5rXn
2OEdtllpyv70d/IgSHRspnoCZ1tA9e92JC7JnThgkiPXICcd225U3x6YtRXVPyUS
AhdFQFAVTt6Fc/Y3xra0ju3rLmA43FhX6cvNsUNqQyb5mfXQdLXKQIL4TxSM1QYA
qo7lvHWHfVv6oIb0KSj3Ts0eVMCRLDWkev+mugfVNVA5rEJE29OAEyADOOkpd/s/
1GbNMXDxfLvAuTksYpEt8cde2ZJBWNyNU5HQ60hGBafR9cp9bLBAMQReFmFI3u4w
upfQbh1Zj7DBxzQjCtA/6ESTuriVXiIoRp+za4lpFFzfRIQNluLRcPy7wKKqTA3k
nSTv0Fvzpa6p17VTKXoQ0aVK6mWOD4h9TRwRCcBvpsasnAcPcBqP+F9eU2gravLV
3VOHj2YX1eNs0hLOTg9wy4Mmht8zyP5cK2oJhtKSujq9qXGCwiCMN8v5eaOVCUEL
HcSbQjEurvxptYyU5gdd9Yy1RJQlnmnQn6pCeksj6yjm07alFLAw9ULU9Cp0XhBi
P4Is6gSz1KAFDuqqeOtfc7B2OcuyJ0TvCEKYPJ/Sw+L1nAG9j5V/Utl5DWFBkpoR
YJkiNZEpIzRC+Q3cOh2Vi8QN6JBVjXS3gLJysLLLbDr6NvHmtobv4avTLuig3wmQ
GqXQwi/KX1ckyvtMV0TKxDf/ZsNFQm0xULOqlcxrSGzceJxtxUr25vpWOLJP6qlq
q2tGJiya+T+/uvaL6vhLUzDitKiPhvDlcmMyiJtoQc/ovgUD1eW+HeN+Y118m2zC
OSQ2PoEoc2XONagTzMxOF2DDa+B3Pa1rSgPuUZAgAm969OgKGuVVOudALxwPUcsl
dieZ44o8xHzC2YGv01tb1R6bOBFnjASdGwFHKLmug852nW7Bxf+sVLIWA7a9rYQM
D/ZOP7P6liJPlVkLfM1iDUR+ECY8nL1ruXqkUn+Q6fQOKbcu13MJr1gC2tYoEwh5
RKHU6BM7Y/Cf8saAUCQYSUfyBCr3lkCNeAQ8Cy/fZsw9CnZ0VN8JDhKPOyIFB1q1
XWyO5/ep9oyRZsNksDrrSrLzUGEQI6AkHW4Az4N42J1svPxVxY7igIo/pQexftcN
FjvLIDQQYizBZVPeLBbGufeW4MCtR/0YOzDAw8OwlJv5yrb58WDyKY3X3S7tFaP4
k7qvL7qKI3TgKEeXFgj4zUawYH6KYL57XlCR38SdF5ss/b8gTBljX+DRh2aVG66y
X/8r7VbCsUTnC7TbF9tadLFMENTdxqr/6AP1Nh3mdvuG/cIeOBUv/SB+LM3pf2Pt
7cqQI5Nh5aTbTZHv/T8d81+Kw+OTau3MSretz51ui6PZ23BV+I+Kgk5B/x7K1qKN
lYtlEYKL8PmWllkileVJQuhQF++Ery4M7D0TkBYwiH6iEAZbS7MqBD7TdIDINo4/
vCJ9IhnZKl+1bzdOfN+mHnwcgcMDUj/D5/jyHQJVbHJqnP1x1aRa9/m6TL4ppZZR
R7EsMi3GRxaoNHwmcUsBMOiioKMwE+vTvIB0C/PcwhYKZ8rYThG7WksRRnjr4L/1
muS7GZt21phKIKrPdbK260jZntjYnjMqDrC1EY3R0/0zb1fGI/5dmrBfSABqEpAU
7ch+ZLQvpJBUzOvrwnUJ8Tw30XnZwUFU0j10C2aDfKnCQUqolhL5Op2rlT7mlmnI
cFUKJxcCsApl25/8aDkb22QuxS2zG7ae6Hn59iaKJz8ZJOZJmt2Gc1U/eiKPVMmu
Z+AJVndKANZ0QNojQ9sO3hFk6TSP5S7xyGHDS7bkmA7CMBs9LPE8uV8Y9YJ/rShv
1KjgixPABxkFRuDt+hsNf3x9jP5785mskMcDOFfjlO2YZatRpQc9v8Ml0NuTyiTj
DuNhTRXgd3fBCkvdXw6T5UdeaJJ+ABeyhrb36xWVYLur/OHeL6DLUMOgNpemkCP8
YfI7fDHm/uMk6iJFgtsyfBhKS3AW9KLNjeFhYPrXvFklJHkgHlurFmZvcv1Flp53
Xd4D508cvmXkCy6uirGT1zoh91RObMg/Ke2cTezWIzC+qg1kGGrwMXSx9K0ao1F2
hpLmzMCjOlUx4ywp+a1tDsu9QkEyCX21IrQn8WGROVRPNqsS/wQmKM2ay92wm0Vw
Bvio1mE7sqApLthrMtwOD9JI9jq23o+hkvFQbsqLUV94BZ9G9r004LnVy6NxiBLM
tNyI6ngVOWvx0XPldQrYAcf6KmSmkaRqnNgjxcJ77sTxmohXYQ5PJUlCkkUxrt/q
Uyajv9OqzfHGzO1fUl6yrJpKZk0MQMJFM2yiCSpXuwxDPq2eitThXMZVHL1KdXVz
YCVWHqfTrKsmVXG+UOF792eTxjgYBhb8pOXN3uXTYj13GoeoGEGG4TdGIr5JBzlz
JtBeB9qQ6JSxzH3B0DCOGHWeUJUbscGHCMO3L4qyERa6+K8L/hk2Zu/GX0rcUada
ovgYb6bCYqR0hrZshvnJMORkGYHJF7QpPRSYIvk0IabobsaWBaLiHq8WnnurEAH+
UVB2TP8NR49hOFpSZZzaL9aPTW91s3J+FaCBgxbr/5YmcMLqyN+crrzePWjJxegU
a0/rm6K7Hs1TRVFJAGKbxkcy0pWlDOep+gFRNQnfZnPnqhS92W3ouoy0iMmHNkn7
2mMtnS9yH3EMsw39d6q9pv8PkvLzcmWimYhcz9NR+TE65cAIM5HQYYTkX2OdI3r+
UKxwj8z/MxOtBNh0ChqrXVHGrlv6+NyDknWOLfO06mHyDo/NeMNP86S4+RBJBxB4
DmjAcfvcAyRtL8adlRpbNYvOob+q+czUQwtXNb+Ud+yI3E5nDMxLf4H18yE8mbL4
Gzf98p5KoWa5B2QTaArpu3+7urnxGQP9c5CvrUp1a81C6p4vNs2e/Gl0gT63xHCS
a7okszRtQITIMc0Li0RtRfn7h4p6d8pvUoymW+pd5s3LceUJNDjNe2qCMSsJBoRR
sw0roILNS6zIFr8SSD+j+QUQyGgoSDjC3vbIb184RQa5J6zvey30IL02OZAvHKTq
7VyWeOLw9VvH7VoBxQj73hA8Qp0GgoXCHMGdxlIngdOU5Ka9tkOahQcTdgpmpm79
I9U2oGmB/O83XAq79R4ys/Tv4oV8WeHGao2oCgqExiigCq5LQXgkX8rE5l93Cq/P
JwYqHFeLcslxSYkpJe5Rniu45y2vEaUdrDvCCOm9YvooYXw2ysdWRyuTZz+M3x3G
Hx7VG66H29h3dqnNrxMCER36N6N8E7AR52hehCgnSIoSbzvzqOjHyL+ggPCWqwvh
bZ/WUJOAB2X2/bBUxmNykjHNfZihySZdRhkqtNb076riXx6thJz9aaJIbu4VjP0Q
5KICzMiM9jjZQWTTIQGEold6CaoXa1eiNAtgZ3Ws7ICcyN6zeMrmAyHM+PoIIpgq
36Jr8HstG56lbGSjEldyQf/3r56cmkuBho2G0hYK6hkGtxUNeXWRU8htAloLJ2/n
utdePJAW59WGQWWLSlqtn5btWhC8yxfqfLYAcyy9sQf5Kms2Y36b3MaHj/A7SRLe
n12/oj3cLKpaVwTt0NBtVslLqpnEkz+YfWMvcCVe8+4zWWXxRq16vu1/MjhqFO3A
wZYPhwHH8mlnCXbQU0EcWYpCvm1wGoYAIW6DmImong8E32IBjRS9XFtKd+bo5cef
21/PB+PbbRaPfkmMF4dKHBqgBvt/OUJEaZkMrs9vA7RUOkdUDUWXoAN4bmu9dr9C
2uHEe/A6jPpfsPl1Kfvgt0/pF7ewgd88tw+jNPz4nn6Tz11E+19aP2xaJa66Xq/7
K0NUQorTFck5Q0XP5mui6eIOOvErClHTzd2Pdv4evqlkh4/81VcW1mpnRFArJN5C
WiIqFAxzdKEA2dEoJxgJLUVk+w2VD5tK0+gL6sdsWtR7IjF926bXUZj68BTcAV1N
Lgd826N1yhx8b/1/8f63g/FSqJ/zHGGTun9F431cTFI0zqYYBla4Zk6NhTupOCGS
p+PR9TVYj1nu+PelLEtfmLPMztW/7Q3mTHxKJ03HUShj5m6dU/kTqq4X38Eh00Ss
6AvCm8JVJxZ/ex9Nx/R6kjUQuCdks2OQ5bYiRCBpy5HYj/JmgTcdn8lpop+3J3dB
ZZE6RRxXMcjueU/10SmS1ntsYfdGPsCCnJSehZwxQnfBj1hGxuKLl2YYAXQRs5bk
imz/i/wpOeB/zisytZYijmxBvaNUDmgRyyhu0GjJwShc0srO/9njkh9Oszo6WC8I
/xDSbhTjvyRc/LgLSrwPA8aqukQ9iTAf8rGsiSTLLdzoA53+qQrxDJIKOVej80nX
Ay2NX7kYYqakC29ThakKhNJKFQLyMHIOqD9c4rB3UKIbl1YUnlD84J4u6H05dRdp
u0pYUUVL81GWCfmwveoDt3K1616YOgdaGxlUDXU3t7/3PQzHlEmK6OQ7JSw0ph8K
wax3QiIIDWqs2k1S96ZfUYW/vCCDmLSX85Ct8qCuORJG9Y23NMBXBid+wXZKyrfW
tQ9HSgz6wSXq/JuCbjTKZk8HcUWcv5dJODehh/jECm6WJAGCJKjWxotv9VhBFeQR
YL+VDLwfyGVrkLnFZzKc5aOz5baQftGbJmDfd2+2MyAC0EaOkOZPhrfLFSXVKwW3
/hMEOe3btr0Q3wkM3iEQUGnsFzqEDS1DcF2+DMXRaYe1C1IO1GROHyeNX1rkjV+a
ztSKQ7rv/+wtQYSiAtLXzjcgBysG6ZFq0B2ld9PNTabrzLtRG5D0o+KuoNSFiLfV
g1j0qQXY0EJYc3KJbEsxJcbCWAFcjRd5LWsGjbAI5Wkl1Bv9My4FwJJ1RkwTPrk9
ZDHBsnFngEgR5aYi4Zc6thgqZ3Z2m+oio0FZr+2RBvJh1qGrJGDJ494l5/a2CucQ
H1eKztWENCzLGq0XqaKYQ7hp9DGH6hHm+0yaOzn7tSKyRHNmYDBk/FD8qJyPt9YE
5z3D2USEzHYCBBDpzmUPFVRrz/VnR8bjVBSJy1xrnr+rXfWTDdPca8bocKPG5M1/
pvtZm01jypIFDT2cDnj8PmEIZFfaUKL5iUbxGpK1fV4a3Egmz2+OWIoHEclfpMuj
RBM+ZYEYF9l7JfAG9AxHPfg5zYU3K9KbixQ70SBSjc40Oy+1hXiD2rPZpJupgiNz
7gijug0D88l7oCz52j05FkkFyTogJvMJoopIuwRTqo8noPJ7DxP1QTgU1qrQn63T
H3uP1Dxa6igt+Tjv5v1w3SU5UC56ndKZIfvYp2oCmCQo5xTeyMd1xa1riUneFBn1
+B5RQsO4BIStItfkFsIqgsvN38bfse07nG1otXJoGCHDZmxt5xpqbASL7HhXDJdL
03Ixk56D6ZY1OVQMMto1B8z6SjbLQ8Ntm9YpOf15UgXVRv2vB6sQJBMqpAP3O2Pc
2wchfxc2yTkWT7YMycTOHO3jsTetefW1kEtKcXT7u8R7/EuAjVGygWnyD47fiDnb
LDxcwXTqtRgMx+aIP3pEEVrv1yPOd1kRcjzLtSyv0FH12o+BhDh8vpiwtAqBO+9g
gToFITIRtNfmhLR5abJ4wGnYNL7SGD6y5UuQfBArEynRqXP8qhF6MAmf6G7E3v64
LaqCr/eWcJYDqJvmcttfRLc2fazJv59IdscpQ2N+JJ1WjmxeSpZggkW1uka6VNY2
hRejZgJiJ7H+46MHbNekCGYtNide/qQFv6ws11hoelcQt9OXArtCrik8myCWSkmE
dGYBa4ECmMzQyPmqmCI8LOdfoqsFEtuA8u95KPbgSQutichIpHbKbdNDrPo5TUHb
JePzQvsA+bqEN8hqD6Dx94OkbfmPDhN3Q7qE5DPOav4pBpKO4cp7H/XdgxFktOaB
xhQYqyEytZqir49xwuEEI/u8zyk4hPKo4zh7DXN7ywllTuaRI6GuiSCyIo3OZKmL
t8dqLCjMai1o3T0vR+74Q3x+zs4MLivr6MbKQuBYWOwvnFzx/ewd+Cg1UKQpZjxw
EQ6EARi0nwYUIXmjWLo5S9XADo0GdVXIx375Y5UP/uGl9u5yEGYgTaVdc0ggBJb/
/mnH+yUJRAt8h6UYxP1kfpn9pwJUhlwG+tOXEVO0gbkgD8+wZORCp6o6wGDYCHQ9
Ntp84GJCDGQO12HZ6Bp2JzayAV268d5h4SnWIqOiZw6pTGnT7cmkUXgI/ZItNdUa
O7NjA36+JsyCxdPmdPDNm1k43ksKnhL57EeEBJHSSOanKHKHU1goYdqd2leNN1ZQ
lA67M+rwnlNYlwMEh7VSaxFj8yAF/dohJdgvTVKyst6yTP3Wlt4KBG8+rfANVMgP
0LMVY5EWizLkZxK0idteETYRIeRRrqJOszDeZTx+xnvt5S/3gmMeVKHYZ0plrEsv
FYUuqEwOtCHsU4BtHnoQblkY5+6aV7u8RqHp5RnhSQQ/7OC086RJ4duRVw3XeNge
iaODfi3U4ypQXTPlnX5Agwm1jUxQRGU1+kEkkVs7r57v7GMDFwubtXCy1JiNLylE
RTjfR+SjzSXBnJbnhCuhNk0i1rxDsx5pvYujwi0X52I1/9q2b5mFMrBdiZ9agqdB
UswYRc8k6QsWrWYEUrJ/voF7FCbBd2ZrsKzI++SpCNGlfHLnPh+xsN1aDc9LOY4Z
O6iJdCAdotclfQrgWKIZIKR2ggGN2bEXPJifu//0Tnoe9KAvQNY52wLLA3ddoQtY
Xpq/I5r9ioPJWgsHmo0rmBR6eGfFxcIwUHsEnBtyq4whIVO6RaSoxd0a4mzwwMQT
aX6x4XTM81xarr/1jHiEM63dME1+SlPMg9geMOcw8DGZaSDCEvXy2YVHTbJDUnV8
AqgJQFpMSB858mJByiANQcyoAdX+b5HqUSmzQ5tfSMGVX7DKGF0qM3S4EH0TWDwb
DH2fGaylfNMhIlRSLB9tr/3lmBZ3NVnASd3Yh83hBfmSeWBQQDWKCiw7OOAq8gyN
FusArCWxRzX9AvEL4EgEDPGl3fNFVMny1NJsnc96SEDev1dISzbo/b9UxIfXUP/D
HTpxjB7URTdDUOnfZkBTw696i0IjSAMXR2+vCRjcntBA47xWwRBrFwjvZAi+PrP4
fMu2p8jRObdd6dPgpwzvNIwLrEHZFnfebrznpAtoR8m86qEbbMaIo9XiyQCqIXx9
Q7DcTvg6aH9GbKn1P7a+VWsGza4xCrM1QG+GoG7BeU8MLky2eI0wN9XwBYqjGpyR
xVL9/w08yP4AFQga84siGIVEvknmlhugeXRgGBaU+6p+Nboa7yzZ/aMcMlvfRdre
yO/2xhpZfxOiS7lcXv09IGwkBmaI7N6Is3gZq6evqnVJYnSa+O4Hf8xZeOLBa0Y3
2wpLRpo0/fXiF8LT3AIm/lCxx6RdzZpICzwi8acnMAgsuslh3QK0ffXD5Ns2vzKJ
/qIouKjE8NOTTVln//ic6IFJ25DHlx8QLDxT/TgtjYC4vrFljD8cB+zEhBtSmbUZ
GiNUaxTKIvXIHhPLxHBHSKmKfKTFNqmuiN/X9v0uhLCCoO+Lre61mUk1+QVQ+NUg
I6SYJGzQocqcM8S1BMdKdyn86IGb/i+ClNFlkV86wDQnD6JE0CXpISie6jIw08wU
vnBRHxFUWAJY7zGadVqYHDEPKeoqo0SxrvUgSOA7X7wjmkxG1I0QbEdTueW8NAeq
DZmtcgca4l3kmxRrueziwwIOV7nH1GxiCFeX1pEZmxl9lMbmn1E5ngNu7TrumzMg
hvem7LaNF4fox9bcaYqj/Ic65kVWVduUuE3Pj7nDvKYHXN1IfXXtyoLcJr256Niw
KdudlJBHqbEyiYlyK3cbDlkOMwC5ga2vt8qbUQbYCRVeM7b9/pjPF82HITQgT54r
rJNqFQRbQcesuGfQAZ9f8T+EyEp0dXFkLFfdku0CRRMlVGDlf3KvqTM0BtfCf1bq
jsq8z0pVIdvCY4a4nt0apJut9e0hyuz6CqbbBqOBWdsuUR+Xj66ld+wYAxp9c4bp
kriOXBv2l9gptDAwpvmusTWDtm6v4+SCm6XCOc+tLLuf6M+njrSAXn3r1b9V8RmJ
yTQu9QHSBv8uG+lIc4jsqQYpEs3aCX3wkJfjUwXDDeFp+Y9+6o8YH24PHj7bZwmd
rr8DCTqwYQfSb/IpMkrsli9RNWEe5hkndolqR8NAjepPr0WV0kAkmvUSdsAU4Rp2
7tV0VTke8Q+awZ6HpvWJKYy16QSZ9mBHopkk4W72U9iGglFf4QHcaF2PK2Y4t9sx
DXY7ukrmD2MH7OpAYFv8PNWemWUWFKJ2zKoRN0idSc1kxxOxYFe+KE/vasskEux9
Em/oWcEnFPpz1NaPpzKa9azDCU2hyZ594FV3qlTbIOmxhKfh+gKgwjqkhhKAnejo
PyXkg2hznaejNQhlHK43sIfoAGvGmJNX27f1JHG5K7TvaAC3ZzFMjeRHcBIWhTI4
Dy1zte+Qm5zSsmnlmIqj0JM+ARTQSMDKaVBuntxMtzDo0ajPOA5MKwQv5ao3r4GY
X3bZYT7zkHtYG/cXnSzCYQWvJWorrTfQMRocbSb+Vk0l4eRbHyMgdbmT64DdRfeE
Rf1yRCjCmhRhbnWjA5hPUzMint80sMCMO745t29BUHdN8LlOglyeRv66xHUOBhYo
fyMUNNp+4j6cfyM+ylNDoVQeJg1koisR19DrzAAiS6WAXD+TKfEg/Z/hQDVSt+kQ
cEp1hRU/Quy77j0xv85QD+qW51rbyRfz7VZozeDfYBOgxAuaWl8Q8yoorRgsOAsI
NGAOBhjAHCgqTlPvhvjdq5dDPE5vP7AU+fftchydiynGEMsBNC9hw0+3X1PNhT/f
3bpWsazLnldgYo7pXG7hnGO9FsQHmNwpJBFOklfWAf/lhXA2mYP7h7KrCnJ4SLrX
2y6elZg38lzS5hJHIU7imJMbBUn2kiYEL1PKy6+iHE+wu6j9DP7Eo7qORnxK2New
2VzRHg3s1J902xH3TYFpQ81nG5w9R2HoBw/tBTBJ7rkNKFGcGTFufYdxt6Io5m46
WpZpzQR7bgUZW31Mqg+XtjG1Rtk+FRIyxP0uPSYd+TGE/g4sYxNoB/FuXWgN7GHr
BUKO9yku5sH4In9HiEChfW33zI1XCU9wFDtBEb+62ZXPXeEXme6rYqECthe4E6gt
eBQk05JEatq/JWAjcosi0epTDed6QjZ6/0Rf07xqPsLwBwgUHAI4H2M4nLdskMzB
uZWEUsnuHygMoAPoGjdFp0RR3I7BgsHbPI2bhX2CHZmekpRuUuz9/uAaZUOb5n1M
ReIn0+VVy4TEHtQ98QGLRndO1f7w+1bHYc6bJXSdhK7RSXpNFrMk/WgXN+9NCs18
5HORHMiZ5UwRFEFIxn7vvs03DObcySg198XgniFC4YveMDVDwWFQywz84AMsa1dU
rALqgJ2t8R/nQJwI82kxtDckQ4Zn+0XeVUOBSnjfZtjiz0oMGkDAd+JNN/mp7oGm
w2KAxNA54VAQKY8BBpIatyL3huOHfW14JLjLMy1HRBfXgJspYNEwE+ECo85zbu0S
DeBUXEiwD5SHuCWF0tApBMtO+xK18t/LAoNQpFjjUTkOtg04gveGZ1OJv/nU1a/E
wrEVNbHE4NE2k9ForNSrXIdQchhIS02X7MhWIz9JTgYPJRuhs5DdVllkeHt0lpR6
NNuO4CCkkIirgjnC1uSB6NzTVFuWNSu2e/AgMkBR9+Y5ugt5zJwSakd1iD9bXdpK
GewvgSPlHW4/2T4LD6lffwtLbPZHOuVil2B3HDYNeEjaalc4MYAZrWxn4qIm4M3p
91bm6s+kQfJQX5AQvGhX8oi6+H/3bWgMLsw3IXvMksGhJvNmSmVgyD/pg47+cd/J
Mg+5wh+a86vQx7cwqTehS0V2TTw9xXy0rvOkYdjIFCljkDq91cojLmQku+Iw0Lz4
AW4UUic1t+15lWn/j+3uhnRYEio2Xizy2Jq+EKpjVb5et/qRKplhy2tazXhP6bIe
eB/TY1FIgfl64/r678+L1e+hRsctZ1VxAgnn8R5C3BxBuhOl7r9BNtA5elIyQLhS
5QmDbHgabzF1hyzZ4vOAd0khLW9Gz+hcKY0Ss2U6Mkhxrj4cTR5T2dLrw5kzjuOS
h33cWPg9uMEwqkVw9mcP96EMBrux3S1QLOtUzUdVekkjqFl3uZjkXSYxnMpAJd17
i+dOH15UarMJxCU9lDT4T2hKNWVbVeTa5pz0yCKDXMOrJcA6TvLz8fCIUI0f23mB
S7wOWK12BY/OVsA+EbmWtwAkSFw1eY8om5mYeuuM9t3IrOmgRvlJ6KIC949NczMQ
SYSHR2MFV/r0jokInAUKk7lIGfY+4S1D3zhvnxkbQDgNNI6YR4MSU9z5p3CFKy+/
zDWTOHwMKxnVqJowlueSJdz/i1OhVbVm+QCUuESyO4p43a4GRR3DAos92YXs63gN
C4FOLfgqA0x5DtNoOOfnpHnEudEedbvgyaqnmMMSy2wPv0+s/im2G8fkZYewnBI4
6kikj7vnDhKvq5ETfpw8eRcznMgzPT2AzpvBWqUf5B08u6aMojQA7hfJB6h7xQq1
1qDfUbhUgPtxsBksvtFfLhR1sQsh1oFneaZYHm5zaEOjQJZUdQMhT+pkFbcWz00W
b7jqcOa2hPZztCoOZLX7BcUEhlUPbz6k3/fst5qy+tTuvOJAGNMISOhmB3xJob73
QS7l4k11x6e18RRQvXvTmqLoTeCED4j2uIuhv8iAo9eex52Scwi4GYWUQBUs15tI
t4NU4H+sHFSPd7ETIjAxcPNIEkYMiO74nwNKm2/PscWlx7oeQ7TInOrf9ZpiXa13
5ZFQcvx7V61RhQ4QQXwmgp22/bhZnFB08RqHhKNRw4GyXNF7PBk+brStiJ5fr26G
GpA+AUNl9yv4pvdfDoYEKS4b42jaoMqMOTdsQ0oze9P6oc4j3KANIXfUMF4qW4Uc
jEKW0SxeZkM5iED2tqWjqyulkyqFYBx76YfGG0Kaq7TYbP5u8v4XxBSwEdz/0Ykw
/7Baka5/AYUnb5OpDce9nVYfqrt+ihxQAROfrk16NSKFTbgPuxCnmsGp4NpFW7gs
YbZ3S4jEVi052DN6X0Pn7NCFnZsKowYEWDQFYXZ7qtf2ubWUzOzlZd7jv4qBbjeD
O+C3t1Yvmfhu0a+VV+RW3mNFWZk8w0LT5oqS/hO4+d7JeEwztyZCkxQ4FQjK95eB
8nLmEl8uFpWKZI5GaS0FXrNIugy3q1r5bqi2xrCyxOTr7Rwee1RA8OJ5t9D3DG14
vLUPqN+KIoq5K+0cNQnIhagYTOZFQl5UQA029FoU63DuJYCy9aYrcfzXUgmbpbwV
WzsDGOprQ/FbTzLEfp0twAE4qzq/pDTtuyS8UCQDTy61lh/ZuLfAOpZ5s2FuRmyy
AelToNt6J6YLHA1D7UEqk6wjstAK4S8L7HlKx9ZKCCuMZlSLrAXiIKA5DWjyl67S
Yk3dbw1VNBiFVrau6dOPiRgdTAmhBGj2ZXcpnr5F+Grv3YgW+zRsonXW7zz6rqe7
NDoBnpRgtURh6HVy+5NIflGXlZWoqhc19zNsk6scnqN/Fav2ObJRJjob9JmE3yKr
EoEtMhux7G4rKDrDLcnq9Vl5G667V7q93nFE60yt3EYpW3xgAH5mokBTOYzfKg87
sBv16DyKQf6Ig09SDSXaavVulfQRtR9adPYWF28TVlqjwFRScxJYjxmGeobDfLwY
uQJFeu3kt8VD4tmmD2ra65tIt3GzmowtlIAoo5YhFZj/6C5OY4S2JlQlYvcbqGMN
TDE9qlTReVapGBsbpryxj149iya5toVsziG7zRiSWJWNYt3YME8cuJSbK9DM1RY+
Onw3TUosk2k8SK4lcG+OjOvCHavoSba0LcBgSVvpoqLCKLoji4RIqDERVRzc0loR
a1X6KvUqvYf3ysOgnM9TKslMQ2RwxDO6cm4nmkPncVyqGuuHJjgmap5SxkplC9vk
gzqPEYLdTmybi9gMYC0wYRUg32l0NS94GYHJ9PDcmNwoLUVHl+yiZ60HjrSqfiQq
1hjBloSHZ9cjIzYZqlS6gkjgE2pTnSbUh4W4+b3Zr0ZHloXr1unxHUl4dt/NOP7S
aDwrv+s6rwnvZ+et3WidgGb0PSxOGJCYvMZhObQrcdwZa0DUetUrJqs0BTHf6nLX
9SSIYG6mYxa7FHD5xsr8yqTONXJsXd45AqmkXoYnjgYk9vvdjCRRIGHs84KQNX5Q
BsQs0YRhodSFGIm2cBA570WtMFmVOR2F39prpI3c2C2y+VEP4kUUn7D3EwxNM7qv
qO+Jp0VVWHFwhC74ge5YXnsX25OEOwEwRAEcnitVrCP+kTTDGN5fTrmd7nf+4r1K
vBoQrbXZYKoxiRnFSSX9eTsB3tc+nviCj8bVKGrsKQqsesKbMvxj9/V+E1MJAcJi
1E3MXU3oK+vdzp69rzti/upl0MdQzGP3pw4xHjFybFkItYqftkHft/v6x8z+QtIw
H2P5uqu+Gf7/hLjhG23ehkEGSkAGsrwxp7liczT8vPnxZHVlYRXtdg1/lQpAtgkE
CoNuxL/gSzQROVpmawSZb/6NGJ6Zi4MJEotNQZVTarLn6dCEmLtm2v2Dw7RZ7RY7
d9MVnUQBDapUy/jpe+wslX22o1thW747SkDigbGByaViEHxlgdRj+2mAg/mBaxav
TgbGxJ9VD3iqbjxUlZvYk678z2XK26GDIBBWK93QjpOolIefAIeeJYCgvih58OkR
FUSOKwmhJlfOfOLdfoNi53JpDvpyTzKfN/+aRfQoM1V+ITpU5YCnzKRxBifphu9s
+9XF/cDlET3vo+AV4hPGnDIyLZ5x3inNvPy2UNHx0GCp8lFt4pzCpHQX87PmzbVc
huZPTr0I8og1b7TFIF3Tis9aI3VLDZ2x0GpiX3RACe7O/3GgUPsR0gQzD7lRKEkv
8Vl0HDsKXRXj4td5cJiI6aapOOSmzT+TpLfsh2PakjTsMzmouM4bdbO5V1xSvFlz
qQ/ZbiwKd7GcMXwvL89YWsKocVHFKvTVIAy3UFflFfj9hl3s5l06D352TXNOOIhy
9CpCEL8G+NPIhA/4u5ndPAVjPuGUwOed4kbcPOzFrWuFYA//fOAl+IIGPPJ3fdcB
Toq/CRoXtIkJkorTKSds3LxroC/u0eUCGUu7/uJ67NRXSigvPVuhxruTdavzhdJn
lrSzWXQjRptTfAgFm4GGUFRWpFXH05YMtSiNuznM0JrqVYnRDn183jLFi6MWgZcp
2Wdhx5bYAj3pvK1UAiUYzAIRi3Mc7NF3UXUQtXcgLlmR0AtJyQw3SCHdW0VHZjxE
yENo4LQiPsxbKKundxUCeSudv+DgpYn//NFaWYWmcbczJYTrwRGAfRL8/8CMXb1c
+L+21xbmH0FOxlAzoDUaNNxfun/eQ+1Zc6ZeE9d6hCYN0FTd4948gLUjJwfumq2R
01Vwd8bjTqxZI9IZ3a2mi3OPaL3n0Fw/6QNPSPor4yrRpSpyCVjpkWNIBUwx/hlb
y84fU0jhYlxIb5Vy/iX24bdbl/FX88w7ITqZMIV/S7miPbZVnYEJWJrMUNd40mPI
kDyjRydPnDewn58au+jefS3QqSR7oZBM+SzV6KHgXBtpW58B8XT7FXXzeXTQGJ1E
RE087mcXiIXKYfndkfm6haSPfMB+oRHTv/zIuyYizBKZjUij91wS5kzccQLIeLig
7qLwi2TWlLcH36IcEnRwfNJcVWn57UB7854uc44+AM3T5XDiOuGJWlN8WpULJl32
WR1vDo6j5Tx+MaF4x9BSjOIUarqWDVcam+GevaYlJ2C+BNs/pLbzHjRqEK5Yx5M+
oIirmAIJ9L+uqX9ews7pmZdNtfBHkRpqALEqn3bAVKXW2qCt0sFGnC7EjSUFw9zC
II3gBIYNMBcKEGAggwaW76Oz3Dwg336sp+FvnGqqoBiQdII/a1vwT+w+Xt28N/Cl
AQAsPUFZ4PP/kH12egoiW4nqXzw5QsyR+Tiu1/lJ1Eb634WslLSeNeceBt4yVqMc
miKufpa6ID7kUy5nc6OD3JB181cCD/UdX6DFbqL4CYrZgsHHyBHdXSzMwMhbyzzq
sqqHrcbySNKmNUVL5JfUqQiZj6aUN9GnerJsGPOApg2jOrzhcQYjrJQWssmHn+9D
3fjwEMQqeS87mOk0wh9LG6XD0E5DLOPv4mxioDx8KJwSPXD1cZrwUltRQXK7lYrb
vPQJhLA2szH2VNYHfqjXWHCMSPlrGRiXoEdtXITUqswZzoQ0t/gVXJ3449sFwM3z
kG95jvCVfItVR9yU8aVE8m5CtnDw/C/xli/Eltum0IYxWCu0PeUfq4fuwa/RQG2X
b0LLzt/3MyZzzAUjKf6NIMIUx1G2MCoLp+uajvnn/gskEuYWXzFhVNx0wywVNm8A
Ze9jPI3Uh3wkBh6935OzLIZUt8HABmjFzJXL3HWPV8S/+zTfFBqNQJAZe8MBDFh8
qjBqiHbCvws1WnBaWSdTrmrmS7wFwH4eHa9Ms33U8ehRaKHVlin8wVcoZfFtpeud
9jSch7xec+SnBqIJbk6Bk+hC0lqi2bQqBxGD3nOTM6/LUAbVSBhjGsldVizijPJW
vs3eKuQXoGVb6ICDEcangKYXW9plOvE3Paja6/zpi0fRaJBSxSp5qYLgUWeB+y6G
o7l0YjWxo/VIODm9c8GRwdvKWWywBPXC4+IzEK6CiW2IZ7jHuIqXWugqyak7YzhM
dl6EdEJqTC8EcDuRVAWU3YZR9Wv0V+zsH3pd9yTzpOWAWOBtlW0R81f0wH/4r+Xk
a61hwHUL6f2/j2AX61bko9KHYG3FHodqudZIf8eZtCZa9kas2H7Ysl/APz1nNolS
1jYUAMR4Rs9MkmmGFcLCpbVnzQJKO3tUvPA0Tuh8V+NiO14FZwTo1VGo0+ZKKSHb
TD+nEnLRP7UGx8xYVUxoJIdb0YsfuygUCyM+/2XYEroq4no4plUXB5ddUshokXn1
we0x4FRuzCxvJSynuSjCXNOX1/OedomG0EXdhNLZZvXYQfaevPUxaIe9KNar04W0
7r3mUsRNWcmY3APYQSSMRUtU+XoqP9loU5ZALHsLXYWzcDYUnC+nuv1rK21ORi8R
B4UTb5CtLQ2dNwkXozVsJYA6ikMg/6J5zr4sCOZpN376yDeNZy3UzmTKTO+hXhbG
MHdYjsfl3hY2qiYh8kfnIw2+vXUgB/1HFfjfnWKDLIcnwAR/Ggsf/Y9Md4H5Wvlb
hWF+xMJfabOWSs0CuEbton/Ip7RBUf0HnkNXvIJjMZKVvNGIkAOx2/6+FaWEF8pd
OpSU9avt14QPHTCq4SYz1W7XG6GxRJ41F+FUvvPe1GoCMe+eEEGtLEaGasuic/3F
0Or5zRGGlh7o/SAftXddVip2C6XE8LDFOaITpozX/uCbj3tyFmX6lvQdaXBoDw4s
hrZJtAt8G+itMZeWt+sUCB7542aJF9eR0Bs31aV/YIstJYnEZddjzeAUgeEuIVur
tprquvVt1+NsqpTSziA0sX28jP2Dx91YKpHIFvXhf+7cnm3ZyU80CTtlXzAY7OR6
y9mkGYnDTnCxMztGYqPoafTubxN/k1mIXfwkVFRBCaIeUgKJYOL7CKkATbLdZgiW
QbbK4pyEQDjnzumsAqCMSRB5U8XcgyWuN47nDmQZem599OmCFL/FH4x6ZiRTW9+u
xCVjZ5vPehDOv2vMW45TLVvU3XPg8oDLmdyAr4IG6DQvVYGj4qNVe8DyerUilxE0
vDnZHLp4PqzuZMVopHC9nNa1AdiLiik6lTQUexduEfolgaVEkAVYxvXAlaOkPAWd
6pW8tpb785tZIdNJ9ZtmAu/dblTWkyN84A/9V95NlWZzIClTumxdk9K90HmWKLUA
ge7/66w8o2O3Wv86nzgB90jtlZn0neuiZ+P1TzPHAo0RshzdCPzFl/YbiUJv/+on
6CkOUMa9OkCAZNheeHKxSS2FiXoTlOzwcFMD4HNle9DHVfaax5E7r84UoIx6tOA8
6DTRmICVTjbitQMx3WJnZrnA1oUF//lyoweMzwHMKLt6REb+eb+WLlKJlpeDEc4u
2WJLFy3cYBjphgXprfMLPFfCcgDLbz0fGpXAbgHe8bFhWyrHHTRkh3oblBFdHvzK
+sejFthjh5Ymqd1vMQSY+61XocnEWGr1XPmjNDuLGvtsJ4YpYW5ynPck+8rFZeff
/IYpwO+S794CgEBhr/Ct/C6bWHe+i31CETw1rfcXv597QpORBtv9IorpMqNi86Mk
SYhZfkBnQ6fOjQynkBzqs9PXPcC+QAJSosm9zGPbB/UBYJYe1GWJTqQ9uGqc2NEr
NYY+BY5u/tzXt4rLuF2IQ0N/pf/mIFep/SGJk9j3dKkSULiNNu9ofBXznfaCpyPZ
u6dSQe67xJy1noOgqXWnQw2vlaAH15xa4HL/vu/I9iWztphuM0kHx4n2O1JxWCtr
ylgZDBLvhb+9IArrNn0h16lnV4M5ekw2K/WNnGx6asjj/25D+fMLISk5HqEOWRST
ogT9QVxwxv5uM802fKzKA1VSU1BAYWhLoSgf8yPNy25fED657kAdhtADkNXu7Gb+
CyJOt89fdFnbv/QVIrerZdzhE88rKt9pNlVmImx3n/V3X+O0+W9zW62mih31iKWv
Ohk4egEmBBRQSJGJ9YRlRw4j74g5iJfa/LkoETBEMoDsd6u5FiY0VDZQqKmq67JW
6Vkj225Tij05Djw6WozQboWSU5SUwKoQPIUcr/yUfS9c7c3rHRoNrXSjr5751glK
9REDCtEovEVUy2qRAaUTrCWJJ7BzfuuMQQMyL/5+NIGsjuiw8vZZfz6+TRzPqTyl
uV4tsxLcZafqQMUq/nw8cstd+mMTCVihWVNmxh1LfDDsifQx2XXRHTlKfR1KoE03
mAb5pBHsBK/18psHbGpXxxkaHjvN7FxyKgKS3LdtWS1iq04IjXkRwjVbQRFuvcjD
NCDpoUbq/ImyB6HoY+zXufXeQByUUVScNMiCiYfTt5mU9ukzQyLJqTODEUJ/vMBZ
Cxl4T/tEedPBq5QLo5kZgrn8AEI/11m+2t+vjWN2K53VmwYhcNhZ5cOliNnOre4g
fvbXcnY2DJb26erqL4Yvc0xdGUomDzr73HjD+HGJoLO/UdQQTUbUc0brhUkyBeBZ
L3UYzQ6u0FsdZV+9tBS8vGuIWnvw1XmDibrYP0GPZDtYZsf2B1GXaqvoIIh05GKf
MAkbeWqALbfoTPvH17o10+//vfzYlMrge/sDcKN1qrpX7BKN/1KLwNJkf9n0xR+O
iUcZyg4JXI1CFG4MvIy2+MPRj9onK/Iq04Uo/VGVBkGpsnX3suq3cdAlRnMDs9s+
hqhXFTb566Y3MR3cm0EmGd728ex5t4qu3XhN2NovdlyGbqXr5DtcJ2Vd/KBsYduV
ajM2Qu16X5JXknKr40zoRgsU8+o0U/rEiBAK/rpAFfQDNvoESapHUe9k1slQSWs/
b3DBtaWP/h3tYQg3RiPi53a018mJXnIuhnXvTHZD7LB2dVXiZqhmPTB1Uvt+E4bL
hE+EcaKTIPyhaeBQApGx0DSlbyTMoxdglBFI6SA6SNQO3OV/n4PRQXyPz1D/UT/1
YL+n8g9pOZdEamCUgU2HuZW2rOoqYM1S//vgWpNtfeaI3907PWwcKgfvKFWI375B
ZjncxcXjniziS4Z+MHktGdJmoDAs1/YfeQ3CEqcJ+Li3f3eZr6hSwC93m5E3CQsB
dzttLiIIZAa9m1G0Fl9ixy0Xg2Ekr4jOG0jV8H0zVdc+5GwQYH9YkfusrknU8z98
0yLIHNBtOwyzfn2AtUWYfXrRHGl9cO+VJsqhWGw9X1dhKxicyhenKBFeCsz8aW/p
I0TdOdHctgaHZATXG9BIwHBFjc4L0CQwtxK2M+1WmN9CqWePTFlWG3qbRM2evmT1
N7MXqh3lOqgJA8Sapal+pdwxeLRMJzw8PM9Zy4iCP3LHNE0xnPnwXseRvAkpVKjk
68E20RFrWdF/OgIpAgl5DzxTUmFNEoD+kmknyyud++1Wl7sbuf4Pnb1etTXkDrSp
tG8mxP2UtlSmdD+npCm7+SP4fQ/myp71mpTysPtUMhgNuKNwmnqAgKEHU2rKNkqM
//cPnFsrFRQgVF/lyPnMIXBJmF030lpGv1nfBmMAfVu+kqzxi/d6Ev6kiSbeunFi
7zTUoqozfp2TU0wtRkmSdR3N0r5rngDDX1HufJ+5k6fHdEaiHPtT7Nt48dE2ZZ88
DVw9yMZWxT+NqnkuYjoRdbmhx3FrEEpo6wl2Jf/uQM4n7TOKI+624ZTZ9nII6D5M
wulorB/JoGZ6znZscfH4/V3SrC5LOnRPU/GifQDmL5Bt4mEx+dGuNqmM51KTjowS
3g7IeePbDd8LjmeTOHp93fZQ64uvwHZKUvcy/ygn9kiPTkiO/TUYf5XnDZZ+2dA9
5SDH8DVTDtVI3lrlSxfONN+v2XhAS9UbEjRHLc9Vb2pY5GIg5wh7VtmwOkNNHVeW
qLDgQX8G015dfX3aiqH9tw6M4dqUPkoBzGAlqTu6HmdLlyjsE4ffuT+pbGcB3pDP
s6vAQin7QEZU0U/9v2alICIhrIprAElIlvUOHYPWDYV+MgdaT/K+oY0NFgGFHOXH
I9gjapGaDxLqhXyHZJhv8v4Jl1KZJoVQeCD19Ee791EI1Hx6IN5AckxzZerITQRV
CiXn83QQptMLMyq04ewRG7LLE7GN3UGrn242T3n+80y7jf/1wmhE1CMVObeFEBlC
InGEqrY4H5DJoumTm2msanueI1wTWnDn7az229Nm5ybF8fwF3hzIUVOBmkZDNW49
QFtcRlWkMfCuNkSz0OqzgnI/G13h71A3yhuwkrMQSRvX2yErZ93bfjIUt3grosW5
X8eLE8fO1aKC4T8Dg/gfPmZ2MjsmU3s7JU4Wnwyy89p6Fw0yd561kWLPnJnhpfsG
IJeTU+Fue4yPmwsZe26mepvXf/X+B06/o7v+zbLvjNc+k2/E2JFBPJUBerRI8AnO
N563PGBsk9i6cp9QMV8a1R0io3DPXqWOiVS5ZYOcMwvlz8MdY8KZm/gGDJgvS9Br
LAK6TmDiMLTFlLl3XKzPY2YKHemAa5r4f0ohcTYk8JxCxh+rR4VmlfGgBwt3Q/3t
RPPKeiCuswGCWKWqwp1Ja7C61s3pF7NC7tZDqulKhR/nF8YramkT3XgJYgQ57PUZ
9RsH1mmClf90XO8qrGqwy6xBUtayZr4rqoX721MDWQI1CqURWGpdmxvbQIoR6A9H
yFrjFbRijKVtn4+gmd6vRu+7ih38Qp1cEO9QEGJvzqtWV26fc4CyHlIWu107Bx9l
J+aWDOpXQoVL1S1huooaHNSE1+pX4GEXjQohycfXXdDM5WmO9O9j9Qc+r7n9BKAh
EhpGWSilprdwcIOhopW1iIQUFnBYpC4d1xNn6PjRzZUWmC5zua91oQgn8PV+N3Ow
4fz03lmeNlHNZh0iV+QHLwF98SpMFq1SmKiQHUlQapuOqg9wPhiw01ncZR4YSpXT
fOplxqoepnfap5GuFRTVjEL5VooDSmtAukaw5maPOGcl2hxTdwu2Hs/qbnknc6uN
YtXHa1kQV/hac3xE+WoUFs8JShTQhJOZzIiB2oXn9LImb3XN8QhNAUy+V4FDytwQ
4oApA5+jII342AKyFUT38JnsEZKi23LBIchQYpzyavSVJqonFP4WPx6WIh4JrTVp
6I6rGSGnX0levec64qEPiErItACkAKI8RnsA1gPyY44U48poIdVtt5zojhszkazl
zNlFY6CVA569xd/tjhGu15OIBm5x4askUVbqZhah9oH6x1FiV8LvqOeRuKyUwLgQ
O9cBvWTg3QpfC0zgP+SWik3qCGKdTCm3poY4RK3JUO2wJehC251BU+/IlI+OWQoZ
7hwxf7l/AitkfDdwzPnAaBZcU82Zcsj15U+GoLo1KDBX5ar2PBORQT/uhrryRw7g
ZwV9Rx3TP+RpHCSl0TS1YsmxFOo9vri8kpVmmCobHo5FJ0DnhXtj2A3nCsZPP+Xd
qaujwF0ozIU/RP8xZALNMt7Ejy8icmrZlTCYgvjTRFQ5rurYzfrsg2ZYQAxfqZpl
5N3TZAfPg/oePiPVSQI2cYwgBBi3MTa8E+VgePRU+Tv+k1Qi6zQml8W9KkAWrZqa
ULyMHUxjXOxsaXvJTGUobRzl5n66UNoNItGg+aNotDSGWy4Wiq9QnxLzDdsTYrOD
T3KTzwtrHex36b5KD6qEtl82fxqLLSbIiuCcFxXbQjAVKUYjE0xsRy+RnnfGTuXB
N+BDnf2rQRs6qP045rnwWaeQh7eZv16fr/b6BYmQqkyf8CCCLGsfqMDQ6n83YJ5W
sGw7rxqNGSVzpcJGYn3ACz3N5c4B1SlcTl1TMQ7ntygDWohp01lvaSm23AB0FI2Z
785vLT+jyjS8AfSzm12hxCTMajOX8F55YVKTkaLg2EM9h8HkdWBtWjH4t8dC+bAF
A3KnW+yxQwEjeV71gIr/yUWxt6oiH3onAchjLRjtYSickYCPGYsbr5Cfj8HVeCtf
red6iDS17EBUYBavUsOfaG/NrzocfzFegtZbl807GJxonad3HBsM4cQGQYq4qA+4
KTHyHjF07P4I5anJtD3NrURFP/+8YhcKQFU+5uoJMiQF5u040MR5CQFv+p1KyIRh
EJkOWtG0bLcj3oDSod9oUroJb105bj3rNFIix7anx+M8htZa1AXJxzy5ZUCZxBf1
hQah5tk1W//nyYtCfDB8Js5z1/GeOFh+pTU+zuIFlMOjduyvhkkCYnmK3gZo9uYk
yhS7CeUZ58hYo/zjVpiNRcXmb9kjNFkuH6tm25sbX6gtM3mnAzpipLjuQLJMB2DI
Vrx1SzjnkChfgQzmY2bVBPBtunVipjubilSuFqiD1UNq26Bj/1ppeJTUSeNpkuzx
4cuxabfnLKcVZ0vvNRzu79SDE44p2B20X4O+nrP/YEsBwAeGSK11O5wQsDuxRKpW
+aq0YNyd0h+mGNg7o8doF/FKUGNhukjrpf383ScLXG7WBDLGESnjF5z0u4Buep27
oEPZ5lQVsG4FcGE+oqAztbGwTjN+Yvqirt7OTYtB/dyqsnMpRvURcPiV8lPQSUDi
8kMrQQflwbIS6GZqnuu/27feXSpD/9MjelQ4uDoqzC+OsyxbV6ImGilUOYzNHLDc
kbSeAyOK8gmEVgpq9XG2PK5g2VrAAQ9vGE6Hg5H92gLldJf6Z6vHTJSgl3uEdF+3
jz0I4+kTcShCYBCtmnsWVJHTlW1Hj6pE+Vd7deI6bUHiAp41peR9eHzW7rG9TOBW
JDZIv4Z1mKZcntVY6e8RtHg+tpRIZwqyYmC5dZ6RAMqm14f4od53lDZ8d9e9kb61
DtABUG/2/bwegBsz4ZDeZawcpy5145BqQvuZSoL+i0qFuhUO9HLbd15Oz4RJQM2o
9dFM1SX6R2Allp1cCcbmF9G8HzebmNq9McGBBzn+9emQzN6W1OQBrRVFFFGArPV0
k0WSfN2Bvv0ZCiO5DieWI2pfU4Ovq/O45U9vilLTjepRl7nMkReHav1d65VchBX8
sxYb0ErIye1NCM24DrVmVZmqnvH24lBiThN6lXl+QQY1Yd2VgAyusTmjOUJ8vzFx
V+emKkpKGWwqZXCAUqZTG1USsXScbSVNaTAueO1JkNq1JEnND1BhEGf/LL00CiAi
x7xmRQodI6Jv/VFvQ7URVLhpl+sqUH3uzOFVeT1KZpForrKcxhURDhVZ/7IVuzJj
uYuVUESjde5lJn7Om+KWMpG/420NSf6ODuZLu+wYNZbMbCJR4CjN9TU3KDq3gI8z
4WDuTCepVhBg1jCfe4FvCXNz9O1yonic8Znp3HLUIeJRZ+k9zPbxd3JCcUUUHhLV
wuNgNdyObcI1yCGq1vUWFFgo8KWKZOpivsBcK0aMiZBqHcv3ODtziwG5CWFAMLjZ
XidL5gPiC5Z1ruBP0DqCjhTsH/uGYDQ9RJj1WLq79K5+TbUG1hOjjCPGgy2ZDb07
IAHcamYvAcOcMnRkZ0FK7S7WhxMgsRwP2Wbx9OFTkbDOMW0AEWRWwevdaYn/2GFf
f+ZdFljcw7HV+adw+m5/zV8m1fmeudXNDNCIy9hUmDhdzWx6uWtHDqem+oD+zIqF
gSSdDTtVIMSCxkbVsvlkRFRBMlwsfW0WOwYrRzceLivghBNcZJRmMF4HH09GWutI
db6XEIGdc3+LxR+u0t1vj7rCEMEs+dPApw+UJryI3ud5q1o0srmImMVBWOAT1k/N
Q4HecD4Zml2aGpvXezG/fqBmq/cl2ijDCcOLh9nkZwNRdgEwypWj3kUcI6PwKSh4
b7jM2/nFd7gYetg73vfpw8gGturWtgkfyUi/+AHCgsUcjHo0WG3lHe6vu5rTnk9V
WiaeYhGxNiDIpon3i1eLMaRnGb70ZzPXLv1BQtIdwUmlSCVrqYhgXYNglN7NCfXQ
qAFl2RVv2fUdwwxc/IMuKdeS9sOATkEjnOO3Kn/fhzX6kvKtaijNnxLIEMue32gL
gq/m5ecmjN94eZOAxbAqREZ3VgJ/oJU8nnkSwvJhjmPMUfLrAqR3dPK7SUOMF7tq
2VRQVnj+Yn4qzmZH4xQumdtTXcD1oI3XSIJsPY8AaFBym7BrMCbPMdUnMlBCK40c
AN5dtVVzIRvD5yjLgbjAPGh59wq2i/PGUxy4AIiFXguWaZ5ZIOKie/j4sW1sG2gw
o5DVdz6ZJ1thBZEqf4wqjNhNyD+nylC0IwEZ+01nzjmMZmT33BbNYMX91Rv1U22X
99QgILDUVlfKtYET0BIL87qFX2Ro7EmI85unJWxR21Osl8eHiQuZbbYVU65lx2Ks
97tO+D5orb5vWCq6af+47w4QgRKJt0leSh8l6QDzai5AboVEbPH6OeHljWMm1RFJ
joNafxGVqX1jnkg3uRD+pc4o7fQYEPEwR7tNOSdciyrFb4Wl2Ve1opIXvZ6f4C9j
Aue9cv/pv9GepNyxS+ny79LH2Vh3136ivuvJEF8oAlnQPG6AkFGTXURhpTOJM7IW
ZZaMeLQ9HQp0A78zdzkkj4dnSmPQV8at8SqHe5OdaWQijurhxkuSt9XeqmhCKPiF
ScCdH/aJn7z5n8UPywQKeL/R+wuGIm2epGlIrnW5qN4TiJMEQZ8OLIa/68lVlLi+
e4LYDnVxaIBV8Lzo63BoYOmsIKaWXEzEZa8v5xonHlJWwh1XRCpOGeNfrNOslakn
RyPfQlSGuU6/565YcPZVSbDJYvHl+cDEIyUvrpfcSAFHQ6RdAkem6e53PiTTkMft
XybS8DhI8TDnyfuEP9HQuE8sSYskdQe3RgiQTfoepBuLkhIbPvfy4lVVulhqHAGZ
Gp62em5IERAOLyRozHRDBoGZ6zMenUqu8k/CpZ/7VpELlPuCRRN91DLGv2P5HVpl
8UuC3PxIi+n53BM6NLTpotkvscovs1oM+nM5RKNMlSmkHYa6Lh04bGX5H2nRQFzQ
EYORhfXdcebe/E4OBmIn3XZ5tnxpxH2KzKnR2w4MPcxFAMAIiogAGINnVe7J7Cxd
saD620XtcOtZxaWUvSAegAV+5cA3SrGGsOT7ea5E9rIvYRHGLVaGf7KgpV/xxq1H
nlX6c9BV8djtYo60Bg9CDIKRzTgVKmz+RYJr6Ej00mce6NrBg8hkpLZjbKDEmOw8
WVM++dBWkmvwdOTHuprDM5p+WDHq4zEXT59jSMxJdM9WMIaP4etCfOzWBcKfkgSe
jVidKT704khkDrCuaCIaY++30+8rngLV3ztx5rdf4mTc4VlmS24llPcQ8s+hfzH/
dy8oQYGtXMzfrzrqdoja2aR/MZxMjCxM3ndn4TiCWwH0ACEnSvAwQ0KT+Hq1EtOt
/CSWBz+3ftD0WyIGAqPqCNCMdBtuut7eREYwicTMSyhZ0ZIIrD7HCuxVL+S4H/i4
QA3dxm1DpmZq8Rc10eMzj5u12sVbUJDirN61atY3NJhy0+F+uFJJA0lp+8hwf4V8
hgmqZL+FKfSP5MWr5s3YibFASVtoJuJ7p1tgZl4gWB4thbhS5I8meoy64pv/CzpG
ygpOz7jHSEDTfeoAhvA2SYvAtu+in0kUA5EsqLv+k9PnqM5zZJpCxbX6809f+OL2
D0eWteAD5TqrNlBQPhyNZtD/z/T4hj1deYUQ42Bk3NEsCAKYurUUjnEQtLxwLlmv
3LGhX3mC1YQvpmL60kmeDn7Dow1DpDVzQC7ekXYs8hCu442eMbc0eadvjjU8I8uW
jAmwCbbPPSgn7D/KQpRNeqKoVIAfPp1nW8MBRPNNMkj7ABb33umtH1Ed053p8YAt
yp3BF37/XGLpoXkZi/n8g8poW2xuHLr314/GWm+qbsCmK7/7BkWpHlIE54UUAikG
L/rJnYTdldvLt+di5+IccifYj9ynN2H9mtlFf5owmZVo/EwaBRT0yJNDCtj10Pto
3YBOwQ8vCoblvYt7l0w1YYAB7wZaYVT1BFwpuCXMpPwg0pYjGmzo5Bd+O505u+Sz
uyOJv2SF9NYbwaEjL5gi4c+05xUfpkuwhoDh5VYiPtkSdKuL5BA379auuhQU9df7
RwD3oR5xg0igWQuk8dCuXe8OgV9zmei5AamYeWl6fHJt0Hvh+RIfB+1KadZlVUpw
pxnGGB3b9XYNm2ntRmUq04jiNukiMFjC+jckPP2fDTBt0FYBAzFLJaVGLIdYOwCV
bGDPkWLYQ1SmGBPQXajwC+nPoQqiUaik+xnziHr8Nko1Zd/zKBeJDiTwFsTNm7SW
iPjJBkBmngf3aYPw24/ELx46eHGBgdcsQV8Pn1wV0n5avsGkz8awp1fkCdmbkoZd
IcDrnmc5ten3nAp4N2ehRZpEhQFtVQqqB0qaOvuO7MILbvaJNP24vhIBYrFmfcZq
SDZ7P9qWs64cHzIX3B3NnAEEzxHCRcXA1+qnJEa7TLYoSyPNGJ/Kw9ac07LNXGrV
oXP52+Lp8FSSx+u79u7iApYHqB1NfX329qFb41Ek4/0N7Q/pcgiQe9d+FDvKOnYC
RoRsbHCpHte/OKN3IxAEZWmDMpYCTyhvcCFF2XW7ZtgrCE1tb8eeWyiqWoK6/HnC
FYJEb+MUQymwIwCTj9swto31X4h1Kl4AKoEy+sworPj4K3PCBd+ZfmHWyzqRgMWC
HKcUEoAnfkv2xgDT7QN8qc0uNrC3Xi5Pn8d5znixviauDrqPBjwldcYhM/MjDhCa
fUFXyl0+F9rsNEEDxRcmj7zKw7OYN49WTLObtLbC8bhtfy8QlVj4GgJrWN/NUV7j
WIuOrp8REDcTAWwTb23jFK7mMjSl7+o/tN5yc3B7F091NcpTvHsHaFwr3HDuAzje
y5teBofDOBFw14MYs2Wkiw8fgOCZ37qEdKTrgt/2ACd7JsyZ0dHf2Bwp6pvkt+dJ
uem+Eo8Ccryvm0kZrSLWHy5RbYTuwLP799JMZtf6UQAiV7weIn1qElxiTRax3p9a
EQySjZSfWMNyq6wuY2TwFmM7Upj4IC2AGuFMvKIQmtDvY8zewxJ/qQXYlJhv5vy8
UIPJHd6TgTSTvVajUwW1zoLgSIR3Rt/fRP1MoxwMeGQwXaxjw2BcmreIWsiYGIgC
f7g7Xz1+GLFLDtimmZ2JkFkr3//oTOmsgDdy2eQjM/mF//IpDEhGMFmESO+ypphN
LMgGA4gSiRKCdO7pwrhCFWjomUUrVWZLFttj/F1DTsR/ueQgF72W4i1Ue+Mhi5Ui
oBIE7yE9XVENpbGq3Ki6hr1T/f6BRhsa7wPUlysSXFd1lUoe6BJDWNhSOxhjftzO
c0t5yle4eKnrVSeVUFbKN70Lfy6O1/Aa49MDdHjKGzrMjFhVNYnugQUE52EW3UhW
QgAa2gvw9sBb5Thj0yL/90yb4SzZX3g0WlYzUBc/TFs1lL7gYg8OQ/HRKCfUZGI/
cZgKO/zZUIhTGee0JyhaVzKCzVb1GWNTrLH3nCI5jIS708TLyeRgInyHgRt6V7M+
1IhWI39yE5h41KpeRDEwxeD35SWG+CmhCwm6FPNcdR231mxOSq8NLrVixZYnSq6Z
Yt19bIxRVwy9RFbiQXN5rCLOPVa08WxhSjVwS9s2Hcc9lHv4bbGdx5gVSREvOCG4
2NiSVCe2os9rcnoO0BtuVTN6nZ6iHloR1FvCXybjyhmEMoQq74WYEg+uyU8TVD1E
8yT4StVxh/iN5PNN+pZ5heHauYFTjKmGlWA6z3t7P6xNiIo13RFv62sQHYvABDCc
j7NgNJWZOJ8G7RfzY4JX3R/+bTf9SaAu24qaxiuDSoS8+b3nXdmFjtEl6+ZncxEy
rl8CYJcatvCna56njdh+SQMkvYurXr3KROm5OBJRCrgf5t3ykvkTYzQYim+od4rJ
gTXXfg2dyOG53DIIuh5y4Fy1hDaezdX6uTdevlq/pkzsnJrlD/sSbujnKhJY6Eo/
mdLAhMdNHC8k2FlbhyJV6ViU7Qhp9m0qOeLBg/55sVS/L24e6H3fpS7QN4XVX6cJ
W4V5P47t9QF6kgt0BeGtrDs9rWAKY5Soh2kEo6S1BXVUmJPV/2C5hAkHulYnvPDv
Kx1Zzq1Uvc9ujv4Y23xJKRSltohA9ttwbUiN63ZZkkigwXpxNsguPv02UW+uzII0
qLp8iCdcVBYo4P7R4QFUZWMu1bTVQUnsM81jG0/+e4nrAlOj8h+/Cruz8QXOUZoS
FtlKFJHutwqMOcSOtEq0Mj9vRmRGNSxcIxVZRlIpTw6JgJiPHclRZ3z7EggVmVFD
xhglyqKR/oh93q2SN6Wr24G2WYBUJSfiS34MtPiK3PWui3ozTqLdsqerJqLGoJhF
6B0FClba8Df7eAi2mAF0/Z/oLQUi8o4lnCxVxBc/HXFdyyEiUBKVu5yV37g4nAOE
7KDjY8RhRDYcuXWQnK9JEcIQTE/9mq1b0VuvhQ2YQd8VT/mqlOt/kl3pFWBnoFVN
ZmKIAb9/MfzygegInvRJIbi1MK1dTLvAquWzKw5cy/zrTqSqsKLiCtW3Qp5bksys
q86SHqH8EdMmYupL/g0AbOqiu+spny9hPD9wozFSemv5Kg8DZzS0tg2BaKGHZG/C
SQ82Nbd1+tyyFfThnv4WFpl82leujrQFcgeeB7m5tlbr/ZAuLtCw+Fe4sgCIojFz
Ad2emd2pqk9IW0LlVGua5gUnvqh/HaukGHKsgaqOQ3nbekbAI9hDjrUyxAhRhsC5
I1CZm7W7Y0dnyHjdwuU0D424V+TKsMab6e9QY5gzoI0fM3wuPzWcNxcg4ThVNqHP
x0GVjGF3ygc0R1kFnhQsFf2LfdTVYs2/gVTPprfYFTJo3bhE/utz8Z7LB3PN2hwa
TDs4OfFpMoBQtO/4uYaSTQcCJfuO3VvnXKmSDucuyJTza/ENP6P7P6AzWOCjOpI5
88yV8gHUPtD1ILfd8kOniRg1joi9Ux3HMM91iCqrpOnCkspUtahTGFWbmlMreehm
UYCR9nC595OyQh0xaP5IoNtgsanV3IeT0PLmPXClw8uMLy2v4J+1kpgkUQkRskmD
/aucbLFQjjYMfl4tGRkmiW8nSrjUrvwcqzgAChh38dqi7FOuaABMLeyjF744bFeq
/xq0xHZFtcgAxi51QZ1PUSlsaqUV5wzhitoeNpsE+vBBcYIjj7n6bxCQCjXhEpNI
/gtw7xXws4juoKfFT5Wvza0XE7TnxAp2fCmMqHFX5JDMveqhi6xo6HDddLQfJ+Zz
gweeDWueW+Jk4RV6vHx0a8R/+5hbuv8MJYN4XiOgYbGGcrJcIaCHTc1d5hiom68W
ugwrD95AGwlGGAIGy2nni4mdxe+vohFxWdpz4a8bR/oahawwxU9n4FoTTUHnR7gX
VnJ9FS8u9FHLvyfQoX9TaIWSnV+8V23BE00hFnLF6OVqHw65HkqJZdQT2DF23zxm
Ll+htfD3KObqI47gB7NRNjmFFcIfihiGdsGy1qiF9+fgWzG9YGXfPXWEL+81O6GK
4EyN9p85+gaPl8KWllRyrbkQ5TrykusuGvnpeW3wgqR8sJD9p+H8ENcVGFJGMh/F
VVM6AiGDV8/NabtdHLPtWRCjjbiodDqfz8gDEhlJZavU6x10tcDzE4ePYeNUCt/h
yQDtLO9bGdXMuY9AtFFzLrY2lsuox6tAJnyGT1o1ww/rPTNutb/WsNyGkg+diJi9
ryP/3NTGI0lnUUxxa8vmqWYUH4+memdZV7SZJWnUr6ACivbeFWgJ8L5an8Ec+Snl
1vMJXPW5ewtJl0IDGpC4kGjv9ISkODtmNtPAGqzoY1Pa5y0LZ48Jee259AAXj1/J
RaEuGyEFjAe2xyj0eeAwAiyhEl3AXQZHG46H2wXn8/oSEUyRcFeKWOV+xRxEbVcx
XFFEB1s9dcM3RHaDIgobY9EOU9S6haPV/Q1D5nYnn25bn88fRdNsxTwEJDPk3L0O
n12fFZ/zRLAjwjQRZSe+Edaddg6jchepm2IGk4yhZqkCdRsVgxfIILAEgWn4sq0z
tRxpMHtaboKANzqkihUIJMNwFvmzQploq4uY8pVbl1TctDt8UZkph+vcCJpr+ajb
nxkpDFvw4eFdmxYi0VeQzpNGEhTOXFEKEReMpZy3pH7zOcaS/U6qtO7uojGEVTcU
Vh38yi7s0qn0CWhs+3o5jMirIBuqUrFypmVdU7Tnn2BZFcDRU84TS7Ja8ASPE2oh
cAKyJXY+gaMu6yRcrnEcI3dUESHmVrSpNRwbn4Z1UhVK7re57q83MUoatI9gaIab
GZR0iy7BZTjs9VEDwlGLwLUMtlJipLOoIzsm4sGNCgbvk867Y4sfL9FQq4L0cUaJ
+Lai2SpWIWj/6OiycSZMGZldIwEwhp6ig3/E01EfGDRY5kUgb6z542WCDUOJ6Fc6
0JfZiXcdeFBLXhKUqYAkq5/QSOjbDlzk+e5z0P3StnzY1X/vWhelA3XdIShvAsMr
CWxYTUJSM2IOob3loN/TbDGYKgoBzCD8vfUbGIvjpMfIum2z5pgDc+EyvtG5Rvlo
c9Etw5sBtMzhKqOoD+EnpwtnARM6hJ0yVA+zhFoc6nHD73e2xigQtEAAEwxBaqgj
WVZG4IKW/p8AIz+GZNsWOm12YfYkJG+FPsEOKk7sNZje2gymnhCvgxM+pnKKqbIO
f7+UhCno0k1Gjgrp0jVykGfJnGi1t1yMbLzKfUdYK7ylu5cNR2uNG2ri/zGpfclZ
PPIOY2XSsWMfw93ZmgwIh047tLjiMnGw2vzs/xGJQkHxYJjTz15ApejLDZbjiaun
Z3g3Eu82z2rQrU5xlPBd/Byv+IMUWSWfqEyP81yEKjsiXr8B99Il1hSldtwgKzRB
YafjR/1yfIah6N8w+GWyNODQl3c5bGcgY0TDr0EfA5MJJdcKDgway2ZgPIcnaaWP
dEzF59FzOyYzLUjeDF3VbgO2oZJDHCPu8wxpD3lyx06BbSjBoOG/acf+cZfMKR3w
OW3yVdByNqX9jEL7Q28cU8qkvW6ewwqtncouwbGdJmTXUnyB11yUZE++uAAoPB+V
Unk+q2UtO3yn21hkifc2AoDEMTXklMB01eSh3jBNJuDW/2iP8kV5WgiqEZIjC9zr
N8O/SMR1rjbftQoQZO4zw+rTwEBUD5u+lcc1YXT+rj7ue/BoUrOFSyza2X1cOeOd
0KEvb0iTMbizV5GZpveYpvYTu/ZVXnwLp1LNTSLmMUQ0MOMgc9KztkAOb0sfOHqp
3YBZSgninNUVomM+Q9439F1TmOmy/CL8wG8BlasiSWYXg4GMkihVOnEM0i/jyEkS
tEVu3SRlgPriawHAWkYwkNQz+RmwPMBorttdDtm279df8UPv9326tOLrCWWf4s/O
u+ImpWftUgvXfTvxFkQJSzbJreiNP5BSNPzxGzPzx9eUluEAqGSHbY8tMOb0TFmg
KKhkFZgnsYcgDxZLpUH4oocHQ3wbKtHqIWDDkSgEAeCqei4rx1v/qDvyvNqOMsQO
VjuIfb0aopSmwgtFlhqWVl1UfYn0h2JQzeBVREK4dYfmFqSbvJRJBIlihlVlSCiA
LnPB6YZc9ox5nsCDMgPAzEaxndEqFf82aMCzrgFjh6ByAIZ0H/wiTlWBNQBNt9su
FDJONk9wudzYG6E5GapW5fP+PHIatKz6QQQ5iqgLXD5MjWaHOffuPw4QVauj88W8
C+GbNOpq6V26Gf9+3HYF+sd3axWT7St5Y3PmwmvHrRInsTWY4dp28jJbFb5M8nAF
yZ4kxz1FRCceDtDfiBg218NcIDc+Zks1Rd/G9BXFCYs8e6Ka7/J16EPrKk/myMdl
CgQAgpl8lT67G8lO23HWJnKs2pcF2iV3p2NLmvMxx8pn2kE6wdJ+K7avEfFfVako
+GW8+3jBexZIij+qXpQOV62S0TsMfkEK0QFOZ9BzxOYLkQeJOrpuWktkYIVZXLtO
ynlBLRQ+YN5OKVciE2VeKYGtT9kwYPS7JMxuyGeLdC8QxCFuJFPRXhKfNVXh8qx2
OcgFrhLA61LSNF2YfCu231CifonR0q41Akk4wqduWEZ5iVOrZ8peiaguuwtqxva7
Ntb/co9w936KiI+PNoViwEQubtzOE5QsnAXYWfmxTvfGM7W8ElANPTNFpXCmmRki
iCIZRCQXep7qCLiFpW1a2wpdSsT3W8rj2HhUG9p7jrvymCAAKyFhTwLdYm1kzmFA
vGgjfKvAItqNL68qzA61sLwwmBikaYGVdJp4hWXWNdVlW67TAbmn/BSX/VyrI8SV
dEcNYEa0YnwrjWGu/1/p8MqeRc1KmmT3FGIGVL8cvkhDXAowqZfHeczhYWx+BHUU
19FTf0JaLe8yB9uNwNcxsAwD//ZgpWe52CfPvpaAcDqeJqaKY5/nVs4leTZvtoAy
vVLDkiRTcV/4zdxf9uoptsliBRwAKx+bTNgnZcXyKmcfkffN3P+OftSk3dFocNBT
kkSgosFlDDv10JsA62WkGZFl1agbuK4IJNR08QevPyq/Ip6zXbp2ThqlksPv6v34
Yau83lHaMSz99WyEMbNBr7nYtUg51PcceY7Gm4c392PKOagDDHM9kGh3qObIDJ0k
RxNUeUbpSLGnEo7+7SadfoOY8Z7Zasw5PtQBHSvRkIcgyBnxV8+jlwcdJzB5/vEV
BkKE4FTBoY/MN6gVoV9dNut9ooYgyxrV72nYB4P5rr9KYQJQdg9koOfMUfm2G64C
vlDBEIVajooW+f71hf+Im2ukH3S6KeYue5j8cLqqtr5y2RPDjhZqDeovzof0RrsR
BJJZPiqaBjwUzZd4G/M6Xc8Snsr9Brrlm1vxmMC/SV68V/AY10nhpgL5bOAxW/TV
KCIEu9fxzO9HR3Eo6L5/EXi/kGtDOFNXOLpBaPgo8HlL7K2mFXR736NhutHF5abM
XXI6KG+H6V1YWk3lItK8a72u1f/+1Lzgn6hGudsZ0M67DJXUZEaA8WeQSIfinM/z
+pl4e4IFF6IBzbvZXdJgzbRwwhsdzCoDuWRngltdBkOlqIP6BqRhXYlIz8rntUts
WjrcnadFoh1XNAjJbfSzfX6wD+i+hKQThwQ3oq17u9maR/rPKhxaREbUsT1nqivY
zM2XDBdGkLJai0jON8/AZlt1oqxvbXwBCeZrtdSGmP8BgICV3JP6YHgJfvYCpsH2
ViUi/3aXtABuQhPIdPnXI/ZeUJVKbvIobewC00R4GGfrqQb9cgVLuhaJDBaJYf8U
ojIRyouCsJvx+PMHKM33apVpVARv2QCLiYEikyYDvGAlsDVVc6bspDf52JRLx7AO
bx0ORFuf5vI9+hTveg7oeghfFZjJQknfbR0WIhKCG477FlrKu3X/YhwkFwU8ZJJY
wUmNPYMk+VU75rlnMwjpqvmwfoVZLFESUey6iWCTaAemWM0eYVK/FXN15E34kPte
eAXX4xRiE5pfYktAWGIumRhb6AQ4pDWRNk/N630R+dkNUenGEM8HFN+9zLq3O3su
fBEOTY9aCr3Ymjzvl6wW1yiNtp596rX2PN1nv3iQxGZFpiK6Ye6Z95w5Qf1ShbeC
WG08oopShiDLaBHAnU8pempCwWOJKiYEZX2qLfDCB5Kws31yYp57c+mZhh3QNYUu
T2AH/x2BdGK/GnZZtogL4iipQbsJbl795U6uFBXK63UkCvrhdwhLPVg9LU3bNBGK
q/QQqa8X3n7QnwcPXiPcpUUjNrCjm8UGmQshViyvuAdV+4fb4DbpLi9VhOhlICzH
zD3wVhBnmSK7+Uql50mPjWomX/Tvw6PsDeluSZFIjljCQjSbnvmHT9nCS9HytDQm
hYdxXas9SnkC4/ipG0iB7OzQ2jo9npR1ZbBGgwDeQwKnOFInxcqh109dXTA9jOvJ
vc1SOZl7WvenNLV/934uk+RhqEtyXDb5oM13FnIX7uab/LFw4clWrHUWIS+b9euc
G/k8HfllKEi0h50Tvey/UlB383xgrL94mGF9rwrmPcsvSamBkliNW2RcMruQyZcn
k6WkOxCH8hf36mJAy9qTmWOX15ILwd3qG6qNnfcshJrse40s5HOg+a9r6T4qFY8e
U45JzFKYuw8rAeEau3VelPUi+6JiZ4xEWnRpcVFZQZnINb4UNhs84El17iHc/fWm
MhalLn4ccA3UjvzcFZgItS35FeJiv/TxpgbTf2JUOR4JmLPHrB920j0Hc5pIdXEi
Vgf7IWPBbP5Nd8ndf3kN3kNOzPb71fWjGjrEi2EU6MDiGNNlrp2Ap+s9jps37iYx
nlYQP0Y+IonlseQLutEpemSro4R1kmE+fETHdLhNGwYQZTpURA1H3XIbp7hpejGC
WlelaFB4am/sBE+ujiIuHCrANIgG6MBy9afLEL3A3CdB3AOwpwhEN9yKwtp8jWLV
Qo6SBtKA3CtSXjFarNSP7wcMwSh0uHWE2Q8Tw4AqbjxT5yibqSyKHYpV8U3M2ufF
HjF6WGZirZFn8TulyBfLOgXwFJ8PdyvixE6XQf0lfKFm0RaPja4B531qzLoidULI
QYv+sfKpnOBgfP6tnk7B02SZYbODuiG+D3EmGe23c0bYKTkF9hYQlbCaAnEwj+gX
WYJAsPNKcdyGT90DfQ/ukhYxPoImd+LzEnfE/gvdeS3M7DUNCWOBOjloNG1JO4x0
mVxk6AtPAphZvIYL/lw5uK3I8bPH5WFwus1zf16HexNrnPIvtglgfyup84hJQ77D
X0NS3wkbxZ+Lztkg9zWLuh6rXsKpZfD7WB6OTBrGngVH+maG0/FmW8Xb1NjbORR9
vB4rL6CoW7NPr9+fQiUAxhuIf/2IdOiO3e5Kgo+D7bgY4tI80M/LXkt9OGKnQ8Qu
fl3vpJsEj7l4pSmjCMo8FQKSVVauybA7/JUYkhkTi3gBhabvI0mXipnxaGWHcLcb
qf+1aB4soAQDp4qzeWVT5cE3IgkZu1rfOL1jtNEht0qdZoZspd1vewLF5gTkq8Gq
ecqFiGKyMcTdzDfECVyy+eBPPW9yzwGo4WnufKERzcMmdjjrXp1PNYYot81XbDnp
iXZ345k7FT7QS1GOMUprHYk4Ky7ccS7L+0sYaIaQcEbD5cMujkx/8FQ9K+/SmvmN
fDHwEjku7cASf9CHCidDnFBaYYG0vRDaIAjaUzoTgCWuUAPR1vHIo4s0Qqrs8TRU
PNeGjhz4beRrIw0TvSXloYWIqwqV6CyGj9bLE4rwR2Hqn33J0PPfp+owwLJV1tei
kDtyGUTRBolWetna2J0+D5tyzJ9lHil8PjeLn1tKyUkmeotDEmGYk4OjonJnxP8u
E1cHcRdauPA+M5IwoKpgkzQVYi1ZTgf7sjS228yW8woDHHigIt5GhfcoS/XLI53R
ejxsx7yMhTmVngkCFwTMOnB2oXQEXvg7phJODU+IcB5LCs0r0YVfxW6nCGGdFjNv
fkijuvYbr04PucfIMNxjKbyGq0nQeJEgRVdAitbyJJxVkgWwQWR9SFlnlzliO1WA
0uyG7Lyv2t0SHRogjyUAgU/E7ecvaAU+Eda953bKyqShrIPUqAIoCxVpAY4PO+iv
mizC+AyJ96lQ9SgJXiHb1Hly9M0QveRXW01siQIppK7QKDG88teguLBPgjbeWW3V
ZfdTTrRD+EOHxCkH3Z4Zqup6nbQEqrLmVC5mwXlaDm09m7o4XOWyeqZ7grPYKXET
QCtOPWkn/Cq3SiYXBzfYXtiGn+/OEUliTVMFzNg66FUNrJBaBs3EizKJlH9mqyQA
pecbdLlIIgvh1UEECNK3Nyi7WhYAw8dGZkYGb1dBE2zC2l7Fw2EHlhcSt8P/m7F9
Rfm6jITi2mgnoKZvJl+0v2f11KAekCK05zNcvasiuexr6flDm/43tTXAgmeMc8y8
xB7Qnv1mHs566bb1g4ulyehANqcVqg9pDPFfvpPCTScVaDcQWeUVWaqjrzSUDl9q
oNWLj8Ri+0Ce/Q9JqDfA5yBTQDUOQGFiwUGvBCasOMHUAMZ1KqqU2wW00/+uLifI
+4WJIRY3NK74tP2OmYc2B6DzCTM7y2z1QeQ21epe1M3sN4KWP1XXzDnALHoPBaPY
YhBB16bP/knfUjAEvp5xYBtcBRAE9fzD+NA8Iqvzen0q/dk0c6+WOFQCYAqowiu8
/8e1QgEJ6I2Yr0GT7EmqZehMIWQcerxOig2EfqNaf37wc7E+ug0bqgtzzCy6QuXo
nJ7SmArpngR7XObhH72jp+WZSqSGbhAziKgLIJl5+LvhVhJhGaWKnvn1dm/td+61
JwZrUKvvvbYwepW8I8tmJezYjDhuupmuN1NTERQII6me/9/5iLk101mTsIEMWjnt
rhfnyKNLLmi8BTk9lihqSWun3PpmGj1ZkQwJWvFCmPP1KABjZch2jIXXFi/1xtSq
FI1VSHbmdbTLmchc1aEyPGn+5TwNrDBIB8P0giTmCOlvHVWhbOOnMGIxDwaAX6Pb
1J3+k9+shsmODHji/gF40VbcefWD8B18GdSmchg6bGqagIP13w+sGgz1S1hRibGO
VvodOwmlqAvIcc2xw1adLEhtap1iEYCE4yw/qmxF4W9IJfKjdsgMzY00CV0UXJ+g
tL16zwB95E4XRCZQipYu9bQI7v2tTu8U7ctOKhL/MipL2lmTJ4cggXmg72FUCJxw
En6atTfjmqgDix0cOzJcnJGbxC9HAOrkea9tJMdVmEkW3Tp6TMDf5L5ZBDhsIwY3
Q99DicUTcqZb8763NJLNpL2eGQ52mCsvmn7h0Id3+e2vtAKytxYLwptHludL8tWO
1ph4cGz4KPGR8fQXXaeUO7ezTy+wSIHWkaaXI96aQpli5beFAkyrZtzgkBh2PYZu
Y5V+9IHaVNi6V/ZDnTPnZhu0wKzkW9DTHh7RchEyXirZ+n90UlbUcphXoFjNGLwy
QQxnH7c3P8JnrCek/rW+JsvcDWBe5IDix4DQ4W27AkmdH7FQyi0uxF9+1T+XptDc
54ahGhhBDibSa7KqmUwmYoetu/3FfEsYvYZy8vj9Av0b5sRppHeil6eKP9uJQJ+4
N/8nJZPTw2mjP7VmcWHZ8erv4A/p5uZJ7itS8yXnV7xKqRxXZ0FPFzr4l+wRH1wq
+qsHdjjiy5GxiMEViKMCCI8JUH3fvUT7JPCYGt/TlkMAPXoe6Q6heoIx7b/rVWuw
F/NeAtvwJqFIP5OuKGWTGe4vc/XDDzWqGyfJwBLIUS1dKt3uCiOeeIoVV1dJ+UoU
v4EFEtRe8bmZtnkg+7RblFRJTXbKyqN7Rv+GSewkvbdx+gk5hzvWYZ6+vQp1pfez
r6tEaaniNWMjHV865KUeEUuK7VIb2t6PTWQPwG2v2sfdDbP31iGVBTPxWjK5zdko
Sfot4BZ8sU5/CJV+G5z+iR/An5WqprMKnRqerbSrHD/uSsTQmBmFUx321F+ag5Vq
cCLJnn6V/YwfAOr+aptaTNl+QKkNO3eEHHswNSzzpsq0W9bBu0oqvMf82INr7Rn2
+C3W3nghmoHeSu0yiLU+GiW6eO7yYyF1oCY70uf33rkbGHiilkW0zO8Va1fMwej9
jnY/oGVWRU/20D2Lxe3R3yW4otgoNTmff6uXm+NcfIpmpkxTA031mPsT+3zCgztk
rS4MqT/5F4Z9WBVCmBt1ceRLkWYhv2ddsgtHrK7mpnJNw1YyoWp8OSdV0CnvSCND
odI83+vBAfQy1vm4IDysnA92uCe5NaI1Yp6U4SOHPf3Ap8pJ5eWSGwXVsx17YcrY
HnIYu6VsbKkxS2oQcpBZg9ysfBvTSww1xywnx3maZEeb5DZlOh+uWLJmWE2bhS+v
NmwcJp7fFk7wr6ZBb8EEQW5uJUhSrsN3dq5pZEPNy0L4UR/vDpmnsTFYE1Iou9yA
77NYhEIaabVywLOamm3sRrjihpNauWDP2QnkmMDdGr/CePdxHryGGKM3GFIg8GzD
iCXXhobQHvKYGmDxGC6QKuTHYnYeWKjijqq6qgjriAY59DkwTljHrjAgsOjPA+1M
rz3f/1dbbw9J2vy1UEcxu+TOARXHBT/olmwXtsPCuT26fsUfP1/hk1/dccbLAda/
b1WRwciP4/A9tqgJLUqXKg1HL+MOspubpnImqpSV6ONr9RFqDTHFNPdO3cM6N7vL
IQNEnQiMsl2NxwmPKS1NfZ0SmQGh1M4rTKzguXr1KXLmP+a3ochXcXzqu6h86hKA
1S9Ns4oxFSnV94AxPnel5u71ZpbytDzjUmVjWW/BuK67aFCVymy9HbNo/us3kDd6
CpoUd04CLuhU/FmlvX1zj8fbsvRekT+dZlxrygHQzBggJVAajpKeOhBoyTspPuDy
WH6NNXi1CG5tmqYNa+Nh8ot/JGmGAw3Gjb6XzToVW9HhMXMdKyHOAk2Q3jTkXHXx
CNyAU0kVU1ADLq7bu6Kk2Wv4/sIXMNFymD7q1mxRZXsX64KLzdaBdv6iwVBqkz1Z
yYTi3Ucng7Ba6ZheW8nPFYK2AGU90+6KSOIvCLn/sxNRFWK9C1Js19xAc0A3PSbN
cftZ7igQtekW2aYbltS3ZA1voxHjULdLpm/eDAJ+QnWVrDSCnSkJ4WIfeq+9yTgf
j2182vkYbJH92TPckB1J28LoZg3IJGWCvGgPZnOgv3azXm0rzyxCNVPMxRFzhcWw
9zQgLQViZQAcxsaJ88GyFGvZ7PxnLMqELle6cDe5JLxXIsboV16sS/71Wx1xqv5l
R+NmMbv/hIGyeKFQKO3DIBFIwMLm1AiuTJld+c/pT4Pn6tNJjht91VafiS3Ipl+O
tIyMHAKxwlMzbd2XvASKDo1/9ueJBV+WqGLLdrYwVq0FW+Iu9gbMxz8+sJYcfVbr
BWno2nQmeR/FNjAQ8klxi5UGAepEAPTDm3khX1MaUOEs7WicATIBb6oxpwEpOvgn
KBmLLgPhAZPHd01MjMaUY1TSHa7cb9kVIOx/CxHQkTrvPcp+CgQZ+B8X5yDYasKA
m47rYQ/bNFAAc3oSW1rAwd/3rACm8VbCy3Dv0J+663bKLkHkm9yxWHDl2DIQkkVd
y4Nj2yHWYLTfaxTwgCkcE3K2GSNg1CxXj1j4domp78w9K9gbBlFDHx0IY5ILuig0
DGGXRWcl9kbNp70j5cb+sPiMyFoC7TYtAPWbG9hJcUjWHBKUi0bRz2RSN9KvqtPO
ruGApReIzuuc6japdEBCUhhZxz8S8bQm6uIixrx939eJc2pjYHgAqRdB9okwFAgV
h9XK3NBc/zx5xdH3zSFDQQmPgsmUsI768MWnIgVGhslbrrJhl5gcJjIZ4oE3/ED2
qTGjlZr8ZKp1p+jVia43kP6qq++jbkeY8pK5GzdQXUH6LcGx2z+tR070K2a5Usdq
QBUb4It3ClqnT2cPfLdc+DXEXxsz3QQzty1RZ86tLzdCqK2B80VbNKvdhUOXA5kp
Dqn6jXlr4yYpPsb+cQhv5CcuOJjCX4Tjr12DrNHBRoMqyJSE4XeLNNSTVFLycnrb
2fD47lrSFPh58me3DBC/8TqEoqWy2pJSRsNUplFwuR1A0sveXOnN5FohPIKL/cbL
CAq95cPbhmXhpdrRpu2lGmJdY4EoQda3IGOgiL5E1ClfwDMeeuc0L4KIkSjXzY3X
aWnqQbB4WVRnUC/l2yQbZdlx6Pnv9UlaU4GdxyQb1RiXEgEp4O6Vsg9jEqiXhtIO
ZLltRnpAIMvBAd/IH7x8SUZelrHpcmNBAXO9ZeGzc1JxFvjDvhIx7No869vt5NrB
XrkI+PswopPHUfmZidlqL7vzG0h6SA/iYCTcD8re9fuk0I6BX/OUTcKIO+uAygaD
noZZL4aPphzHMOtdxsIPCqtHjKfkpm3On1MF6tRgXTADN9rhiEB/b6wjipLtISDt
NJhN9p7t631VUcRnQ11KyBp5LQfKRppD1LXiG8isNrVVtG5qaVsmGUDczK+upCZq
y6YLdnKn6II24nWNN8AaAttUCDXSDUoqIpuYOtkag1pkgWnORL7WXHBoUaf/kD3k
eSs/r9yMUhqLNvpITY9J1RdI4C+OzgQJv0hR1NTJONrzut09XZH96CbVk6fiHGE3
Q8PRUpfCFTQazR8e8HRQxwJkOo4wE1mf6Eai1sfiHWrw2eSoRcwRgZPSXVFvrVHN
dn6AQnWaRuf5ywWMHd040znZ5PCW3UFUDvYkOHtnAmuTH3H0UmpeD+HpKqdKqXnr
sAJIMYBi9ENQZcvm0Ehc9EXoiIm/5F12Ch069T8myE45R6MTAg9eHh9pnb7TXpAq
nxCOMbp7vSpZPHz9jnwmwzZW8KgDoZWXMu7nFaRie5/G6c0yno3airxpysUR70Q6
U6dcppDrskAn5/PlmaRYGVw0LpEz4TkVi72QbW+/qDGZk1/NRrRKqBz9l+MlE5lX
aGvm61egQ09nQk5yvLsSzKbZGelyL3qvpPyOp+ihj+py4ByL959k/5M3pFGrcEo2
9NsgbrZCubCVBXQTetbCYN9q9FnBL48kPwU9rFYKEt3PJt2yVlNvi1bSV1Ce3QYx
joyh3Jt6YlwCbG0Gc2EcvQS0OgQXHNyyixjht/OdOhYjkBeRmaxxVCxtZt8/Ds5T
gkCnL8BNWBFrWB7MTrFHl2Q8uuGg0uN3dtFsVnybI6tEE3Cxjr5uRD/6jRKSO0G4
I6Ez4dtLzI0imDdrTNVhSebeeIu4NtRzu32SNYgkNiZrmo1vQhPEyb6YDbLp4pIH
w0Dp1jRDOdL6yHQB5S30bPionjVx1qq7hWxR4N9cyn0ZvH78v6tnHiRt5n/gTaB2
cfVWNVZRcYMw86ZJVRIz+MlcWaMskQuDquXWo5q2I2rn6ESQO7hNRFntDdCyV+/c
+EWStswQfK73/LoEcBKNwLU2rsl0BnZUdc7U1ZaW8S3XAtrgVPJwGUBZErtuc1BN
PvXpu/aFGHVyg4v2y20OQynQK24dcfVN7hMBJhb2xPHiBHtxWOD5uwUj/DvykWAN
hC6v0plKx/0H1tyMOa6mgstYVCPISwx+C4jr2EhPufsWhlfrCen3vnJeEZf30jUu
bKG2suogqWdAdRtE0bpSM8Qgk+sCxam3A8ngmfTiiuqXHo6r327LjqH8cf6li3eZ
e/VP2EUbJlmuzlhrjm0gyar7vptGsbL1W7WfhTvQkJjuKZiOEraOX2o+t+reKs11
B5+CLeTQY3J+M6nFZTmh2htrfk6kALcV5YYxfQnZThivrqAuR1siRV61R4YZ5W+O
uxGQNTuLiDWrrgW9eYvhkmlR+JIxXAHtoSsjp1d5Am+jw31roIk9C1FQp09x773q
iAs6K9yxiTkMwEqVRrR9/5Qk5C2DyF4i71iIbvBb57FWCw+bEtFN9+eKGFtmdUSe
VvRGhCeEwg+MIirKZPZ+brJUYREnV9Od+npJYAiP1GjPRzMKzQdi8Q1VSDQr8UlC
lNl8FFHZxLquXV/lp9doFo2R/yk+iuaWxB8rwGSOWxbVuYyVzu6apqqxkVgoOZ98
LP3e94cGUETF3RZsfxe3GOku0XAeNCT3XbOJG5BmX/bp4mlS3k/IkLvVKmtpUMRl
LkvV3egVxSorYMqEUQMrUeAExAsCOSXB9gDf+5W3TT3SilAYD67p4nTjHgs0HpK/
q4tMB3KAYn1mFTD1XMemW0lK8M4RkWVjeVbjLQazbY+YkQZLYzOF00Y9bKwPA3t3
SuT0JOVdZJ0wlCDNzaQ7B0u/n8hWLgzXofbEVMY3izdHLAYwwZmQD0fENnr6FKwR
UBLUJOXpDbvdaB5bzmiZEbkA5tK95LAM+EnWeEQbiqhRQtvhoG23t2mISotVKptr
oROjgtriKvmvSbVEzntvfV1tUlvTBLwW1rpwU3SKArSD9Ge1q5K1BF/md4Zf4Ljm
gnKhCRCDEMqHyvqJKw89X2mm2S09uLJmVBrVMrBqExlW1Qy65nxGY7lXgS0rBVrg
qIKtp2zBKTDjNfqKp/rMbSafzwj22oInMhoSepOv7eb5Ny4Yd2Av4/3MOzO9072F
1kS9xThWgpyRfaFi5n9ggyEkCllNnCl/cxQ9KRV40gZRR+CGkoTyESNVyjm16DLf
Tqt7wo+9gE9AdNQ20fGkJD1HXOd2JrtClnP7iRoFOnEsZoQ7chW67YKuCp83Mohu
BhbH5yuFOu3I0dyCWyJzUAxEFBByA/MMIcgE0wtAvBbpoMUpG9MAM8u1P6Fnw7yf
jLtOd3IIh1snwMD12Gr17Jl4NIejv9+BNRUsi52zSCIYTXzUnjzPpLpQFI5l8Zcz
ua1hE85J/Qyk5UDcGmtirJiZZi7Zc9w1dafbAy2EOouJRjcZa9kUwFgrwglD7KrZ
sQdyoiNcAQQ9rS+eleYQ7wltbv6+IvAcucASoYerqt7mY/TE0ehcztst4PoeVupI
pN7Iucx0nCmrXE8ikkysKrebN+2Y37IDcSkj51kxHs5EA7gW/6p1fvM6lXGDu3az
5Q1FraaWcYRICB3GHLJkPr2pDFVLyWJwQfxDNR38hfHAzBamQAGJRjA3xylqlotF
nbR/5R2lAcEdKI7GIqGlQ+kvD04D4WTG3W/1PtOHHprohsFeB+X7gWcH21kM5Gay
ZzvU8rZYhQTaZ2jLMTI7DgzEcXwOzxJNLqiQrjM1oKLPUvCAdcUhKRIMoZbV/imC
Ul0w322l8J8VaLXw5uv7Pqjn3jB/66bcOucMfv/cUuExQA1Dd5ZAhIoosIQDEQal
k6tKyglkMZhFlvXwFk5vy2FWCLi+WuTflYzpHe67TnBuGS2hBuUPA8/eoqpTpi60
n6EArZbRj4Iq5jYaWTe3V9gedV+rjWngE8xP8/V2MMOF+7dXak//U2zLyDfx3sfX
cQfapGdhUFCe/By8iWaJHSieVSi5jZCYQ0PUw9MeuXjsDsNcu0zyM9nCdt8MelJU
R51hjmIAcnBTLF1WE5EDnP3f0OW58gVNB7yeGZhB8nFBxDazLGpOO8iMPoIPsM1k
B8TSJN5C9/zKqnPZJoKHck2HLhz66lYyNZbCsJX9+ukIpV7z75rJQru6POdGsoKK
nI0wKXHGR4py+K1yEPjFcJaXeMsKZo0kbLRcdW4HJs4Xk+/rFCh+YSF3l8c90m7G
2rFml8ijGJwhW/GCIWWRI3PO8Y4az32DkdIj3PuZ9e6ql27vt8v1xrmU2y9No9j3
diD2oNUJX533XrgefS1k86oiDjVQ1s3IHPm8/3gtFLw4gl6G6Dyc2riNCjCKzguc
kcb1hDmc+dbfV94QihKhi2PkGgBbptbK1EVo5M27ivKw6CSywZxfMEON/hoGILH7
iAktqfYInFBsRp6XKmAogo2xlpO3oYZw45GtH5aq/tb2tVxUXGZnrZEKeZFFGvo4
6X2QeuK8mwBMMwpWx2c65gDvxQ5t8slBXj9LgC2Q4DcU7peW7JWbtuE1X1lFoXAs
6q3S9ZMZkpbKaPH52xjMtyQthsyNnq6bKrja/sgkspf4XpUrlr7ccWWzHmCpmSxI
mLjJ+Fl8u7WLRPSaSjCy1bvhkHet9fDbFZCQu9TC2O61exOYOrWvixZxK+X1Z/W7
EsTY+CmYrbfTEOzuHS9bdCsZk1582X9mHpN92WOvyvVX0J7LW0Nulv3MImkHrOl8
yxF84ZOdXJFQeeenvMFJVGssVKS8yBnAugO2m9n874TwHeyDs/tFGb4ivPpoyU8O
Xo/yLBlAcmVyc0D+byDLsyyTglceWVLDb4byUPFt1E5P66RgJHj+roib9ATTYpOc
5gL+O24mnHt6ETKnUP/1lBC9Zg9nyTsk6J1vEcELV41qWGuEckgmplTNmBit8CIB
R1Z1b8E/JOk6r+MbrlzEVwbliW/g0Q3FVYNz1TF9eL4cdulDr88UqXxcWSS+HVFG
YeGs65pkH1Cv+WteQ8ti1C1TQOd1Q+9KB+GgXkv8zLym4AA4xtAw96eFnoKiVMga
AWxKOoaWlfcZ/3LOhHW+KrkBb+G+sr8Vu4Zof4e87UA9U4Oqf01pOjeoPsHaVJh1
bPZ3bFdI7KwXRzfWpRjWHDSqXiWmPxqTAGb2eBYVpx/4nQoF37B4SMfE5RosehsY
Dpu9Pu7aqOa8Qww3Fn0kWBR/ScEVPsVYdxhpAROhhpevqfsCwcG4IhzGvyO0ACBi
E2QluYw9nRiVbtoxZqbhshhgLz4vBeuFGAuBSbaHSWHnb7XCI18cJRMLpYx3qb/b
RqyAqFa0CDBKrMlKjSvpd+eIZ/rb8x/SF5e8Td6rbONOQ12z/b6wEQfit7nWZzUt
Mv5sg29jh1jeyCqtr7lEM7FkV6ndkkKloi5DCkYXEmsjDT4f586KB9XpOBw55pAb
LF355FFe+CIJoP+5N7RuVyB3D4jo8qXtzRXlzcyAw6YgA3dO5Uqc1/ZVJsTUsRW5
pz+A8+r1lwVq9P5RWDWa65M4p/WNVAugzzErmuR7cvo8ZOFhHGDSBCg4DGXajTND
78r5KI3uteWBcIyeEmcELsT+6+Th0vzl6khzlOtxXfjkYUuXU5rxzIw11iU8B9BR
GXSbNpbwYj0uPF3cDRvvtZU1sgfZb022BXctui0iOoaPzWODYbnqIjhc57VWAU6A
BMHlyPD2Hmka5SGcqD/Ln6MxncOz4z0fjuNsQJrduc1RQps6zuOhPMrPFMGFdskK
rwk2Ooa4n7LRvryteJJgw4eP0g5aigKpGh3ps5fbVLga/xKO4ciK5fegD0s9nNEf
O31n4Mi/3ZPD9Onv6neASf2utyEmn8xGVLHMk/5FIZOesjKKPdyg2y76VkDh5x7m
7oYtwrDlfC1rDQdVGX0bGTfNJL+VNIw82EOxnntOQvnUbVHbVKkiG4rG45BlY8aO
vEXqxEiGbPJ573Wxj1HpMDkJm3z/NMmP4lesw0rtZJfO5k+5vyxVkJpl8aphf9NH
HmhLjlC2wwY33s9mSAyu/TxmleCQCloAlEeHR5iiDtnaj4W/ShEAXMRAvGJ1SVJR
QR+8qcZyLsoKWN2V501HCA1RjbQXqnSBDU8ct7nnPm57iJMEtT2GErpetkbcnTd7
LfbLTUbeJsYQdCW38fCqzExn7TW/cASveJGo5plTA6uLAFlVDJA74YfyuPpfYams
KZbahvsHa4UQmhE2wrIjHnYdqJHJsrEUagnOUb3ohyEzNJzzoc40B3xwqW7RXF58
nXcosm/iOXCbXocxh9k9lAzM/3Kc5BV1C6DdubOI0cGMsM8cc0LeCkS3x1fRMxqy
/Fg/zrz9lMxIxUpGc8vHJR6zdc5r8i10rIfV6gVUgLAX9mcEfsSXspZ/QTL1nNgh
mI2dreyCGqlcpxeZ5NIe/8x+Xw+s1y7mrLqf1bSbO944hyLUNoKa6PeOnwgW8oXG
n9AiiHtJgqAZnC/k1mIfS/c2o26d0eX8frkvNNHENTB5bnlp49Ed/PirUSH7vdoA
xfYvPW6UwhcsIowswjwu55sPUCqSypG5PGcCa3Cq4ci3oCSBovtvCTJQowGClX2j
JIVhaUqhH3jUhPebgHJfasSY1SMLZ+TiZOuitcyF1l2zB77N4aSOeSVcjfgJ5pIA
ZYYrVfaC0BGe3o2SXeI2LypDIDUx5w3FTqY556el8jKSYXjifVyJ2V9vkICJ7Mz2
ulDEKPBml9wzwQ67z5Y9TU05fv5C4Aam/OyJS2CWjyROo+SJI1nrOAQ3hieetCps
ec5QN0D+LQBkd9mPMBDraTuSeioo3BD0dcguABvGUsh5MOvQSGd9dti7LCXFGTkQ
LO9zF5VqWZ9NFUpp9JqTJQt5/+xv5+hezMaHgWOnYCxUu5xCvZp2kBrwJ0o/9shB
1vY8CbGn24CuZmHZV8VJzlXQf2tqHNngTlLUBBzLB26rJVB1MmXzlz3nZ6A3gNNh
EXWP8dAXl9Mz1lhAHTiPfT75Qc7+P8K/2Lde3zH8OWWHdrEq31RUFJvltAlj32i/
1Mm/pxDH5EPhfUi0BQE70GJlsjuZj7HG1ztJM4C9tH1Y9zzRT27DBGdE+bjq7DK2
+x6PN/LcdOemgNvxAJvtLy8LI02zK3r7soUtkkjt0aJ4lw4qCCA66zEPmK0koBoC
pVWzT9L6+C/sCtH/3mdOVfnFKeWMtfa3m+f3opUKjdxZ/007bzFtfxk2neul0AdG
ZykgVeAV4UxsRgZYxZy3LP12FOMOl06/N7PijI/0EVnuobbSFHCYsQrNQIoI64hx
HvIJ+oN5eCB0qb43H2kDCTl35dAvm0lU0Yx9idch9gXVbT+p4cklTAcZUy11Q1x8
R727sprLUesqHlZwdL947J+RIrXDQZhefC4nVTL+cx4z7lNWp2D3dHng73tjKzvI
uk0CzNx9vP6AOSur7vjutapXfBh2dWmbAtLdegujIf+LOVAdsI2zw0lhV48rXLOQ
p6Omkdhiut1+2uYUXsw11Qt+NolR7yrxKBU9Z7K4lT2DMU8ky4DvdqObQmkrqYqA
SnVjaVvmnLyaHjD4vlPfCQz7OZoPvHab7brfrXn2tfzxv+qPn2qYFpOVl67rwk3Y
3MoOO6lRQRTYuE2lld9vrxzjhErQkL91m/QO7Hk4FINh+W5kC2thaGfyVptJW1pb
58jj1vO23xTz2wYXlcrmg2l3XPmBsJDj/r6QqRuWb59W+XCW4eM5VwgtHAwWDLge
z2m5yE5VPNNI1AZr/UD8jVMGVOn55MbdNzfO1m61Eqk5dauhPfPGneh916Rh96JD
An6Sa+KBXY6ZbVfZDcDqd96wfL8FF4SAOc8/sloJYswVZLakwBC3Bsz0TSfeVdTN
b9w44Om3CQB9jgO58sm8xHxx+ohnUhYTYV4sQRtNFr2BkPh5GrkSKDIg5lv8JwLF
SYv7u/f3hBrKj8HwgCUAa9T99vtNNux6MsfbEiieZEcB+AoMYkH5AGBVbCLhiH3f
hDx7edDafLsvB8yrned1QOI2iuxjZF6DMUT/zLVvWRtZmKpzAIzfNt6f5mzFKQHU
5MK94QPm9ybl2R95VBVrrDtUDCurVXgWcOwLQK77bz4VtgBR4zlHa5HKHumXIKp7
o3RpARm1WW8C0D4YF2lf5Y1Au0F0kcZsqkQ5g1W/KJg7NjMOL46O0vYC+ptsZ5D0
4l43QFc5apiHBh5hAgyJGL4OKOQ9SbOrwt3MAEbiOIBRLKEFbRi3ht7vVhn0dGVt
UG7PMBCO94vksB4uePqVxXvM8TAd/faal9vD3/qVjdIxF+smlndZnDbdZoL+9MfG
vZ6n9hhnhNutg3sdzySg0YawTLhA1oJTc06yUGXvhdm9Nyid/Hm2nw4qucQqr9Ni
stnx77LoVG1sIK4Bx1rKqtdoLApXaniSXYVAWdxbMkHOd3FaY7DGi6GWAKMpeUEG
xu8oE2Fu8Zi4QU+5YVWwI41MYYHgYQgB571oxU+BUbiazEWIbqDVHsFA4CFeImwU
USW82JvoAGusS1pv4IlrobpK0n94j5bfceDzFE3EeRZ8Dw3okJvWqV2LoODbXGmH
XBnK9qk4ZvlIHoCNCTMRPDv4aFjDRfLCIHnVvSKWAhVIHAv3MQSgAxgLTcGqmn0M
LErl7ZHyzzqES7htkZNowvd0pfIWFpnV/FGqoGHTDoxt78E81qdlkGgNF8y237pm
xFfJrF8O+9lkHmUdb7pSUIZHr1m1aLmkBT267jTDL0qD23FSLX4BtZHvxQLPgJE9
Qj13FqZ8V9zAvHwoP4+yAmK5nYG/RqS16AVhWRcC49EpVwLbyTCytALxX5tTK3kr
Hs/RGx2KK7SQalzQTjVgSMfGgQnpv4zYwS58AxCoVYc699rFKOO4cNBq/RrzI/WZ
sspW+ZtrZL+ijcbvEg5XRZcGRukLwxXTwlNEwOSY8J3ydqgRpdjPguAf6hO5iWQ3
FH5/AoQn2PLaUIOoqeIxcF6n5vArmK5bbmrtgbj0ncyL9CBBeUIzVcVemyWZtF7q
guOXyymzkMmOKWg6BkPuYrh+IaHH6yYf08M7SR04dV2A5by70fOdemIzlULDQ3SY
NQSIeOHQutHZUV+pZ/W9szumJtbLKjPqRVGoJ/vyMQs/jeZSzAa5fZrxPkuO7ywp
Q0jK/aE8aFRQdDeRCdh2o8HpE1IgnUrGJFJZVp4vjqC5Jwg6LXQjg0se9bcRTNsU
SO+crGa0aBTqLL3hMl0J/0MXQX33B0boh+9chpKVu/ifFme0d9Y2wAHHeZBSzIXP
YdnK/lTa634L9y7vG0ERaF8RCFCWIsl7l8PZXDchdm/B7XFwiFv9MJ0/szcdBAyA
0TMEl7WQriAc7WLRAMAGd/zeXpPzQqw2+8gFIpXyrMxpBiTp7a8gQw5u7lg3xJ+B
EIVu/Kcua5QWk8aZ/mlnwQD2ROK50PRIAp0lJFneYd0qDLrgdUySaefwO+woRfRP
OPtWOL8x/2bYJq5FeVf6fOvwpZXKSa8i/h8Ign8JhFetSnxU7mws38lO7lNmFnxn
LrJTzyb4bQu3rQ9rUPWWUHTUrnh9SyLTxAca3Aw8tEHVXEltjDUT2XlhOZHxgTJH
3PelHvIQCgIeLFJ4HYa+X0ujC2pj6Ka6xc8IzpV0Ffv8ZpCo9qQOaBqcgfUjJJdg
9RgpTmlV/S5tnYZ8jsx/oD+qyVNXMNoD/hRCD2vadDeNHrQ2p8d6z7X2k1cBR2wm
SDxzw7uoCJS2IIOlcsJATbfzzmaMsZeFG/SGbxJLYIRSwwzScvwQGmCrfEAPFlqH
ynjbuqUOauFsrmh736gcq5K6hxljqGrXrSdZ1tK8j3cThYD7hANIjM0baUzecFW3
Lg+iJTAoOKr1TguatKNh1lkoj7lV7kMZKBnSB/0vpdN6fzs/1uJw9iefzpPz4yXD
n0UD0sq2GT1+5xyIF2JlAe2fRjqOFFWcu53+EgRS0AP68vgu80rVfMXZrTmGdhKn
cC8fkjssrubGgCIkNlJ4ClMUuVS6UkmhCRdMQeSW72ZT9RNBytHvHOQhgfTDMsqy
gTQ1u05L9vvIQDR+ZrS61FbWQkmUNY3kdNtGhVLGlgzgsnVVSVlpabnkYV/l5Nk5
Egj5NCtdhv+opLzcyYRhq/dk8m/ZzsYkDwiXLbgH8GbCZZ7YDEB3CmvrMc3jmkeK
xwRIx82xJ7X7tLyKU7iw5GrlrnnT6qUSh0p/JuGFFXQYopdwn7qKKTbH/L6GeavH
+b8drf7MO4V5CDY6sk2NZjafdW9CbTjYj95Vr2HoIi0eC2eewXOE2gYjLUraKC2K
VWrGp3J4thW5sLmVsU13Yjz2jbOWtN0uBLZ2zU9sT80Mb/NFjiZQQAr4R0ak9eYx
d08QCm+i+34EFWN/pnNr2Sq6GTgE68EHqj8o2TCqtr0LEpMtbk3tqBNKz5HPVLNs
cdCM3zy582NECWxUwSvrJJH/q6TUmlUkMRhAlKlsmMTBHcEybJCVxh6CYkpPcoB+
Fo0Vb1myRMwQVNLnuQDvAVN+k6KnxFEE6e5m1tiP99/V6feyR47WZ32ni7LxLYa9
DWE8EO3HtrcOwuIyNQHBoLiAOaopdpPAOEVh4H0WYDrpjBQNnbPo6Vq1rwsNhj5z
kvYzuV+C1FY7c+f8Tv7fdc4Fk+0vmvgTrkHjFxrKNJAVr5KIuZbo37BS1H/+1A3R
R9X7eclJ1MT4lkl+aIx9oarQFcn98lAh96FcUfvAAeXSTpuXPJ7m8HjQebng0Res
rFRwc0xGaosgtwwEZEDnMrgzdM2jpDzS8R223dgh64wpZmNfYsjtKgXvbgqjNaKz
vNhoClrv+oNwD+XjS3UcDXy/HtBTsicgxpsqBrZ8WU5tQcv8cJwECo12Nwd4KcoR
MiT7pZ7l3LbvcGl/W9hPPz237FsyR/BmecuHNrcow4JIef0CK0wBBLKeVU4F8z55
nU9I36hNTSDjDBxCof5N7i2dPnOjHrN+RKW58JJmagqZFgUsbqKTTa6N2G7xk83+
RDncz5ljw6FALOTkkdGychWVs5apZNrO7cXbACMUwHqwrE6m2nzxS+6r760R0pZX
WpNo8B2Uq4EePy/P93T3zkmKz+LrWTYYWE+J8YDSjjOQ4FBsuW6L1XIngHq8FpZZ
bOS6OjWa64P0i4v7izzeWk4B3Yp89wj97y8sUSdV+UhMi/zMtaQyBtVS12n4TmTE
nTLMCfbY76T18d93n+4/e1OzmEnemhuAPFIGWvCgrfznuwA+hxdnHUURs5mZJqa5
3C042d5MO4V42AMhz93i84EwCQCMuZJzpmFx0EdsfIm9BRgKehAHN27xVFmsd9y8
r++hLdoFPioodE5zWZf3+TzvxxKp2dqrOLCZ2u5FW8/v3WrnuqS4NKubAXlkYy7n
KWoONoOX+ppQCccgK+NRuhI4nmXVmdPl7gVVkCOuDkPGYr8B/cwWsO+a0AwDY0oe
jbNI0G0tyaMl7Le8l1tiW6936oAvGmKvWr+7ScbHfTbLZUmWClPmhFDB+U9Hc4ez
BCcfiI79w5sXl2D/aqmjOl8hudQAbppuJMXQXOPpwQaN/yub8a8n7Hk5/pYnqolr
ujPdOg/9Jhe0mzCQ7YMfWhjg7lqs4F4HypcjzxKAUjHQK3JZ68KaY1SnAbxtqET8
63XkytrtXXDEoFBevSPrO3z7ZPToj1RFiEpnkfKDAETKHIxgIzoVwJXF5B/VX1FK
eYGmTkqH5JYn0EDvjuLbZAri9dxfNqqcZ6josgvO818tG5wKuaAi8xuXN8lzYxI6
57TYGZYSymRMlOfqHfb8sgw0ljSq2xlcpYsHZAS8rDj3ZNd7epkfg6BNuajHovfo
T2/IdZ+kDUmSO0sunZwGKT3eVmfnI/CF6sUGE8WAxrGFsHmJaowIiK2f1gNre0+r
b3piece8Ep4mRb+BbLPWjueJZPm8z8VICtVSwGyGepaGKwoXAdrWUpGpBxcZDk+D
C4ct7bRLASutS5aW5LDvU9A8Uv3YEmnlYsmD0QXuFyuJKQDjSxIZTeWD5qusKhzp
e109eRbEM1rxhy31Dpx65QBIqlO+JcieDCmBUz63oXWJMm1TcnirCsuZHGBJRZ4h
0YvIbrUzFsjbN9JnxtWdsrrVrxkX0DL8G0b/h6X/A7qqqG7N82ydLLhFdNit417T
D03onxL7xwfFabI/dgodN7zO8KuXvMTo/Re55qX6s6ZYpQG2A6XQlwfppjqT3u0p
kiFnEUIPOM+wnHIZYbjV4jO3qyB+rdPvMLv+DcPS86ta1IBWdchsI9Rnw4Nd8oXi
Jgn+TXcxU7GXwHO3ej56NySE1MxK9hqB60QXxQXsEMkH7LBFBr3h+Xo6fQCzzjnf
uanhJpT6smfdJb/jaFStRjonK2vJ59EmlBmb5nSTMKYAzA09/TMfl8VSYqJtEwO6
bvGWUZMrX9V+si4LvVKj/N1kU7eub6HPw6aeF7wdmBhlDvCrhLSP0FY0WX5ElWh7
U2YXyKBehs/ip8tNZkR3V+/S+oPyXcnjgjDGd6skZVaVgv4Lom33CfMJbU329a/k
3mSpPHib2p3jBWgDa5lxvLYeTHdYZV0AQTm1o5mWPHiRRolwJN0/YQ27WCs3Gtnz
2e+1XzuY0hYpFoHhdLgo0xzz0rpvmVoR0NM5N6ii2PNOfs8LHnEj/iFtaLCexxt8
VuNIc1CrFKdXgY3m3pa3p3rN5WB4ycoGlDo9oNmC2rrRL2aMahuZl51ovLXKzVmj
iLgpqsEOI+XIJ9lEqJDXRh4kXhdIIWtLdpSJcmCjHeuBrI1ZErZTWnBzh3FGM1tI
Cq7MM/N/WyuOdfuEfiPkGGgXNWwCrS4/9VHpsODVthSUdipETTuBpbkNvoiKUCEw
PB5dHIp/0LBnYBBDkIIWUCIh7vYIgDk91lq/kqCgKukQvQVhHO4b9hBBvANsWPfP
mS/7pTfLTMpXXg64BlC7f4yQ6KPnkDpLUuGCIPlHTBByOD7ITFL8fGtvDlnulnqw
icXNYFfa7bt4ld1gSny3vZr6woEFrd8Q9dl9c5r37VFojULpeFrGbRaMwCcLoX/X
OSZLAEhhUJemHpJjuNcHFFmoMjb1WLSDwqGeWIl3vT7vjk+4nSY/IvbInaeSU+/w
Uw8pDqMSf54H/3WGhwE0/dcEs9KYCf6almciHqJBNmGeIPsDu65Ezjngjzc1up3g
hkAjhAjv+qMxY/SNXxSkmHMvQFb01lj1PaPV/FKwLQL3peIo3QaI7PPgLOoqp8AV
Mpu1snXBN6YHwZxxA6X9UMvstvWrBa3cTHECo/zV9Dc2aHNoID3GlmKOC8MTVlEe
xM/UZ0mgfxlDmv0h2JsEw0Q0FSlX3bdNtk91vCObNI8m7dHkZWukLwLN9FuhAJwU
yZUqtnWGlafrcV+vOaXA+epqlkWVOsXpYDOPzo4CzZN5emCKqex4xPwMg8w/BlbU
+StYiU0Y63RvA2DHX3OmEEfZihu3lBKo8zMaBpKXEKGX2ylRDGlWreboJaOwxJsN
an9s3lN3V9HC3v/mXSYIU7W7QxRMoE0oLQc5by/8JHG5e0pZZH3zFsUXXWR1WxPT
VVeYhwrp+MHIAgkyhbOfh8KcXLCTo6lIKOaIxOcHTYzR1rilfDM4k4BQDmAb21Xn
umdc3V8i/EYzaLptxh6/2f4s3MGtPNHfC1bW1J245NosxbbwsKgTP+a/d0SXwJPP
RwVkq8Wd5AanZcrPNjinxP0bbDoany5RygLBYDWN6QrEVVgY6y/zCISaQCWmb4Ec
mTIJWU/fQ8r+FK7FCtHD0y8RS7eCWdY2HF7TXrPw8ZVDF8FAFNggoOWGtcNob1I5
WitZpN4gZYtgpes1js7GypDurW9obnqjAHveP5Ceqt11Rgm6ZLBPMN+nFLBLBrFu
X/PD+FoofbvyeZRKDduiAdH11E5LMwT7GQUampHWxdy63ZovYXQ4o4BvH4oKwk4U
W6MEQWgfiVcnkEUN86edVRNHFrkwyChcKssxXypzfO9JfKZ+bNSHzQJtUDbCakjD
WK1vzG93bW3rilnh5hlk6bkhwhWtt69AoZZGCmM0/kZytafTAd0X+TTQwhae0HJb
fLRbFL/H/qF3zz6UcUpE8v7+haRnTM9MmD2IcKApt0TaxjcFgYnFrQSMPz36RTat
NyvoIAJ5ZhWPfX3+jsLCNc+57tZoggl9sdk6vdbgWSRVmBU+FSpWVl0izpHNxmUv
yF8UUzVt8Tyw3NuVRlH6cQKPY2Mi1SRp4Hn8hOrA19JfeGORmgDApfdZN2Tc6dLQ
7davX2yKHrdSgURhjbqIISNMrC2CVLGXAXRlJniAvQTZTbGWoxY4gzeiI5wtFPZ5
kU2nCcYjNjPQ5N7Rd9HxQl0ImOA2amcy9U+e981R5hk7vZ3kpGzoVCZPTMK9Y0C3
qf9tDj54owoepx5nyrblyKhYgnaFKQeYKMvKgZBT2gweqdYWVr3Y+VrT5dTDDhCo
sy2bpFn5ltw+weh6df9JtFr5HGgCcJXxVcRD/ofNpNlFDlKbuTEkLkgIX/cDRXr0
vFiekwmA1ax7744A5vnhiS501XTSNtGrkMhp7jaH88IFHangpZA2pF9tuDPRHnuh
CGPrWSx2lypSeB21TW8AAtXSc3vRMonSOjsAGFSW7ZuwmfoEhKPvGGcyeqhSgP3B
/ic14mczo45fl6n/1etKEnyl53Vn2XAyRP4MTXZqufqbZ1kEVOI1fsxIPybycw+s
SpU+I32Qf0oshOth3dMlpNLR1Xd+Pwy61szopgnCT9OjBKMVO1RSAbov4mAVzGGm
8qADQWL81mtPd6Sz6uJ4Xqzv6hpYeD2YiLnsKC/MtbznU7QHtskovxhaHPXXH/zD
iUSqYUKfwJqIvNB17+z6egI0XzJnqhgv2y5IuzEGBZzxOaLQnCwL0jPe1hUeyF9G
m6j8Lchm1uckEjay0EkTbGV/RXDu6CfvjbeS2raunSLFqVkdCGlBJy1BWuaMmOy3
QHgt+zi6vr6S0UxCQa6fudiIe5sum34ND5Cn0Ou8v2BUjvGvZLuPTfLmlKEyKRXG
+rNRRtMdWN676w5Q1+H6YS6K7mITBH417TDmHgdHXPutPNZczZ6mId1JqljvYkJA
6dg3dELknY97N3Hn4diA71qEQU/XFOLB9AfYAiMuxYRg4HrVOrT3TGc5sQlkrhKr
79qZyij1lyDKm4ZEXjgAxDVHsHZ+O8CI77oVAV04sEoLXpPuK8j5YLDc+iFvNtKt
/WTUjy6NO8tNMK+MXjWTCmoIhqYS4Bvtcx9UadWGKpmYDrE4fP2GgyOK2DrPwIB+
j/sPZjIfJGV754QVIrW5xzcbN+h6K+ZlIBal0Vzbq/iQ9ORf13aaXP89/gJI86Zu
BeARFao6oCFIxU4Ssf6CypAlt+ftUQhCVbKwryKJ6c4d6e5mcFJhVjHaoZEAK3aE
SehPSZ5Q+CctImV8NcLyZHqg2e78UiyDQnVT20KXd2Tdn783e/Qm8T02xQHHcp0Q
n903VOjVwUE3eYdl2GjqaeaY+qgp0WiWjp6fmLvsc6efMLmjuQGcL/2n8sQoY7I4
8XZZCx4TMMkQHDePmotl0BXDhjqpn5bvoOz3YhzLjHItGDnhl1MP9PfWVXA0FXdk
y/VDVsBws4QupqcRv/DtpXPveZlPDJGe5nE2dfds5qGjzd/Nea0sEuEJaAD4M2T0
rWSgywORgQJWyVPEHpdaFTWIfMa30Kla/42Sr9O/KjIbFmcIQr//hp1/S1ZYQTCR
NWlMXNiw59ZiAkApViC18cCHVx2/XpKb0jga8iqBiC/Av63oVf9aLDA/l8E0gUfa
3fvuNoHly4QdzReLzeZjOVY+V0eBCSw8lqiUKWy3c4Xqvn/5tqHpj6jECibj2aDN
WiJIBSIWNRDZ8V3v4Ny9hi5NbdVAVMQvpZ3eHyjWJuSMZQDqn2g4QAngj0z/9ALN
MmjR0FY3oxoYvZpQ7FJfUEnLYO1AI+yg4OXkD+9lOzEzhyTRSuV3GHLxjWhemyOs
R40mLrkNUqCTJOdCiIjqD5c5iKIkzOSkSsw4C2Hg48CZKperoOOYE7ayYykVd0fs
GOOdmOtVNiFSE510lH4n1+2afnh4ldVDiOLj77pGxWCDAG9ZNYYUjS70818nhy41
wWUZ7qxoMX5nrIok7eoAFLAzBFHDal0Fav7RR7hWuhAsqnp0fZhrBv5RnfZOmTC0
VSJCianYb7wvDUVPzA47vkWGLQyG7xVm60vMB6deKEgB1iRXs7NvaR2jDpv/S3da
IUzfXebtfvVf9lIOzd+JNoIBsG94l1kLHm3MRbACCIvUroWL1mzs7qQSaddxFgRy
b+pf7HSkclcjzdxEc5Z7UGQPCdHYsQ1N2wwJY3C7ECta34TkPsqYrYmOHwLz3Lkp
tPSIWsYgTBReckeP5kX7YZ7S20HhVJ5Cucih7XYNXv4CdoBHbCnLr4If1pdE+l/W
ORSedGJ/Lpcyyf/WNgQhzoSaq2cwyozIdol1YXkmfzK0+0DdasdIbg+FMYpC+xG6
VogGCVWpgyTsgY7ylWqlCKMiTcMD5+Rpb4NLACSJSgQljaVuiS5GMTK/x+0dh59q
EqJrwpcPRUmjSfbDWlWdkX24N+TIS4VMdDlIcrPEaquwsJQ+fIK4l/07Qug2wFib
K3/HkFdCaOxsPLfTiw5I71aiGgrWspJ3eouo69gHRbR7/MYliKgexX2oA5p3ydzt
+zvIfahxvNSAwyWqRbyV6KWOtNe7VEhzr6hAPSronzneqeERHhwNytzunlegbUCq
qL2V1RAlzswr7kDeowjkLS5e4hvP1I5XYw2fnvz6dPB9pAz/CVaxkyXwGZKbyHun
TO7S8J7FseLMtY6I9Wj1MRL+ipiq58CWvd/KFl+jo0zwI2ksRJbwd74B0jjc/TLi
3HbRRCF1YgmD3iHQbe7Db2ZrAQRjBTa1HwcbB+rAK/TO9xsHOQauyUNZtsFDdiVC
yPk5SVJEJpsq4Es/2ExcCobogB0lkRQ28IbaaQcGijSmC1CHkUKyyh4YJ+6geHXv
1XlG2UlDJXg4VMfZb0+WLtlc12DutbPe7zghqaUDj/dynuCSt6f0bKxctClXnqgv
Rd4aT+QaqEGt8RVWgCpCzVTs27Q7Eg63PxqlzOxIk7x6EknSYS2cp0DQS087KIgQ
DT0wcUERY1ZaOVsbI1XB1oeErFzcyAt8C+eTB+7U5uRSLPAnjMKh6+zgwXtXUBUQ
0wREyxLGDhWbOc7xuP+p4RJpAUCIkVvrc1r4R/FDHVbIE0kCQg6krKNOeFA32K25
5DEXDI9WdPqXo7QcL1qtrNloiDZ0Ru+9HSQglx4ZipvjZqRI7T9V4iV+xtLcRpKh
SiIW6PlHz2dwqjlRg6KYzVDPGyYBkildwN5m1dZxEla44fihhQQuK22+2pD6wNaK
z4MS2D8JvGp2ITmS1xId0iUwolqfYohXeMFeArRKJZq1Oo2FkUlWqPRGTxvKnzD/
nEKWXEv8IfQq/+r3/6LmE8OyMF0LUk2tgQXIIlCecsJ4n3gO57KYOE/F4BvN2cpK
LOmx6cUHxH6ECl7KwN4eySKAAZ3n5etXGQkS/EmFhRkm4TArHXKd/lduLQj0utEi
zNIi8ZzyUFkhXSdTPGkQzwuE0zwLR9ndr8ssaU4jPph7AnJ5Mk6uQ7mYmdXTkQja
N/okTKcbyFYJQKmlyywqUY18Ct8WZYU0h1M/z7g+CjnTdvL+V/x84oXPWmlmQxa4
e9cPuWA1ASQoVp3TNWOBYADJDYHZwpgZRVn9GusEBXWwWpTyGrObw3RQPbiOs4aI
C3YokjsMlcuyN6CI8VY7Smixtm/D2N/1nzKjs0kBnRTUqJQF13zTUBSniR7Uuds6
If8tXScTPz9tfG28ZYVi+F7NwRT3L1Ba+MJ82q6dG+0vzljYE0F7ENa9okPdHAFk
CP3EQdEHjtPJZIeug6VY1aEfpIyVbW2qezZCtcoG2MK0t9TyyABWea2UljO2QqSQ
paru4Ve1/dshc0htB9h9rYCPcB7usK8K7kQcq1dcuyZYHDtoRAYMwpZlS3BnHyqB
vHp2/XpiZst2ffda8EcORcYvvpv3pj+ldlsw0yAAbQqrTmOh5avkKXxEfQmPZyE+
GsguXKPIF9k9s7fn//9YLKRGbYvDI4E4KH4CQ1vcZKm6XXI2qVurxcOaw1o0ztUx
hciZGS5FMOmeaOeY94+Hjh4IxweNbsUT7RjMJDikdzjh4pJRfppOgkEu6/gj+I53
v1GqcMsZn3TRUiTI4T/GeJvWxB1Vc6VCUigsEtfVt4dS8qudEYHZB0Dk9fHs8EOb
Kt7fTdPenxL1pfeCJiHTqSiVfZJrZAD19vaSDgLfR1+HlPqMR0D+uweR/MMSW/1e
GqRzD5FiLWWUbYmOX7sFx4zX+JJLKmgFvlDmqjbwOv7qeUR5PBQRXt2wExG610ZS
UbD5WPCjmSEW+29bS0g0I/OXk7l6h/gpKJd6wUXa+NyQJZdVmW/G19aZaJQezRqE
Lkd61WyunC9ha+LiX4ivlKXBYAkq16vrnxAOxX5OqJKRTyXiJwhySvAj4dimwtKb
k6A98f3sh4UbeU4DNZ6NjqPEx8b55wF2YmCShpysUWFV1qSeXHeiea3WV+Yiwfbm
gRs2FlhLCfsTi4qamURCn1fuPtQcGKhx3jp3HdN2UpJASs7R/SSNgYT5n21suamG
vNfp28QOaVw1ilUwFe/BRpm5wLsmspGZWpaUlWWHV3Mutj6RI0EtgzbeN/LJ9l8G
FlQ50JZ57+y16AXB0WKKDnSCmmx13O1/f17Z3UyhOtD0dXpOURFafMdxfGsBdkbE
1kPfjoF6//s21HhfhaBCi+E/8c42YZkVMuI+58DwZSwLgbRgoIvOdxFpgmjDcBs9
X6oZAl5gDXBJMqAD3YM/hiwKfdRvMEQJ2gNEx8MsZWNgV8Az72YC38prz9dcB0RE
7+CTLqfs91cf78fBSJvfi0JXtKdYkYacCogerprSovXu9FLK7kXNAnuWt7JbwV2A
7zUETBIJo6uPr9RcEtwhzMUPFz1AU16cNMAo5NmTBCb69Xntxhn7FO2pqDRgv1kU
k6DIlyU8o7UuMqbvLDWdyozuN6iOEc6z2jrQcggUug7hLgiyYbHpMXSGpuJtt8+H
9p95QWeZOlA2NS4Z/pdhGkq/QVOz5lGpubPeNh9p744T9++G/G+2fc0k3QGOSXU+
0JIGmp7MQncc9ISSMHJQNc/nIycVzg3th7d4/Ht9j9IvB4xDNTSra+j5bxXQ7UV6
znSsCcqwmaxeojf8sWPyGGncsLAE+kJLmvYnmo8ydDuEvvCwx0cFnMaxzuKE41qa
fptD6r1KQJegwHbRW41Dny2kIgHA7g51gN1mKmw/QUtlRYnERO6R5/ccaMWgP1MM
8XkY2Qj0dPse/dllqQ8TvwOuKk6zE18PPxk6UWvneKBARRYZOFp9Q6NEYrLGP/BH
HKfHhvLHVDHCKGsSGcu/Al8U/l00i4C9z0iyuxY0lWvy63McHFZnNULV2h6lnB8b
yQ8lcWzSKkwBvAqQVpnptCFk97K16oOUCzk9ozpH1JCwp+NtWh/ewqrMu8piFmP1
yv/bdzF94gUJwr+EdpM3sZz2T3bt6p6fmSerMZKkkb/MGezMe7SkJqcEsXy3BPwl
RqxyZ5lUOO/5mJAGJR5SSF+BznEBWEFcGuQyOXbnyzUF+t7r7z2Ajv0jbYDahvm7
/ogAeaE+svRkNQMpbo5WxEWLDqXzuqLs76AhcySZ6qyRYOA+oGcYVOiB49bcWcna
pLlYl01UmbLB8GT/YhGHmnCkJ2ai8y6Wo8gYqDUdo9BMFXqT3jLnYxTUDQfT+Fce
d039uSM+LLi3nheH5hLK4D3rZ7EckDXtXBXzSUiMkTkC13wgWJR3YtIoOgPnPvNT
eg7VTZvaPqlSOve7yvyClrnkYkz5VTfIJy7IbpxiEYIz4q01q3o6kuaJxgg9W/oW
14L9E7X+HhZ8trolXLU4trDGbVdujo4Y5cw1v+ON6d7O6NabnkdLa5F1XoY1soF6
8r2caJjbHASxAYqZqlAt3yf5rV9ZcAruf3u9TMv+zdll5NDgo13qvU1U4HT4WZ8i
G8RxSCqS2g0qYWZL9b90QoNdiKsyUqRes5jlpG6OFFCHBrKQ5dv3MafTN+FqiY/l
bRvIeMAhhPkRaMiOBZZEe96KStVeEYS0z6npDB/NXHgaDDmTAi2RT0cXQck/AgrZ
2AqgjtdvrQVxclhcjanWIeSqWezL2s/bLbCgiselnRAj7wpNKO7JeOGiMEWcpFsA
+FELGWx6fggC2VsoFF+MtrV9/qFC75NG4SRQC/iYsNX3KmX/Y53ZDbDP6h2fi4TQ
CqPOrdUmRIwBhUEs4CVWUuLNYlvEL8gFv2M8/kOLwCGXfYJKcyVg9obIolHrKliT
wHS/UcbiDaL77nzeZpdJwmzjXVgc8mPMIp7gs5FUcQO0uhfwymadg895TShUfMHv
eqoSNGQdg4PkjtEMeW+Ds6s3m1v5/fH9UrJl7BoQsSwLFdTI2LT0SZomq5upV1AL
MdbrLiBcNtvOsVy8t5l9Ol87CebhoMTmrKum4XunxOO8vK3OLEGyOXjKqiwWDB6T
re5MI5n/ausSKgbiscwAKYl0gGwHoCLaV4EG5t4cZK9C3sa0qBzHtwJmXoX9rs+X
6pAS9d96t9rlerug8gvz+qZA4Fmc/mlnvpnLm5Kj2orbEVk14gC7Scv/foaaVDhD
IGxlYHVPRj2I+QSlBo1raO7GE+njp14Je18w6v3e90R0mbGxkahtH8E/IYaX08f8
Wu0tJWs+Glw7DnhS2oIuKTyelP2N5e+E9iWjSl4NV7Z9q9bat4umIjZtrApqDaRH
Uqgb9/Ck0e118Mbp7ODm4f1cWpiLxHdbKAWeMJ9dVnvDrMBYOBMPPYajHzGz6R+B
8k50TCVZJrLV4N0bwmxbzjCjiauNUfuTDlbMMTupmElOpue92WThMaByGXUuPKXW
Vl99nK5+JYfjtWxWTQrbhwWp3nLZ5zmT+otpvyfmbf/Z0ReRXiDr/DF6BcZ52ivq
tMUeiNxzG/hm0ZqOOiYg9wM/qjMZYdC+sEBpNmQJz7cfCGMoeeGwce/skV5VlR3L
++H87zEUdEbGdxbeCPmp7JgQ/RDSkmseg3/he1/SD6mPz8oi0wAWGEJHIEqBf3zI
EkukbXYMcE1Rx4fVWZYhJUkyIAopLrKX/fgxN8h8rq6i3B017SMt+yWa3DDE5w+Z
tR331D01DOtLY/+4GZ0COOdTFavn6BeBrGhK1IRTDWfri3MAWvFsswGxpw+fHv6s
KStA6Zm9LBOKEFDwRnEo8BeFhpM/Fac2ofFJoO19UVpBbKx1esO5rupoYHs2h5GO
J8dZUI9ef2AfbZvhMBm1iDEqESPSBIAMozCPawyJgAnTICVZ1rRPUSI3f2qxbKP9
9AKjzWEAgzQl88+8LLySNUHWo3JaOTrRK716cHTjn1Qh1oYME/obK1U0dGqfBG2e
DPZ4s5FGB3g0vaONimFNSZjoAh11MA+r6pUKS6uOJ+t3UtcoyfdrEFy7lBZmBwC0
bgdPkcknU2m4EntYimY4E8RtJ8hD88SuZyYWbapSRSkVAXUxj9qCSEZtcACvYb/p
/3oiH3W6mblIv2hSX/PmLdCtuXmj8lXy86dbOLrHMv+ed+P0q12pe2dK1SK+cLnZ
kIK/YDXT3iguX/SH34BVr17n+1o1dvyzul7wUVXEQwMadMsvjxqbnrjZPxyKthAC
5mlgwhhDrEooNIu5DAuUds1MqTVrpThjocHmVA96MRUpUFuP0sH7AtkhBFUW8qk9
mc3+TsKfxiPRAYTm2Du6U7Cv6OoZ13C/ke8euQWiE0ScfF64YFGrvv+YSh8jvgJ2
yN6tFW1H1wdJOoiN5o5DSkEubz6/aEq8XclgLHmBYmnWqJYReQxN9RNhy2yKjl5D
BiA/8rThQtgcNyQ/QtZo2iM/0piib+dTFYBGZo7747hi+JspH/M0EEhn9aoZlLbM
F61JN9HqR8KX6CmSi5yjsmFRJNSIMvrr73nOlcLRrm/Nia3IJF8hZ7bZlXvPzRJt
ixs234Q58wtjKa5dpw3vo92MvKiuqFT2FnGaMbVDdrp7/b9EftmjPDrLAAHOeSLF
a+j5w9QqgqOina6A93sdXby/+q+3tS5O2Lgq8l+zIn0OQuqKrvCWsohTtiXMT6P3
tmY8XzytuMS3jJEt/EVQc8YBb44GpSS/u2wfexO40yzq6cTAvULSifkqiaTMinLF
Fp5d0kAKReH5M7b1GZuTu07qDQUpkSyLim3gs6ZCtrek4P11J6nn3sxy49R1XjIn
eDPsHqeSRaX4J66VDl33p3SmZx8Wwa6h5/Ip28WJpUFd3LRlNS6XCIxpx6AYdgQS
JwVTv81yRzvKCNvDefeFrBe9kCm30bgAqzA2pVK5C+GgFeykhf/gXlLEFz04P+l0
7nqDTFCD25f16BNwN8cCl2Mtp4cSfGFc0w99qhhSeoSxGX72nLgb2eSu7DTvL7vI
aNZb1ZB933bxs5z7t9P5TZS31Yn1xeARAd+kMaaNpyGdGujueT0ZR2eMN4nPGHyZ
y8G+I1uOPhaDgh0rCK8wc5vn7WH1FD3q8rSBF2buK3mrndhWLD1yzg07eh0nclFo
07NLUcC3WRY3Gwq/1SuKp//evBkX/ayTCsX006l5DIph+IH046peynK194vgE3F/
LHXpA77HdlrYMQSJCQJ9BFq6fxLs2unCA4Zul8v39/RYwo+cBPxDb/P89yiV9pdA
dRc/kIC0yYALm5L9tf+0yZwbNJcHrbjzpnpaiwqdCQaMFXG71yFPAdqTGlFLBdhN
mvDfrZMfca1Olfh6fEaSzqEAwf2bQFSLvsoVWbZR3BkvVrU0zaWgiHSKYfTwIFd3
d2ouWnXFUxIWUyNwh7iuFG6PjuzM1/AQm1IJJRwI5ddFxkixVtxIEgXTJG4k41yF
OOdHL37NQvPNu92Qsc0wb2fq1x9NjnecDJ2nAacJIWR1d4gP01Hy8GuKRupboECd
bO1soGT+s7oRwmdcch2VpxtQ/CQeswc8jOIamqLjXleeU4Dpw4t9dzzWJU2pYziW
61Hlw7QJwzctidx/LaLrjn44Cq1p0TxgJsuA+dxCstzd+3muWMeIuvkDnLlr/2T1
eUWMNDpPkPr60mlgdMa2v5eiG1Jq0TwUjFgjCMXJQFK9BQ0Vj7KsCScpUTV5c8yG
EA94s0RJiKPVLOJkzW5O/Y9QIr4xvuk+y8LhadPLeO51waYO7BZf+Y3OybB+7SX1
ef9Ra35s8I23Ud6cNLNWqNaHuARv6OkoRT7QuRbQnWHfvLPoYpYNPKTCwjk+nzRo
dhZE3QMlx47XXXPSi1QDQ5IPDyAuZzQgJNHtvoLVUGhUnnQDpJ3hnverQni758we
dkSg9OiiWrsrVUeRFjwX9SVUhtggZHtli3SMIxNWP3z8T0wVq7h+hGeXK5wTbMbl
pPUdMD/BTMF92Mji+ZdMzJnpEDDHY+BIQ8qiMZ7yZvFMpHKkUgSt1ZwVH4DopOEG
6u1g4pOBdTTRSdisQbCXJhgdICB29EWteQPYGmjcj/yTtMRUpIoJQjEDUKapsE24
bTRnC7YEXqCgDMMz0ngSEdCfAxelOAKifAKNK5MmoH9e+3Vpz55Od1oNLGa2LFHu
9zmbySoHn7ht9+PshuAZrJE0rHVeR96ErV9NAlJkZnGfboBUJGeDn4bIF+t4MzVd
1ijhjXFBez5zmiav8fcE/PIgQ7yxj/c+oNpftiv9S1lCeyggwrA/650ziWCYgMtY
Zzg9AJQW2x+FGZNbxrROSXNzbFA2dsYVga/9yepQ5bcKrdW1XR6qwO3mf1vVXrGP
dc7lAlD6sBUaSf53yoPmUzgjqNSpwj8qRjG6QJW81WHC9d428N8nVuHFDjr4PHSc
0c+slButvnLKk2RDt85b0ZLPiJbLZSjeU5F/8OiIbmDFMtHnSXZFStDu+JUI4DGO
5fwTdoQKtMjB9lfR1P2+HxAqRKfjsPrJPcMhKDsoR8w5JXv8t7x5bAlBsoY8wFVx
ZjmbbSopl5omi+JR40vGOnidfwfYne0DUGGoDo/ydO7OamCwoHn+56vGKCg3xHqn
29+iTf+Ulnh86AtnQKw9cqXgeNgUKuUaCcOev/I/+T5C2u7/pFCR0iX7ACLl2Vwx
St68UuBIPRAUNZd+2kPbO43LA9Iezkb35zQ3EK/dihFhpRy3CFcyzDXtWNYqKKtb
UY0BfPucMo1z8btuy1XuDv04UZ832DBSk3JNuT1gK88JXyMU8PdxfmDs7v38VIEQ
zHTv5y0WyJngrBfTHVcrfNEJGGHMPbg6+esw0ARcETIJJT5xIW6RrnJDqCGQ5TJ/
9SE+mPrv4N6suf7pxmgMd5mObbM06nsgj8VFD31d5exhLpRxJ+JME1smnzxdi4f9
6gO2h0oeiJLRi0twN9Xnlg3RapbAGtSI89UOnrdPvhxu8fEZMoaHC29hJbetTh1j
FATfj6LILsyf84kg8WP8uSC8GOKF+vYl3sjVpzwvzixsNHDZQtd9OGHlRcqUOHzo
3ftFGU4Y1cKAyfOrhpXIiEsnsthAhfu419493b7AogH2zSgV9i0hlsRIrfYn7Pxa
hI+kb9/DvauojGwziyxecOfKm3JOmmILp4v5393pb6k38LBWhrZQUzzt92/aWEfr
fRBzLYPc9KJuiibXTXHrkcvNwtaYfonuVOYMDrgo7iOgNT2aMbsGWoLr6ovG1IPK
Y6NMn8o8xdYOSykd7MgEq/cD2fn7SGLlAuZ0eWxGygPT3aVBRqqM8bxwYJCTLbe8
WSQEZxNbO+bArPJCnFQMS7QuRGeelT9huuOmob21G3vMiyrZC9Ie88MmhTd+RP85
dhCJblY1GdEgi8YQwIIxNrNXSt2NAIwGI+87zhVVenp3LM+Qh3whJjH1Ogps4HMH
AxVQNS1DEpON2x+1RbhNKH2KWvslAicHchnEan3ktApD9LKYyXjcq4EYZH1KK9F9
qMtrS+KCQWZnCMjDKcrH4TcnoijElvvUhAePRwTmThA8ObQxn6UBto4jzQPhFD09
NJE2pnyPOpis48+znWroiJ7hB0DirmRQoRY0ksMPoipgpidEEPZDXZZS6aUEZFRe
r9cK8fEJRalFgBpfZnb94qtluhIFSCfVfBem3439cHYFSmTHFkA5dPuCLKk/MeZv
pMNkT2ndS8XDtvo66p9ZlSP52CPIyXQmU8Ux7QUvyl7jsjIVvnkfnuNTjuQMOcMB
meO65Abx63u3Z2ZdLwGvn+/Q5+NOse1ROkGkFUpMystYAFityLOmqk7/LgvQFRGz
M5Oc6kW9IGSAmudGcPqLfLVkNjsk5vJ198qbC6uZhHQVpQB9H9QZMyWXs7f9iYP3
5ThBTWE6Nr249RpFAYr5dvibPNWqumJ9goGc9poP5cWN2BsWKScOwhov3K95llQN
jbaiR3hTymZxRyvVGUOAM0rdo0b0v7qwh9btMCrRrl+nhHfbYmrbG0+kQk02U6f7
SEuHr+/5993h/KDVzjaEW4pJaQCd43VslVhw+HwOj6TwdjfWK0YRauCOZ8xGWqml
ZpqrwMiBP0GlmL4K4z6LGCicwd/ZCQfia7m38GXhQMstY7P2v/qDksrY1aqJn0LB
gGdDQ11MNTK0PbKMV/+gsFUTkqCyHa9hXRlIoeuxEYm3jDyMKtE8e5Gqhf+eGTrN
4RVZkNDjIZ6QBfvMiNJPCcPF1U6P7fJlHcN7URZ7dg/GIcnjojuUo1y5vJnp01MM
gbZ7z2GwWa1n9LI+71BnPZP/V7YwW/NsfGNqBa1gOtq3oL6oM2DZVUqzZopBC4JK
KKcRcKUeekkUhD1zKcMBxyewuVnjYUl6B2Z9RIiErhWl4N2M5Edxc0v1ly9PHtb7
l7OKHwIHv2yG3UsAWt6CbTZtNMEEOibIzKcwZp8X2vuJE5yFjP37LJOQsKGc3xkk
OJbSck2eUNRjgo/AU7llZcniM5369nbfH+N3FTaO43s2h98PEaqzmoYpNQvE7/jL
wkpwb1rNveL8bxvXCnAGBJtfsywcsed4Ya5NRlS72MwSI6IA7czcaQokBnHQhRJ6
aYJNImc2oaEexEa6nsqscqFmaLp4SYM9e5IydOBgWB6lgpzThVSAux69NxMW4qxG
5sbG5w0b8M1eQj473VOdNf3eW1fCFNH4DSWdfP+LEDiW5KBSn5Re3OXW6lh3yqoC
yhHB32fsH9zlvK8lqPhRzQZKbosyHHnRU0k+5SkdTk8KjI5bmR6eSybB9+dgs4RH
EX76RZC0MOGZMklfSDe1dB0p6a07c/KJAxDMsZG8KOIZiylXefDyEYMxAilUwFgT
oMyB2zdIAxSiJiBhtka0MrgZX8FlTd8qfcua6BH6cogHRdySQfTGuPgiYcXVwYgi
d2zB+Dm84K1y2XR1xfeBJOoPJWYcNY5hw4iRU+hApg0LVUlDZmpztivfRFVpCDXb
U0fYq/xCNjI6efWs/TErRFqAXfI/KqlOAk22Tl8Z+DJ8/4ruBSjSYL3hsZl8HoQd
xEHuF4liIitPymch74SRSag+SyahbFKQIvpt+woBS1bpg/oTliCHzbeA6+V4jaPk
WkEL2Wk+L+X0u4Ca+k4CsIbhfUOXzHD2+7SjpBcuFjmVTXl2MLUoJN/gmEhDItQO
2W9YUJuHM9afUsXoD5G5LUwA8tNcvEmm3TDQki83rTwEz1wMveNnmdLCyVZ8KDF9
ixW9ytM4VjWhst3I2q4uDU/AvqqMZF0BYZjxh5djmOfV2Rzx43DeNlxwt7Gl0KEb
UiAQ8C/9uTB31AunfNcJq+jthpkTMoIWQ8gGMLtHDsiQi1ERMuovEBrpZrxCHijd
ifIl0Sfg+50gpDF9iE0dDQQ6qY6FtcrKl3zdQYhZGoLwpE5s48GjT5nvuXLYMzcn
OEzgT0tGS85EYNvbPDIpyIc+tyXD0uep87txFZYF/E8YG9/n/TF3J15u3xapxOdc
9ZRhnKG9iZCBcYkL0+S8QJwYQCMiWX6IUElDyHqxuxvBWSxYLmc1zt7ibbraOG5J
E2WY4y70NLIwfc7CrGBmzCrHPSXKWnQfNTIiIGxWZZ0pou4Xh3B9DIe0hlBiimoS
xbMaGYztSA9H6Ul6APwP4bJXEiwH+L/oIUlAcfeu6RdoF3xsnJYuHxirPqYg8szl
pa106Fr6LmeClhxKqCJsf7zUHdvgW0l3UOYOfzIbs+ZQUkvR1l0pfBisYEp1s+Hk
xeO7pm1+TdPnwKetlY8Yy5waIXmqUifZbY3fwvwdB6t+3nvLOTIiBWPZSVvcrbvq
rnJjMNHtlYDrnZ7r94OvTKwrHMgMXnk69dmLNPjRZLMdN3RaUVHmuqX4bgutgzpl
9qpxKMgSBExvjYZb2l4XvrtvJmaAVSFYOZZ/6+wZ2Xqn0AQtg5zMjx20EL+xZXe0
BUtRTDWrRDy3JXQdB5oSLCm2QNMylF647jgOmOi7mV6UoDOtCYujgu0LzGHvzf87
wTr/UqeCYMjrn03Py7td52h8w7VyKprNqWkcLhdCIdhJBuAQ1FkDTZvR+ZhjxIvU
to0WG8BkkcGTWvqIrMRNCcC0dFsoMRFddZCu9KAB+lNL3o1OefIAIovxAA0bj6ZO
4YjKRNZVUA83zCPV/mNVIiEUmRpBbuUQFx73SlA/ip0FzGG24FoFWrjYRWUzxOQK
4so2LP0MqVl2nKZwmfbQH+ZoL6Rz3F6duttQf4IfTLTxQFmBjFj9SRYc3X6ELvZf
DBnXmfHNY5E2G/0iC9faNc40auFNZcV6jjhF16h3eD2M3kza16fGC2HsMeGhZJUJ
oDp524Bbf47AEmcpAS0QBXceYofYuhxv1oZC4RckwH25mDrwyZqr90ea9jG88P/r
Yv6ekyk9Q5mDoPgMxYeW+h3CRepZCK0gcu40VUP/Q89YWoyXCbv7Q4GvWoUmOLL9
o5UK8c48RD1mN3IKjFdbKX7fDylxaYNo6FYY7D7GrbPrA9W5ZGKybWofsNVrN5pB
PvG15lObG5AVJx2y7mhYC13ZDMG7E+WeXthPWwVw2TF5zdpm4Q0oug9jHiM6Fi7A
05QPZBihlDK50TfQByeEUeCJCavTPUupe3MO4gInhVuzndMu0kteVBF7tlVPdbtF
DUuTGP8hKQZLkssK4Cw+suSqD7vgHu5l9gSSpP7Tloits9TXYiP249iMu4HgaLmX
9wD1GLAt2HHfqnY+KQgX9qrk2Gjti600S5XJJo7SU066g72rBC2CpifhKhmzs7sJ
2jhLZo38KDfjLyum2qlMPjN+ShY+daJrKht/mR/vKw9rL3Rrakp3lgxaVb+gnsfQ
9WDZ6taX0UsFF8P3LOSJIR0avq9kWtfeArQLSbHHpJWUR3k5h5IQcOudTpWrf8nG
4T5tIKQ8H6/aV+siQfCWrdUjNhHPsxH8YgrLy4SrrN1myHjU6hQTP9BjaPZjPfid
Zm5OpBFuhyWuWsYR4ype3jqBd8ySZkJrRRfww2DFjdjQHNvWNseSy53F7VL/+c2f
mTuLxSAOvuWsRGLOC/asMS8MH5TZ1IobtJ629sDXSf7VylnGrNyWdTlZPFw8YUkB
CE9f5+yySjPGgCdnvly6T/R8LvpTFNO9bda0N6CiutmdsRydUASEGO1mONcZjhyQ
K4ZjrckzBjsZ42Xjx34P3XoPIZkSYsqoDVoTmvxcjlSsQF9lmRpXc7MpuQr+RRcD
tnRFckv7Uh+5qK7i5uvD+okyZI/eLOwQ39BOQEEWjbIh7ARYQdrUhVMIIirYO7Ab
ABhZOLr3/cSc3FKZWP8iyrCDb9ZkW8RDPN+hUmIxfeqfRAzD5UV6SRnG1TGUoDP1
YqlMLNIJBKgx8Qk5ieOUVkB0JRlgw8BZKuDlqwgIA463Heq/Y5kDm5ObVrAWbVlh
e/vhsp4jkaDxrVuFwK016IEV6fQqPLD3u6PGCbXfQxJRHOwOkV4G3FBryZAebdN7
JeCEDqPtTDerNswDo80rfEW8LspB+qJSxUIhHoykdJVjV8fFFU20TqGO8vKUpvPl
BxPCCWQYOaZYtyW9KiSC9pLZykRMr4Tf9a6LrFzdqZt0tl7TOlcEUxtQEQJMfo/K
6pqKSxTeVvz5Kzb7UzfUAWdXJnmZXYVeCnT1QWbkhhtX4HrEa1Tk3+83LX8uqTtB
vheojw5h2igMIWR7Mvhge3uTYDyLkp9DEFFUSS2g7J4tEB6WiI8TO1NN0JDhdLVe
kSjVQXWUdBjG8+e+1zhy93rVevaS3Fq9XXcgMjDa/zh4k/UVArjQTi00smOjzlcT
uY/wpkKY5LB4PhwfHUfEmXv198YndeIOxkq23If7zSh1K3G1QHRfE/ttRWWvW8XE
tz4UslSuFVanIZAldUz9P7pUIue0/ytnjyNo3hzkfM0y1FVI5KZvZWAk0aJqTEFe
vhn8/krZxIAcZfr/LLnnbzpQGUVXqSF7y5tfQY4MWBGJAm1GkAEn936XvswBKe78
/ATwHP1SCLTJfEEWXwVaApT47LfYXjSedaBWKKWakrcQkhciI/62M5vXbU36w9i4
vYH/P+FHCP8vGLxdkDq8PhaZmuDuZ3TUhnBbghBFQeMpKcvnaWR5wsee10CMuAqR
7kuWqE0AKR65GzIYZMkwmkFLyH3Wjj3+Ru18pPVth8FgA2edIyGQXSpVkSjvEKZ+
OL0ebgsiOU971N+NN9LYLx7mOuyVHQX+i+eSAsB1jdxCjWn80d3LLxM4dxBPw1LK
VUTEBjd8aNIXIGaaabwrDPmmnnxxX7lvuHB8wom0CdsgYOY/7DEzXFZnjS8GcIKz
ZV94RxKGEWPw19F4b64K3J1w0Z31GBsMCgWtL1ORrKr3Ml0w6Mur4gMVl2eeeUzB
wSOsJZHpfXOSrQ3+O/gffPHdEkgXF+196aqvLmO/KTvThDC63PRPxOHUTXDnxWcE
Vn8ayzZb78xDsNead3M1VCtWJ7ZZcmuUe1R0sCDYmUbMuHckW9E7xTF7cihcQTr2
GE98Q1kf0bfLvUygSzGl6oRX1iI9UXNhv+TtR74RhcRH4Fh3GXCroWYOQzfKfeFR
Yaxis1yLPCOck/EJNVGyYMnrqT+Ckd++KP2xAXGAMajeDJFXw2kPDGh8KPUzTtkY
V9Y/UipeZ3hpCKNMTXxEZGCzRkvzVDYywYqSfEpXO/BAHis3YHuZf1pThbVk3+WI
H4njm9aYxt64hV634brvW2dh42jhS5DaN4x/Y8CzNiwNOc2stu1Z7IuEqsT1KhfJ
uPIQpbb8vLyGVqNIKZWuCMmnPnH4As8Ue6JI9nSFDgD0Wg5ImCO8KUUfiSzcuIEc
75T3JY9JedaBz1M+QnJqlcg0Js+tEHEV1xVxY9LRYuBJd7ANIHeUHeSY1UrBaG3H
0di8TW5FgrnMU4WVgkw2JqCBy3ojlSiV9hu30kxlQ6+k87Ja0bj3MHZtt9MQ+/u3
fc0OYKsbVQ03pRkAfFtXLubaZMngEpgniNlwcb+mG2hzkaa5jE2n4p7do2L4iP1G
GtOpVOUDHLUVseqx4y3owRR+C4de+807Cl+cECUQ5GiUcavQQFhLthfLqlEW0We9
IsIGsJalE55nuRfO8TbSMRWJxOKZ70pxaEQPJlR7KAVpEDBDp7AWkqjOd0TZUF5L
RswwNto9P8szcnighmE6QcpF9FDYww1bdCUoaolEzi0L6YqwmLE2/M2d0Yhdy3rp
xFi15j7DRLJn0yYbzWz3yv+fy2dpYah5/BsaGP+PMGK+2+BS0Mxzd4oNJ+LYPvWJ
0atAE/oMOq9v3+JL3zgqM/Fb42ESK/exoadg97BMrAcCc4VQB18GQsfwrZylLxJs
HJhAPcnv32+PdhagzzSwzr+t6bFnfiguv3xs1Y/X7kBpMNHzBNbo2q6qr8s7Tp4/
ppjRlamrABnnbwstaA9tCK8hyJTZfJcHWyeu2FAnfFgGJWmC6aKaEEB2k7rR7jb5
ic0pZl4V89/T172SEvzDgsiw7itcr58zKKxMUgK+YC4CP3mBS+u1WActwCF6wwgP
lwNSp//5LLQIAAzkWvYc0AKiyh0HTwtIqqIimkYb41MkoGCnZLAy6ndiiQX/z/pi
C+OudfH96s7YgO2WNd3SUj0AU/Mk7wHMSO7EPl4KS4LIqU2SkTBhwKbqVgR0tGBa
1xF9aR4BBs2cgVOaJe49PUlZOQD2Qm5AZcMJ/aKIXhZCJvgDv9HBaoMrJaAaZr2m
7Imt4zy2wh2V2QRtkSPm/WproGTn8aukQjtAuiCNXM41a4F7uSQJPhFL3ORZNmCa
IzTIQYn8MaB4TlJ6Alyr8OB9n5w63YX2B09ea3pCpP8/t/lRTU/5UFiVaSmVGLpF
b2Lsm3mY+p/KZ3gcyECAdEudNhMIY7hakrnWvTucFvTBjvrXNqUxyNhvNoW6Tl7E
pPvbNMnse8/tlbbrE8Q+lHE2GLQIi+30YbTbHgUON9Kdw4zn8sWKnYNw2Oe4dI9W
LvcrTXZaXuDAKk80rE/Efh89FiIcsozAA1NYcwqKcsEv/V6Y41b/lRs0frDSJYtx
GVEG65B++2Aq3RR/BMjd+2mIewBfhKV8fm884SHt4s8LaaLM9s3GRxy4UZrFksSv
nvUYaLhxyd1ReKZMXYQbmUutSnRmJoDveCbDDSLCBVG/ZEN64cG+mmgTRcPvjs+7
9tf9T9OvZWkDQDFcT60hqxsrcUu8EvM97+IozQRx6zrRHV1RHKUbGMHxtwDOFON1
+jlrS2rWIxfpIex9mJ/CcLKDybjq/l4CXwk+n0UuC8yykPKWRUrIWqg0OfvXaKVY
C/r+wY0OtgKWNBYEbTgQHq7SSLglErLz/vKmpuezj/kjRoKQt9wNlIIoI4clk2Ld
rZ1voPbmfcKXi1G0GOKRtg0omdx5W0TkaJuzv8yZpmghQrCFuSQMD79raBsdObzD
zP2w5DHurzjcWUjILq2dulOXsmCYcxb16tmPCTNt9cfxWHJTKK3iBfj23jqrI2Ux
6J0pfTo54LbQbPalNQ8ON9OEIwW+W89ZloQEOFLW5qmE0A1ErVysHTf2FpNNdNH8
FVEJujUhP6cgJ7UZhYvYbtbr8+Qx0XFHZC8n6v4u+HSXmUTL7ZZa0tq5+Zhk2nAo
2F9862XCMwr0nexjNxrZ/hr/iIfImp2Q0751ir8W39+qzXlQzQCBMVnl5b8oNUHZ
qzFLTSfcAgfl/2B0vHO3hqoCTdCWxtsE8hhUxo+7wkoEFVoVGP1PjPwdEy2InCGt
kKb/L6t2V7ld1GOgI/sXdG8SDJgM4g/mnHL2h+CPWnDNGtDJIsxl+GkVAEXIO8/P
d61/UoEP6lwFuK3dR7cOLOmKg0LFmjMHTYpt4Koy0WHA3c3Q8xkHtErR/R0yoFXZ
4EIhT3ncVvYSkqCHbiP5N1INTRkO+0WIhT+U+QlCavW8Yh6RZfvr9DNzxOCcNH/A
FN67CHS9sJLAI3lZchOzpb99/fyIib6kY4x8BVSXWcT2a9RNj7pLQgvUZL2GS2i1
9N2foNTkgu1gfTe2IPYAaweyf4t5sOLGNAY0npxAoKXOf6e4jqGxkJLj3E3BcLfY
tYFGlP6VjSrHporm4LmAU54faazZ9wVZE+C4aCuHIhC+bRIpQJmHDWlG99WYMLgJ
s7+VT7DyjyFqtnbRlys6zE1W6SfS4wd9k4VdgINuSUl1jZEwzSXwBqAZS0kp1QFc
80GRiL7ZGtW/gkgk1eKGWgoXZDPIns3AfefRZj+qZeKqQ0R2Yp+3pmQRwJvcEJpz
NClFiXbixIk5OP+BOMAxU1h/mFbSFKtoIwl+TA2tA067YNhaqsTHtRPSdCzpFQ86
u0PtkKjd4PZPD/NVhV0N0FDMJGsTlMr+ICOTqvRKDvDDM125o4HNhubbxrtj46av
NNbmADqBnXc2ut10GsdW+JLJSbwdeRtD63jR+jbKv4ysQ4UCXZfL6Ov7XQ89eMVm
Oa1iMn/BihDnZvqhQ43rqPc/nQfzmr1I/it2fCRVdtcXILHTya0JY/HAE03JBNEf
1NURfcCmTkYJrp7Eba6igtLJWSZ06gmIRGbSQ/IpTgD4mQHebzG0O/eXu3I8HiHs
q5dCoavr6gQp0R9h+Du0zP/s/jSe5EJa3/zmhojF95c3RfKjQRXJQ3AV6kBHOIML
QO2z9gKGo/G5mGXxWN38/RyT4Z+A3+LGNyCazkr8MWZqpVRP9JuoAkStr0qtmC1+
toRE6Yiy7Lbq0l54hNt0SfABChcu+Nb7h8sMr2TME7T4UT02RX97p09DILQgLgus
jT+sQrHmsAeJcBF4D/A9vqJjwL1Pxr5Jql00Rj146gY7nc9IoNhTP7cbgGsraHNh
kJjVH5gpr0EKow3VxVsJVxn4ymk9n871hRvSbXRovA9Bzx90oqZo7E/0id+VEM2r
e4czVMLjm8fG6xv9alFKeBxbeGD5IukGAT3Ub2WC7Rrjod6taN1pDztZOD0R0TbQ
FhqtRlvsqEL47QOqM9ywg2xu7uzinkLagYMT8vEobyQP+/SxLfypYq7xH+q1kUZu
DiEQLExkM2zSKLwJevvBXiw9pVwlU+VW8tpWx0HDLa0FCi4yQUKTZtOP+cEKNdqA
tZOlgx3HIdHzXfL0tw5IAf5S/rI411fpAVCni5TCGG7ZXDnp1KnBfi/6dZ4ghI8S
llvgImioYapNIyASGkqJs8LSkHzBg6PNNHIuvpiQASm6PPpCfnBc3XlfnBl+5ZvD
JKEUgWo2UtrHWpbpHewxegepFW/e4OBES4RNDghOw2m0kiQbse+QGk9YFC3mRJEs
++8FRk/UMVWhgtdCGdPfSh8AUUDeId4SuKICYR4t18+Y+HM9NrcafgVw6K3TBaIe
9C3DXmwChQa2JVRiYAvkfgCbrrEs1qokK5rHpCghcDxVeVsM3TCwuXuS18UCNl9I
9O7bl4e5RD3cCbXvpAf6BFGHeG/wNFe2nUQPs7govkYabcGTCK1QBHWfW9ogXxi1
n9QMnGeIacfhk2on4piwQ/oaae4wgIZeKxpqmFWagE7norOqnrEkfgGjW67SOT/7
EGQ6O8hl4nEyPYg5Nl7FLBIRT4wdOJZ9Y7pcsGCM59pKbuvf9gY6h4+NQOpdjY/O
oPecugp2u9dyphaSyInfJasK1PHfRr+MP3x7sLqOYOqJO66OLyOhrKKZ1+wCfwqu
VXtrWoGpQFGlsIXfcNtNW3ABIWl6C2kXeWRM+6VujpdDq9sDnEptUGBrSAzTL331
MRTg2SK5lts8k1esltmq9/zsVkSqUGNNibzpSBG5f/dn2uD64KzGlugMm+PAxdSW
XcKX4UzIkcpYEdqGAJ6uSXfdS10Vfh9BoxmCBJJKG4MjcSVFMxDLUJZH8jym6TZz
iWNDm9BBjGnx27cnVPCrAb8v29rc4P9MhY+4UmFrETpCADq8/XgK0OW+/1gKeV4m
LyWE9LKpu/xhfWS81vDzLLtcVucw28HIOGiH9R1Wh9KCPh+CA+DmeErvrLHE3Bts
XwDdaXoRPhTbLQxz1b9mAXSYRkyba54G/C/1gCgv0pZnl5d31B4ndosFINHKyxti
9SXoYakkf/WLbSOMyT+LkOGvFuiyX61E/LtGoyCoDM/cv2jPW/m60prW2tFUrwxJ
nvB4PQzV2OaoMXFsHVC1AAcXValGgck4tjYkGd9FT4x0zNcqLQQ73fvhxvTc3F2M
/l+MqROe42n8g53GV8QXqsomWN71ZMWjMX5pXdegJ9LLYEOeA5MWGhO4cD3Mq4GQ
c3BQet0TRwaOBX4IxLrCS5MvRXj0kaxfZiVPhhkmTB8D8Z92ubDrkySAjf5/PP0T
LWx8D9dZIi71QoB+TGbKYXfGlBeeTyeE9EFKlzXcCTlVTl26EbdbSWrZotepznTi
CvxHEBjqCjkhGC1G1dGOGrvY47ddJPC5ZCm/OYEBeiSqQLQ4yZOH0TwditKB/gWL
01k1cJAXSWfYuOF7dRmOfXKi8Dw9cp4PrLkxFiI75uR6lYIqFGV2jMzabhBHi5RM
4sG1UTFP33CDmyMf5mM457kshKvyzsPOnqSXrwVsAD0l//QdFb7AfsnMERgQS2f3
RcJsc053uh2GUv4Hz380k3w7ID63IBTCzjaSq1+4+4bOgWA/GYS0vvdd3k/uw8wM
yUGSlIdD7UnGtk9dTpYLX2/g3IIEXzwnwi5wK7V+tUoKbnHINbpKbNFcf5kkYd6T
9rK6DPHF14nK131Ve0EZzes4eB7+796XPAnE+ouXTjMj4Rq8WUDQANvooQ7MhzLO
KordZbvtt7lquI6InLy9zNgl8z2FUKXOwjlDyq3sxJGvRfU/IH23kKYrG+Xyu9uB
vtqrodtxkH+c/5hkrHa1hr5ukkx5kYvbTVE4Z+dANGh5DQnZRc5Bdf6FjdHJ6Ymg
H2QTW48OocV6w9ESpaZemPeQQNFB+0ODrYBQk6ByrXN0DkjIqBQfie+cp6yHCuaM
zUDqvMz0KYIhbA4vOjXYN9zsaN+qRxZsgNJ6AKHqlenjFoV0FJUw69I8x7qUc4N/
X02mgXoHc3y42MzfeUJTyT/nXl7xR+PxFNPa8Xy+DsCMXYCt/uogcxfx9cyp0oF0
KQCJajhHgYSjhxeezztOKmmVetfFIu/AwA3ngr5cKdfxWvz14D6cNN6lLnh77MHR
L6dCGyIC8zGhB/8/rtoDWJKVJVPKU56gtpFGIzhj0OIuD+4tIaFyxzJpcNarO5jt
YoLR/PNG25/c2eDReRm8WANTrbbctidcVuge562utT5rwImXgec6AJ+oBNTNNpCA
VaQQoKNFbbUaT9Iy4xestCyFIPy87M88BlmJxcCu5kOFOHPCBM+zzsphTphJvmYt
32HLl2p4p/q5nAtr8BvpYGBymraXTBg0wbEOEku+BlTZLpONNJJ7TPHe6Vz2NsSC
uL5uWsfUrpKhB25g5S3XxklWGt9xq9SeWInZIfoYsZVJrEQ5SJHATUbZkFXYkoKz
B9W+FsaZbs6b7GiZ5s09jQnWHrOtLtcbt/fo7zp29P2tYXOS75AUNqR2vQIYC9l3
0yZIzdQ/ikf5WnTOydlcEK2jGVetTWhshQUFna9opshMKK+V15VJ2JP1waZP094f
uqynsHxSk+VRv78zsWTjRI2H1Dl2CYOtDx6+85c2KJbh01ZPhQUWRPBQ5UOeOD3D
lo2ue68/swIc1+6lCosy9C4r1q39+crc26D7dmWsd5rs70bOomONONW89CMATYdt
oO337VsK85YnROj9heeTM4NHPSJ+i/Bgc0iquM/bk5FNKjV25BGI+XEh+UxA5Ydr
VZUz1t9NqNXvywTpms7zruHA7XlGF6HCDr1UXZu3hk/g2PsH1nddaOgTO52n4Nm6
AYU7Xc8cdYVK3lCeOiSA1vJkAP02yQHjIWKjckgePzOpvsNQTZE4oCLFVZkuIxAT
BOfi1dL+FUrnfiG+ryBYqNjWZfJZ7bRa+uu0MrV6bgWwlP9Z3cOOaijvjtirH+W3
ys3u7PNVKPnhEWXJl6+07+NyUya7vRG07ZGuVkPJGVuxNdwNb83XMMntUmZ6FeJ3
8wO/lhZ4i1nhzDKG3m5F8Kz9b1N+uJfMgE2L5LFYkOs3/nJMSeoxl/6dW1FIsxbN
yWjxPBeVNJmG+avPDlnoTkn2IfjNo+uRLiCerxrlXC+u39HJ62U+hf7RQ79FnWPP
sBD395XrvKtEbiOHQfXtWj5+f4mLYMZona1Wo7aJT2cUADhZBKZrq7dJohFR1CTA
v/j0YiO8OEsVa6zcOUEdWBQd2seuCv8rt/lZ0H/pABvPOZz0TyPQFAzpFQhrGAHo
ChSQHFPSeMiaWNskRlw3L2mRFTvw+LunlcudKDWEG6WH1jKRXsb5QL/OtpDni/DE
iMOPVzmAdESfCujy4mhRyVd0lwiNPL6bOTU45K7OE1c9E5h3cr/O/YibOxblXxDm
R4vAOyXaNv37jgu/vyNryG4e8H5U0U8Al6Xf5wv0J1TaBxhh4pRGeiEaHzIARENh
Bp8tbBKveQziXD9ks4s1/qqAd7rbDVBt5fxW+SH5QhWzvq2F6/T+xopdSebWHY3I
e2Rp7UaoYIMzuNnxT6qwRrKACDxb5+4qHcpLnLb1hsLiIrLLTSbwc3X5Veo069Ih
5ffSJCW1DZRiaBV1R/sjVZTEfbahKR3Fjhso2WxC1Hr7iRa49RoTZ26HnCgiwFLf
MvdeSCtfSTicNQq95ZV9F4mKfrhkZURI/NLd+yudCCLj24KQ+r6fVfwnKSYVKfUV
WPkD4NbgebpZHxetZgTQXqtzKWAEjyK2XGOXEwEfm5ZPNGTuMgsuNkh0FdDbW9Oe
auoG4lQe8L38nia0tnvM3qcMq2gBlYajM7a05WmAOx4CKQR/KrdlZ4VEY22kigbu
vMMdl+JlLnP7VG1bNTVN/CNuYmSY04PBDmFcR16OmFvg5Md7qeeRsDnikTBumU7u
BGZDmw5irIG0uhRE+ojab5ZRx3F35qcXbO53BF5FBPit1I3ySjDXhRsjYHQwzWij
GnSJMy0tl9sRoYb58jW5QIaFgdzZ0S24oYqYncHkOw5+StXgQqzvl9BHq9H3ZeL2
32SKy7qZ42Dn8sPagRZRBo5daruasuC54hqIS4p4GqTiFd1VD/WxbibehlTPdx8Z
X7OVwsJ7HsEeNkvAExkWlE1gP/479CqF1ieGa5+nVYc89SLQz8QiuxfqqnsmkXou
Mj4rXgfrFXJvkiAJ9N7rwa+pJoZyCHWqCxUk5cbvLGMk6Rc9FKBAuBDWVw1Qaw1o
HvDE99gakoU4o9/1KZFspfTjbH8vADgSrk/fjfiguQ2yP/by5wAGFfkv6cCSjc0V
4UxOTCMiOZmXM0CoQg0FBXsbjJXb4MppK3M5XtKQIMHlumOtwfjVuCAGmdVQ1IZb
7FJfBuPWYi7qT+4iIjysYlBodHvjAA3iQYADtD/XYPDsfZnWQZueojLH/vGIZlrU
1ZOyuO0F8gPQNGnXM4w6XyPebnl9sJ3I0f1gG3e21uu4jOSWUqOEu6E/3RtR2EwH
FzG6Dxbyk+sRlUSaYFr+wp11yXLjB8n1wTc2k0A9Ej7Ph1dNPuQQJGvLbc/8HqAm
8Vrj8tjKBGU6/StzdLpPAxHoVfiZ//+/A1S38A5oIdNisvVy1nQ4k73KslnSDtPs
zBHp1Yl2Cvnc5RhXtixrIHfQ9BxVw1T+cPDVoMZh5EKqSZUs1/vPBUVsHwDewMYY
ftja9qEUoVsM1qqvGIeq4V4VFsINrY0YFeXb2jMYHL/Xgu4ZdDGAa13bS9iXb4KM
z1StjAAUYABIyNWm6EmLTxHCuBtR4wdybPfmi4i+mJZ/dz52kV7dm6dOGERYfAXD
0J0BUZ9qY1GISGr4rVYsMWJqGgL9PJkyADbYR/xsHkCBkX5iROGAwRVweuGimU+S
NDbtFNU68PBHLpMI9vMqSPMWuKwgN9SFhZdysEcj/sHGE6JZB9ESH5h2VvCqaYY3
DtcZms0kQrjj9RPSdAp6q7hUNg16zOo39NAKqmUG9Ewj/Z0+wzGVT/QRJUcVuThV
I9cVCfHRjNvRFmlSlzpNsbQ+q+UqLhaGJTGmjxrlrCgxk5cReTsDPiHgGLQVJr9o
+UhV19wppwBeg1zBujkem7D3AxYA88fRvnXJwSqCsrwKMPXkMRoBoEsSUfIJyxiV
fsbnw+wY2wcBULvSe0Rs4yDOdF6alyCVaD5QaOEocvk+w6oucEtySj1k9lqFNH3h
7G4fR9TkYTfUBmvG16+Ki6mugFCIkDXp28OyZDoi4J8GDLaGb41K0YN/r5oG6wXJ
840r2AS9GD0VKaGqzzt41k5fWsFdBQ/ubqj/stzNDBWTJjYydnKsfaempAAcEK0t
cTjd34GlSR8cOWEhDedDEkuEGZpi01mpnwGPHTjr1X+iR+zUAH1knOwjd1ePwGXF
Om2lQhDR8X65orU/7hy3jfJj8E/J1dwHSpIvqR4tgCq7yL+clj2pFEYE6N0ge6bf
zoL19Q6BpYWStQiXx0++c6+jegylYr1Kklf3s6spjDQ30p7iLTIGLlCDW6cIXVDR
Od/GON/v2JQ4l8kL79VQuF/IqB0Gbxar8Kav88QENvNeRsukn5HtXREtDJbVm0y8
nCkAGRgtKAwpBSU9l9Ti7ufJTnn1ec13md0DUB62H40cTcCwMRjbCiLOfS68yZDG
r7iFW+0Ggvx59AOyj2TEGRE8cY41OmoPEgXzGFRXNUS+0Scc/27TEPpAEkRFWpt6
XJ+jCLfwVjZ1Vy/TDEqXflkUTeyZ6l/Lris/vRPjGtzO8j2oSkgRHBDgYrpi+JTB
vUXtNMl0w068YZ3Kvuc4OuRyijmNU4dFo2bAyPlBA0zdzG6XkvsNNRe2AoepymA0
qHBdBrwVBTkNy83xbV3Rpz662zJcQ+92IPFy1r9dhGEvh3suXf2oeHvs1rGrvbCS
mvozSLZuitwGzy32NELmANLnwx9Bl/58wlhyF0t1V863d8yN0EIo3JvUcYwpuWle
05PbPXWMLSgLZ7ol32K6NEqLEQFd+s+lBW3dDOJsr2Ds06+Aj4lwulUQWZ/zggk8
xjaKnlXfyn0IhFcALHfhHfD9gEHwOlcrhEDvJYY2RmkjhHLfIgvV1xriLXbNoVoR
NGtlknYwyRa2M7jl6JgjthyjASxEjj6P01bMIOnQVOhoGxkfXQkhPRQTBLQ3240l
Or0sPRwcIq8aVN8/NfRkt6J+k6EhhHLrufMYsOD7uz6nNNpQNLz0Pkgp/9BEnY83
wndcSv7bmWv1yBymLCeIWob9F8sKxmP3YuenFH4v9iWtY9LRkYk5AJBmBBiZU6wn
9cF4mpAxTiPY8Yu0/aRdNHl/mZGNmJlELFYUfLcVu7qysMjnDoc/07Ljx2ydimfm
wmYYx8XsmN698tqpJpf9zusnaHHn9pKy4cw6/LJ9pFtUk2SQNjDYHdRIBNoIZtPB
dRqSZCYqx2fIS5eekE/Vd+uMSmSdFQ3U5WoCmbcQf7DrzF1U9OIyEBoDEMfi3O/P
2g4CdutDrQsQRzKK0PJQncQI2zITbnpMmEarRqV+Wce6wkwu+UHDPO7v4okYSu+/
lu/uJAznMWlD73XEQXgYCmy9/qxyzlLulPNflpHIWdZL6h0Ko+CxqzE641ZGraFy
b4MI9SBsBK1hN1Top5eUrhnALi+GRjWbLRNDiayrezQrsBrbl3RBWz64mi/1QuVu
6aAIDB+cXjWtOEMdPV9gZBkReMOuAXCpSa6pB/grZpdLU0845L0PcVusQmGL3xPX
0ZyBTluO8kyjr6hUAAQ29CW8VaLIyiY2WoXi4qcDbABPJvhXBq1XkKfppN5NFVQo
FBVSVPsEM1EzcVqSJamtmd6tirOhGluMHr8XYz5cKkZny3+ozhuDH576YjBasqrg
s/PrI1TA9m535pDjImwTofV+Qd6SVHbYMqph221htqdzqPJDa+zQvfjPEpMcwTxv
ET5VUXG9oj8prj1SgQ/0zCKKVrzTG7huXiO+liaWQaOkJIGIQLYVtcr45BKS79sY
lU7H9HDwJ++urm8JETspnyMu4Voi+tNA2YGRZ7qOVWw0CW7DF9a1ro9PPoY4Zivl
Nmv3zwdtU715GXyWbj5+uRlB7WTejX9ahl3/V8EHvpI+wkwlx0joYI/kJYAuraGh
TrxI1MDlNp+NuuwlkcOaQsOvQ0hRSJ6sX5IYq0evp+Ntemfh5z86AZnLmlLTxB6w
ZbHGNcd/Q6HmSdddjbJ0hNndBYgBXi+TzwjnoGIn0aDdggneLUyE4UgbAoqO/kaZ
DPVzoIz3Crz9VxMxR+dgHUMqAdcyuH1onzMdMIyZxm+WAVV1NnKulPNUK23CI/rJ
QvqI6WDYdyrsX+17HczshsczHcrQ9HiJuSKnCMdZBxfox3hfUxXLqkBl7bkXvGxe
Fj2ouoBUYHmPYu7MJ+xen1tWFIs1NRER+OkCMEB9USU+S3bYDWmesX0RIdet7Hmz
t51SvHzQHGyPNPT5VjsOB2tr9que45kS6jVBXUoy//qjuZkjNU43+jWgGuNM52+z
8ycvtVH/EW/3B35Eyu/ZKS4eRAsz/WRmuQkvxr2qombvr/nEDr9zHsoc/Ph/CwiF
he7mrbw8U0yLKJ9Zo92zoEUiUPkpycIhOIV9yTm130kd8sQHRx7xQLehgavdNCLg
NF2fQ6O3ImXpRF7LEKnXQT/5HzIi8fcazUoLRh9wsHHzZGKwAywngkDCPOKIJHo4
3ETEOnsuax+1rGHaSZBlj7/bnBD9MlYl3ZJTyraJKDY6eRSCy2iXg1ll327lPatt
DCOQt1V2nEfq3DCtl4Zo/eHKK05gNYcZSxrfe38zCgFsymvW2ok7Bca/P9vvMgHL
3R5BU658RopN5sJYO0aayc9KjGMtxHA/5r+KFRBXaPlppwE4LV1K9qBuhCznhXG6
DhoxTAK+GDp6ApeMW3RzCgmo7lqshybgoV0g9zM+5VmVyNIn0SbiwpjulSEAemDt
pVhPcG1CTAjjqlBlGfsuymymyo+PAsApTaZWBrqYnwNBwZ6VayCOGkilu1W8Nok+
FaBxO/TwVejkfC9uBGKM8MsFTTO4Pvn5CPVaZqlEfHZZaenuGRu85OILsoteoOGI
Bfu4xUiKAYZFu/uQq+GV/N4gDvh82gPvOipc6e9/+ihqSFJOhBgXnYytKiypwYnr
MettAUWtmNbdLQzXdvFndkWU8K2IRWD/NNLA6+DEMazdQ4+CsAxjpRkENlFPplVB
rK+EyGxfy5Cj80ot0jBZEn1SFr8vzCuIYd/nf3AdRPCfeXY1l2tZ2B2UK6szKqf6
j8vXeg0F1X8ihvUQLWOr9cH3d9fl8mus97Ck86maMzhrYiVDfOeVF14yOUBZa1ir
o532BBEOIXoThJiJHy4BTOcko+0+/XOym5tBnc66O3ypVf58z0d0Vb50FDUd51NS
jkoJoF/xu10xBEnHMMTgecunTD2nW6e++uF8I/6FMN/hIj6uDtm1c7N+uwH6b0dZ
nVtY2JGZDqUSeCDvRNs77f1zU88J3Y9zhAZhfmJVSsF5UgEgj2pUun3IKw1Ko8ys
cVV2HM1tnmS+OTqudkwpsCTgK3QLyl7eu51s5StGsJSxh+XWg9pFG8cIID3/N727
q2D9KPeCNIFflEzb6qcQkyfmTcTaPo7CkNwWWIhFs7VGWxQ1yB099CuziLKZNTKu
WrD6h6kqu0M4BOpc4LXDxnyQC8oAQ4ZZNzoVhYx/RSZjZMdmVssVQEFGK4eX6iwE
GVMqOu4Gi0J53ojkKyW4X7+P9kHXdn9+DVoEpirWARMZXJRTz+F3DXQAwQfek3f9
O2zj5/dz6zUmY+UDVz2p/YSNwhcdbivohipbHxLNXbUraiwY3x4Qv4JwVhs5X/yL
32453m75SXssu02Akw3/x/GywgE4HOkNmOnAs3erQ9spLQRuNWlHUikChtVeF+ik
GBY3fywGwsD3ZVTVHRgoo2DGV+EsBYggVr/+fLf0OGpVff+P6pJ1tsdYd9oOJ4VF
KRJpaecHW8QVPQvK7hTY/johTBEqRuYbX2dFeRKWgZTkZZSfH5HEbd/vvKn9pPw1
bq6rlgXvWVVJDfhqkNAiIkdgucWVM+psyGToRbeW0rRKXfu7kTmzT2Phq8bPgg4l
gk6jRzXLW3qxjOwV/dIwO8+hN/7M/CKqgggKjqe/Uy6D0HusSy3qYooxnzSKENrG
XlsaXVwJI2B2IQv9vRR/aDPpR4R4YlT31dckcsOywjoNoBm+pln++HN0WTAcwks1
huNKC0eln/ZPXaLJJ1qYZ/lPfmeeebYrmS/eQj3AkTtR76YDDitrUONWadIPF3M8
LeWxfyez/C7/WNDXiEDBgwhaT8OKuesrzdxn7Cj1GL1bjCA3aa8F/PzSpwrTcxP4
bMybg3LEZ0zEMTdkDEp+MH99dzafnwtAPAZRvAGiUhRqeQO/j7toFx10olBO9gw3
smc1/UyLLg5uB1Ur4ZrnBtkOjkdqohAGclpxTenFnCQvgc0tsKl4LVlqCcz9pkje
PGVp25gvGwXPSrb7+PZoSDrusHHo6PiJVwAvvt3R6CI7LT1DDt3SuMsAEKzUJLls
AmcPyZXsb7DNc3TqfhJvWYxn5y4rQtfkrkMFnv/B/Bp16tFWpRH1hIXU+d0hE0El
munc7aGxtF3vutP6gpWXo8U2EPbHf2KB5lfg0nqO4xjbORNcdFSpAS5zEwam5rfZ
`pragma protect end_protected
