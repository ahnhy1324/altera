// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
lWoytpc3cPusPsJ4OOSBlGGxdVLJMjAkhQwXks8Rr4ipUTwf1iMkR2ibNnLhIEb0aIgV+a4mdnqy
mfXRDTrVDhl/QAgrV+AL7PKN9isXUn6KVm72ZzkFIzlng0PVrzlADYQ1I101DJ6d24CISInxXt0N
ybBWxcv+EOJiHL5ksc0CpiLc01ytd1Lnihk8cJJgzu0cjdMBve3xlp0rD90YDzAz7BPF7wZrWXbu
uJngHwpkymkQxGYzaSRZU/Hl5REhHIHZ7PCgGqfr5HcPU3kaWszfDgSTWchzIRVeOajV6DBTZGNZ
+8tGFigwg4e284UiaE9swa4IpJgSf4TC8kdZbg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Tjlngbpbcs6KjX0vxryxdzPGTOKQ2VYg/PvBQIl9/jBZxxFgjE402/Z4kImf3X54OFuhzJpThRcg
+Muy4mOTpDwGYUEdNqmO/a0WecQOdfMJ2KrtOm/fG0VAMUJDipFKrqov/jq8RVXJZvQuiO1uejPw
yiJ9SFfidCKP+F538/PhPG7p7K8OYD5bHhKQ3O7cW4/YjSsc0vgqZAWYdWEIGqKGlTXQmim/0vie
eAXTlzDqIlP7ufSrN2uuVKC5TNf5/G1eeW6MDNewEKEwuqKVeBr8n9fxVqnANCABtsNUY75ZZNWb
5yycTfep5aJ3XpOvNEfPerV8TRqkk1LteY+ayN6ElSC3NeBZSR+ZnzzTbrL9rYMlYcW9KvnJ9Z0C
rYfSoNCcMaXIS52hFiI3ptn62yPKU4VAN/1LG4RCLCy5gKc5WnzUsHVn1rLBUtdpLwrC3YZJCz30
DXG40sIYupWioNB14Ybbp8dSinOhtBcU81Km1mMlFk8tn62UTyJ4sF+5YCBqQCOjMSmxkWlOfz3d
Gc9IzJNvhtRalPG5TxGqu34q755EkxDqd2y871dTmx07l5KihEYeFpcyN0I46CyPvFdgF3PRBEsP
kmn5YkvoAjI/XzgdPUrR7TO0SKs6L0SWpxTUkvzxNYi9omQdC1WjxeibSH9Jk3GH+HLiiZmhIZ+4
ePFx2h0maPw24P4eZc/tX+1PG/cMrV9XC9rVrLRBFQvFbjKNp35Zr2rsPVk+kfnnt2xLUKGIXsgi
NkT6DheqvWkwdwn9CslMmuPFvMkwuYUE+h6n8dPEN6hlrE4atNjk9N5n0Sh6Jp3ZC4wbcLflmeBf
krqoYJePb6fNauON7FDRDqA2ODU/zP9EEE9W5NaRPzyDTOM+iqjXbJ8X1VHfUdeei2u76wzlBqNk
LA042KdCk06e+YlED/zekLwILh115TCyAQsFGX2Q4aoge1TE+rMNLK9k7d4pMSsg0UuNj7uXvsGp
QaDVZU/YrnHrYiSnDzfYxC5yT14yXVS5VQQTa8YQg1qeKKlpzYKflSyI2I82O5tBr9pLF7hKx6dC
SzBKblxt52BsIlfJY8fsqPW9N7q9usNY57uEpVekLuY1XIIGc0CUnoBAfRlgifZR1ba0n10It/uo
+A4TtjtURnOPSf7wwm+/yxCbStbmDtw8SK/y5IjkY/U6cRpKn4u2L8VcuM5hWCFTsMrVNOSLgB0O
jtHRHt32+RxbUADo6XcpPbLv+4VDYNTgL+zixFgGbk62HaNkcR+PuAPknGPAuDQdvCMQ/B45ecVG
Wpzti3GNHoBUXEZZY3TFCKS+nTxqUO+dKLZoh/ocD4zJXDyn6O2wMa7Oy653GTiXf93/FZgSKlh6
LECNQiAN0qKvPiGPAnawUtiwy+QR73yuJAt4Le+mn+qdH8BK6muDdl7fw6/h9m0uhTU4lXxKLb0F
jJKBFUWoF3R4RE5ICdIp8dPTpzZrX+VSmMa+HxS6JA90l6Zmp0pNoJnF5pScLaKjugZ4AS39zUVR
82uIaWgWcwukGRLAyScEVN2SopgkArMLz4V+883FtoWsUGuNbOjpXRIzFseWQAf/oFfYkGEFb92d
kw5Nk0YDMgyyZCm6Jj3I6Aba6d426jTsqnzA3aP2oG7vUuugxZkr3sli/reH9rUvOHszyXY4i2E5
jROEA5FDdqzKfinhRMMT8KE6/YfRaa4eg7JNNtmYjJ3+ufInhsgtFfzZbMlJiXezvCGtst9qJVge
q68lzKHlbRpTnKO2uR8cCfnDgfdHi99+M0dyviRGoM4gnATXgE06QL9xkMNWFkfg/TPPxH2px0o+
UkOPHKezsPxymmaN8514DC2v2B6EKBSdp3Qxg0vFxvQ9wAPGDuCV2oRXYBkJAjt+UOpvzxcYBS7f
3BRBE89OPmq6LZfhdIJ+eOqmwqxE9c4o9tudeRyjSC9/ouEsA87bISPyspiYtKL0klr8MPz2hYoO
vPJiCDuj64ec5JOFditioTCjlg8Dfg+UuaYgZhGdMbdIeAzNkFeEfLP8yCokyIW2aOEnjg10xbvD
+oMHEStazvn83nN6o+oUmyB7rMjCtGoN5mBoRvGFgcZiUcNiPT8NVOUug5h2iIjL/K4t5ytURrrg
Q6ibUBkDdAgeLaPMIdhBSJ54DwWF8ubp1cRv57WcZRo1U4tKCdjvw8VLw6tTk3MgWAODS2Bt6HhT
hwmv1UW6N2eky62QNCTk7Kf2xyPfih3fEsuNhUDtElZKqWu38pL696uPVp70ZRl8vrO27YTtdj3s
z1VNvd6EGpRRWdq0vvWNn7FpFSo0nu24v1owTrvhSJOGv7Dk92ajv79XBsOW/leDFEfuT5P9o7Jd
h2jOz+cBLN6ZdOaWbrqAvDvL/nJwU20yDPfOWum6wgw6p6VO73gqKdp4XiOPE4WwoXHNI+JooJKI
DewwqhRRXt5lc+fJPDIx3X8nKDs8yI+e6qIxIE7BVAG6NpgM/xUNggOhA3Kvkl6pmR8hc1fOVUrt
bjrpq3DdSIaYWP763oBIxEWVthEQI2asXSxVoge5/FK8RvN5sBiKHgcCy5i5s6eiOSPj+YISHbjC
cEnDcSLelJ4JxIIEEDvBbBvjvIzojHGWPOi0EjtMWe/SqsN2oM38ytpymdH7ljT2r7D3AoCo0nej
0Z4rTbAgFgr9v/aYVXfU6fzQla5UKrFzH0W2ky0h0zU1fxoLawugIIy92Y5RMRb+VvTFivX6m+tk
QoDUuqVli6BL2vH9j7oi+kzSsV68Zvz6ggsgXuWVrttVc2fKaoTQxAtg6TMYRv8c+0pNy5Ie3A7O
CWHQNCQ4HsQ4I85I9dVMKLAWdatTe2PEBYhQ8MvhLO+GGDkbRRsscdF9XFwEvxsI9nSDGgQmIHAj
3YaD0MbW/X8djAoUrxLY8wJ+hDUm7SbLLyFT7J420d6S1Y+NK7spKPZuaxqJ6mpKWD9cg/FMZwXR
7EPB+Bn9DvkvPGvauA/YT/t6Y0m/gH/Ilvp/8YLTh58pzgckfKgGeITqy48wb+xI/LePig4c8IQH
T+Fj7LNBKZTr6jEQvqFOXH+TG0tCHTWE5In66E7wqTzbKNA1Yj3DKvnCf4K8qMafT1LAWs89btyq
tlorriFkjgc8wR2mqAPqGW5LrPojl2IUA8BYa+vcaM4GaUTTGdOWV5ttJOIqCbSfyFSaXUiBQ5Pg
vjkQkxFCrATAIGhudkrhasRCJvVief36KWuHNRmOM2yBaMgpyV0rnP4FSNDpWHQmFDtgNfo7hPVA
/glw2ASfabVLUuxjIeIsJsDp+EAo7udvy3ppUgkffAAO9Uu5OiEiWHWGuXcyOn4qMqJJyCPsYvbQ
0S1PUZNWBT0ZJqpldk5U/3W/alU9lgvEuW5BnzyBOfIAB6k/RvcMo8pz3zbmIWTj/hD08oF5gsyk
zaJdO2+lxZHkd15CEJHcnyWMVSB7uQS/O0jgIOBhfCMHmPTmbw7vR4zSW5ORb1uAEBxeJu2FB6e3
9c9xuY6yG+rF9sL7S7v6w13CTzEHaOs29tvfeRoqqArj1T0cAB4cCHVN0xKMxPBjx0kZFL6qVou8
Nl8x3TTA3Zl4vNUmoAMup2Wz/x5MirMb9unSKEhNVNG/Vk/0q/xkbHHwumYlcW3x4tA+nEyKVaeg
XaeaVFav6vdAbHvZBn1IEzM6ppptbyYQ2Dmf+KCjYFKUK4GGOEukrsOSiT6wXqGXNmcRHmfPMfrC
zUTZY/RDG262OmI5i3rZFm7hh95Zs7yy2aWxbLd7mgvu5UaBCHbFeHj9IzWvwGzt7ug18OfWyYYB
l/SRf25N9I5scGrG18Ond9Ca2LCaSEET0ygjgCYqN9uuEjUAcOx+RQDxAssJDZdnyYd1/kPqzz7a
ebb4QvwZFxLu1S+bOYDETGwXiRqqkr5LsGW4HdOpiVv0mQFL+j7EsoIu+3O9UIH24eIyC4LZCTU3
x04HCS3eLpA+yAmqjKGqe9XU3OOOKpkEVAzbNA/+wEE1f6bp8vJJkFgvsXSTQ03Sfi3o3X9/crP0
QGL1KNMzP2uIwFFoEaQMrHauX3qfvxRYrmn4y4PLMhIkq4cxUWpZTEoNMGNyZ4CzxsPIlkwj/cL2
y8GM0YUXlgBYf8ZZlF18xpX4BgNeo26gtmgUh4Ws07cUFz0n3cW1UTJj5vYC/mFd5Wbs3IVtD1Uh
k07JO3F61+dLneJmyqe8SVrNfmReIWVgsMDmeW6WYYcnzi4RkOGxpFilqmkIUIr++HGWrnteHhUh
Iu0tUXXAs74pynqZHNHWLaCiJ36+1EyIsVqFuSEd5EQrr3P4z7peE1TKmNg8BmR5EbbOqIbO2f8i
XlYMIjTxURMeCQIqSqlWj2q9ZZdvcaS0nCLT4dRaKmbe0pG7AQUaYsKEyil/Shm2udEM2dDTtPoG
P01x+yzS2Bcldchk/sMLQaDOSN96wzHidgvlPDi+IdvK9drMC8kLG8SoH5QUKxUYdveel7khspUu
LNcDcwse7d53ywoeygbiKDqxJI6h+JfqyfRPM8LeV2+bWi0h8BjJyDDxiuvAE450/Nhn7o5Z/PPZ
9CMuJ1NuZ5qUB8yGFey4kR/sxl6xWhrtTewcG7p80w+AvgAwND43iJEKhY/BhhxAAbS004Yj8NrC
WB6kL4dfpxLJmkQaaMIOO5o5ATDDnR+ydHesNswZkpLffbjV8O9OYPdXx6xPlQDIrBiMI8QIb8XR
nw0OHp4X21ljlGGJtvLdD82haGF8lL2Zui6pvpjh3GP3SpOE0JFv+5WYgH8+Fhi73e5iXBwlqMbH
vzFoih9RYYCCqaG9vUbomY8Ekendqz5eHWgNG2V4Z9slc0XvJtE4KDV2vej7amY42shSonehizyg
2idd6ZCuXT9ssolgrcZQlE/P1PxVt9t2IDX77OBkoI4G5CN1KHrNOD1yXUT5DiFQ+A2J2rEYSmIZ
MOIYrJusQJK1M6dGn3RlfqF4vFnqopcGHlMeer/q+N0G7nNB4P4vwN2RQNnS7bGgLSkxfawsfnNU
EvlOgZ4ZxXhOlUb3p2yD1o8+Aezh+465vCTov6THBX65nL+VG58l2RlDq1B+CkhEclc3p8SqH5id
q+thBW6zkuqmhZuR0Msu8E79WDDkjmVAVdOGSp23z6Tp5cqQL6c1vErZPnGL9lts7Nk05CG3EMcx
1Fo91/cbX5nkziJLd16Jc2d/KwRtqFFWUvVz//qOoS9Vf8qQD9hbP+duRZJBpjAodoY4pfnfBH9H
PRuH37TWGA0p3u1x2aUqN/T5HDxYcBIRd8PR5QV6re0245BxenrhXWM8VCpcc0wj+fndAhezhQ9t
kLP84i8pfAkAzW86mDcMtccgbqIsejTUyHNokhCzg6y0fsVgiTrjK7EpSccDn8AiK3DqWzCTfm9l
KqFd2c2dTZ01K2FnMnkYcg40to6bY/LfpOE7+tOHcDcj5VcqDIqOb9tOPXy9zNDzy4QwCOzNzsmA
dZbRMsU4BEcbBcfgMSP1zEi5IgiL3HAkF+5cjxWbPO64/wocWuEy+o9m0qVw2i4dXJnE0a2AYvUf
8Ude//4Ye77FCY8OXEnbcIRulwUvBBZyD4A7whVLSfvmV2728dXD3k+5kMVwDA2ojp2Bh7VGDWj2
v2csWlV/dBsyCjk+aMPnBHpG0K/o2pNbz0Z5Dx80j1Roc2iQekNvjvg7Urq/ql310bHJlFzxNwpN
g6xagnP6XStpIGSscIO9DD3AhEqXuhRqMjBN1Zt2H+RvsJMvcNXhYphW9GqyKMmR6I/OWcM4q27g
HCQMlarHUWN41lEz45b6IYuHDo7kLTCLx9THi3hogODdLYMxn3/l0SupmCtLKePu5aJFjRvx/QZp
v5b/Bq2P+Yf1SnUfDOUVJMMNk756NVqCUNJaElG9LJBNm3jlXxLkc8g0Y/9qY7C1f7ZPsOsTVE8X
r+0WKH2mN+V3R/Ausjp+BgidlTJt4ctosArZFQBSJl9dIW15FUnfjbJeTAsv+AuDr2KceqFFHPyw
kYptC2mfE8lstpOC6XvEWlsdZ96H1ZNg5MvIP/ExUr9P7lKVYXMgyLYmn4Z6Jo3B9zIH7/51nMkB
TdJr83YU4Plm0tGthheeBNVW7xmbQQMjkErljf32U7sgZvR1R2UnNo+vDxFiD1b03LMwKrwm2lsx
rOQPhiFDsiy+fHQhqOABS/rTIRxW55z9SWq6HJmbqGKaDdm1+btqGJNF8Y8DPqdt2R83zdojcMPO
kT/fqwachFixGdV3XOl86oVK5/BlDKT8bIy1RqODkEdGzNQ/cwWjpQ5vrvAQivJ+/055mf5qdEaw
uJ8X1V5/mCkfk+SCU2tOMnlesPqrBb6NW92ABigX99+fGkf+CLCHSf6PjUzOnJrsQSHAZWM1D4Ge
7tyRJVj/ICuiDb/kDLx0AlWXjRi+uW+ZmxUkTuXHwVAHUmGcMzrbvHsH49eRSI9dW83xDn2L25/r
kT+0ZXmWbCw8oi36ltF6NNVpVj/5fnnm5rXJcAHwgXiatRRiS1W4utnhXPAifEayraNrn6ySY0Hf
jpGBVEjWFAnPDg8lgUrn9RbWk2aX+bsutrZ9E9yFnKl/aAfTxr0L8RwtkueAK3I2LoZXIDYmCU65
D8aXDJAbqh7mY6pB8Qi+WPJbH3EqPGxdk9/GQl5u8s4fyACBwn6SND1HX6DEGAhEXZPs7Lgwdj7L
d1AJXpFi4KnFRTuScHhRan0/w/3NhR7ziP/ALxF0D2SeK8rlm37k4EY3n2uUevGhThPa947DR2LB
Owmed/XXUiOmckDu230NARkgg9J+uaN9gOAMXTNJ0iuOLkJ6G0+0D6g4hJ6uYTzE3vMtNcYciIMf
Na8Up4V9HbkoY56JfQXQxdrlLCTbC+vpx7Qr6+ofzJ7DXXP0GdWpl7KQXsaK+mwYFBv9OMM7ZK1S
Prcv6nl49fyC6NevXS2AhJo0+abhCNOBfvYvrQ7dBOnyXDmROYp8BsGC2VzxMA2SG8tM4kFC2vTH
S1SYZ42u3ioQb5eMgCR1EmIJQbt3Dp/vH+DCslupyQV9A6PlNw8iz8iAoGP3UPVmZG9t9RoHSeLT
jG3k+UEgqa26F9SI0rQJA1brfV6p0DTsbR0QdR5Ap6jd2Wn0n3gBHDLY/zWw26mzQrxog0yHV/SO
fye8mwYBv91amPoWZ6jTuAug2REp10U5SpZ9Kk7oHnZBbJ6kYr9QODHCafV8J1mooqsa2yRjoG3s
CW+7nfyJDwDbnL7I8PLnSLa2+UoVOxuYtJKy5yNsGkvZCQwg+gq+u4iefcovC7Uk/+EukWmB1qEw
Yu5gJdXdz7LIpCF1BqmlqLcAXQrwnD9BnuXBxFoWleR5iun2499+zkpTEr+Zs5MAS5lSNnLkRd5i
SllH/oU0mOM4K1GcWIZE0Qdl2y3vCSXzjtiYOBG0k7tZt1LPlRzvlqrNw4lkX7tH4SMBF3HQyO3w
hAPu+Gmw9WvlUq+aOimXa57HzfOEawPGqZy6w+I2LlF2OEq4DnlvKDL2K9Z0hHw+Xk+qtB0lZpQl
X2SLg7wLZHFV9g2//kFq7jkRg3dVMxddsg993yBe6NAXW0xuYAZ2qMedwE1pZOhLyhFXbDFf5Rib
sPGIcawPo6BmlBLctn7cDb5CrF2RxnYhQVM9XzNpB/vgvUvNMyjtoOXijZwLMjuPh7CQyBAuuOdW
YmvFVLGVOzyMFF8skXWaiAG+C47do/RPvMyc9U7nS4+tRKhbm8cZFZ3WDAdmtV1464zoE7qZd+sU
Oo8b94pfWEpDn91nEvyRWtB+oNhxAt/f6LzCVI8dWTuTr0aCe+d1HPsK5nu1+X22NjyK4Xlx/vjz
4QaUOFH9weQ62K5nfT2OBn8bsOSmzpwjyAytksoyIF6ULSx6BkiNoVksArWv5B1ZeosTv2bZZRpZ
4Ef6pu8VqkrKiJM8pL4fGl8O/z9s8w4ee2x+v5QnduvNvoYR7sZld9mtdP2rSkNYuP2fUb6MPjNi
ZXuPnuIIvrPCkpuvoTPwago0FptfbKOJdu75IU9IYEWL/X1BfR7V5lwhLpzp4Ng0TS7RVlBNE+Du
SoxWTinL7tDYTuVP5jy1bFuzFPGsYqLaIiOlxlN0FQupg80CipV5pzM1jMF5kZWM7EICrkhkNKox
Q4hffXSrFM4kgsQrtNF94HPShDXhv6OUaplqFnyunb9LW9ftM6FhdbY6nSZW46pDxUub0ROO2fdD
UppYHjJBgEhB2MjsKcqkNpTSdneS+my5SBfoIMVLJouBawSaM9cQdSRCJ13NjAo/J8W7GarTFp8A
Rqy5nR+4tZsso3U7KDDZtBFvv1+IN9l0B7nDDjAinVpXOdmPa2Zx0b8RUr6zvtlWbjeLXhGxeWMJ
R8DM5vudeDqjsGtypKeGm6iBObau2yv+47QJ8hcNt4rnPEfIwX2cqMo1GNyuC9DTSfDhvQS/uEZV
GHlfmnjVLeQdad7mzvvK5ufGVz0ratIUZbBQZNiGo+IV8d1WfCjWLmB5xV+WldlCyIlpXpOC7KYn
fFyUB6X4i4ebwNIe36sxZNvAkPCoyxLx/xMOojYN2K5Rj8jZeGqleeUjLKcqAWn6vDi1xMYRMjD2
DxOX9xVLP2p5y1L2o4qWEZRiGuRT4WyFYB+pU+3Q+nCWqCMkmeAAp1UquBM9yXVwUqoVc6qHakAa
TH38rXCfARQpLNSpq70Psr2sVno+2qRk7vxWPr/GOulc84+YA/QZ17iFuMERnBU2xPgQwK3TdUEA
baDu4iXWaNrULBG2TTkq6kaC2j9zovggJBFm28HQK10xteKKHxpF3SUsnoiQTDJqiwOXTMBUlaUk
CGXp7o3D2b+PWo1YF9DAGzxhyzO2Kpn6DYgXuEFWsv9/ShDSNiVBx17O3LWbDnjGH2swdws5WExZ
8P+5dl1JDUupuDQDGsRmGH9sG+1/yRqQILdevYohIOFc2Hrg4C6g8cr/ETmFsdBqiyEoF/F+xUp4
4Huy9TxBPj4thz2Alf1nqlA/AI7/R020cXHjUFMk4OSyhu15qs0wZUAmjrMzBZZdouXOXVbhRJSi
k84hMhSJQEPUQmkiik6U2uHBLM5Rh9wXw9sRWHP+gRvBogrDNyoKeZaCXDsmcUopaVsn0zahAPRX
EJ3h/lutVhyQjs9S/TkUqY8qcJbZ9jN+4i2o8baUh7s9n9J8DCOT8GDIvcGYx5GfBISgKm2kMCGx
oiRj1u9CSQ61hd7TzDz/L+fvfjmDOuT7xNE1mnp/jICkK6O46pbfIddknsFRvBLQlgfj112tDhJb
4OkGvMnIGc3QjuhDtO6LpwVmD2rxpknehSVHgL09FFHSGfbOOkPLpANx9knoQ7hhd0De+pVzXZSA
ePRabpgdrXP1W1V/OQslJdAxpI1oyp/SkJ5SwgLY7NuAU8jKQ8ifnUP4zb+qCbMw77CLk11vkyZu
WRieJHiE7zm6Esr+NZ2vP+g1+j/GvYixfriSjSkPvgiovVWEjhWXFi9Ix3jWJUmHCCv/WQTt999v
mwy4wZ2k3OvYjb9KFcZemmdYS3/xhoR+Dyrar9fCsoztEYM2tUrbXM+WzP9g9YsNcDphvDUBFmzf
lkLfZxgtIzZfIA6OIUI5LPrO0ld+qQ2OWWc6JvyFP8i1eBh/DSkx96BZeUn39xM3fYvToVqS2gi1
7XFDxroO0sFk756JB20oiYOx6BrxmGZ77jpDqMiAj8AOpH30HeI6YrNZu2FPXPiISoLigeS0/jQD
tVmppMs4l4N+HAfv0hSN1DFNKhky+EPkLIJHaUsSZfv5OhRVim6R++dODkBCailNngQZwcaSjR5F
MOtb5/q62hgvlCLFi5OSMaEhXAQqJsHcjSDRZRHYhXR7xpbVaOqZ2s8oG6o7JdaYuBEhfIDiHQ+5
QUMnhrhoHDlYH+LBi/z4UF+vDjMntV4XYCcmZWrv5PJVMp5fG+dH2snOQwOjBhyxtBTSPJ/xweyG
OyJ/+exs8oijtvD50bU09ZxbhyDZmhaHhwE7qgiGYoauZ45hhG2JfCJopPeKDBZAzzewfxe8/GaP
z01Lw6fRNAG3p5HPk2Kc/8Kq0VEJEOrn1N1Zc5Fg+clC9rOhpRpFSuGn4kBMdCdcy+CZCa2UwI+J
Q4S+cwnWJFoLDBJCQ/IARlYXyvVSKcMcqCb2qTn8LKHuvsk938s68aLinM2as8/nifpBZz1BAWWq
3zdoxS9KtIEul1Wb3/tIwsCjWsO903i4OpCsvC001mv1eJGifCYkmMnPMtns6fzWJhbWPskE3sHL
CsZ9ySqGaS3aCnNsxIIzpaXCDR6DHJ1vHG9gq/kTGZIZRqeX9P1uU1bl0VfbMaVtUBsnfKr0+7A2
CWqhOctMje+sBtTnKS+7X3gijUY8LSmEq1FEEkdxKpRDmZKhYxQ1Vc/OUWsRTP+8iIVkyyqve4LK
m8Lj9onxcw9pTts1upd470J61+ne2zijOb6Sl5ZS9FtcZTPUaxsLgy9l1ZA2Td3LceJcnltS00Nz
GS6RseUZjriifAX9h0HBgV9Mmi3DTQqnMYIdvnfiLisB/jsW17kGo+CESpE9Z/OueZPaOzN1FbO1
RzRBvY1ny4Edq7iSGoWrAsIAWtoMj/81ePi6ykTD272SJSBNNPQEuo9EzTXDexvOZf5cL7dFXGML
+rofLbQi64WXK1GMO9XgshbAmGfo38XkXOnu+Fa8TALM3iNmESaJm/NTe2RAjT1dJcrWuOiIG44J
pyoUM0nDq2s9LG4CdVOPt8r6HfUFuQMC+kIbmN4ZGJPW4+mCb+7Z4XOW+oGmcthrZ2FYgW+E9JCG
hNjpF1v5G+huPB6x4R4Q9ATLRIYbogQYzYChiS3+DzDLiy7MQziZ2EEBSHTr33TMHyGigy6sJyxQ
gv4FfvljLcoW4OTV1n0RoC+k+/s7IJ9zfUFl7TTYkvKwiGCMMyh+iL6BIgwCeD7TIBtCIrBKSiQF
MhzA5jY02Len/g34no3uQXwxjIbvDsfurXcIpEO2/MV3uiBVy9kaGVF4lHPIKu5kYU0833RZNMc/
gZ7Pj3a6Ur1WqNfAzmzMY3QR04kWFjldOJR0PkqQz3P/v3CIlk7sVmR+CrUTq5A2z3r+TnaP4QyS
c21qmp/ofF5bwQpZSEgEBWq8NSXL57mSFRG6v2Ldz/x6GlR7H9DAma9ZbtLzqY7/sAhG0A/GFMAN
0gNFNZ9mbAzDE/cAr4A5pxPqzGj6xRx4+291y8yocHzX8HLeUOQIPm9S5tt+04TZoXmxjiUFntSm
NFbfQ8rRv9fwLj6HgnSI1UgBflP92O/UrAKXAczI7dMWwHh1zLg11e0xVbVuIcV/jfPapAZBnzms
25vuy8QSkewunHGbr/2BORh2wxkx0oV6SNVdUIeqVAaBLUjtlKJ6P25Iad2t6JZ/CdaajrRUsT7P
tcv9H+DW+iN2NE+/Ksntqe+SXDkjF9YeF+6kDQRtn/2XniiCnz7mm6oZoG5C3kCMbArdXVoRfdQw
7zmqN/hlIpyBhljoy09AZxG6TDh5sJyLox+N6599sde2YrJYs6LbDjE/Zu9WC2T3nubje8mAqZxv
1jxh3TB1EO0dEr28eaUhiGYuzHYQgMFzaW98tnqtE7rke1c+gPdEfgtmbSW1kt04WRRkeYvMvJpj
jistYwp8neEUezogQQnylP7hTD2mxjB7QybSJ/aIZKAH7bEG9PlDCc2Q3Dv1v6sBBJa7s9rF4WOd
UlVbQmbFBUSptN0YT2bVetGHi4YzSWbLoWCvGqvKkr+4gP0LPGsFQXg0Ykun+vw6VMS8bezZqnU+
xEGozXFn27SFVKcLtuCnAaxlAQZquZzDK2ihUI9rtg7hMKB2FFuqL4FJznSsHFOQT9b+oPOCAvVC
KooR9Frgq3DwHCibQqKbNeZOLx7XW3xPi8/SesIHuFr3SVP2si8QzhWLjsLYtH0EwXdbX3Bqphdk
YpLiqJNPRliEuBPQMXSTicgovDwsD+rE86ZSVYw54GEFyeCOYlcf8JRD+xYd780cM/WEMaZ6BMjd
/gE37uwXEsFaJNyQ4BxysyOIKCrmrADjChtx4iDWLP3JdUcUMMqf78yjo452pCG2Tcp/DtduA2q/
QVT2JIjTUZtehg+dcfd+uxzD2cqyHHHUnlSFAYkNScK51ywOVMMzDJV5qLv9+zB62tIxlGVHlB8Z
XSoVFbsga8G80JlKT4rUB0SNyR/AdAyso/zTYBCaT8qbAmKcGyHGJwX/y66miPHX8t3kb4kzxpCE
RJmbgZ88t43lFpKADfDUuuB58XJTGm4lKRqaQ1PytYLufH1xYzcn1S9bE+emKmxFZQHfLhcpTZoD
4D7ujtraji2Ee9w+jvU=
`pragma protect end_protected
