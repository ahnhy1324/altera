// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
l0FKhphswtAi5/y31Yt/Fux3b5cGyxw+OX76KGrxx5xuyOvYG46QU1usuP/eCQ09iLySa+wL8V1o
4DhQYqEx1daB4N/+MyyBGh+MyLVUzZTvgceAPhYuidoa8YJmW7yFA4gCKviAYSkZ253hf9JaoqjK
iHO//UeQpqeZNsX8M7b6aXXAW8V44zDeOf7kKZwFdUQR9BR+1Iw3SyXbVLDDeBRaMw6XjgQ35c8/
psPlvnjmy9N/V+y6ZO+HGHSWhsVSUXv8tK/EleBZMVprBkPY+tDX8od1wAV8lb3wlLhrNvPRYgAN
w5ptiJUWrnG0R9TN4M3CSrqOZ1/1AvYEINskgg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
rj/7mIPrLzNVdWb6cB4XnJUuSKsMGFlHZXWTetgvsYgrLQI56Gl9hFJDpSY4KjO//QOsZjjvf+3U
2UmeU3IqQ6jplNm4OX/5cmLq/mqCDb2upyITms42RP4+tfD4Xs8fgnk5aArw7BkWK+zJbLr+PO3V
EaLcNJXTcWJFL7J0kZS33zbD3l/4c1aeAm0R1Rslf+UZph0SSFDTXWuK6gds5cLBRge+d5U5YVuS
N3O6+BLgyVHTBGW2dsQf+aoaGTBwhSA25Qqp8hKMOY697qujyBkr/c5ZZfHSR57XL8+7t3rX4WPY
/IvNa6/222NkdF5gSyB1bSf9F4pu3ypET/JGFjdOK016ZtRhJhN981l+ySkJhqQoOz3xC5AW4u8r
x10iPavKV1WZEbO4HVb/HnnNzvt8bstgb1+1a+qnCFIvdJJgDZ8QALZOr36Mda7wsbFcWFTQ8ZnZ
UgX3je6lBStVIUH6cfUeU1W/RjN/lg3Pt+YqsoX4l7ZR7AUOGmW+E21DWlNfy5FihKpd1rUiNxAx
4eNyMt/MuYV7ucWxb8sP59T2hpqKd5axtPScAbSzvTFdHwlQ11uAyCPKtPviRfTu0ufMbu+/Q7eq
c0A3NKpBMUln00Z5cT4H4NjEU2aGKYu/80xVae9kmmzJtoICmrkgzeSh9IXvUa/EYQL6SqwAZ7dz
aOhRd4nUWJ5ya35yna3swJ2adE3xAVblYwex7fXSMlHclSC0XKWcOjqkI9c/f4RXy/TF8K+aavtW
V/YSQsWNAWsWUwY4h2B+FsDUsWEMyXPj+gdLLEAJL8NI29PZqeugSfEdOrM7ZmbByhe4usVMZiml
eyEtX3K3nLwRDHb/ZFmLhxxmvr+E25/tXtA0IGGo/+Y2+jHBqTW5Di9A3GasqfrjWH0j6zU7pOq7
zRwTOwLr/6/2niJQ5bIVFt4e5EFdZ3XKpF4XhVN6+a1MPmtHxIayJR2+yP0W3gXY6rqDnni97oUd
gkuYqhw9Bijy6sZFlRzsMdUSTywT7tDnUjEW9Z+QHTnu2K+NK7eJqamaPq8lXO4aSngP5tRCfbDz
o44jeg3HHIq+ndsQbZOAkATJTvl38D+hjxGXUFX7PLJtvfZ2sljMiysPv6V1xRrqmOXArd5T6NXg
P8WMjkASvkwzB8Hepnn+lQlKyWWpINdhXF6uUtm9VIMGNNjbxDJtinZQmoYnFJIfeBaq1fuUlcwM
HBAu/O53wDmRW710BYH0PH4dGuJb6OvjfFvZxS3WncK9Wc1Mo2iZzo/3SoVSG8taLMjm7EoX7JRa
LeQmWdjX3k2sNv/xe7o4LDrwq0hMVLFqqL5DAcnpeVipC8dTN1ZQputZkiDedTE4dMF1TN0T+tGj
zdJf0xR7MvQ7op6Uom5WfTa+GYBT4l4SsWV+55ExL5U1xOU/njzgVKQCYr4S3Op3oqbKpkrFKj9i
nEzr4Fm2pQTU74BWswpRk8QsPMcQbNnKFQHuQqjeelCm1ZkBGCJy+Lhf/60mMdusolsE1tskY5TN
hpqTV6CQTU6Yu0Kr1W8+Ccs4noZGfBGTzcBuIZfYg5leB/TcqM+2DNtms/xDUvFnE6JpVXkUNzgA
PsNvgaoMtcr8DcOa0W52IvpEuBFSgZXWuG5UI0AmVicxydugn+ae2WMixI8RRetgGaCenM7eAaLZ
O/arf7tnPt0klUP0NvLYIAXAnDY79ShYGm4+5Axd0TA+0kPROu94dxZUUVYySvH+D5I+HcrSugJ1
/grwim1kCfmc1TcHfbUcLWCHSmzGhhSxIcpWYIb5vkyeuqcENvkX/08f22VucraN9DagHSEoSSMY
7QIGgIzV6PaEqSzrgJWGor7O+KGh+WLQsCCkVyIZXM7elGg52rPHIHz9XmYX6Yeer4m0dwXoKFzN
eLi9itCrQAaybc1mkU/d8KVqYar2eky67dCiNr31QhHSaoG4T19UOlV+4oAMuA31dJiJq/e1ivGD
wzaeL/PEL7SdcQFQQabLPVBPJ5crovbJYGMj00m2RKvO0uOmaELnFNGUZhTVr/SuCCva/M+cWG5/
cyg0C2xDrqS8XuUvThnQhIUdZKFmOff5+SQ+dUpjwc+gpt+AvPJH8gNjMRN9CB8ZidAdSvlaMose
jShZhgx7+zN6rrjdpOM9EtoWDbDnzeDM47r4uIxz8MGKFK3cVKLaxJTQM9uk8raSslkRDQ5M93/K
fsR7r9+d4Dy6sYDsV8AB6gDQDLe0a7zdvjtUMnhqyBNkcGRVdBvhsez0yz62rPGl6K5lQXTU5w1L
d/qmYYEvl5mmNEHVSSqnnFZ3gRjMtDwrUq4GTmGIRBI32PuiJ8afzHT0dVEZglbJvBjgySBFZ8Og
9htgZOoZxxKiyNz3gSJhZtcqQKCfbw+BwJfyzqj+p8mePIdRE6XQQEoHDfbfLoVSYZGzrLv5Wrzf
mimITv8dXTKiE+zgwgUPyvMkM2/JmSZoyprCeLKyOincWXShVxvFBk0ZYRNKpZa4Gw6Q/nJkAFK7
JKKWImfrbuxBdLuJrq5c3Bf4WZqScANRVCWh1s7rF2S7PgbHN7JakUyinrFGBvlpBYUyTCclzoW0
L162nVJ7s+8VFyMAZTAgOVS66F8tP3i9olWCSo+4fZTT5WteYFS9T0iQM+mAro77e3Q3Ka4bWUDX
x5wc9WHGTyfx+J82BUYmjDhcmkJus25oKL9Ey8CjonShQWtjrp9bwW8OlPH2N/F5eqXAAX6pa81V
tUqrPA1SNlgiRndkS6rWDf+lq79qtoqy3v7JwoM0QAiNzXxKMFRJBFEqce4Kp4kGc29LbHyJ6T84
4Gce8QZuLngltZGBL2wEw8vF5t7YGiMzHigTOakcw4z/L0GwdoKZRzgzXjosH+XGLET9O5kILNJI
sSGvLtl/UvSMPOsYZu0Wjip07d3ncb5tj6og08x1JX1RpM9LDBocYvoTcmSYZ7hpu0ANVoQU4BRW
LtahXRRo63QCe1hz2cxS1MAQXB1dVHi2gf2sXTui4o2Q+XOxMHj5gax2+PBUGAiIB+zvUVLovqBt
jYpH0VnjPKC8b4eDuxSJzZgZeclflSRNpD7IOAcX/m5YXhpQ9a/vlpYsJ1hkDWf1dCjzUa8pI2Fn
dYBM/HzvclhYBt4lKdATItYvmWcaQAHi+HyZC9XidpfDUi5K9ANT2g4q5ualsLsmNN5ssdDqqyQz
r5WJQYpEv1a+fJCo2EhDpcCQ0Gzsj+Fm/U9d6qBnDnyzQv9KJRtyIt+GZ5G4sPJWxpsqcjIY7Mje
/onXpL+qsZI1qpQzoDPqf8KoAL2hdOznadZYcfjn3CsdXq+cv7XxOjXUWKKdsRUewmFmbqUZeztg
JJBg61WJfBQXtCuPpKOnanutE5IsmAMxiTYasx2zO8L9/vUUN7FNAPOGBawYR4wc0ajCP8sNueGl
OzkdQPNAI0XR0RIRO3dF6epXY5/xvUiCYVsp57KagZtYLhjlxQ4RBa+4fn1hejoIGkJQcJGyuKQH
QAbEkcF7RXvqFAmZNKlMBV2mTArwaoQoDw2IDDmTdDOOROBAemFzbUH1tuKk7/Cx+oXXYzNh0Alt
odICErlpBeEyGfU9HFm5XpW5G15xCKE7+T0PwK5x8+7nOybvyQ5mvzUptZ612XshpWbRyRahqueg
HnHeyaG0PLIL00A48WeKO1KeokSTewzmQj/SLB12Py2YeaelHa3OxTS9POhm8jwXxea5ivByOw+p
D7FpM5SZQxUQLW91Ka5XdnZ6/yoI5q9MnyMrihGfLfA/4qntk0hWtiKOaoYW+l/6Xiajx6vfWnQv
8gIQM/pfzxa7ZiqwfElNcNnyn9g85QF8QuWpi+ChsYzu7PXpuF3JkitcmPmfTzCp4dwm4qlThBqw
abFdSwKyf0J1RufghTvb0p7ylctShX90Uor714REy0Ilt6usFb7UUzdmk+ePlxxfABqzGQ9tmcLO
XLl+etHcGPyN+uvG6xF3ufDrBY894D7GnXY3PyGwIm2H7j2NoeqeWodtehOKNx8PcGeq8Ochm5Hm
ns/XCjqi7ijUcOAIlNY/inQa2gS3rATisbGH8Jj06nG2WKwbkbux+hXt2EciTcZMapaUsP/g8Nc9
w5KY7bpVjODEAnMaDQa59oZ3hvRUM8vnHgPXE+ZfBqzp+TPjcbE32QBYUaNCUfbpV6bTmC/MWNMy
G6f9VuSh9qSsHXEkkYiFgcfF3AUL4P+pTpoDzhDP60eE50h2JtoSjCel9+ym6KIPTSC95fiMOPO/
+p391qdbBTMmVVBDRF9oC3fyWZLYotaTiIqhGlZYblrLG7KN0CgUFaImEYXMjJETPS8YMEK9U6ea
OX495lexW9EturEMh2QgC3VEt8KBWeq4dJsmGsFWrk4gTqwR7rGYM+0yUJ3m4MvEd7GxmrUSKvnr
qts9wc9CxV04PQPm7buQEoBQuQDQYGO7eQz92DBpU8cX4vWHSkwSfZx0RLpRWQ6WiXwS88mYE6y8
xNB2bLJTYkicRDNWaqL8xo4LoU32PLFyavdUQ75v/qw2rQiBX+rH9JLxYIuVevMcjMPwbL/v/hnn
q6tC58gmU72H8G0UFB7QmEdfQYQExLY6YcCj2RJt08Ax+C83RuiZV4m2S6KyE421Ewok9BbRmliw
b3oFdCu/WDJJ20V+ObUsbMiIX93/W8Qiy4Lx8WGUd13xFudXCe1Rj3k7Xex7cgd229J6rbsaACDa
+oou++ZjPdofcJ1WOzVtsR5NC8BKWDbyp6VWGmMg5MSPeehBAHF+gWronl0OCKYXbZppZJyytvDP
QahaMaf6y/oFgKVep1tg4rctOq/51CR8Cu34nJGSVjU/k05zRVKmS8DmX2fhmEr4EsmuwmWudOGo
Dkakt5UsX0PQGdkiBJ9Dam+ADbwWlG2aZJyWTNNbET0LOBPq6thIZE2wzmryfbJeegEbW5FPIJGM
C/aIVhSRSYRddjNJKiOu0O1E85USLNjhknbLLTzS/vzXXLtkUjyQxnbqXFBT2u+rCP4edDlZLlPI
ut7zPSAChnDGX6ZTnUMLJdEDo2AwQE/3JDa1LNwad93fuMNmugTrkGA22dpLDRIheinbK3BRmpyn
f8m6vwKzUdm/s2HAnAJvxGPZRK0fFpp8kYObyZCXZX7v+j+Rh2UzStm8YvWCdzsasGcIQVEtlxZT
Pq5zudwLPYatUpZWAvkoXMrs10LqyOHICXhBRIQDgNEqlrvVKJhon41jFAFWYYdtmzqSH/9MGfY2
fJdEu7EgcGxqYH+8zi57/C9MrFhUmASfuKwyO7XcgxsxSz7ScO7H61466sA1Zhb73l892sdFXQth
2tQXBMIEzaW+61pfBVg/wNxC2n95YCAxSn9F1HQwBDRj5WgyXpChJTSdOYnta3hlgZt9nGReKXvv
JI2tjEUC4fNuI9BGsoazwIfXYGXpKrjUg9iiyXel3g/K/Of94KSemCf0a4HRVukWCwFh1PbRABdl
s1zp+8ZEGewGzlEpvIi/kh5TeA0QNGeaCxJXS2cMtoHQJuvqkg0xl8DfqRIn+egO6S3uGJjpq2hW
0gLnS/tqa27LG+VIiTVflcwaWAPs90jGtOh50OTVFLN7JHbs/Arl6NFXAEHIo5WmgnuPTiNJ6FyD
s9RmmBeA9YMrQv3GF6yQL8V10JueXYunxSScQmzRyRGX7g4XnY5n14fv7Le6rra5bJHf/xG4stvm
+pTEXoFDenaS04LQUtOmrV3Cjq9D2nl/dkE1orhUELTZ/orNftcFDDQ9eB/UBzeuxCahC8cTryjJ
JsX4vdHH5RPMa/Yw4AXFrvwMR2LKH84Z6ZPJeFXWuUQUDfvFautsNsSBuCjUkUr/xNcV4VFmLVzI
TvEcPCui8f6Q5FxjnnU2HufQzvKokrXzp0R5ZWI3Wx5iDY0UlHnta39b0ZzI5FPI+PKIWp5rfLfi
im8sl9wM5eI16U9Kh9I/C7RS0E92qldfIcCSAuJerppwKpP/31v8pYhJLYGx1QsackpbaBAn2dp3
BJNE9y58IWblhpJFuirXbE2S1r1lNGTqaIOFIppmlGN6tZ5hL1Dp3z+ybFibVNY3NnNQTm9W+/wG
cSQDnjLRNEA7PCmrvS/Su7KQU4dyIn7cs2qZ6TlXkL9XmpkJNsbvOqxRd2wAyF3cqfsXu2BQAsA4
DksC770Hhg89ZKkkF8X7yH0Za4M6v7eg4mXrLMpniCTHOW/WuZNzCmRbBrwdTxIMsEsluvIWyk5y
s+4Avd6hgVaU+hjFvMeuE7GlBK1A072lffDbEs6LjMlxxUCb2FChPLI+5zdKQNw5IUzZiAL9WxKb
xwlbjIZ/dm7klaWnWI/l/fmJxvfRWFmPCBKD6gJXLtWxwhG9nY36Ard1G/945T92GKDkYMiFqOul
sCM7g9CjgTnLzKYZYOHDA1YzhI0E7tj1pEp/m4ZdjFI6d0nel2xV8qiOcq/kiZfzVicrxB5wc61v
HKtKtRkWuRSYm1sQtsr+jIeLGRJHx11kNb60SRyhvdgtGYwkZSFMpwlnIX6O1ubHLCljYcdkoVbK
b72i8BdecfumY/bm9mgJlReLulaQHDHq3AxRNYvK7tW1wr9CurTbqezNYmjJ0CYnkvqoWAPdl/+f
jeMYRrQ2JgrnftQVkCo8Yxwb5R0H9uM/SQY0kjkQgLVcBfWJ49S+FUcwf3Unp1kduC13sFlJSy/a
bMICDimBbtDsXFoGI4p4F5Cf53xmOZWssvgfweI/aUhYpa08wzbgOly+RHw8+v0t1uEf+q7PTRBC
BUMmUHgWR36s80nzX6/I7x4s8lQcdAOlw2DS7Rooua12PkY0+eMIZKtD2upIrSucj5boXaRM8/zW
gQ0PdTc5yeQbUc+sivghBuSPOGRi4lyCLAFSHivBhtsIXkz/KxoKV2zKklBEVj9K5BB4Lqwjm3vT
dVD3Ziv5RocplK1vt/ymRY+tNngWCPalskeuA60uuQVZU00LERYPKL/4X0BKO6/IpUPaKg/evMN+
QR7uAeru8ZFTsw6Ic6SJc4C2fvMzy+SvORapMvGYMiTTTyNtsHeriKLoBgpso/e8FLgDOXcGWynz
ZPceiZDcTmOID3jNhsHffl3c62AU5MFN22prPVT62XUt0YNEESyLNd5uQ1wpmUqYmYJPWSkBLm/O
EbnmQ1U4vsSEMGU8pgM0nqIpquuZ7A9/drq3OX3Vxu03zgK+ULNJvH8dBMowWvymEADCsUaBHDkI
u6FJkaRc9sMs8hiIHzBnRwiKCFpbmztwjvoxY1VCdcM9+Ch8o4cciVtrxLx/Cw58zVPAiwbvI+XS
IldgLXodWfQ0UO7NvDPowjVGrVzcoug8SdKoyDtdMSaHSxjXzz2asLUPbSGXgoNmI7ea+2tYf2Xl
gcNBumIwH9YdrESxZ+YEjhuf0xjG3AEjzebRDdnAZPdNAgFBYe4XVL7YT7LE3mINm8qR6WIll26R
TLnfnjQb6wDkSC6/SuzkeSsZ5BjGdE2nkPE+PoCtCF0sTXCR8kqMKdgA3zY2Xtxf9mebG7X0RjS8
YEOE6/ITziBje4qodvBxyyM4kaXo8iqeEtoM80lK7sPTHTJ2/YpPQmYkAglndu9Ccl7FMybZInJ/
tvcH8uw1MEZGb3FYcjERJMuELCZVwxJOzDpHu94kQX9RDmhNG6L1CBovhFRRxcKFCMqN877KHtPu
B4C2yXrW4SML2Xwy9N9IHGtZ+vUNWNWwATjJhUMeyhIizGvBLIL8VNjdZ3k2t3p9TrQM+HfI4J6b
mNSsWsDeIruqneFI1EVy2pJ0rzzpK5yMTYUdjssUGv1bH7Zn9O9Uyj2wfjFtKs5w5CWMB8+NfSD8
m4WkYgAUSUwOLwgCOTlxfQh8M8CGBYQvy/VnYnpsA4RsA1SMUyGnMQU05cy2hKxvYUwlKeSnafHq
exYhqMNIHnCwM6wHVqiUQ9abaTkTRHLi/ReXKuD/QbwAYF3NCzo4CsauNsBvgESZtaPSQUQCiaMY
9TDL2FoITp9Gv4y4+mU4fSpEKrdDEAGdUhetAjrL1qbaAdXquxnQ9hpvoFJK9/aCkfOqeznT4EkN
v0azwf4QBueT0ys5GwiTv3JP0kybr8z3s2FP3vDN4g7qxMyOTC2ZSf0tEyZ1WZWplwUMXL1Qd5AS
FjQ/xg5SjiEZcPkahFn8vATNj3EyRussmLokr6XN/ahyvtG0tTDNVy8OqzbMMKpQYfv6fklF0Y7L
LRlYGIz/Vy/w57pc2D6HXwZMs/1uJCwmIQtLQcO7ug7XO35CKesiPGS4aMuC6rz+PJw//x8K9E6J
+IZissQ2LudLfP7vuVxKZ/7oEWFZTkyFOpDqVAVZ0Y8nCB9jbnWIAqbpUTEpYwqFWM/Kud24O8S0
01hD34wSfbu3tP73ujBvYeH7BcTO/ZNZXWXErTpc8EudDS+robGaINCAyjeCdgVpQ7FAEY62p5zv
VdM/HFXhqv2++ATNwVW1Rxs8TpMBj2khzT7ljflDfja0kKTxmGpY/qvlbIzC5YpPzJEqLKREa2rx
Haqqv8mgaZySbx4YVUL5inXQD3xON+kIV18ebbsLLt1jrS05kQx9QYrPY1mrR7ZHOvSAn0cSCT/+
z4iEyJJia/cTXWysKee+am2g6RSwVEZhvZ15nqScYVfH2KvU/ofHrqOf0gUfGkhF2vW6xZ6lNoF+
nMt0IGtZLCHQ341V8i57HCb0TzhM1UvVtnbEkPSx1JAZSSrTVol+5hykjz83JZXHnHiM6CzLIoas
FD83bUDrDvePitaZy8SvkOR/TO4lj2JFWSIwSPSX28S8HBaa46YAzdrJ+HsN4aOr9hPXA9ck9p6o
NKm/118yj1D0WXlUdh2xHZscBUol8XbH6v1ooBKAJ5nzWZjbJo/JGxsXPFhmLZH1oWsdJu0/NTv6
3aD1+NujEwXoEdsOM0UjHiUMfPMLIa7LbbJw2GW+XBBwwUK1sBJxDDLvFQIxPMjJWA/EHoiyLC2F
sQYGIF6nbFBNuU+xiHx4U1iWIoh4clfnGMWdshJNs9MM8tjWvcjxzOhL6qUDqoORw2IJtXAIhqwY
MMAFaKDg1PHtHElF/ruTBY1UkTukn8GhP4DRcbF/Cc4yFdbAVDQHJ9ls17MgmRMTWb8jMdmHknRP
zqr1iLwyVL+i92uNuao/8CwI/+VSNeuODRmgQjApK6HbVIaqZXZ5vektayOtkjQ0wwLsedSv/7Db
QXek4ZbKkxbu0q+zZGwo+74jIcn1hvbp+ANgN8NOY/C91XEviUYGbbZU5dIryVRyq1uJAoFR8Z6Q
yx2BvUAu8Bte5iJKytBCzvnYdG/cmtcTasTZy5N6syWgUtLHyhW8hF0aBxuYsrQ1dKZNUATcGUjw
9YP90w8LqqIN+5GZHNfrV461LcmYk4rrqh1LQCj3dMzuhPGYB5XIy2W7/kCA/mgpYYAD90lCKHUR
6tyQOAIHMdXyScgmXQI/zNsfvmj1D5Ptk+8b+RkmcPnjB13NTEOkmnQXRGgGwiAWY8lF9jB40rlA
HALoERBMmUsb2zhbmBcIbZI13vNakZ8nUiZmlSH+frkcCP+KmpUs0QQ3GafsgjFsy1TFk4EAt9oN
fNfkOJ7VVTyjgdnNannusLXWOC2PlU5sEkuJul95zbwcjIuipgCZ5RFS3IC5RNC6ww6DRGRM6Hoi
+zJADV4ZoLGf3K54c4lYD2g98rrhCSB5F4Qm4t4l7tpcnIQsVEB3xezGLYV8A/gqe3ZpM8W+ci97
rcoVNSTx9180n8PnsiRPSh1OBqLbe2wiORFWb3PD0mJ+8auwl/AWISPU45cBgDtUSTgiLry+jbPv
ZD00JppoAXWJl5zEsatozaqhMiZ9hrqx4PEJ61pCvywlY3NR96LAPrseZJla/SOhrx/WUPlnWcL0
h43GpTRuQtQjnyD8anbJ9mAcmag9y0bIL9zwvjz7+0T9dTCGtSHrx9MJORKhwr9SKXMNqHPsZdfZ
cM0avJUJQnklfXKfeUxdhvbF6TnTO2wbEQG/gvx1lR57wUWJAbs6KXPgxWv/SqvMhgIwV80IZdej
Ba0obnHbBvD8rCJSd/RUCYLrZmiZJyBIT6paeSvfkwt/o3ZcoolgTqj4/Deessuyg+aHnKLcE8yc
xqWt461o42apG6ioiaCSfvRuh1tXlOZzHRFeB14t4Citq7hK57hbSbyZUbSNK6Nt4Jq42gVvs6c5
7brJUnSmwpVVduMGy8D7z4p20m0/E+MWM0PA9DLcZdy7dXzQVhV+c7VQNekwVui1fKXvVMuIjYLI
nIh8TjHHuC7nhdWfhzIBl0e4QwGRkfhrcxZWsyt0uHjiJQ0xifIVOuLb+qe57BIsupfa6AdfLUoR
9AKZn77jZ5uJvLvCO2UBEDq2Che+8X7GfDMjkNT1XdRVh3WuATBWvqcfuWTJMwll9uHhmXjU55fS
8rvkLQvUNlcyaJ34VkqM3ENZlMqAvLfyWrpcGg8F2vsZrKf24qg8G2QIQMqTpxuYv7qDADx96OsR
ClCRBhmu6sEq8S0/NZqw2HLxb718zrBMpLy2U05n4Wdw0Amz5aHqAMrmtSwtbGiAdMkLs/o8V6ut
+FFVRmlVwCUnNYnoMvWrAhvzPwoX0DvxVKiZPu5lKCsoFeaVcb52+ViuV0z26us9LRvamgfJ0WXv
032tRkF+HP+pmGVxjNMvZoyxZYUSQqemamZ58Wyn5z8I0XLA2D+X36276RaHnPB8bXrFmp/xQHsV
puQxbQK6PVziy4qxuyq0hUpZiLMXhNbUijYYgmgR2yB2MzLunXdYv9ZQ0cIWYSny/1uqoUDL0810
XnR6F1C2wohd/lhkumg19DGWg90OJYIwo/mEe0/R490+ewd/dH3ym9t9helNld6WX4SHKcquOgkC
VrHOHGqkAssDgIGJkJGD2Ehske6u/AXzYASBzmveKtcdgpf532uMOAe0V2R3b8Sv2yrPYudc5arw
GT6sLR2q/oxJDHxkrPhO2GrCaV8stD5YAVFiKVeO6H4L6pb2fRu61byqLFpvizvUU6KAnippDPyA
OBAYSCCR/ZT5OwMC1FC1NAjyhVXoMoi7b3fNLdo8IaM6rwceUoVe+W9rqtB5hEaFskzURaGW0neV
M6jBX7H4Lj6011qnGszPM2SQLaflWVsViBaGJ1rIH9pN58Y051i34aJCPrstBHJIBTm65+w5Mej2
EuehHEkAj5DQ0fjAXPLNI0Ss+F9UZtVc9PK3G+rsFqOnFtS9ifwtUHHj4Ph4U2vX61Kp7WI2cH0C
YNrckh1o2u08+a1r+EhtOu7qtRiS0iB+mGOJntftLX64BNXvGRo6N/CpqlND5RpQQD9aC6iivBMG
Fwnlk2O2/p2yGcwlpYi5n/RNRtgeZ10Xlfe/QE9vtBYrEzEk7I5oeW+um2JloXOEI9GtjkYPvzJq
XIzd2i03XfNmhKt2nlh60H6oroAtNgJOb/wd0t8ELTkEM/YOMyRbRG7SO9YoDKeiYqKaM399+BRk
L6TJ3lobzCt8TdCrKgH+IYf78m8euIIDOQIeKiwV5ko/cOFzz/444GuUgPxJA3T4cenOT+1AsCIX
gXIUU/1Avf0qtCQ+sJzm+VBNAqTNPhstglkCPqWJWye6VWLQGfD0HExIsvEW8bFDRduUeov8kKTA
NlPcD0NLCJ/fTYa6Arz94MUWvUVTuDrKpY9892Q9oujSJEgGJypz1/PyaJE1eIWS0P9xjO0pkV7P
j5NxIDtzIfu9A/Pl8AEgUPIJRpk68pYH7uIfROLiiOOhjlIXIxFy19L018KWXyDvxUEE0jFUYjDk
2yJh1I3WOMHdMnxBnHFSjWzTA5GidJRY4p1rZ/FtUglIiLHEVVn6gpOCdHzPZWTkjAbQThAUgwm6
WltIctuzQRL+fLeuVWGzZSiAzgsawEwVFP9ZQdavyP7+trzZdPDYrEIO8XZ4QZuAm1siPZ8r6Q7U
h9hWVcHr1Vjy3cRkILchmDwSSDldMvK13S/ErUA6R7VjjCclFjE8DTaBHaVAMvRrEj8GaXvGW63D
jerVBizBpqCVNRKACu3LHZXXzCFKGjTPEQgcUlV58TweZZgI3QLBE4I3d5UCxUUGY15uHNDBgGwC
53GfUNPeJknFQRiABjH0gcOxOJoDK9s2W9zVh94dhcOm+fjRJzpshrIj9BQiDo6mnQqLR/u1Y482
2hvv0ORW6qazx0iRpfL1eZfWtUEDq/Fw7BUKET5mRPTpY5xrkWwuIL/vhXWHup9RG3jZrtsPmIbE
Vysd/2AjtK0Mjpizy++E9sx+hKPsG1fs95SD5R0yBiAgtgJp6yU5fSaMWCv33TV8zpPBPbZV7QLV
OrDKZKX4xQ5Zy+JaNEHzLCzptPLQDWTNzbkvcDNv/PJQ5OhPNtrCYM3DhKrBXg0FKEgXSZasc4nw
r/ymDKAtsCzpkcvu+E4hMZj2AnNh+qPrHTNO2ke+rvByD+r3NnVdGfpy2THEJCpfsACwkPwN/shF
01IO7l+jFgFCurBqTRb1dfq9zJaIPEo8MsJJfFlHun4CWFqL9ePJ4wbXoXN8yNOG44rEwhCDE6TV
byN36ZwDLGTMedtUceYNbYNnRe6ikYrKsFOxN5nS/W1zlwnm4N8VGmQ9aXUuGbIU5hqTIfbSzDD9
TqVRwvd9cLVzS8mEhILeEm0kLgfL5n7cIta/b5+QA/drWzWEGLvoBCpyo+P48Wp2EMcyolBLkGZs
P2SCpZn8YwU/oRs3n0ggyjI+Y1d9TRjB8DyV2YuWI159rnoeyCORZFnoBB2AXZqpmYhxZB1iLPlR
H8g1D9CC0abmM5OHnC7OOfyGDrRIdIASeCBKN8597XFurrxE4udZ0sOxxAfxBaxwo/mnCKkmz/7k
m/MgxgEmIkQ15GHZwKegznBgikNaN/PWQPXmoDDtRvtbzRALPvxr8xCi/BmT56dvhNftbcyTt3r7
W8qeu7Oqxvy0wo5DGzrOs6bS+IHt+hXttyri4yRXWMVxdET8rjs1iM5JLREM76ofdT+aVJMpqCmp
wJJ8hOHPBWKgnhQ89McBBa2wYDgWBcpFN5aaUyfnkd1vD8p9810krvDjpAYjYBkUBE5kEqgeAzX1
y1VoF3Z4eDToZkLzh+0gRn8QuSJ2Yo5G7Z8aE8kUelPHWQt8JgosO63SYY6l+NyXyp2ANMINrEE/
Z/8Sg7LL8HbMcNib/3yRkVThp5VXVc2t594MDciCFUAIuJxtdkV49yj63/CObNgphXqlJ2hNQ7Yl
ksZojJEIWtZ+TKoFKvZxAwiPxFDujgLg8ijzMZo0Do5CxpcBQBEYqaGvV5tgHyY0NULeE+aG2fzO
YwzSfyN+Y9Wxg+gMKFpl0SJHHEbiOi0fFsXlUfLkQZARckzvqJS7SqZSp3uZ5HAg89KKdX9FnO7t
fGxTcWcLrYuiQpfDxWn5rISJIggu4wbo2pHmiExD69TpEkb2SDYU0gvbNWG6wmpgDsQ3LHJIqt4r
2jmfiOki6KTmbgOeJILtrNrOQWuo09Lr/1lBG7FHlO7RPrCY0PMA+2UqMV/wvUuQs2AtSH/gTIlF
yqwvL4WJWpJub95KSBjLOI+2ofTz1iorxy1kKY0DjfSUMU3z7TlD7SD5Fm6FYWNr4G+slekdu4GV
wYS+muL6M9sPG5Ff6rlloEYLOLi/f1mDsCiXMlZxZwQ2RsjBgRorVW7iF4RHwWmkfWkk/DpyNRrX
6K013WGbg4sOadY3B4AaOcPh0SP4BYVFsfrJXk3P+fN57m7VzdWlOBoscBzYols6ZnRF1qjtpyo/
g9Y5etIu6HCRIvCAzpCafya5DQfrn4YZlH+CeETpPkUBgr26fS7RXh5PDZ6cprqEA265HHw18Oz1
aDnBEBqIhb6bPzBQgP1fBby7mUum8iYW8i9pIZsGDIchDSAmCKzD2UQ5rEuKkBCPXdMQJi4j9Fba
If1i8Ygh4jXGGQrUraIbAHVOtlEExfnT+xRVfPn4rcd3vEiagq84wtAgzsV1u5qujy9yVXe6RNWq
XbfP+ml4CmuW8VDiEy1eHbKrtR7Njh86bkKKzRFasqazIn8TUTE773JdkJJfk4mJvTUV5F425vzI
Vqgb01xNlbO+GQv3k7iaqPtoQCwGKJPo8ROHuPHwiXUcXsqNrHv7CvHd0loN65tgRr8PvOgOzJ/0
fxEfnNc0tYDyFNFTY9W1nAma/nEqS4ADan6uEIOvVAVg3GqOZiqNfcLrLjcMtnyq/AIuS/FVMNyV
njW02nMxleb3quwxU856CSo7HLaKxTSmK9UqMTlZHi4Ilug4XunDMrul2u5swRoCWQGQE1wDyPYM
pWgKM3Np7AlIir9MwwoSjGdxLfS2nliG00SoBG/iCQ3OmuzhXreteNyByVKOMcnia7kO+IkLR6D4
fyjrK3XdGL8YUmQkQxfKB7icfwy88eisSkmW9V/6SZQAmoXTMIGDWORCv4ZEMm43t4RB+oWxvjtN
hvqTeIzZc1IwFoTnIuvYJG5U4tEjChG0Cue2N56N+lxOwLjs+CTSLsmMnDD40/wnWUcJALVCOE3k
mrP3DSMGTK7XThdhgcoufEKk8Y/eJTVBMiY1aZcqaG3V82s/z5EFb0k+7Kd02IvoSqBHfaME1v66
k9Qyt4IU85f30iuERm3HNFkzW9KJVDt6Mc34HyPmqKQvF0wDwlaYQZh1AVsYULLxC990BU50aqKf
KTTrqvmndUw+BXjFxs9WAiKu0wZHsb54llbsdy+28XoPZOTYGxLm5wOb2UOO0J2mdsrAB4oGCnX2
yD5S60l0wSmeCf4aYAbSWVMSInbVk98CSO8S0Zf65g27n0Ko7FuHf39EQVeq3WvkgfU3FG0ZxD2M
jmGSbhpED/C3yckoOMWvGyQFlIetC7xy6Hyr6BJwsbPjrVmu3sPSj3aBZ/e4H0zRoAM8NkkZ/5jM
1iPtr6449+cW1vcpMKKa9V9ieMAiDYMSioS2Pg+Fi4l3CsmrWuJgw8sVPCouur1TOi860OW+qYWf
JSBYm9WXqmUJhP74jvN70esSGpgqcKQyxGyIChjTmahNIi3THQmmMWB4y2uLhyLckZUzYlox5i56
G+X9OmpA8ex8m1D4dU8cG3nsl/TImwMXpNxQxdvYU8ppSclgEDxptB2sXOCsK2F1PzcG2JRmnw8X
cdQq9dX2PbyT/h0osNn9lXj0/CRjS3HCaW8XZNd3wekwlR98AHyBEmZzumBMdN/hq/0JqxEztPbG
WkJgQbyrOlCIuaud2KCcdeJmt+uD1fN4iYbrWRxEipLUC2Wfetp3ZWfkIJ6hktSMtZeGupyyWirn
Y2wI9duHoPCnCIMT1hoeISKbxifI+7UqWnzns1siIugCndwxlav9oSbRzvVBrFBJZmn6/qtokikO
F9vstbl6zuIsIBVSlnDW3dN21kBSNkuHf//lu91SSnS7XLUv2RLH+tzBbWlDA+/fDGuKCJ5LBBLP
hJqfwVh9BYmhInV/OkcgW9HFMVvew238Ri2VqT3PL7jBGvDGesZVwrbqXR/CWOQkG/tMDbjAbLnn
sA/EFcCl4foQpKKM4CnKmk1efuuAciE+6YmbCQFPs1GfYwmIL2JkTFL9J+IinRyjjNDu80xCyomY
hRkWbLq4CcSbQ5zrSaSvhsCLpc+mcDmSoro0qD1bb+HvBgPztN6DSa2G1w1X/1qSoOAViFoS0Mu0
N+dZlsU+Q09BFHLo+CQW72h0rVEU9IsPPf9dTrslwOYbMBN5bx00EJJhzxoBJeyelR4ou/2442lJ
035aEZIobnKN6O6N3KdytPqvcy4o7FLyjCHk37W9lj0GGsla9k7zae4ugLUfTEqsvjuy80lZILKV
0qpjFWnYt/qETjXspvZgYJFKvFhhCal8roF5YGbsBUo5vrCSp67Z5FuILKlip+7EZYyxnGjC59MP
0GVlmQVq2wx10G74bObq0UKP/xiHJnPNvDEGTpciBkci8g6D8dYf4vBqw+whozffw6Z0rPvqOJXZ
EOpvg3p3LsyO2TXuIgRTH85Oikzwh5wOornHNkuNK7u1t5SM2xrhTyKhDQUis+Q785Ugid4stDhH
Khos0M1zvQ8laSriFLOpKHpTr+pgjf7/wC96sGWfSkSgSnmGK0LzCnJzQnxoEf3oa7EQMSOdNmEO
ZmsfD3s//5RYlo6R2ozCvThkorTvJuDtqdWQCUWKxklTJ0rXnW+ARNQp9Mu+GZfGpg9BjRQrxQ5k
5HLSYK0v7QQr+m/zU1Q+QiSnvP+YdicrLDS/1LjPzge6LxBm2QiyES/4B9YoGjYgYoVrY40evCwv
InJR0z2PEEZMQHcNcsp2ZPH2YHurx34bYdoYZFz7q3vcsLmnm3eyIQFXAdpEX9Ox/qsD6jXiV9ea
lJ2zF97G7B0FFNdZNKaYJDiHPRD7/8tB5Iyp3VJUOk9hejDD7gKA3wQBT8h0FYnaojFkLxM989ST
TRrIPkhbIWNDsrW8mKeuce4INuGHIo1+IYb8bXqoa0+PNspWlbCIjhny09/pUpCKJYCp0SRs0YAl
UahV1m+YIjOYkl6NWORueOjoEdpIY2EgJBnsyRN6/+x/GP1TZAQcDg5dx4PXSisgTs8dHmhrgCgc
f9gWD8pEKrNgIkdxOgsvo2xAnU9c5HkI7I56HPPxMUnGG/3HDStvzfeLyER6aWhuJ4CUDK+M1tiV
f5iTd38jYVEvTrfOIUa/UCSJ5tAbsTPAHUeadLJCxZ27txoFnvdqw7BDl53E29+DYvtYBBNj6CpU
qVCTZ64C8L0tUoMg457I3aTaI/Yqg12dg6vIys2C95/jDi/7eGKscairba3uLV7SROf5AS2GMrSc
hnlxw3y7aWozMjqYCQzcmHkH5xgJ3qB1YPxnXx0IXY5IX9bmUAIAWD1sjO19F8Zz0SCak47APkUQ
xXAl1WIL92bwry0V3TwtSDXfPk+BjPyOufPESmuVEeo8rZwDWyPfdgGST66RL+9/lttGAtmvHWH0
P6bMqFsqPcq9vqnjvt78MLznzveW+Q+PToZXv8t0ppBUIS7Dnw8bfGW1ejd8rhXz3OP1KIfmJI6A
GU9nBUrFDn0XvmkQKInneezHRm2AF+1mGQ9B7dEVZAm52T10wqLllpL16v7N9pf2DICh7X+v8MOQ
7HROptqtWsQ9ZDnFQzsK+KNuoeWeGg9CVq1DsEQojE2AsBcuNr4TgAFlLKkqK6q5hWLWeuzzVIFP
4Nkgpqi9bQJdFi69v5gv2fUcukx4reUKLpgnawSpsoYrCg5JS5u8/lbruITyJf3Rle1C2wMf++gq
emE0rCs3wPI1K2MxDFO9q0PCCG4CCokQHyDo332NKv0JA6H6n+jVUlRc21Go9ZhvNtCFVhgD3vHw
pGq+CtaLOJYOlYKP241VbEIDPbFp84RZNkvyYGjZtSbJud38l7T2WGY+DW5trd/U1EtQlDjZVNnY
QnPvN0mLMrR6ThC1SSvtHAAStWesw3opihhcM0Sr5HalF32WcqiM7jn5I7bvqSkkxU8h+x9aabkT
K5pq/6Ao7Mam95RFz1qPukeiCmOE58DhMuKvVwL+ixhQkptR3lctaVjOiDNsqVUIvyPxv8Uugiia
SS2zeyAHDYwONe9M/eidpNrtq9FpAA5l+jixY33LTzwiO3+ul4eZD+V0n/36dZf/lbKVVxQygBqp
rpL2kY18UZSRXLUttkwVj2bzVnDuV7hGcJWOM2L+ybaS26erg4GMEqxUIEaZo/OpUUYMI6uoWC9k
LKlOzK2Nq1kmjnnSjYKrXRyGiwa1MYIlvz+aeacBO4hT9XXPuSjgzc/BjhFvf1ahR1tW2gxw6Kmj
a6N8cJTVB8D8YtCWhBz9oe1JZtHuiPQMhB7a6MgQGKmnc3s+tsnOBiF2hUUDmqAL4LRbHb4gnOQO
H8eFQSG6Jf+JrQyszYFH1gHtXf3CTTU4AIVhs6dkQxrHazjj6kH/xzlFm8aFlky7MxGFEH0v61in
F8mKtlVjYstfzJLuVE0f+4GBq9zaIIpuesRcp6cDEyXebwPvdrgAYXFhns0Be2UTegsfD9G0raPh
pHCBRYEA9fw8fSyxBGaQLkdldgYHuL9TgEO0OdWrwbLfFtau+mxEIWUE9Wy9mx0uOwq6vJdNukW8
rer2at4F7v9Trnyy0MbeqHqc0dFupp90KwkNP7ZxzG+adJRF+T+CuPg6/+5Fb8TB1VOfNQeLQoxc
A53osMNKf0TFbXxzkSwBqghVLqoV3ptaUNRE3lsJo2ON3N6bGPqM2uI07KSCTpjgFvx74SgIqMLN
j4LHvr/MFUulDCcs9uVaOHukWw4jhvC5vG8aJtBj2Gfk/1R+E1e0zYQGsckWsrpK6+PBhtJTQSrR
6VJqh8wqmQ6c5hNBjphQ5pb8BL+qzu/SPa08w4Rw3yQCc1hu33oKpK1gxbzVKDQBp+Ohv5bpzW0J
4wqimlqbimZ1FipRXCSb9sNmJktGgskn9NbTYpLRezP/rKEofpwnxAdbRSMA+mIyj3NiJ5f/O52J
XOHddWZ/FKanOA1x5QB/ZsK9e6L36AoIsPJPvPiSYSYNNXrybMODaaPH9pFr3w8OqMMhMr6M5167
EbwcLs5vgBaBEk4ZH3y/noDlaY9msCPEH9oGnP8b4NvkyIevcJ4IL4lD6mCgM8sFNRzh2Yt0ZJAc
PWWHwdwXz725skOMzLgQn/GQJ/udv3VIcNr21KzigUsebZj/6vpwdLTWG3vCbemIdtMtSEzPOKRp
t2k87zj+mtCwQ8o+IeSGUtNrM8Rjsu867Ps1jjbCvMQEELuSvmgReK4WM0Nto2DFGuFN6za83O/V
ptIZBuYyx44PO6HvoM8H+cpc3nU3gpcnfesyrjEDKz+KAaUA/RG7V2QhmafWlq9BpDTQeHy4cPMo
HgGiCmbNrgUgX/7kahKYZTp3WafCfVDvn8zbGWerVKosWoHWEw9gLOhFhyBrsCQx2ll0X6pL5O1X
7kO3Jcd27FjJ8Vf/wTnE/NrgiZdsLSxQQPpOexDyyuRDnTHqySv65efa+Wumzwz+XcTJ478QjaOb
1I63zavMUGPPG6EXy1MCr8Qvp3uub3labcboU9hsJQR11hhJTl5OrxY47t4RiP38ubBuwjHcU2Ht
ZfM7lue4wywfe48Cw2mac0h9FBwmDT9mc9hKZ1u0J9vA5/ekyFrVkUylLsS/9rVyfupGwkiO1ftw
oPOOc0fUwRpxq/ao4lyBYxP0HyhQnKuUovTKZf7O2OM+01FgfSvmfFJmNGjwufe3j1MU0uFFBm9m
CxjZA1V7Wfnnnthkjnzd+ak5CiUVigiJ+XPwgZ22sjtx16V9/grBsviDVIdJ9CqrBVvLVjiUqobC
ps5Ol8+8owC/RaywWBbRBPWizYt8+apyFsBnJ5wkVZUBAbt7plDy6ux7vWN9V/88Y6GZRyQeFuQB
qLmzT1txJlSMHgoeczrVk7vjbgwqH6n/D2LZzpH0YR0Z+bDJBMhKd5tn21+ygX5vseJQxCfohsVw
RrvKLykVyt1HavTOZ+rKNAIzdM2pSwB4/PapDhlQrq8ui8H0k86O34KOAmBa8uQPGvWIjrJoZFkM
/c3gYCqR8ZCCJYiKEfUs5sYCU7VYAvzv9Qx27ZYKtANVKxUgRI5KUyC3WOfKT4ClTgvCdehRH72f
2lSEk27QNNco4tsoVHIzMJZoXjKbHownvbC/1Kh4mbcOhm0YF/cz4rBZulbtLyBtQK5UuQwJoJyf
R+j14n7lK6YDpfVtWM1jKu1kO83/PZ2sOdEh7pej1SKHo2zJm98haE2cK0VqHnMMjYW52KRSRJRP
96HheItkQy/GS7JzSJEWNhl0MrKNJ7OJM52NCkzgrxX3MWKo0q8cV3L+gNMv041QHKg/5BaWBCYO
smsEGes7frDlf6lk93GIQy9aZ+ToX9zwm5N5973PSpa70/bFLsSbs0HNb32kjQ+po5Cbl6rTiUk4
o8gB7bMHxj18Z43sa9cHfTv3OsMr/4hQzzp1uVWtZO4+hEqifuD9Adr1wXphQ6373qKl/Jn6n+Xu
3idr2g1Nnd0PYNXeDSzOjl1vP8IQW8wz4rayMKy4c6s1a9gb1LUSGd9Xw6aeH/dZo8sZN8ITp45G
9DM7QwGxYLt+yH+ONeWIv3pvyHXN4NW4KNaqRsGA4RLCv3iErJ1kd7XmEObUunArl6788kLpm+42
eC4jWRveGFNIQoYBtuJwkjMc97isYz5PeqZiutS26vM5TtrMVlGfVWzOjJHGTz6qS2GLpn4roe9b
vYZCJZ+vbgP3EiQgv8BkjAUxUL1QAQxUEV6e5ZCe9Q6POW3PeigtizeH6DYxD4BhPjS5kqfTU11z
BiWzjheIVMgW4adKXE/Wq/caOj+phSm292MqoQ6bbdbm3ZXpwJ+NabKiIKYUPSK4ZHM7xL95mClq
iPSWm0gM7tKqD/XpsjcDgHSjkWZoRcrrD1esxoe8rAgWdUq5tFANzMJaotoGrK8fywLcSKxRgVux
II5Kgr9SNzDTzbRt6/73biigXQudGdf5q+sy1+0vNeyoj8UhRUJ3hIRwkvJlUdvg9ggowWjdPdts
PoIC7paU1o4nfUzRluYTAiBe7Ux8bn3QcnalhkqiV3qMw1lfOrdL6bSSQrRJAyElcFqYdIFTmvkH
Qrc5xq3Gamvch7N+hsP0UPCq9Pd+UYgqlWZX9zOx/1DXE3yEQazcfA0NFdhy7LxA+hTmAjiJOIML
PJ447Gz1o/lwVTbKuOiN7nVOWskeOk3DA7mrzoEsB/q8JdoeOEEmVKpHAcBro2AAbjN+Z+qSKkqN
aDsIZVvkKiEOdzSryOHj50IHfd4Oe86JViF4zcTZxiHiTGTGwgCfJLEi2KDbjE/ip//dv5fGXtzu
aDFsd/ABtIyEXNMsZfcQLAKYCK9ywU8LE+iyRg7TrDIYEaSE7p8BmnPsuXFefK9Gc6ZhHS2qqPu6
46Xa3QmdNeLtj2/3nFOB//eYTvsIcwZBe+6dYdfxDfKXQ2rRUnVILZ8v0ScqRDRqaYoiQCn0dewl
dRc7f8DhM5NJMuvqmx0HzFnwFYOrqEMfSzcutpF31T+pfSGlJdFCnOMLOF5lGFichoOhDOOYuDaU
tQ1hqBauiJwHT0SXKo3D92WuJh4cS3dyU2yTCrgYuvX9utY8g6b2SWfER+0gv6o6TlH+UETqElZH
+lXV521W0VVE5ebx2SEhz+2yRFqrPLtF1iWwmHtAZRC9+isWQYHs3RdvZwfTOGhSINkOB2fqngPP
LUArukIhWoTUidFIXqZtMbWCA1HL8F2Py8EDOrNAevphBAa057hqrndky+uDyv4TzPwdAKdsTUuq
cvCgGNOv9B8M3HZz9Rx2JzjUlam4Pw7w4lATbbpFF7nTOixmscurZQN1gT6JLzkvmapViKcgudbo
8a4WEMtqiY+YiEob5Ipq+vrsj26UCtuUropr2bGcBHLs+ZoFCta6TsZeR8nsD5QUJqhoPFXJ1oc7
QBTQZtth2wySC2s6XSzO2RUg7pXOhxGU7s8t/s/yKcZstu0ppe13QlE9vvK9EUoDobpKDoKdolAO
ZSRdxu4sYLgyG8ocWSljc/fNn9ufKtT+d63mASrIAMKlbPgTGPXvxV3o2O8WGB+KOyahIP6upWMo
yZ4051KP1Dniuk5eI2nH2w9+rpwqrZDEBpoluT0MEy7yqCvoPQjQGbPMywiMIy+A7rCaxMXo1T4O
WQ4718wlvIt+9aHmxFgWZ4aMZBk5DqDOzSqM8+bQpph/kWX88H+GrSDZpQjI61knFUnwsPdYOXdU
5VzU5EXvDOB1NnqUvtHec8746fm8FZlgxBnNjk5+M1YL2uJk8sk/sY5w1cBWx90rilEldzo+9aaK
TqNNufuBmM+3gKj9Xp2KniViA+nP9ic1D3USOEU46iP0a6inhiuMW8Z08PJr4rbAmRbzUjoD0Tu/
FoW42G1dQRobHqhVP/6oOSvL55nW11XzymGXBduKDJljT/19cdtgCJpMFSMMA2IB//SQDx7jSQVK
StdcyOzZYFBsKrJbdeQFKEuY7K6NoHsKus0eWhU1qfLsS37dC1EVjFMYAgM9KE3hTu4qxUl+7rCO
YUbHMcY/a9HtsJPwRKhNc3y5b5HFd6PPG2hirUeUXOtRjwIN6fEjvxYrSOst8D2esjDhEkQ7nFSp
6HuAc6MG+FU4ratYEuOn4JroUPIIDTneYDcOg4wU5vWhMp3cmFkwMP/usB2C3+KQIR724MXM2HLi
25mSX2+JShEA339D8cZlHQhh4MQeyJdO/1U/hTVqG6k0h8RHQjYYwg/MvB7psBUdXnHXvx/Qjrqa
/Mdja+JMZDzaaMn+en6PJX+bDt/Cr1b0f7rOm0ng9xamKKQj98Pn2aqEwv3QafyqDKMhm5eWNb/d
2MHkw0RBG07ClJ9dQ+EHYfrlvVLbAft84hfo7XsUMrN6T1mA0QTseBtCmi5bsvfphy+1qkrvEi8I
Eb7K+Ya0/wr/sB5FKWQyTXUGaX9NFV/82p2OLNR16BflBXCZRRm21gaQ4MJrB9vbXpFKZ6CeHLBU
PxtbWnNpoL5VSvYzlIOaAS+ZTNhw3/XMoUH/wBioecHa53b/Neh2hS7zoUvyScI95ZIN5Z4hzD88
IA8nBeqLvdpzxFttns4BTFz09U/KlxXQuItLVYP309sruld8fzCEWp+7qw5VjJwxgVf7F4UHU3Ws
xf3HMfITr2fBwZcepLPSA04suGdvbcQPIgaeu1GE2d5sWne5rWYuFs6XDnWXlCJYiQmZMOwG+jur
dfnL1A0t2n9/P+vwEPFHDrZKHQGsvb1hl05U3zqzVyOUecrbIFxYs680NTysW0wWg1QF/hLTI8WH
r8WiSTnfWMt+QHwADwBXZqo7UT911hwVac3TGJAvLxIEU5M1IMnTmb7xwzysH6qLE13nVqKngQYw
vwNgYGIk/rCQTAKqO7vUZb1K7rdtxv5YtKWCvsvo59yvykoGw7Cdt86gsAGGP2PqQCMQ2Yu6Geqz
jCDJvzPtPMExlxcycj6PAdzOBStHlcZJ/7bvAEVUNznBL4MP1k3p+kM4yrdo1zIz+05lGh0jXt75
crI9AeEwaMckEYTO3wVIoSS+s4uFNQtYCuzCV1fvG47Bqym9DxE1ey24YpemwrGpHyYMHP+TRWje
AAqgUSyZ2x8grEPAnoy8vP0tU0tojyQ7SHfyzgeuMZb5/hpRm6xsiMP7x6/IvpS0tVJ7KjBiwF/I
egKFJ5XHcPQLPumekyUN3daMbJu5GBMRajQ1xxqfEJ8v9ZFjGVxsdFFGn/UH2yUZgMHM0bW3SCMH
b40ZS0zFy1XfZ2ZpF5/+QSOXJQnKMT/nICmStKBWdd7Atw4zCmtGcAeZdGPOINd+R9Hdk6V51dk6
9GCfRcGNMcyONcbGPpqzZHpHMBuI8fmonawMP3h6yNu9wcVf6dZxGWHLS7m3jv26or+IvAc/Nju1
7rIKg70JOLMwDzznKy4KD5S6YZ6ebMiFEXeYW3zbxQmkkkfDpsHGTZcAA4zV+E65n6+uvTkArEeA
VfvYvhvBgnPxdkaY5P76soSdqoWWWmIaipvvuX7Ft6la1zu/tTKqeR5PwBOHSyV4PQRQQuazYzjb
3Rr/G8+IUHxDVUg+NlRnfAJk2hCNN1RElCJAxt7/Q9lcy/Qqq6GPZkfcKB04pYJdSPoq5uvVtPpM
RTDA+eZvcYjZTe8rQoa0F6XGJ7+u9TDJsnMvvQFyQDywzeWo+IME12ljb+BktVxC6cxBZvXjxNfm
W5MCm6xWj7hvGy8C1XBrf5/EOdE1mwDB+B2yWs5yRvCdv8qYWEhwEOc+OKVqjkL+WJ3Vx500v46k
mmFJNCPH1O+FNVSXzcPJu9/gKnM25AQ/I1ANUg1l9PZmzH+bo6eBSpJ5BDNv1jcqF3Vx1EhFzYFG
bqdjvUmzLRBQPWdm4BTUswmChGw3O/JjOKB5XxkiWxs2FJVOb2pjTUdj2EvoLiG/c5jkmV9Yfrec
S59v4SPwn5DYN+6FnmVEqXnUljP0LG6zuZDnwfFEJbnu7SLUm+zSCu48EkY34vcQbVBgwZPVbjg/
ZlP9tkStHRYc72BWKI60wdiz8YFUOp3/qAzPlM8QBIK5BsmUeTQ4K24UTH1sVVCgPS659yq8DTtT
kpw/9uU+yoht250Ltzj6ymIqKEQmui0k6f0wSOPR9ktoRL301pzo3HmU+w==
`pragma protect end_protected
