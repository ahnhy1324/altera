// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fwDJbbWYefGrcwNyFei26dQkXwRs51SeyHEZvpdsydy4rjIffrufPBmU/PdNEGnK
fKIuUx7NDwsh2w0AKQk5458g8iJEhAKAvGhcy6h3pJ+epIYBN1pJ/1mz0S/goquV
vWIPNXpkyDFxMhV2fF6/391wwEYPvQvEPaysw3ia5kI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 88992)
/DvVRYKGmrDofUi3+T68wPLIxgrU/+tQclUqseWykcjidlWml0HkArT3HoU0LXQ0
hKFH6zwKWQQSuTdZPIp9AiZRaKA+4zMss7sypNfeLnCaXZyTQfzgAZjPxt4z3xNx
aQOn4HDL6mK71JihWos7LKY25rYcoHz+kiF/utVBPIYXeQirYWDago3/vL9v5a5Z
Uncx58/5X7Ldp/fYcqeLkU5+EyXUXOmvCoS0vIRQlbh8rRvsVkJPa7PciLJlqfgy
60YJBeyl6hkfgwds1veJYO4zndqgvhbCr/Jc5zEqa5Pr7JB0GnG12SZUjR2I9Krm
I1Cun73rtdN3tf3cKWt5seGqFqRa690BIp0gLQFPgmlOiIdgGKMQWVQvttOalXA2
0be9vqTWmoZo6qF4nImCs1R5lvaiKkhr5gZ/2BQSa66SlqtvLZVzQtFG1oEm5sjR
rDUW0VHsUZtLiRyIMKoKsQY7EJwytUihHdeYKByShrBz24fVrdPedk2e1HOw9dMJ
HaL305XrDEcmtxHFheUCMa5HWEAPKFMK07b3cWlxcGpw4h0isKWd6pQYttyFXwg2
LlYKdfujXQ0UXdgs/OpBPd5b9yJzUsj4Xta10OuWVdfoHbxnvCAnF0yGfT+ny9uB
RAGUiDGU/brCbkGfUE60N4EaDYeyhOtIAwdjahneApCG8XfgVckuNsG8XOPMAOc6
o5nTQG8kPBo8xb+yZdPoZgd+n9o52M9QpotjJ/C8XtTaJcnAzUhh/d0rw3IW9nBn
vqHLRo5rfCyZecFpNewHud3vtsq5Umwcp9YMiWrUVoz3PoWr3UcGcUe23KtD9CEQ
bVCSGjm78219MZIJrUvNF1TojoBtzDeMoMAvb1TSXu2S8bgQUcJhYm/WsqTlWZNC
W80KIQdviXpeICGBFnCWEo1Sq9PdF5rkV08XMaszDmHwj0S3H+gEqey1wKFgvQRS
33GBHb3ikIHj8WcMHLa5ZaNWXI0qq+nqcXHXO0QPoXBKsXpEhLVdCVpH/DxQ+/Jh
rXYewRF/lZX8zMsO9A6y/0Tl+A9YOP5UONKvfSsJCILi/cEXnbqVpq93a8yJlwpr
6IiiWHto2HI6G+6Wo6icgp3Dj9GVVQHuv8ptsSihevqdXQj0SuZPb9mSWRdS9vNP
wx+MN6f8aZSIHtCV6WFgPbfZ3EU4w+MOcnSNByiTpWQwizWkFEdMbnuuIA7cfET3
ST6nh8vOZ7HRf/EbHnrXsnSODVihtN1gAkvj8ENto0Lyb6ZluGogoJq75mMbO8Kb
r6le9XGb4MixXmHq7ZzcfIy/7LTOyII3Q833ow/diAw728AE9lMe2rh9Q0AJ4MiX
Uqo2VLOteSdmhVcnY+4mspH8ak7Msm/SR1605IeuDS3QAPEv7N/ePcOexMMva21w
I/aD80sb4Xa6jKhtQV3fLz3FxCg5AOXYnNsSrAFP/Ov07jrt9g5lCl75oj6dj1xZ
PXwxTNVD4AmpdALFNR46x3M+iu1A/DMNfaAmoKRUbQlngIXhqK/tG/16f/4r+Eoh
ItwojT5GSQpFyX1TD6UEU7X2PG5YuKCdCrgaehrfWWRKVnUc7IhKs0cgElWuvTf/
TG4mGGIQHGDaAddg7hFq61KllvJTNL1+EWCeJe2i/3C6Y4gQJG1keO15m7i0h30u
t5Yk0/p61eX22FXRo+JLYsVrXco1ggghTo/QuDfu2fLHMojq3Ev5FitCS+F1/IPx
dT+ObcFIzadTwa/fmr2an/anZHQsRf/pKUuvOMSpJ3NB1lC8LOsPkuANCrTh8r/3
NsHcgwe2057Eq4gK4fzGORZYtFEjS4D9EjfAWB7Z/9rRrLYBPfRmGBFn6WsgyIcU
x1V7Hf5Kl8LTIIKdkCQduHM5/8f+DyAL66UpjizXneEXa9LMXM8E4kdZzbiWKM+m
ibZXbmgEtre6oSJCjmAfM+XL/BpMu4Jillr1ZumVBK7zr/PygjP9ZRS7kPsgt3hx
DLh4jk1nIFG7LF8RKK1f62qV4LxarSpNcjdWc3mqRSxWShwPbP0cECPFEleGv9oE
w4ExNKFv8iO9wPoyGQZNJc2KTmCIo/LzrzlcgsFAaDcBM53X52IWsf0ZwLCIkFFI
0Iu1dSO8tP714QUqzZMkD/rtz9H4SVbClu66+vRxucj1dSzwRIHL3Kf566jNykcj
xcAq5B22CbzbWLSHXh8kXmOMNanD/rbQb+imUwZRNFQ4IsjzTHILa7TMho9YJCU0
+M9YaGEnTRhz6FQFKrWfgmuH5ZbQ39qCdm0b2B9oG7TvmN5yLEuu05evHbw5KEaq
hoAjQgHGtUmgyLeqTAHCIknhWG+9SYyJKeXQ9GTbX8sb67fijFa3sbMWfI9cqZw3
z0WLOO/ajDkqqIyv02LIk3WIWuMJ2bQ+GpNCyzBNXt9/t9LZ3E/cBYl064xfZSX0
0pVmpWCBxyB1TRbI64eDdJOSNjaaxFhMU0F+3ATFmP6/XpzKYPzyOKicnUtFxZzM
mrsoECRRFATobbVTUy5iE8bIpykGIZuedw+4lu+XRWLRc6L81h35AngnwluYMhpF
RQi0T7aRmJXOT33mEOX0X8cJ2MXuXTjTmZVkLtONYeA9+OTFj8/tmmIjGVDDGEnj
37wtaRRXbYdhY6YGlmIgxvhWwyS41ZBFWx9FZWsq6C5EIlrYZUu0xn7ioSn+EC0R
/atd0vse+yyQUDcmP1mtViiqU3axn3PKHhNrz/c5iWo7VJcxn9RFa96ifNYTLpyo
F1Z5dqtHbrG0TyHbDL2OnGB5Xeau5NpTxTJkua7yZFLF0I43pIQ7vDbLwJdk3yTG
qV46PkLvRqVdlQo/Rtf/4PEQFCKgSc2r+hnyGgRlHxuZW70UaqiaCeUQd2HeB+id
6OhOFn4A3uL7HT2P4lasj+AOFJ5zoPVsEZyTQ0863UXcXkfujYz/SGIiLb5gb6uR
JMCz6+zAWn8esFJfz9hgEYC60+5C0vQtZoLMTLAcN5VsKabeMU7ot/qY0YTYHFd8
sqEMjOZcUjs18wmD1Qu16wV9HVePHw2wT4ZsV8TSQSils4sAAwn7aAto3Uh+p2GI
rmybwBoz76goH4LAgrZkD5lOYZpANOeqoCG0Z9bSkTqA08RUiW2rzSSe6AEULZDX
NO4PTonCIb3Db7fhuP85TUTB14gt73wEHJ+wynkMqjYhCKJXPL8NO4Kujy5eyksY
JVSdirdJOexQhQ2fIfFsRcfAV2oYa4iLBxlWpsGk07tQ9eXRtl8v/ARWkLgolMyo
lCZyaOqn+V/qasK8B/N1lajWCFzkpA5TXDtWrvH5M5va2GbcIricq46kJ75SYlzD
o+DxxXISJwn95fjjmRq9K5vijbSDBWECerJMqp+sdLwm7W2sRq5ol9dhnVaR2fuj
kmpbGrTZy0DAz6jo1hNTZkkLbfMBCo8iFcNxnBkKh+hwiG0vyY2wqjdmhhorVRv/
VlAj3xBY1KOSMPCLUFZY1DD/Ejj0BfIPX1C7EXrBR9g1aGoRgs5w2On/nmNPxZYd
RzRs8VwgG5iLo9GLU22zbDLuBLrCWbIIbnvFOK1Ab/uDCIGvQOue3/RJM8iguNd4
sLPmeBm8VyxN15VXnS5Jk585Q/AbJhD2WynAT/x8DX9Wn299mydLZtl1HNnXRRbC
rcUepkLIDtiAmgvz3M0XqnT47JiOCKuFOzwJL+xZ6XJdtFOaRwxncVXk58m64c5o
8E0Uz0flHJSax5g5UsN4HuDlSKjIlOzCwIYHBUb1w58/cahCGqrcpcbfKg9et/Ke
5ciFCN79JZv54P/27vNTA/2HFatQOoNSGmUWu11fJtnwDCfi+aE62kQ0DByFujZM
D2Pfhu6FDZQaDfZHT+Wa8b76QDIYuvgiJrwkLh0N9iH1P7f9dk3qlPKPVN4EMwiy
7dag9db/fMAWUe0EZ7o3//AHjwPDmiqDNHyvA36s3jGHrNnApt+jfUTBARn5McN5
wk7ulPNmax9NTLsJsUdpMYUPuLb9HbgxhU9CC0tSG0lKXlFdebzAubSSfyl/HOa+
Lfy7K8zzCYoxGsJrUAcJuVob4yCwFrVF3bxnMuHaNzIKadRHhXef2/sOqz3KEdYS
CVC5XbPWDaEyRbwm6/jWdZ0ssad0g2oXAcm5+7zRxYR6qPPkQvZvsffgnN39nbge
nhtxMd+WxBDnJFFyugexAfTVbNqS6Iq5jEPEWNVUsvtD4FoLF+DeRoO5QJIGF82h
uw629aA8WRuZjZ6IP2J+XuNZFbUeHuGFlP/v5eRt9JNbbFYcuO1veBK4sgWhtiVP
bD+LRy+zIcz36yZSnzcsr8kbN7vCwKAAjpH7Weos1J3InU7kS7nIBfXtIi3ClV5Y
2Tnz8jzRd8GqpGZ2c1OhdNoaMTsK2QAit9Twyq+ZpyvuPbmF+19ErAf8yyviTGpY
uq/pvOYEWV9p+29GhdWL9gzW9r884BdvaSbl+dHMWQ4A9UHbRApcyNM4Oarvr9vb
B0ZKEU2upva5ztxXGSuzb2DULmq5QftrXSXVNfxQL6aQdy2R38IO6nDXLqvAr+3H
2k75LLmXbdzblRosbDUn/PfUHVboR7oT7X2boT2lKDw04uRAy26wpeyVjCD9ZyTq
lw2Crt2dU4F70cjEz6rliU8E4EWs/ZDHmqWVN+5nz6cn8Cmbgn+eEhQTEvLS/u04
j8jX0cCWiQO0fBB5qx2pxA3haJ8pqvIbEKdU+NRUPssDrOCnZq3GTuU/Th4GOCK+
mSaG/S11vb2wxWp8xKhGXESFjDEDRCHr9vGv0Aj9VdlLDNjQ7No6P5Y6fEkGQQ4c
0oWDBm6S25P09v7b6WZgdBxVbskN7eTranfWwlTMcXiD5fFWPZ0AK7NEUTUVyaDY
p2NQyPqASkiDiFlqmhIVNQfTVN/NTt9z0+8PDSd0MK3Mdiu36QrVHfN9iuFxIGvj
D7A/cP9E7kc3XDzgthcBhJlOMT+CBmskShqx95nUObIqjuFrGwZBwdOmpXmE258E
j88TZ58l0T5rC5x48lYLYQXeVTQQc8SSHOaGYlzOrEbPI+NDYvushESUVurz+9fD
wJRyNl8MT/Db9gKQAp2qeIuAChMloEu96nRtfbutQZSnBtKHTMyoHPhYAhoR9r4F
nFZh2tuk2kFEpsSkN0KnLJQjwGJRx7nzZugLVQsQLpouGGJeiG0HtPO5Hb4T7H+v
vlUe1k94/v24ZZf78scMc5xNsGMsMtiNeUbJwOnfi6vxeM46u51JP5zHQYw2AHyn
sXuBOvBtLM5J0LKZQ0Uh1gWDrQGMCybMF20VpioeiDD32/cIvjBZNouk4/8nufqQ
9ornKkF7r5vUtmlhHIA+LiIqfsmkhaswb/Z4hV1/NSSFcYwmIb2rNijyy41SpNtv
J5NBSI5kwoH7seGNONHkLRPHRn5GvsqfoH/5vRYx8p49a+X4VwUBtiY0ZBZ1Uw/6
npl15dh2q2N3yTJH32mnyh4E3sp62YluIh5uHtVaHvNhrleT1WsVJ1K0RCCs8GQH
xv1/4Jll+c4LppGntxL5Ig9C/Ivu+8W5zgxbAsZGBq8+ACmqb54xF2ElRsXqLb3b
HjczZu3uOIHGDF/jOcuxhfbW8RYgyRNl09p/zZPqSb9EHbxfnQS2I9tUetriugLD
fsFhA9ZdkECY5QInfeVNPoYbGeH38TaudkBcAS66960NQHOFrsowCct5itLSbiXK
r/KvJralFw7x5rzpv6dd7r176hQFk42Ve/bweUplGVpZPIRCj97uqzQbQJni8Opj
H1g1fLHFx93tlgDdcIb6ed3+5heVQqWjsLNSyzabnHtvx9feM/aptIbvSNrumBkN
e5410eo1Q29VmcJ8GuJGd2qqU7THcUt5ua09WKUeAJFeyviu52DE8mdeVLDhNeQ0
F4rOQqWn5aTygzgkcppUzrZwjG+0GrGZlRvOOV6Ck4PuYe7zX7zMmL1XZE2U6BkT
9tolrW9RlER0dJ6W6KZ6uAtPNbBF0qYjpDFB/gIhmmI8UygvsAcTFVhBGTL2m51j
TNPmiq1jqiMEFYfk7yujS4xx6aQWWuUr4Fa7zKS7hliwMsCxkExWbfgKBe3ahDwQ
YckPiOvwAMoGDJ69u7vHaiSWF9DaG2DkT/C+QNBz4wezBbE4TUlUOsRingWZkJ8V
LS5AMMMNnyi0r7qQz5dmC/UiL9dQbk80v+c/i2r/PgecLVdHq/qHcvIOMFzShuon
pl8KK88Aoyh87GYYXonqAQzhc7DnIrMhXFd6vIrn0k1oWBKc2B9TKWVL+1Hh6Eeu
SLnea+z4Z8NjOxaAf3FPWnmoX8iZ1xNaoO/XchCnwH+/ct8DIlu+08RpgNkBRo+f
6IsrWl73uDLMVmSnHjOUC5H9yMsJ5xiVOtl3lXs2MAbN+qTbnBPyvuPmYmsFEtMZ
2g4FOp/e0NG35Rz5rBwm/Ag1dZGzm7X/F+Gd495c7j6h7XuT9s0dWSH79MtLYhBZ
CNe3lRkW5HspkbPZsl2I4WUlSsO6W1CqIGj2QrX/pKXSd29/7sp6zRrCrk0zwGzD
bwmwFasBDI0Owv3/wsRqniaeI9+33yNk0xV14SZEkWE9sOxHhg4LA1kITNyVfOLL
NGc7xxFRkQf2N+x7PCFA00D6cYUqKNmqTZelUwKvMeDFZh8NVdLaUytz7YMh5tRZ
G6LkB7hFmCUhSUsKhxpk4TkJwmuc6FT+w0G/vXOGav9Gk/1iVIYpOxRYon9T9fC9
ME6LRnSgrWxczwWvjwVCwN7DacsNn2G29Nn7QkFC1VRqEZfAzf3sy40FWHP61Y/R
1D4mGnl7f2bJjyMUjRzyjpEqy1ASA/HN39RzV4vywe1xk1NyBdiGFn97ygra+Xzl
Qk/lVwCn1lEp9bxW7zarV32030CMG7vmcTDXYS0xnFWLtY8qT+BueatLWQjSlFFp
kMon/lOTkmQdNzDw5aNULB/y6aqHDawYJ/A/4WvANsgc33LGg0quWDmZD26pv2FJ
67CjFG3N2f1KMU2vvDlgBY26NAn6lEN3f2AUuCnZXMpj2AH/MMSw1DHDZwzfjhfI
KQEJR7J2W9+WSzrKCH6Vfb9x8PLLn1rBXJ9Q2Ok4Z555ywIF1iX3s2wnSdZ3OjBH
Pf3Wl3cBRikaCQBZLwl+yEqCCuhVJb+byInLFkia4iCpIx2xS6JRXkM0GaXmjuwv
LVKQ9tTEDXiWisFu1JVtr7MTY47t+4/5Kt8YzN+30c2OPU9crPKkkluOS8R8K1gK
oB8Z+gZtetKoXO1zQVQw8zcNFifnsNGfZrl05frIyCOnpjSLQ8XibHreX/sYlJbc
9OZ8s9HJHqjyOOIlHVGBFn5AvM5cCt7bba0/ceI6lI1YRWiUJ/ktsGjNBfke2X1H
x4FTyW0xisZnW45ps6069gUzLnvO0QfQbCAQ2JBY1p9mMREOMAIlcdX363ETp3M1
xu/Gr29Iy/yyUhxh2njOMUEmfZtpdyLOP3gOxMMoYG9/j1g511Ixhmg9YFo6Tbgu
/zrZn2P7mqEBietvLIxYxV5rtftlPU82jG3YzbnaJYhhr2r3Ka/FqwbE5wyMmkIt
QC9sNCoTmBnUdSJ55toKzPxw8zhok4Z0EYG/PsjgIqyRd+jOwXRUL4L6KQu24HY0
2VwSIZoLDAt/7FXYiHNtdoNcACQaV53Jr+KGiJSPtO4LPf3VPRF48JPacpQ9kXxz
iMpf01iNjkRw5VlbQGBdjffUWKZcucPQm2AyCno2kaa/Gd+IUR2F2+/ydznBP/YH
UJVNNIQ7J89kCoqx34OOnFvwF3iG94aV0C820yGIcYMR5J+cWhZRux465qAvizrS
6hnXTVKGdLK44Kl6z0O02t76BFJ6p3DThRY1yjwdNS0/bz4fLEtFAx1wjVuTan38
2xXAyzva94FUTbF43jgoHRKYuAwfrd3YkktIu+H7TOsIx4WdSdhBviUqc0YUFcl/
OMqGI+kJjOgU+ouS2BnDFPp73qlIjV7F3zL9RbuFwi1walD3KUyd/D/+QXTBh9xE
3E9HLpL/YhsERVyAdcXbJ6Qo98xYAsE4GLfcpS/RtNoKcvDa7F920qcWriy+Wtg1
oqkKPonxmI09j/d8Yj4eThViNCFaAopnVH1mlvczLmr9D4yVZ4viy4jFXxu0Z1cb
sTPXy0FvmGxxAnjm8zsKPBjt7jxVL8uIpp00avzjVGp6qNlnYO7cqpjxNVoYAoqq
qwlwv1zEtw0LR/nzC4CZaihruU8Qb5Z66TB3GDcLxu7H+FJ9lGa0aIXq8sID8j8y
zpeZlnwbIKvzc5l4rCmvaVqSWj2jqIltQiYTP2x4ACdHVEGKHy+lcCB9cTRBHNqG
H4PPWYns9DAI1fxPFZdKtahUDHeNyl9oQ9cPPawhxIoLPGW25/SYPdSD3f6I8AER
1or3g/VZp2/XdcebePT356hlPV/IEfegliBGZDUN8YMy70OLJAqSNZVCzrZLDxhT
iSKtb7OleWu6KlQFpaOBuybI9VOaeTpeu/3yFjBe166jAN10X76uE6e5b1qXL3tL
gUbMTB2ADb7jX2qnFKev+CUqR6/4m+on1m6eFdy4EEuKw9Z/7p/py6n9bnYwxawr
+j2NL/4241SGE2utkMvADZTBHbeh1g+2uqFEr71ieqhHokahe8WcVL1nztSH11QM
mtkZoabITRjbRM+soaBON1F/hgY1XRnb+vEoO6XsGVKqPzGiJd2DRVwcT4VdXtJy
KSqOduFm1akfk9luCBNiVQD5WqqGbTofE/Zd1uniPhvhLOQdwyt32CITG19v/bjY
jSsOs7JMaWrDKa5WTZpOo889YkNicwpsJmMoX8kwu3Up9f5G0SS/HBhZRCU+sKXI
+WUD3wF1OyRfZdeUqsO/XrZoPFWq0uI0uxYMxzYciB3GxvPPkjD4eyjbxhcbP47e
0hsZOnJ08TEy9/SzOpQPtq3bFPY12QVGD0IanPpVA++kfunzV4+Wt8/IqjZCwAEz
LmiOo74uC3J2j82chHEyml4oWxxDVQmSBNJBE4DueweCWqlvMHNxe/RgU0m7ehsS
NdKJVsf3XzqJpGUyCv4ZHFMaJME/OBPkkNFs2Dzkmkn8ga6YaVhy7Lgp/cN5FyC0
CUb50cMW1+67TSS+5GjMNXgkUtgwJLVelpXYEeqNc0wiHaHlb4KRQMy0DYkJtMTw
55evWw6TKC8ui1RyZt9zu9NeLEw+C475Z8csuLB0zFIisTiswW54Pi/lghT5Wf1n
g92ue6BcejVMzarv0kEerP4AclyRgu/iVSxv5aLVj7yrYUKL7+XQYSGG9NwygouI
xYp3Z6wXyHK02l/N4qNl5XqllVLrvdXSEHSosrlY4bkwAR+0qHWcugF3hH7uGXG6
MEMatsQG5h9NeS0LA9R3A2Ie/vRBzYWWB46qzZ1F4NkLJ9ccnQpo6DYc91glUrUX
wOr4MSj12UP6yGjfF5ZiDeNVfXEDeamhObtpeNZsVB/EopB+r/VqvmrgHtr6XcxF
ddEXqlyO+fXrbQMuv32pUXY6HUAQvcXes2+XoOHhp+B4FutufD+PBw0VJt7ZQnaK
nMg6t5KlTNLOCAdoUqZ0s4pzJbJh0Kwr/qik/GNYePUSKmv5hD7gyRNf4zGDFjqq
ley8e4oLoY2KM66PSHoEOT5Q5z0XcBvAJLcG9lbkWRHF6e6MC8CNwvFYxPsk/AFR
BMsDCa2zIwrqbOkDw8/rt5vI/Wq7Z+BMYmdT2vcmFssWK21Ohw7Qbvj11A5/ofJK
SpuooF+CltUDYfqmctIs80W+YGhCJiI4OW253ji3NG2A0ujVfJt+CtUEwT96o108
r2YBl8qrASaZq/Si7VSeQehxEClqbP875ScmJ0K1VZ2wReNwLAWBeCWeSCi//3+s
stKQUfqFuueUH7rAjXiwgeK4XhOf7q5Jdpv0UTaLWP+Bw4kkEbgsNz77A4k/1irt
kqCtbaqqf/CCf6Tpbwksg2uLgSlF1l3L2Lt6fAH0Z1mAgMa/gfWkkoW5CUT4QK6G
2XSjTSrs+v+xcgzn2QQnVqKyqjOj2dGJ+H68lZr7/50b9GEIWI73cTNENGPSYpSQ
eNaJwN3iVcLh9bP4ZilZ950y/aPCQrikC64Byhx8TAkZWg8Qe0TrCu+4h8cUqTZo
k1s24VGMYeyEV0bRR+mSqBJsvXBkz1x1VBNBV6nJQX15hgTvqq/qJSCY3mb9wg/R
5BUwiSeWO4sKDAlv/M62VQPli0IEmmFymRErdQVYt/wcUCwPLVut5TvnrXoeyJAP
A2JRBLN7yEvAXGUAIoPy9pPUPDkz4roHQDmlJcte+VzNeNr1i5dW8wAzNqfnEPIZ
zagVFvsrPxl4zaK45AhRBDCFkhUWGRDFsU4zHvdKPXD0e1YOhTe9wBDvO34wL93X
dOq67W5yvE23QiCxqjhlB/JjMWiGjGWVgqIw85VOliDTuJalkDkLvt3gGlEmt1iD
tafR+2YW2X8PqTHPnnu6hm9kOW6LDqtbnd/Hh8NB3o8YeNa7KtrrswvTUSMzV7XC
dL6ScvaFGNQNAL+1xDLnrlm/y8gQP7uMTJ15ptd33Nna7US0MGOw02WLcQpfNwH2
hxPRReega+3jzHsqSd9zefYcG/p4OTLav0AYBozz2sAlZ8whFFN0PsfACF7ms6ub
b5utjpIO/UA4aoIW+JrhMg0fh6sQGLmiOQobmGLfJtQXidqtXzgE/rqso6H2JEJQ
bo3GlZjDx4TcQotOmQ9PF1yWlFSKoHJQmVYmC2VO4IHu60keqKlwxOFYxxznb+yL
n7pC3IYJ7Q87LbKNlHBDy8XWnu0ViOcmVL4kBqdMtUdcH9stzBytw23u//nZSWf+
2PkFmczzPWh5jJBR6C2j6bSZmnzQczoXDJu4dlOkKeu756y0RR9A8Uk5AV71l6wk
VnEVKcpguSIOvPfYOnd8/KwirKxpsmThnvl3P8J9E1F4vCn7BFuYiURp8QlhOnR8
6Fktmzx2ZhH/FvXP5SLas1yF0/bm48O5h8AAyA418zZV99gAPaSbe7UlIIORcW3H
xBqbbA64IryxyJO4M7e/+cxDTR1pABwPN8j7m0qUVEuiYmvpiyV4Yie+T3GIJLiH
WVpGlIDMvCjpLk9p29eJZkuJbguJUf4HnEGYyYPtX0AxZpvSnUxTwTTup12JqnA5
9hneB2GOFQ1MD8dP8vRKPcIiKjLnDCyqsMCOWj7g8t5B/rJBnh6JHPyRxXj24egK
KozkJLrlbZfd1fDMOBbYlQlEZBnvNIQMXpIVvvo844gYz5yANYERnkQ6eg78juVr
hyS21U3k6iBW5K+AJaCoXWw9dKZKRu6W2GKrcIBPIUZzsTfurxPZlzCb77OOr46E
igCMEGgc8eJIdNmwo/NguClqPD0GV+1vrARq424yDE1okZRV1l+vx5PXZxClYnEd
ZZzr89uh8qAV+zM4BpDxMLKwprhsOCPwSbAe2G9wFHFOw8D0I0nQWZAqTD6PK9CG
VvVVoxFuFklZLbIa6Ee0zNPCC+yyzXx4y/4zZ4a0d7pxtVljpsVs/H5O3ziHlXNr
BCd/oenrBPVqlDt8l4v8XQ73it1uQM9CW0QnDK+m+viUoonVz1Px4JcB+vVEVWo+
wFUIKq334VOicKK4KZKSo1FbHYCsRW2Hi4JK6ui5HnN93gUJD0aNsg6EDZbQ78Ut
LasDXjnE7s0uiI5Ai8Bpgvkv08VrZEadJZ2bTFVNI/AiyhferTs4cMnXWdvgob52
FS//vhidv+ehOtUz+R/84i8zqWA+PpGQvggFlSCaV0TK7VeXXycW1tivk8dRRomc
fzL4hI8+izB22P2oQnq3KQua536mKJ2AJtW4TXY4H/trIRBl2zhnCNnN1S7GFdgi
TcBz6RSNhD7Y+vsLf3gYUC3cXU2oD7zCeC5KMv7u3Hb9sTgaolnCKVeoZDvQZKNS
z12e9p9tMczMTC3RFR11tDUCmNxfq9zIRoRVie6LnfNaSisgVQMfvNhEXpDa791b
w4a/4RIQr+SAJv60NG3SXpIH8w9pW3A90ej/WorOvrFeIr13eb9wVp7xu1NtB8DM
CE0W50wQtXi/78+LJ1wFW44RZc88a8ScQpdae5K5/bvypBKGC3XiWMFLH4he4k1d
t4/4lAdAUxrzDP5oeRksIrnlWACb7pfhDXMNba5zmKK9ZfjRdaFtH+QdJXpdUrMC
ZZMZNYV7fjqajkKLf6W4GynMiLSCV04arQ+yYXfgu3p8wJ5pIN5blqBU1UWuCWN7
K/M5dSXGbLyS21+DOpeEsOR6UQmHdqBu8AMgRVw+/pD5NndHEKEmKXDw0cdHAJiQ
z54cCHiYyo7dS4qm4UvqsIOfHI4dZX+C95eB+zpUiJZ2MyyAnyryvZ+NCyYxKVMI
Rb1wGZi654puIfZF11z1M+w6MCTOjeZAu/QwsoGcXXEcSlR2a6LMOHh0jrSYFhyp
as/+yOrENGdrQ66oDtgtS+JHIHifLKWY0w4Md82/DrRLV4BJl9mq3gHNebcbzEqE
xUpNHywIG49UbykzpVjuFOYALiy0H769qZSb3jtQ4PGtwHxZU1ZJ+2ckgNlUhRL9
rPg5MCRG8trW4Yw3wx/fGYpxOgmSz2Hzpz56IVbXRmFDxxlNyo5JUcSQCHK5mIA2
b6YOYiqQjrvmfAyCp/KOLgeyWV8BdLi6VQ5FoBBEPM0PJR5xa4SWEwk3sXmGcyna
4Sv7uVGerN/7sTeVShzspTl3q0MTlmBgXfime6NDhH73YXIuYPS5heuJLz/RrLbw
x5FdPZBM0zfcqdOj9cDogZAmV1Q7TKL4XAwRBsvLuXWsGJLqErXTb4L1fPt9WR3v
CSxMy28k9eCK1rOfTPIubp7HTXfamWGu4OteHzFCswgZqA14XGoZccIE0qbJZ6F/
TAuEB5zwyGQRaviHJcw1SiXuBpATpB90qon69Gnw2MiyEcqbs/iVtoegyvKAwjOd
wpKJ/fhj70JkWzFWYBTnq+ziNAYuNDo/2ugnpPgLnSopSPcOlpeXmFN2Dq/qX7+g
JMtGZb+ef7qUEEhtgal4bksiD7eMKoKLmCCHf1ldgjPGNRhKPWZtqjqCs9XP+ZnA
Nk3HC/o1PPqaiMnL/3Hqg6VSDe8zCC8iUSq7MtaN0rjVuovXCgTpobqp1VvJLzab
oO9scMtWmoYycKuXodrEcq98E8spbfP3Z+x7uEnawybFgP9lMhy8IjVVjJaol7GX
BZOi68V3X0OoVHq09E1Kf/OAPOftnmUD3nqxTmnZGK24HS3oK9YBtPu/rEvL0638
/kbmNMVJV2C2XPOx8ixtqq1YF2oqF9ICYrv7OFjtkCAF1RZM62zAvuigRMUUEXNz
xuls+qfFJz8tl/hxbKVv7DiwQ2vqv690xqDZRnogUMiUtW9+xwOknHsgos0kyXCp
ZOkfff328eJjFNerJnQKQpFYJU5sghi+XIQppVVgAv1Eom6Pb6c3gx360DWQ66Ax
7q38YdBciyRg77JzqELbfmZdlY3FTKsMKAMY5IQX24Pi5tyLPfQYKUagWt5hNBAp
qoyhqHKciwDs5oImWUmVgkO0L4XUb0mdN+MtRTFFaD0NUJFhqdffuQdreFbILNT8
uVNlSsHvul1Y+irKYYZD7Z84/IHJbRnU3Xjd/Pwx7yIUKThHF2J6mrbxjMl6r8d7
iww8Mr26WKBdhB/Q2qI1nY5IkIFzFE6QdTSTM1JbeN4D+++FLh9M5aO7wfC/OFZY
Vn7YfXwyu7OQWde0+draCuXRly/HBF1bLbarAQIy51B5i4v1ieuCcEQgFSHm9MCu
DjAnz8yQnF7dPUsCE6xtpjdLrhgzFVSGBHGoSi+cygBzfaYeIIB0Wt/d7dbi6TsT
UaDGWG+5/S0hp/qx1gJh0jyGfe1mwxh+dSdiD1sjG8n/LpiIMWCE9mOK4v+fMGfe
yb1lmjkVa8JnIMf1CSABQC6N0JzR0T9816hnhNp6jhPKbXhNmb2waT44ZmqBi5QN
ggl4tKzXTSzjAnGvPJiSPsf+CCK90FiwiqNdQ7hM+qTbLl218MYvEV/iFdipb30e
QJabxw45NbcVyK9HoIrrn/CmC36vWOfmzwFtXtAbol9hmkrXad9fmfH8c9RgPf2Q
fD6yLS/nBo9qrtmFCASwZkuQTT7XsXzt5cxExnLZJjcGaKQB9wMz4V0r7k1AmnMA
9nwXUkVQ0/WUcF1WljaaoIbUt0P46eGNQkRXfJpvCK4aNHwLO/GxSCIx2uT9T3w1
tISRY+wDoDE4j8f0chJ/zDSs5HXZtrlKaFRBnOyjoj2lurpfCMc/Jisza6a7cXAX
3cxcfFmDYghA4QEiCFgj3yG9XEtM1gwevb4SPNJp87QBsPngJz65dmU+9tg/wQfy
mOiLkDnYbLoUsZM8TO3bfb8/l6yX3XdUJ8+WOaoa7APN55i2RYbV2+9PqRCUf8A0
l43hmOILyMUSZFTwKF8osZBOsKMHOILu5xIoPOifAUFSgDsapGpFFXlEwJ6WvIRC
BQhKv88abHJAfSpS+IxhQMcj2rQJVukT9fGm8N8RLfCMNEgG2Aagwy0/k29bCMUD
6YkmYZHA/yHvyAcfvByMzoLWZOIFvvOzWmP9fxvAoWoyW1/RVP7wJdVaDoR8PX9z
WS6wEJSO+YQMnHoNxPHrnwpCdNy8heit7vmJf2eZoM2OE8NSlnI2TtT8NS0AiRZf
tKcHX/JGgq79WcUGCX5j8j/H6AXmCu87WqHFAxZawh4byYPFr/hiTlAgFGxWgLuI
RCF7GF2tCJtJExr5czHustyaWnmy5ZZ0lc+53kVSAN6N75PLCWr3TvATtawQo3Gp
KCpRjOBmeAEpyRS9epC+AzeKxIkLr6uMFuMMtiHwO2VYBdR7kKB/IXoof+Dv75zp
1gw32UGj9LdhWTdeZKmnlEeI98gjsDG+yGDeH8VA0pAa0dtWGLILaELm6cDWOago
VubcyHOE6lfCrrhb6cBq2J2H5o1U6EukwaKCFD4fRqmkciwYBmV9/ISBhXRgxXh/
OZ0EsPXz71vrQNG3cUbLBGbzVvzme6A7Ow3k3EUbswG5CwzwcxsefEyATeBuMEXZ
3IkCVzXljXDWJjFLfIFetoxRUFL9YLg1hm1WIiMl+nyasnjssr8/HsFKXb4kCoGb
ldOpXgz2l4VoQHd/ygBy27+VobSGLUREJc3UbyyiJKHbr6LuH5VdATOzRfUtckUA
TKbZl4j/3lgnOmW5CiUvgSa4neCbgTqoFaTImnmgL+jgqwJtPontv7G5scuG63nQ
TcC+zL0zgG1wL2gKl6llOX7APtoJFeOhv7quC7nNcuhZSYRie3UpOi4dvgsgzCde
VXcNKqu4KXJvQRvic8Ua1xkrnvYMD02U1Qk0DWQT2ZVM23ggpCdHMUr1p1rAbZrx
V3ned1cyVgDSqZ2DUvOxwCuKkKuIjbk+nVqYpxwDu6mlMd20tc7lpR/N4bFNLX7C
zifhUSca26ZrRWSlJX/BFi73hJbabc0hrTdSSLdNqIQYGSNYtllTTIjIyU7CmzJg
6I7PwMaGSzVaCsPNleKAOjcb9Up4VnlN8DbOfrc84YhX38a/OquydwMU9EFdyPLQ
N4Sq+xSj0PBeqZAOpCIjWU3lsarJ62aPQ1lvUOlgPZfvNMVYEpUawHsfSn7+Cf9A
pvK5xc52nwzo+gSiezCgjxjBtLoPHR+6OwVZtzi/BoymcsojELLvua4tr/OpVcoP
2OolDmtuiB80cpsWa9J4my5oSdUslJ/WfbUsI7yBnhgWRgfsI5aaj18dsGP0cDDo
yot6Nd4g7H14B+Z34oBHkef9Hmy9xfshXL/KBfYQF8uBn7WtwL14Vi8vOpVNtap+
7pJ4e7TDIEKtEgwj8WGrNuUNeQL/jfNeKICm03g0zcXKgaydTUTSI5n256Nc+ve8
WPJ0JBRKvAcFwC9JQLNALnnWZL4XSQYQoeNPvGyyWjFH9Z7V5pZMRw+0XSWpEW4a
rqwtah8B1Q0gosD65nlvI6e9OPB7rkCCRrOKwjkUKn4b2DPVhBA6i7hVWz1hbqoR
doK2T5R0ieQrLkRYt9ju4s8yNlCp1qIzbHdasIiqgH/wUWVKUZiUJeyp559IdDYq
1mOArg+Q5yz+8CmBBS47oeGNsiWkP9q+4BEmnQybnGjI/ilmwZYXdmv+799rFshS
6+MoH6Gcz2n6asHM0w14PBxHUdMEGKOFkWPcSEJmbo6RkpwEerfn0cKik3wQVkrm
mMoPWuxXeKseXBbwXpQLSZ05IpGnCf4QNUImUPS5alDq7toe/NUxRgSxSAhuklIb
/8HTx10f12h16pBDpvaWONNil5+f91GZt7BV5QcURPe4xGygeh/x8WtynjD/YgWM
j5iYA+T6WkD8IOg+smIxUuI2cO79mXF3olBrn8w0yMKVTg5YUZXCPVuQDmyTnt2f
3yX7l+AngTzhnObjejrLnKygqAa13WiZ435eFTPQvDLu6VZMwisVS7l0YqZnuCsN
GopOlWEn0VHzshkFXUFlxjoTVmvi2NglNaXwIZld4K3jAEZf2/iz55hV9WMfobJ1
Wr/+8XPlf00i1eSbniS+SvX07ZWC3wW4yi4hlvWNTcRuD7Af1Kir4pryGr3HPriT
NvB5Bg5MvN0OCd6ITv07TXfBchjSysEZyhD5fy+CvWnbgK99oeF6GGcrkabJkdfs
Ty6PtXtrNbKL2T6CShwDJuD1cQiORwvC59V1cQmf0KTYgStACWXcvZAExiqxWUeg
5B4PfuM8DN9BeAGJHEFiK4tpjm+pmPqxCA2XDCJGuuk7PHzh9bIarqNE9lPm/+N7
l/Hxa4hLg19Tp6U1NHE8QX4ezZsQ+3Uq7RcqQNQjXbsx5vvMJDMLwHF7pNkQmRPd
MtnYuJCcW99dK9UHwMfHkM9pKU/eLDolm0v6bMWLT84XHKZpbmUHpdzkSX+gUz0L
n1DEzaOxSEosWGI6urrhhfjZl2SjHOcBno+ZhFz6CzrDB5iIrTyyXkiYrcAlE8pD
YjeX0gnlbTTH7a90v5awCKJ463Pmd/Ppwk9WeAkI6IMDCTGcpmAb258U39hSP2zC
2ojbzT+h4qURiyotjjZO0ahGQWdd/yW1VcU2K1x9+S/rEDmjXRoF1j8jUc8iBe7C
rshfb5oV01iXX1z890gHNr3PZKl6iAi7E+uKhqmwl+JqOdyrseTzJsjyDxjGAAoV
jFwfma8V9vGHVoP/SdRgN8E1oDrbpiOD0BvzU3zpKyIufWDFPEZtdKZeRDR/Ve+6
o8/6p8FNhzLX27ZFI8veLfVNyxB7YqavBAh8SKNkfMtYAWzH66e7/W42JWLzqjOq
0q+10mUJWMBGN2gjS+/XeacoBPTGt/Ldl3ADbwxr++TmZqyP/6d/Am8y4Jj8YDJk
FuqxAcOGCKeJ4DwdptNAxgLriwHlo+9zew1vjPktVX3Ffp9m8dOWnEE7Xb8RiEKq
Iv5WYBZRLLG8uFXZjYE68KoeTOzfY1TsA14GvKyG1ZfYG0FUKb8GI4aajSatjjeA
Vpu49FxOtvW8rY2LSzdvLKjnfjc7uLN2edGKpc8em6cOQ2DebiyGOUsn2zqfec2F
wGclPllUZueauvJqYdJTdnHvO8EmUS2xqfcHW+qREAKB+dWPlcMblzsjU9UuJJ7P
M7RixBsiWUfYCOhkif/rSvLzAghL3ZH0ZclPlLr2HfH+PP82kdrXAdD1EwAGHjyN
5fB52c+t1J/2590sI4zoh2Y3ag13RSLHEiq1lXXKHgaoX7IgH9JsUxInZlZ5LnIE
VpxViCM9TQ+8bv08zCZr/ZWS6Ip3FSbK202RhnFvqMRCJv+EGf4Zkevn5KCwuhbs
xmq+qOGuqARzdWQAhc9qHIdUXgjPNwg6P/qxVEfF+fmEAoKa/0uvOLEDKvcnMq3Y
ZECeO9SS3HQun2jr458TsBnLvc79i3GvNsi5UkF31GMxdfGcwTlplsbgZWCBUHK+
TeuNEO1S3u4wb+kjnkx0/A3DfbhZPN3KFuklV44rnbULbkHMZCLyaOV0iym1m/kU
9bNbHgVsXAPSRtrVCNAYmRGzMpsNB2zOkzi+FPYxCP/TTJ7vEq16g14UUzhnG+21
TV0dqXSQeF2PJ4OjR7VukqNs0z4376QjGwSUkUSS3IbSGs11xDd+AOcrkBcB9Mjx
hUX0xQ9CeWGHu4sg+mlFWrwQhvIPuJFSm2wPlpZEdbpJjITrXelTjr2UAr8ki1JR
5i/SyfIIcEoJz31mo9BcYNcr0yazphz7bKz9GFHatlCje1i3lct0nAR0GQ8qX5v3
KxtuhcT3hcMEJylIWUk2G/PXFD2T8aAFm0pYzoq6Sn9irPv4UWdE4uaPXRDEjSMW
jpx19r2ecWLY5Afqxtl2CZ2unRR9boyJQua5130jFeYfDpcHNtbkgQPRi+m5RbpK
bT7oF84sAc03OoIRUkA4vfvX31fYV5d1AK54E+EPPp99WIGAjcV8fZ5grqIY5Mpl
buxhVLOBOz5Q1dBBXI2P1HdviZVVqGy7sR3cjdL+a7Oo+4ujDx5ltD0ygRq29Eda
phTk2+onTY2gwWbFtXxvKaTq/NyJU0a554vn0f8c+08yAkhWcDF6NDokvSaiYwbI
CZSWt+Q/km4iGf5DGukHc9nnBuLuywDmqcJWcD50IVulEDkhes1sZhCncm1HB3ZV
nTvbbWqgLuWdEEH0lrA+D2OCCPKwm5qHpVN/NudOfO6HTHPF/0K6o2d3d5XQ4n7b
1m0EBXebI2mK1QEA3JyM4GVq+kNEI5dyoP2z/KtbSJ+RZqc05EnBVJQnLsbkdnZN
HqDmA1Ip7M9F6wmWgnCJHTctwrWx11eVYS6hPFlIaxwuEH849e56HRPKu+Pd0mC/
6BMeb7T2yymXe7zSbI4/ypLmG0mNZnsZaTUb4ss4f+WkSETc81TWLWo4QRIlJQ3T
if2SmZPxCE59phyOoLIqZPUQa6sx8T3pKBNLLQTl42XapW5nngbDH44iNW3e4gvz
87dn/zsJJKOiRmVcVD3RJ2KYC0RFLqYH8V2bcBuJkaHWSuqLbPK4mwbcqEOzLxIy
aHfNOpEodIaagO0xJfRwY6pWPI2eKM36A7xXGyPcMfSx/kI3BKPrn0Az8o0qy3Xa
zx6ijWwti1LusV0xBHsVtT/WhALKZ9rMdynLgMnLWhhsz21o8NhRhBFhVrbgAgBP
/opQWmTT4SGweVL94z7Qzlq1NenEgP/rvt2dadWYx4X2qANS4KUBnD8zxH6+TD67
48+5mELM+skAE/fU+U/VP4XSHQBTRQAg1Vm7z1MMR8AQ2dekerFWom9t/Y4Qb9r7
K8mcgncwLQAiX2VsKrLzLP3FwKSPiie5igW8JwhK2/XT2GQmAxcFgf1Jk8WKmZGY
aAjgnM8zGQ8VoizyAcIyQY8AtsJ6ODj4khOZRX/gPzGHYMAhU4c28cwq5Qyt7S3v
6TLrRfTg5LmCJ3uUO5X3n7UR7uYZaQLewChhbmyFquL3PRRwLdSwFS+zvxBV+UPg
PdvLUfsCY03rSaEbkyPDhwb7ZM8peQAVu7/WvJBvXORERLOTjTxearAolA/LI0AV
e2fv8wn0EHdPRFIOvQoSY5aGiedscJDVyqy1X/pTTt2Jlqf6LqgbanUl5T+z1bVA
c9QcM0ehlYXL6fw5bsEhCdLg7FV5n7s12KX7k/9/WLNCNHhptK3O0Sq/h70pluXz
ZjstWRQ+d82OLYA/kCxvb6/NjpMkx+K0Kaavpnyq54cKTatCIgt7tjlzktZBHCKe
CR/3/L0Px7OWYHd2qWGLQfSaCMyL9zT4fbsxk64ESbHPewyFyhJjWv0J4MLLoRD1
7aXw9Kg7Jujf/lEtpDo/Tmx8EAHDu4SnUv/dIbw09mSkuENUvExbTWQv7jiNPTyd
53pxgCFkTkEp56pMQq/Rob0N6YVvzxsgZTOUCvhYs9whIjdgFoMA5ZIMXWX4Bewm
L7lPd7XUOOkit/OQnCr84WMDdwcKf0Lo6OWyqyBAxRNZuPGnt0rGS+JJ5rzgq5Ov
pApY614itVwiBIo/aP20X5twcbw4JvHEDOKLhkt0ZyfwpcNYDlhtSkTOqd8p+TKa
P45n4awYukBOMfTL660iy0nX4xu/w0zYrVyTzC3zVWv5N9JKYTBe0Fyiq26AmQOj
phHaWqypMyVbTk/vIaTEXZPv0/RkFqkrBJ1VebKpDt1OrboD31mKQ4uud48t2fFr
8hlMIclHWWTQw7E7rd+HNLma5EqKQ+HmoMGt3VgU+YC/irEPu9dfNwop7s+F6240
Du4em3HmK47j3X3VWslvxfpt0vBZ5kAQRR/qUaQs8co2cnULEobpmgaonDZMGLiJ
EV/+WLpXsFX5Z149vSTK55+F0U9Vl4Lt0dxjQazVPGcjK0ujdKwjW9As01niVIz7
5eO/v+sc2VfxmIT864GY1MwQrXPdVLUuaWhIEKKMyZRcdH7/i4yhE5z1OMeBlUXE
f1nSO1h9p6Dw2bARmy7caZG+dT4BdSTg4v97TzyDltZrHteonIj1AbhYWBNKsBXq
vDntdnVYNyjmAdUBao/+5tCK+LFit9rCeN3h3jgvCQ0HUMol9/67HxWRlx5FB98/
EtrAo6yCCnGRlMWFGtXm2VinAme+xZWDyqfRNH762mpfuGk/MnksavrS5UfUCMCg
Alp4arV4e6Q19HUVNuOYDEbgyo2D14sgBSSALcd6TYgZuHxdd+gNKT5ZhZzBFyJ2
EJNQaJ/bSDrti9ZC0xj3JBRNjbhJyPd/XdtiKevZg/v5CvAtEz8gKC7rMV2BTKdt
MZZVA3SUnagsodK7hmc5Dni4K1j2iTlnnfqXteiX1sL1K/JR9kAHdfk2yrAWiluL
EOwttIFJ9xDF5LwUFR6GFD/PYTReTEAw6r2/dw4lx1qBD+I0R+bgpzO36/kDzm8A
lzA5sOvaYJZnt2TuwouCFIBDK61EiKLaUVJAKJ8LzT13cm9VVGUEMTBwCRizow/l
d6eid/XPhdHfMLSqC7gqI6JPMVpFbaUv5JwGkfP6chxUiGF4Ge5wNzi6UfD9nBim
4RjC+UxMgy30eO77/uzRe48j8EtmUJzGknxk0BsbKMvydBXr/LMrZsjuyimq79/n
3ekDnLUPygsWWJvIzPYmO27qZBxwe4FDi/kZsRPJWXGSYQlXFHD5kYWhjeYHJZHO
HaX6e56lW657BqhcLzy0yvl8Z8x/4+w91AKS12eJBCH0HWwW2TjI1gJupUTx18OA
6pa78njzldQ2xQLwlcuhNPhFC5OFFxSSyuU1nM+MCkMfw65LeaIL7KKVgAUs4CbG
tYkAcWgiUvFUJxkj63tNyAafKcngmy/qSDFTk1QOzPiIdCib0qnBpWW72S0nGEHz
egZEDK/gLV+5Liwfq9/Hw3num91/28d5Ss6JF3QIW/H20LulyOCRnKKO255FcKDE
4YrHdydxtw5igNGEo8bd7VDxkSfjzxKFdI+0Int5uE6eC5U5DijTnXzqSqsMixj6
izSlXtkYfzbcGagEVP/tvkBjwp2gOQqujn3ySt2hKnUPDjc8M8fkcv0FIrwi7Ysk
xKzJnqOPOyWUQcmroOJQwR98gyjgV4MDVxrKhWWQhqWWlXgEiimQC7zdbmvFZ2K6
iyWbxO5PnUZqh3/TUAP7ZCs/E0/D5Ht+Qcb5aR/M0JIF2JH27d5faFq83iw8V+sf
IkZ8n3GD/iUPVck8qd+TvIpVdXhk/cmEFbHzncXcbNM//rBuDCLPxbeJqa3VHdfn
wUcEerEW654g9J4BjJ3HEagcccBK6233vWGBzoKNGOI9Fu3S/hPAYrYlsrkhd+tq
B1D/QF6sxbjQwnpR2/QcLgH4v4RQoldAg7kcrBL+mSZtgw+Q4e2j8GrqsPFdxSO7
qRgLj6t1KJ+tzAM0LAiowm8CVot//Nbadeo2ssMU9+6h6I5ty3t1GtK7/wLlAakS
HoFJdWrd0/raUSkaePa8qOiVTzZ1YgP+hGd9iuF5rVwXDNayxaPWLQM3xr2GfoPP
Ci2dKK8cE8vtytXwyMExYpC906JWRxYTkR323MYQX86+SQWw1U4dsQk6ggEw/zbO
InWkBQZiyTkdj+z7CWI0qjdyvPBSQPEkAEiwjzt/qZB765YBcvDsG5543tUneTtg
CBpJFwCEDzeUfi359L5v39pEKy8DalMF+kL3maBrwQ3iNf9523n/JITsGn6Q9WkL
BfssEgyFlqVhU4dp6w9tl151srOj+/HRZvwRl+//DPxss17kXYuNULpKcVazlzwR
V6Gb28QO5bQPJJa8mDEhY2OzgX2x0wFBI5tk+v5klyG9P0Zfnz8M4l+e58qoT2Iy
z3S6MgNIgq7oqFIMeS7iiyZ2shQyXDpfcRSUuHfUYRLbHRja+6P46TD+maMVtX1C
j7hQ+mL57C25jLLBrNq2HAzwl3pRPBZDHWG4YXMcDg0uFuw2S0gTkGwQCzlZQEtM
w2D55arQrpshPIDSBWTs9Npfsdm+xJz0x2/qVV5KrPVbTNw4BPm9w0bX+YlrrHKm
O9znSAk+RUE93SSwKtBX4n8aceiMDGe8VPBnVuqfQmtRpPVOAGp8rr4+0X6yMlpb
rclcYcAiABsvj1H2HkSsX5n4Qs1dxVYUxOaQMKhY7l2xkOhACJcMy1JlTd6tlO5P
2BA7E96OIWWLtc1AX97misw3dXz2+65eUpYxfMdTnskNw7LLjhZ9TSl0FRqzjCYU
acHNyyKnCqIkGIhDMPNTbLpdSouD9frRI7Jhqe+HroLwGa4Rc/P0o9PgPwMaS8i9
IZ36DiR6m+ep7dsWpePMjNSzmqnRbOyQsWZvi6fdJwTZqTSDiBtT1RsO7iGQjdg4
6xMzkplngtiMK6B8bfElX7zIaJfFlHwoqQ2p8sF4tFKk/lh5MTtwbWRFBKvBK4AX
tHEjz/qwDSm1x3r9LWu7GAubULStxb7a1iDMzEZ2wcpnC4yl5/413U/DuvuKIyfW
vFn+6UWbdJr0HNOmO80CFUanKxyvp+/8+ZUnKFk2AuCAsBWOU7T9YuqpMKZ+2O81
7HS3D/xjaQo+g3YQv1znycM2hoZ5UuDD0k6vEw8OYzxUnJzIsc0GxqJaZEp7zjjW
SlecbtetuveejN1PpWHJmxknfaBFYiAkzd15br4ly86CM1xUbe4VX568d7Owjlzu
a5Anf7kHNd8nSkWAxN1vWJT7ccqsWmOtPdqmxlX5NGFUXW0Uque16fh2PieX5Rui
8lVdSZkfRfLwLSF7O6YngeJgc59nQGuRfs4ueSY4WlqBSEOJSJqfP6BJ8XV/mc7f
Aoj/yKKtS3UBG5z6FLjOn9O4W4QpHSEQ/MDnku7qSbmWd2FG7CO/f/9vXEw5Bkr2
1BmNIm1WmrR0R1GD2BsXjj9XttLPjGYMpAkCd9bHprsAzP1cmx+JQXfUAhFSWkcM
LedY8/Smy0YmiFxhF6opuYIiAq3r/ue3qhFoEWe2uPeZL0y1FvWRmBIqb3NDz16l
Bz63YbG2OS4y3I6d9GfVJb4jDUMIObl6+BVZ7+G/uWm4wiuRUQAn4gaVByMVaJjU
2FJqryQvyIg6mJXT3AhrF/MXjD3PDz+ZMFx0ieHgGv33++Dz01i83qMfugo3YCoq
jm0croWG6mxPGYSe2JpaUuh2rEINrRUUunQ00teLE+PCqaKjur8Ivzwwycwg/HAj
XzJm9MHtpXwUOHZuhZ/+WdOCcwPNa5jhicdahzA+qxThF+LN2JJqJiXHfgyQFhH6
lvNrNaZYenlFNOAANCEbAf/5+v7NVxhaoZgauNtFsImDTVg/EnshZK7bAJQF+JUn
oZz3GcCpiTaf3LEu4sD31c90dhTyInyTbakN2YWvSNEVD4/vlNQycpma0ajhgBIL
TqstfaWrnTcETI50mOnDoLNVAPLZfvmGdLq7f+lCXTAVGLJpjQ+KQgAJELHOPfZv
31POIINyz7kZXOllwkpTpepsamzTNcBqCtNCnwU+3qJxra8z/87G5n56HQRushCf
B2/uUmhffbGiaLjY/89Kr1ZLQK6J53GWzaqDayPy2APWFEEFpuXLbuUCmUvOn8DD
31KQutG0YzIWy6jsmv9JwMfVEtL2z9FH9dXn3BJ1xACrTK2af39EkABeE6UKv9Az
2pGJcmkkiGiuqyknAXxnTkkdkl1xG6wqDISowHMQaJhuem29lbODEiVGIgApCV8N
XR5vo7P5vwBGdrpep4jOj4qcCqYjnkhRDlB2MmR6F9od1p5tzds0IkMc6pNfcmIa
A7NXWyP1c17Wf0wn9aLANPOmw+n1KnjBFqAW/7pmAoeUe0MJxBZ+rhAk0gETlXjD
sQzZLrV3yrR+sqZyXqJkuWz36eW8b5dFe1M1sF7fldaZw4nnxH07n667CX18okYx
eedDm82B8cjENaJXHAuVXKUXEQucxNw/eIbyEb9+I95PoqibZrjLih91QnTLrPrk
V3rokKoCDTomC78jwRRxkiBlQUCrSiHCYQDYaTwF66bS2/4yZpxklcpIjgXZFGd6
97/LVKRAGAhysaggr3Ax5+X3isHkQL04KQdi2sFws8MIcvGre3KZVroW/Nwmn8WY
pdYevnU+cg9rFRI1yLRhTFqLj+kn1rZcHzJ5Ll6bByoWuW835/tA5r8vD9ZTH3zg
GaspIO7szx0Y8UZLWe3KALagPlE3cFZu/WeI/By72+y5/nLwQC/fm/5Yq5CyK4E4
44nuU2vemSiciy4gVf//s3GvCEjkh1mWyIHKuTtBYi7JViVHSFeJ8XWiI/+npmVG
IAZo31r0TT4jVrtOXMrSppD7+QbUDHAWz+SpS8jMMXIdfCcLWqsVgyX6VYVfok9i
8JmuXVKavMofBOD0mo5yKUyhQvRM0hiXY9Cbf+0pciLRcplyi7uQftJujixgqTlq
DDswKp6L/0L0/y+3zoP9pmXFdjL3VSUbP8k95Q4M2/C/jS7h5yZcoIBTqlZlmdU6
WRZoG6An7S+g/So91T9v2EA9eRP3QFSejhbrRWzs0wGzE8Jfo0F9wpNL17xtBzuD
Z0Km2p914LCOb69IpQ80CTp1aTtwST5CPdAlhVaSgON01BRC+wlmFClZiBoayqKa
IB978clUys8SIb/EUa7HTXlj7wgF/498USg9YgaRCwcep1P+4eUZcgdEt7uOixYF
Wa0zhIZyzfV1qcvdb41bSoADdG4sGK3h3Gq8b/hXiBU8OIpZNy97ctpXWC44HpY/
BkLztWjFbtpCfAC6MuuI3b2Qi6vuWfqlhsI/tF5IXBiSgBEbNxuJOUWN+LDZVmD5
xElGiTAhYICZosJbc0bu3FofjRhva7VkeK/jncBqpDDMgaoqmxVmYr9AdxIpW3KC
qWfIo7XPhRkR8Tvb9I8m2EUmuMeAy1gi5RKGcnHYTrzwaxIWiGsktbrEDJk9kdUU
E7i9wmniBkYqqsO2kpKdqq4pQbJbfc5Q5PIX8+WylpNByP0oecYeaIeYtXPYpWJV
bDjtJk0SHth6YQZu1QBkBaH0zgWsNaQe4nOgcnVnM5lpxiu+2D1ouZ234uZtQMYw
3NYe2T4yLr0GldIV63BV54WS9cpQeq0aNi158l0CJR3bdWpyYevGHI65gongIynL
7HSwkeFmwSyUcBQkkOUC/lNC737QV2yoyDLR8h0a8V5Y5IASj2KD9fBxKuympQno
oq6sKlsrO0WlhffA6sbPpQxr3Z+rFo9WXhRtEf01+Hx1uzKt6gPuZ73d7B1R2HJV
NbKrs5ud3uj8Iw90i7ZH3mkEqn6ZJFHhuIElCHMmhzR5CViOEGBFc6+V7uEmScGI
U6o7QRYuTHe51hByMZ3zzj5Z4JJMZagCRqROgKgRcgPktuMlqiQ/ECQFbW+ZTdae
EgmV+lahGN9Kru1V2Uv3EqbbnCokvPXOvnGpEbaiBzmhdCIK7a3DJC/hE30p5p/1
3SEhiUjKu7VKZtyXQzidA++cAp/Kfw4mLFDLUZ1p28FrzQnPwSndOSH9j5UKkbLP
m1NmilVutSZy0ePyGZc/mshJuFva1Wh39ehfvi5E2E95Us3yx/vldLU9wi5XcJl/
85X7bn5ITfPjE2QyYagPCHBSj+B3Ka0LwelA2ZA24wj2cY7bNvxgm3xAXS7iELwx
7MWVuvuVCM+3KE6+T82IVb7yD29v6TVY856uN8YyrCmJrtRNV4dDS3tcdxG67CO7
Sqiu41wuVKeAZBH0bUUGcMMCvySALiRvT7BWStRNtZszj1XS8uVXJOinae8yvz+5
8d4vFVpNbJmUpiQjpCvbk+ggvRETt0rbOy029KquFKZz20gGD0CmO5URAnah+/bx
9G+XHgVee6em8SaR23xaUMhfpN2EuvdklNQaOsCeQNTJDhiIrgBCW1Er/VDOayhL
DSY1YlltwhO8vVhrv71sHO7r+bQlNKrTXYs61uy6OVTOhVBf3rcPIVqrywPwWinK
90qthrXXn83VaxRPTOcBVt5ZO+wUEZpKUEu9J9nd0rxutL3R3pW1OyQOyqETfsIZ
G7YEpSh1jbPe9ni1XVa4aguwSBgu5+pNP6j1kiKBxX5AtUkJ01TkF1EWM9tai3i0
gR+jjOC0K7E/gjqFTyvt0D9JqW2/m/pQIJiUh1cKQWYOacPyvVobNRbHRRjiX3mK
dMujpvRoBXoQQdyHZkNwMqdpi22Qbrqud4ZclC1OacRDE+xcNTVIZRNWhyFsDYjn
RggyjhlD1L5A9npbEFwq3wFuR7adJQ56JDIjnTJZcJ1NVa80+BoES7KcMmD+1DKg
+K22KH049uVMHjFg/6Ek42lfNxIaNT0nPNrj4zOtKGbJwxOmF06MOlWChglltVxI
Q/UCzqHIEMuzjvkgOC0UtATJJiM5eqHKCznHGjYugAWWH0hJ0Mb+SGatq40HJ+92
oKk28Gt18qKp45Wxk27s+KP7q1WrjXWHNErQNm8W6hGnG+aQvs6sVYfoiI7OMZno
0SqpKURZe/1Qu/jX2TSveh/ivxqLrLAc3vbfIY464IuFYZE/dqK9fqUZRg1JP7EY
6227jCD5Ehl4J0iL13qfoNqn7bOwlDFDOYJZdmZAo5VUY55u1HK3tBhRQrll3MD7
Z3vrLgB+V4uRN/KpVqIXhWyMpzEzPqYSftrYQ33a4VFQ7FNrf4/dR78spPWZBBeO
eXlZ2baNd6QuJ1CT+T9XVXIm4hURC7JSJTNWBQ1xFyNgkEU4inBPjRljtzxoKxTN
3bE53l5LxMlQOSoir0fV7Cvrcb+UJ0gLHYPKpZK1rydHtEAmUaTKtouSO9o+PHEi
WW6Q32UTL+oTscdzb+RiG99vkwrbN0Kpv266Fdn+Gc250Pp0KhfT9N1Cpe8MH3Om
nmAAgrENxqnGSePevcIFHmHu1SaT6jHptZ1ifr6PdMiAvaXVPia/NOI7wqx/RVFf
hySjD7zce1uuvHSZDHmtYx0S5OhNajLfcHUuuMqoJ/aVyG5C4SmffWu8tUBmGW+x
l8zsIYYnPCJzOLq3YXY7+oPX0oC9JXw+gBd1KCsMpuu72K5a9Dy5MMyeHFEp4PpH
aAayHGkUtY/dyBQR5UR24Sqh81jo9uCD8GrSy0oxjiHJi2o7nJECthEBUro7XPWK
4dsRXezsmo7XYfmaKL+Pf/3ZMog2OBdBMFaI21bLhZPHHTj4dCFLmOr3w2CzuK3o
UgNi3Ts1ZBcQjP8n39MjYvQHNAts3QZ+pfgQN7pmuHmf40PSzw7+WQylHSVREow5
mOz1V5kR3QPQtYtuMAdpq28cJZIRwIZpmU/0RCZWNM5hop5QUdLg8mRz5Qv1PdBq
FzhH7hKemTOyKa0+gWjWc9mqsvFlw9SwJVKztS+NaNV0O11V++SPNf7vXVHWGSZz
AIcH5Clwr/eaaUSdMUHmodNnMc4iVxPfhoSauSxDh6oik9s0c4wxvzs/18QcUrL4
x5Ac7km6wwNBSZf5W7saFJb1qNWrZ8V0LzGPZE/Rlisl3iZLNK/vrLf9u/LSjnBv
zSvuQEq9qY4mZc4SZBxNPhyXn7xzOTALn1rhgC/093Sa4GTESgbZnUaq8Te3zzw+
SHZue3lSbpiIweo1Oo678Z4c362Xml0LV5PGHLn0PJNCCZRqqGXYmNZvr7PIORTo
gO+Kp9ItxOusAo7rOso9VE8LQutItxkE4Of6dGg1v+e/Mj8G9s6dObi8fxZufQfM
fipAUsfJzNVzxzGxabPK7q2gC/RTxOBk/bqZWe0vRFiJuhwhWU+hGmMsVsTZrn2F
vT4er2SPo00q9AqzxzteVTGXxEPcEi9oYWnx0aFxQfKeukTYvOV1glZsGpIjV/Yp
Ukd5T7FBZOzkp5e0ViXqEsxHuL0Qkaxaga+ptG35lj1WeaWpVLM5rfZUwZ+5fcqP
6FN5GENJVQQfjjjV/r6ajd3orPU86tQDaileaKu5L2MKOMGwGIUwBRTOK0wSSKgi
e8f2xYeA/EepTYQW7sH8qmHfgnb5hctIfpPyJesUmr5kW6BsppYrJ2OF5YIckEgS
NoOqboiztNv5TF2dv+G0I8FrLUQSAGxTBNCGZ0eP/aQFgNb5spsVY2jaP8GW8PT9
2rtBGwUvap7bKcV7vJr0qRJcC4ttvCL9jYOW9ZK/JuOsSE3k/rVXAHrWMeopNCD3
7QXiNAgd/l6PJisRUmxrteREUZAZfmf65SYLbz3UNfIwcnbNygm+OSHMusZgX0hA
dS2x9Yxzj72k/hzySf9sNN2HHvo7cKh4xYD21VqeTNIkgmpkX2t8Y5O+1Hy2qoYa
s/2FSuwc0NSZJI77e5aNzB/dqJrddmfHsdfPizyr5jzL6paI3+QmITqqMI9ueWRV
CfDYIvzUWWMeKjOEI/QoV6zVYkkn3ZinIc3dYcn/MJetEq3k8VxMXst74Xohp50D
diO6K+XmZQQZFa+0vUJCioR1eQNN08AoFrzGOF+i9rSKBLRZ3hjKV1we4Dqd2AIc
h0ROCibX1rLL6ZZUz11ndRRI0rZFStr0/rx7TmINxahAqtqvysq0Yp1V2gYuKgpz
HItxfCzfYC2PQBP+c7jF+M4+Nf9je4FUbhXK2k62Hu0qo+82nCVXJ4tXX4Nv3cVK
i7GaZcjqwLiEtU7YGqunzMLzcaDghFRUQAvyUaaoa4AeAj+HZ45G7zbHiC0DF1Ju
vRD1SfCaTZXQErAC0AxUvH9ZCP03o051mEa0Pfo8nACUT2zztaPmfkLqHqzHFssJ
v656q2Ll5ovj5OXCv5jqaA6JTlbIV3UKF3iRNmOarG7LCpV2JG+LH8HXs/TmkumR
NZdeJ9UJVzvjYE9+IfJOT3F5mXRKjJykLKlhUzC9ivf2MPY3fsWv5fKpnT0538gP
7xs0Yg8ywk/5TLChNv6sddR1cCjIM5afLOvMRr9WTf/X+cTmG4HWIV7G/MHLPY1D
MQSqb4UfeIqNaVj97mK/sSCeZpAT8Y2xDWDIAg+HTrp/UY6HnK1ZRxpvB9tEsJnz
WTM5BxiJRPj6CTIE1+tAQxLIvY6ORwWMRQ/ysq4UDaj2rM0DLu3E7+Ph7gf+sPUw
hkAVSj6ZLvK61sEht1QZEDcim4jpnJ87xnhzfzBQWwTpf+rR5wTN5y3vmtmi7Ii5
+fq2xCkdomxurzWQNFnT7BQazJo0HpEWHSIcsAtFwymyWcRgLZX4WhXiwjr5We3a
SJgQiSD4IuuP5XKzEoZuFrACzWgxr08S3kXCChGf0Ezps/qgey79gosJeJ0Lwaqd
e4R3tTgfRrfSsBF5zU0qGveyuEBQHQEpP0/pE479g44R+ndnh713lF8t/MZEWEwV
K6Emk9Iy65ejETas8/AAn1BUAzsAaTMhJTU7YXNg2yGkJbOOxsX3Iu8vEXgTsUrC
CBy9lZBwK80JlX8PySu/kKN4MRWhHyTRbV8QHNjfVZtWkstg0KI+4NKWEDzD96Jb
l4oOrVCPW/8Nm9zephi9SmXYZFFbS1fNILmbylYmgLKD7ulG6bNy8S9+jNWW+TZu
bcn5gQO4mKhJGsHoeKp5Z9CWPPBSHj5wS7DoEFpL8JAhpnPuZ3ps8N9kxeZ6K3OJ
T0kCtjBH8PidpTCUsYmShDMWmRdvt8drJEkTTpIKTmUrGGhrooXtYnumKTk5NBqU
vDIW+JsibOC6l4bB/GFa75G77hEM4twsA+NFl/bRZcpLXX3xgcfyaNSPgjS5qUFK
4HoVIKG8lcRaB2fe870Lf4KstAgqyFFANXo8ldvNSX+zkoEHJj+2D4MiTfv1unZs
5F1I17IWE3UpAEwNrJy5mG4kUGfZsRPk0ftV0gw17alUvgwVQoCBHiiDpXAk+qBh
/iK9iR4btXRK6AiIjwb1J30hTjP53HXY/WElFrUPX2qSEOnE3xcSlWy1mBqeUl6X
W3hG5STOP6NxyQqV/+LMsxoYuQw6fSvu2A9l7YQ7JtEH1bnH0SdQ+swwkExTKD8v
jIp3X73bs0r1Mcf9d0d7aVl0PoFGeGWAis3S1RfpXBTf05/byLeosWiiZmAHtva1
CCet6SQ5uqwe0iBp3t6TjQllVQipoK0y82Zxye3kROav2HGXuY6Sdc8hSEYgh4qt
P30LXq21VlZCYZ+cVa4/n8hj+uaLhfI49jbee7fRHomnyWuou1fxhxWI5VacflYn
gj4ypCXYeWjQEpgofll3d6qXfmDpvApEhAny3FfcbkAHBLKVTBWnipzmqp2W3hz8
pRZfBtHdzlW37OXBbFSGxxLoO6jSlj8vQ8P4j1ik4Ifw/qvmPXo2aEy2e8J/OEsD
CgS2be7/1XJBTnLEVdobYxs8LtBns3nWq90PEphRBLJaMS3aDb0VNz0N35CFgIrL
gVu/c38b6DaQzhF4c5w16qrXrHsH86cWrfmrQPfRmOqlKN7bLmTSdDzg3u8mC5Jb
E4jOkRT9v5QKfsKOaR7c5U81A80deD6L2mlUyuhyj1bz5UwhLfZtIv1G6e94a9Cf
K4ZUnXCjrzTG4j7g5UMzxqptnzUqbV6pXPQQ16mshouREe01jp69ALOMinbAo9LG
nFjcU5Y2Pb1+49sZhOfhBhfz3JjhTqiYYrYZX+3GVLdhTXGF+/UX9PkJpbAboJUa
a+sWCkE+fYhDrLC32diaLBVqKRYpsr0QSbaK4z7uZZIutUYowA4U1Q69YVl7ryIk
VgsgIrIIhZEY5P+KG/buhflJ3vD3wpI4MXshXEwUWNMc7vaNmlGL0PIpaGm/Lzt3
hddzFgLYkcuY8+GkjivNEL1lURd9C3s2aTvOrTf+atbPUURbAyJTIGdX5Qhciaos
hQpcKUsvCBUAAVvWtq/69iKgMQicIJqOMLeqsUmr5fkUbUn8O98DztxnKgND0k1G
4YyUzlc8cKXJeAjYHCZfig7bONpE38vD8M9JTiNKWWAcOR683G/WeG8yuwGaYUeh
+YjdzPJkijqxDm+Rzt73ntrcmwfxRVefj2l0IGWoo6ABqcLNXnor1q5VK7YL8RHc
Hf88DfuZ7uSHjH/9Coz0ltrzWppsTllst97ciNfjdFieyAykxcLAG82TDLknmZsi
1xl3WLQaKnpBdz0r+mMrFoukT4dbr4a5Allss51zryKye8gQI2LzaXrk+h0UoY0j
VeMp+MRAcF2aN3Scph2/hSI0iq4SVJSir//DLFfvQTf37qUs0Ce+ZRBSKx+3kEp2
Xj9Rr1X6VOlUEmjQ5UtcuAh9zMgR5EXx4/Kw6xS6/j4vHVw6m6hPFnRiBCKSG3oq
Z5My1ZwYl503m/p4dkvU5ztVOjw79H8F7it1HZSd2K4XMheY2nqgn4eiVieW3mUc
jXPnLi/7HlZLiQ2894cpcYDCtMqtD3cMUPGy5K/mfxj8AjJpL/n81/Xr9z/rvm2s
WKZaFi+mlLZ0n1AkMQsUhHsKvEjQprb+/7NuXHep0wIxO/R9Vznnv6NXY6p8rMCr
vVmyZf0jxMSc/Tx9MB1OswKOK5W6EJKJan55NqZGlpIQrWggbRtyrhg81Z0kO7Fh
ZUUgZPGvR6IGfFjkVvQChxdPCt++0al7k+2zbTJ7u1uMnAtV5q9vTCQfPvG6suQi
uVdER5mpCcidsvsPNQJrl0I8LpHpYygPA6QDZPgoKIu6qme455QhSPSUJx7BQAyt
f80RJWYzUDNOQ3ShGsMpdq5yUq+A99Yw49uJlm51O/vq/s9YkYEN2J8KJZQR3Z6D
IqHMlbBd4UVM6TAKI4xSWKc5rz122eUomJE6urq+2G8KVNUFflXt4KRXgK3zkvgp
6SXnd8kIEb6lLvMeWnA0BkJ+l5FdoW3n2hGybAKPvGtr/IhJGgd9UIU1H+BDHx32
Qaho6rfD03XZ3g6Rs/EKw0tkrUHz3wTQDohRnrlb7I6hpzpd/kHydpmpF0FqVls+
Kamj4tzxwsJXLfOUl0+TY8nyd0b/nGDgkIVCX8Gr4TckDfTvF3h/SGHcSE9TTyeD
gwbOsQTAjKw91FR/jMcEXL0kslgcM9C0MQKuueWIfnboK4QRYLxIjifvBrBRFNrq
pG9HvpBaXlpgLjJj1XjFv+LRFyua0ZtCtADaDjWaEbSTqh4SYW9JuWneT3vwnoSc
O2teXbluRyPdG5Mw7UERbjRK+W8fdYm1nBGifNINyDliyEv6SHOf4Ua36/Q0IKmH
2DOSya9Xzcl5d+OS0D5YblZU1sSiVWJZz/lToimbz/2JZlzhRwu/bwesIw1u0skE
cY5vgRz6nUuIrFHbwaRVdjDCreioOmAbxNMvnu1A0r6sWn9pqHh5ejv8xlXuKCwF
xfzNbJPLxATg92IWwcCu4W0BeBw7dTCMWHW1HTJNLaV78Wpr2+PA1jNnuhsZt1X2
Y/bwLWdUib2tAXINTZ9xGIl9/FC6A81VyFgB2pjFVFvXXWyHne4UhBmh4A34k9Oi
WEZEotjG7ih8kOyC9vP6vzTdYtQ8XmoFlJUM4x1wJv9RNrFtSACIo/vAMyBBRDXq
z4JpIZEuVnyWcej0Sne9ZBA187q3tqz+OCanr/K0PhWYyEqIg5gZpI237YhWragF
RPzn/a5fLu90ddNDK7aNkG9XlpMCNex9YYgQaPf40fNuUL0beap99RPOas6xczEB
9T97Y8JAS7n/izwISkl9SSWpptvTs6CNow27G6YhkEQ8pgOlj9MKbmcaRdM74gOR
rtKdMFjQyT64PKs2Iova0K/505IL7W7rTHwl3sfWVw34aEGT4ul7XjK3Hioq3pbG
Psa4Z5cbDglcrfOuHMl0N1QPySBPayj/o/V2szSz/tSA6GvPtt5CgdMM3csnlVjU
UzJYOft7hE1JgU/uUewht4nlRkrSOxOOsYpFfJjA2HNqkcxU2WhB+2gb06/rpY77
pnZU2QZDrLtvvRVmfUQ1UzqWuIRPEWNX+k/eRd93wHxmqEYtUffFlhyb9p6fAV2s
W4DLHTfWWz271hW2V8uIn1OH6Cqy+VYW00KRdfIscVWCxZm3AqUOdpTHV+br1+VT
gWbTR1hGtMkvTWCIasBEAh7fSAZBSll0UFPiSOSl4V1Tv81cNA+hSe9LZk4FrSzv
abbK6ObSHAK6nQxuxz8ymy/Omm4Qs0gSNiwvRk4+L1S2DcgqMd55x3GDDc3IDXgs
Hybc3S+GnsZNcmY8j88XhNjFT5z7rjGjLyT1B14YzEy3QNch1yovJG92Jl42MSM0
XxC5LjIQTDhh69VchRswdS/aGIxkUyau40uBHJUbCnlu+Q65+EwwDJyBgqxzCp2d
xkT9Tb3wKbtnPiagyr4PsQwx+UrVMVTuqQThFHJqwfo+SzKWchsqIuIQnWt/n1Zo
v3mvORgQwh2iAqmkqAuRTqWVU9LXgqqrWLocCENLeD9+j1wjCjj4Zs4GgSdcZeZZ
/oMFm/DGyxmnXTnqj5BSyNFD/W1wFag3IuYI8VJNAoiBk0yZoa5QyjzAsGTUvCOf
zIOEADe0nlmCLLgB7q7pzRwjWD6IlJx640BGP0C8lIumoXD6HX9gTpmcgphG1AuA
HHF+2Qvf3ZHmX1HeBrzKJB5LnkTczSKtEiqXr4wyQ/fxDdOdIQtP7Ys5peVXxy6e
dzHFYJdug0kPR60ZN9el0PRpAc81Qn5T3Wjo61owQs6rCV7ix6xaQB1Qttvfl1RL
71JuGDZW3S7K2rUkXXE9jgXx8lztEibvUUL9aA82Lz1lKs80eTUeAd1XJYZaB12s
spliHFC0nFNobjRrRuHUxl2m5/6KO3GzbK9bD8MHOI/F0GOooxcYBccOM0F9jw7y
pLumqu23JUTZip+mYdLMKuOBqMpBNr6yCdIxOPjcTV+wVd39ovQJ0ubMAYKEUd3e
xSaFz8sNja+Fr+f7bn6YM4O4790oMsFLr+wAjH5aVdSmgyeXCpm6fXJeAwsY5lgf
QZkIzOsg7Q3Kqp+nH3YOGp5J49YNV5OM2EJthzPeK0mKGaS3PU4+9lOxRZDctbKz
WLc1kVEE19/iuX0ZxJq1hbLChS/Gg8gUxZ7I4lDD4Z8Y8CiZlu69ZGh2qxi0DHKN
uhiqCi/7hd7lKsyszQAGJja1MqfPEfLCLgB7j1tqONDoNhR6DFCmnsNQjP4o7bMW
bNhG9mcjfO0bN1XuS3OmOSsJZ4cYM0BJoUR5PCBFFql/hg67Jkv02MphBr+6fxhL
BAihoeqHIurlQ+AgEdAhh4yOkikr5vbDx118cri1C0OYmVk/c+qvqRV9AdAQSZDq
5vtnsw8guJiXLrlahsfvUp4963TUqxuZHVN2RwnHhDWcbyOIXqbQRF+zgnL+TmmZ
eed5PvMCzEXjpaoYBBJlKOHUUfAqfDq2eF9ry++tQtk2Or1HWGnRrB/3hKBYSsgB
N5Wxad6ltDBydyVn3E10rt8RQb2pUgGFn0/fW4UWdbihfawsNsheXhegQWtbQ7hE
nRSYzJQZVa0EmIgy+CW7i2c3C+yv9pYl+K5REsujgzvgBCg3Ld0SIJZIT+fXHFkJ
du395pUfW2Bfj1y9YJAgQFout1L63RABHwV04Q1cQn82b5HqN9W5SZDMXcnC401U
8pdMkgcGFcvyaMQnkbQzrSz+yU/mVc+q1fI8yk0CWnlvroDNZYfqmthoW7Wo9Kpz
RYdBSs4PpQ+oWNPkdH2OkmZSCeV5XJ5hiBRm4Aqz3lVM3sjDMTcUt/RfaDikk+VJ
yPNCNXTPpyyzFXfZyoQ7DcV/BvDjK/Z53/BJDf1PwRc1brFiHhGY6EF9es+1qNrr
UGn/mV1/R7TX+tstD36Ka2EoJpoBWPiq7HFj/ahQGQzABOQUFxOXRUnlOivkUnmJ
EgLMFSLVPuGm/5Xi9LuODWNs+vIFd7ktHTNiX69RpJh090E0zsUJq+OdUu2FCogQ
s4AAClR69OVQsklp/9yzM/U2GyoO2RXO67dLYwHP5glA4O9II894cRfMAPsP32jy
wb3C9R4aqd2coI3FTX+J5KFD8pxwUch2TGZdTQk/zIgjXddzD1Ymb9iwILxQnTZ1
Tw1B70PLvcIvEsFH4Ojk4vIlkIbtEQhauFC63Raf719IZmcxjMQi627+Fial6bhS
a4V3Q+DcxZt9We07uvzEYIeGwRmNrMkN+z7vRk/3QzNUoNCmgyOrVmGtOz3a/h08
TXevt/Gw5JwIAOr2/8AmjgTtqS0l9d+DcP6StUgnGU3o5ZUr2fY2VswrvlV/VDX1
XtC16qlq7kNCr79Y9fi2IZmf+WYpmejqLwrYaHvFTSZvDYdZ/J/R9xLCEziOQR1e
ZxC/HB370drfPy+V4RI0uo0BLSAi9eXcPMJh/Hdvfy0dxonFO1X7xQOnxknoqjoj
BGi2QujUmYlLeOcVIujZeU2UO0XnUCCFAw93zrZqQhuXGSc2xxrxzO3XekATLNyO
oh1BPhZyQGnuMbN00rYCoruhrXFAfoSgDQ2PLIc4ErjnvwMtWb6TrzfThwhyjVqg
WwxUSW44Tu+XMPbjH0oTCrV937XEYo2JutFLWhV5Pszd29RSPVegr4fMruR0XEDQ
q24sceOUTCVIEJkxYzHZdQF2gIXfkNfv3GXHC8db3CgBzd5YHsxnbgukp7txIJRr
Chxrtmjg5k3nct9mEEjT/vAl5Cu2iErQ+qgyWjz+hZuYgORFDCY2TT9uaRQsNzDg
EogKk7WHxHkWR570wLT9BjVbiBgTNQQkBdtgAfMNXDtmXt47+nuRiLv83/7fARAH
0AW4RZAp9ByEZKB7dECmwRy+aY/PRHvHPW+mV7So2O2+j24OnkzwbtAVyp56TlHM
1xcv1HVBWfYLUWDqO1atNhC5iGj78Vdg+gX/sZ/swtjg6oNTZt4kAl9qXN9dlPdv
7wCv1heftnlLScqU18TKNlR0h2a502L2HSUJaeAr7sURAblgM2a9RTUWwSnNr5tk
XiVEmnhHqtnn/5hHybxzemzqEuen0hfX25OKwglWtK9IfDPyMzW3HLPIMsOPgxY/
vaNZsyfVlT92fit1y6zadywVfcfz3zLzIGi+of16Uu1PtFdQBEjruautuka7vBM5
wXcYZWQU92/ksGCOWqGha1cgKFPqTfuE/+9cVbvRCZTqUpCyBS6mMjiC7oW7rOa8
EmR0h8oi3CyvjdT9ucdiP6z6Oqa4xuHf1LFCzm4dUVpS3tVR500G4XCYtwo+cilp
OD5l49pGNcv/lPNKV9vO0VYe//qlHTb1mhG771PEX+kh6rBUvcDEI5zBXYcwrjTW
MmaWp7Rbu3PY1q750anoV4g+Sjh2tVoFLKMojXHOiUX9UD00GbZ/Ms1vG6/1Gmlj
/izNWGo8BmQty/9zkcOr1iE4yi2jXtaKOYiq2jibkI9kJcZHPqaiB7GZhewiYTS5
0cpe2UKdPTc6+aFgvgmF2yDcxUIy7cSyKRZftJ2CLn2nfjgKWCb7raSTXTqlPdzZ
Vsdvw22smYdWRDoLJH4GMCqx8r0lhBlmDwPS4MXyzk57DHHht3ZIFkBv+esyVR6q
g+qY4TnQjburOPDpG+mO9syUhEQdt3u6VomN4y65DoRSjzH8SukiLP5yCLWTrHzd
/mZFHlNMBR6atexO6LKf3zCzdWzFz/SgHVp4x9vp+FtTehIhERsyjOVADYISIwez
hEM1olzz+2Ox9QfgKLN6jZhbYZrTDXsc4r+Jloj8Vry3sWD39rRfPGwKkfujG3me
AUNownetzoyoRjohiWuVghkLKeEzvlUWjwGGYtCrNXEHlySEk9ce/AMIDUYC4tdo
0HhEoKWsfld6dRE4lnbt9WvZOXCWNVFTY7GiNZoemYPy8H2XmEb5H4/Ukxf6Howe
TlxQ2uPhIOKbSW1YrB9lD0uysFSn4TIUzNl9DgwQzkW5pUy1FKyirnOYDmylXiGb
pwjlGs94QNpM30SdnZ9GWEGr2wb3MO8DUqbQRwNdsc1Kvq62vXraNvoWQ4zjEZhy
SLhMVuBAHhE7gEdytqDgjZ+SJe9RNlYmfUSRYEI74UJX8CSg3j4M4jow5RKR5aBO
eRI+j9rvPvsuJz5YRBzw2RjJR6+BJYAvNpBVjLnT5tyEoafHGRu9/QFb5tJ1Fb7X
uxtCbKP6HzPQDljRf8Qhq2I2QsVFm1FgxGWz+DCYlv4AE03R/kztkK6ncFhMiMM/
yw5gxRpZFIX6S+EDoIiUDVibWJDclEU9lk1CvdSZD5KcEA49eqQZWxTBQ6FQrfRy
WH9YVPfgx6Nysr/qNnyJLJRvPQHLImv+VGmjUAX63y1vjm4xTnzfcoWTf0MbYqtS
Ba5fQb00+8QItHaPMoKi1Jakk8QiXQ0s7OsBcqraILTzQB6xwKtC5QpMujyN+rS0
pdb1x43EPIx7eTbp8kWXq0UzKUx9GnumbbIO8DGHX8P2iE7/9MNTen3gannJKXDm
l8KUYQ/pA/jTzaOC09rikiRCOSTp2v8gTU8usJvr//fgNKGEouBPhEE1NK0qx6u/
+LWa3s/vegKEjijTOIR5vwh8kTX9lHRjDqc9buNS2+TGAjYVTjngYUUrfMZJ+M9q
xMw6ISzaBygZZbRWvJvRdJB/AxNePqKEXYzwhD07Tlk+OxOBhQEoH4+DDiJAEPBs
aurOyRVk1+Y3AhINIdgns5hEXM5C7t1BGEHCkNLo2oon9dYtd56lIIpU4YdQjE6j
63V5gBpa+C10kOfXA64khUITTz508msxg5kYg/kfiD50dy8Hzdln5VFQn04+SE4U
b062/10SyuPCKhDA6oNpFYgp46pZ86J/Zfg68qny8PKuQNdbavtCy97OaIOd/JwS
aRfUEtJ11ZPyBKTkIcs3H4Wi65L10/9qriGR96bC9YqiqFkLs4EZ46fEbqp66gtX
hKI+dOmYqbz6Na9KZi8MqgyAM0kNr0DUTxBVJmpqYF8+9ikLo0swKodpy90dUnWT
Obd59CCOBE0L+RnQm25KynlFN1yT5yoIeBXRDzrBf0KGXCnevS1lhdR2CEh4vYqc
qGBN71dIz7tB0d/8uOyamNu7K2hqvT51rXeZqUw1xd5kTawkz/tpr1BERWotrlYA
vi6VkPa4qaGjzdzcuYF4bU4hDEG8O19HkXrnwSoF4Wdg5CLup6pwBj6TcbbmjtqM
0Vs4loFVbgUbB1Tjh95z1D/ACG7ai1c94gLDLPSg5u41ZRnHBrM3GzMaNUDKqSGL
VJ48auZXMTCcW5dKp08i75Kc/ame100Zeu4XbJZmBSrs42eoTSAdUamEVMr9Wt3w
BrHdCbE27pWsS1TRqwkLtXnsdSA5Lwc3n+BiydG2lTVZCjZEYT08Kc+okHPW6Y6y
Ls6N/xtweCxDTM2eU2Dls/Ma82FQunxSe8RLiti2yNz+n3SpprJj3cetQPnfR2GZ
8vz+UiaVSUuad64AvcqgRQxonrzPuVbuTc8V1+9itq4cfAECVH1DO41EP9rtM7B9
KDUfPhdYSsn4BGXKha2fjspDAv8CmbFzXfkWKhirWhVWvvOtXGWVGL0FniWpF9Rm
flfXQU2chq531cEZVjc71CBEa1GdQfwosjaAh5BuBvyX5+8rQVz1aNNx1JyQyS8r
H/pEhvS74Ny3apPd2sfRREDdBZs6snMjTpn/6yqY4UmH41ECDGUqxvf4pmYnbpXF
+qPRVhbXgNly/SFCoFuOyqIqiJKZLznjFdA28LHLq5jRN9+GhHWLP6H0MmfTJDN+
lgC1BzuLt5/tMVRuu4G86qNf/ctCR5i74nTmYwqZpCs9qtCrbCzEM4hDdG4XBwdr
FvUHYmjmc4Hs91OIWWPFNNWgyE3B00F5M7RLzhnEDZW4wL2PXO91We2bNsQ84jBJ
uRFSGPZG3DX0L9IFarLszuYbYvG/uW7GB4E/pkiZlCUiadm748F3yrgS+UOyhy5V
+BmMGMjSa1AcOTY8+1DYNnd8xVKmuKPHTz/TVv9NPHnLhEueuhGaYuXHpxdfNWwq
zffcBVCrQ0sKaMZcub5rvFop0oMfRZDvWuhYFsnf+gNdH7L34jtvzDnbyEk9wzmW
GfduEBsG6MP0kDCSULtdk+zJcnwXfnpPd4JUeejRFAPNeYsZMz8VdU5SUZHTvd5C
55gRYpwIQbc5ZMlz4h3hKtDLdXHJVoeT+3Z7vzCg/p1UysoQElV3EEFoYdYWA+iH
PO02spY3MRik2a7YJxwNbY9z39I7tJG4rVPqX78dIx5UU1VwFqfUm0XLKZLh9MDK
Qtl3RsBXJ5+fL9qnhYjWsgKs+ALGen6hZ8dkqieXsVnMWk03pKjzQTsfZ7EAJSr3
nJUF3MYcrNXLz5ATHaDRk58nhN3YH8PV45CPBATxJdpFpB22/PLAy1I7plOFPFSb
jHuWcsAgQ9dciYF6B6SNzBs4Rxyz0HuhMSF0pVDmuvAnxM+MBgJq2S8mw78b0jWu
yBQS16/hoMNdL3Bg359QPg+lzGucrQGcRkFQjvFy7zBUF2Kn+brSSDtoWP34DCaq
g+Ct5Z3LqcF5kPpC5EiQ1ySPwlOuHJRLJoKiqNUw4HudF+/L5euLk4eq6KS83dTc
7HNHeOuCELd1YtHpF2mh2Lvw2VeqC4/ou4miiok06J+p269NKo7Q9/htfQBtzklB
58vVkxbTQgJyQWvVYTj9DFmmWKQJ6lsIwfzqtqjmyLclKczqwn2M+yPoo46IWQlS
5uG4AAd4fIQVTexZtbYSZXnUDFE5o9biYhMWXVKl0pGtjH1Oxkp+34w8ViKQEzjG
9z3FhrOgYaf81KVUgm9qlMhE1U2fuqINdSNqrJdk5GoTExEaK4pEDde7SXwWCVtp
VhQhsNqi4cSaeHgJ4v8s6f+xmRgAnh/7N4Bkfy0YGEpj0a8afJbCoO/GI+6LTlE8
9MGFZJusE3aFzTQBc4LLllQ+0bAPGHkORo9/jGD0BFPxlVr27geNbWvZmdDNdFiZ
WOrpbhjuAZ7Td0TgBCj/+JTE3zLRfj860BnR4E2wDq7knHK5uaBdbGkDJndhp/OK
Hykhyw8u5J31nDy97lFcfzuePbzGodd8cPCpIWIqz6/yqfQEoXR8KuLwQapSnrx8
AMvrkXnjgseYMP93PSetSQBiPHhQtQe3ttjtVOj3bD40JaPyGcefsl7Q+Gg+g5RX
C+uXwT37u5vge09ldNWbg93P9oAtOJD83mFkF3FmNrSqZfQso/G/9NlEz4LfXQpA
OemMAudbzWNCibVMX2E+LKVnXiCy2wkmL/ngPGxil09TLVCmYHNxAPdhVJFjix1/
tzHKnkGAB7L97+nblnO+lyzBE3Up0IihzcWrd1hOcu4lZx3WBaCHcUdoe3EY+pHG
JUa+f6fspeTUhpLWJGWlLkUHwUJ5glQi9HqAKRd29T/mdAhUqd5OLwqsQuxGksmz
5Tu6ukXLfu/QpSzJ2q1j4o77D8gntYKKI8Jr8hMnMJzcL71Q5vZY5/hUr/trkW/A
pACnTqK8luFYJ42THwmNERuVS/WBf5BRdL1iEZs82MWr3imdhSzrA53Hfc+pO3Nu
HUvz+0Zq/PK1LXB5pIbQhPcsE82rIQx8fUxKWT64tiauBrqXroeEZNhga9drAiBs
1IyLTgGUa6n+CreMxI2OQcm5HopLQohZZvqDEqYaNq0OLVQmoSlY7pCINgUgodwi
5vdJBm559hiLwLlGEV0XaZ9vJ6E334oPEZwgWwaPxC+vVgiht1H7hK9XerCa/RD9
geRuH/nB5FkO0Cz7nvzzcRZsOwehegZLDUuUYC6OsyuFn48nXSBtnf7aNDWUvMMr
TTv8fCDovOaIFFo5in8u62ghMF0f1E2MbO+FJs7K17WWyBamavWVkaqVZjUTaQsR
7PxIXinMbTRY1vLqHZSPKNWf1J99jV5lI0uVCCNMyfJJAg5vSDaGrnvUdWyJksnd
aXGthAz5J5hnQ0DGSR7ad/dvYZ3byfqi6SFXw3hZ32RKwSfz1z6D/gfkz8UA23lQ
A8IvD6jkWdQMTRMk9+PGL2KYn+X8InBTi6XjVdj/CsaWyGep4Ugfb1cUwpQ+EGH2
XMXbE6VPeqOF9Uo3haucMwcEil9zclmFWSu6Bwn0ItRRa1XrBG/DP5cjrCX19lX7
ISHYZtdDyQ/XhBrLq7aLvV4Vstq6fGsE8GkGMAs/PNO/o8K4ODRfu5MN7yJxCckg
ogaIBa9b8PlTK8aEvyiZctaOUqvHuu90KQEJMenuzr0dCMYAynLhVEMSiFjo6lFQ
zK0AlzfsiBMFH8XlOXlsltpJSzqrhwfpJbbXaZwW2qzJH933BxYI1HyuqTYA+6O0
A5MWZj9DcIxYYrDna/uM5kERCRkLY6xaqUVgD2QS3nHdCteIkTNzEsurWeuk62l7
BeK6PgxrWotTLYZueNM1Mc6qsY+1Jl6gScWDChMRPaXSjaM1011WcsPHluNC4DEh
AGNHcZTGinZ379FV2MfVjHaRBVxwcAbOavdnRQaig4y3Q5RCl7ATsZuGplQ5nKlB
HhcSZTR2GsjncutNN5dEiG5OMn15+z9phigokS4xNe1mycfjnHFDImS2gxJ4FPQD
0g3aJgpHvqr/15X8P0eSY0jN7rsQ+aOqizmN0qmZwvGPAA5yF5yKqpvcy3R8k6rt
JxPFbWwiaVK1sU7/AMnYzqALBm+CSVzHLF1y2M8JpouWspAX2KfI1k8LPD1Po9Yv
LrZ2LB3Yls/g6HKiADdBJ/6Mn0wt/g4nGZVh2vdgVwmMB7s3Bb6gaWe48Af7LFEI
6J4o35H0IeCMj6mGzs7URCYWaGGrpQ7phWzoE3JIuiHQ0rNQ78GrCtjYvOO9VdHX
zEdCoCgTY44eyeaZktTCFvivduJA0nezIlhNi51kMKRX2RbobdrezOYznh6QCRb2
1rGbbxapmBBStp6y8CQmz+sGK1JtNo330X/b86F7NdfR0aCO9p5gscN9yo2G054i
MEq9QAEduOpCa30VNVBo2b+Hdh2tu2nOIzuRWI3+JYIQjyElA8IrUmqYhQ5CLTrE
SRJqaqMHjG1Pn42uISc2WiFSJHyLEEMhPqNqs5CH12CcKyWaNPBnTyLNt96fRbMe
oQIputueBifN5h7g9cDf53u2ognswbklGHRKjrGQAm8Cw7DkElWscbRo3oD6u4t4
oZKacquW5RHR5uAzZr62H9w4TZa2qQnN3JZ0C9d2rxJAVP8T/qrn5HLPQvooEGna
YJ12GcuiROn4IvxqTH34sW/I3DnArcPdei4F4n5aWIBYuIEyvPPQC22zybaM0oJh
+SgYanlDSnD3tdmtNCc1ABiBX/+UnMuVTScEQwDCM5k+DwqRIY65C8tH5sG3vjdq
2u8F/xGT2VHEt7MIjS+ZQG4dabu2ZJn/PJzORRTFdZCxvMwcQOwEhiuW/OkrFVOk
WjaE2jlIGI4PmqmQjus0jlJxhI7vN1TubGmuU8LIA5Izb2PlX0HbxRwpDr2rzRyA
uwjXxrg0UsHdky2n4bXNQQ/uL2LPQJ9DsRzfJ9Ux4VJgqmpc2pU/Mt1P14oyA4WR
5q6MxV20vu3El0zoQ3tbm6IKbVbc7LyfNEPOWSFMBaJYreO1jmymDFkDysUs/iLn
s55guV/nxzwwDpuXNd9zhVAd1T/r4uOcC514xobMrh3QlnTXbUffytjwUyDtG33l
yabC4WPz0P4pZZfnNAy4q0Skp4Ky9Ipr3HgAgZ8jMM+EfMwNU9zSJIzCeijqCLLT
BDQsL/N4YbFNxkQAr00TR1vvy6WRJLChDlqzDiQCXzTF6RxiEoMShqLVsaDzF/DA
7NiRDHZXRE94Vk2A3kWs/X6+LFWW3yE4H1vT3GYfGVtU9jYVk9867/jnsn+23upt
CyB6/i/hMU+5RBLMWZFxh/CsIJxeELKeb057BdIxr4hcFgvCh7nDIZyms2qYBgio
UVQEx9VSMo4aRBwJSbcIk5NwPSaaFjbFbhY7rkANpjaOQ96RXerJI/jA+hxfBG0N
3r+Ocuo+fwPnMzMEoo7M0id8KfKmmX46AnfQSTXz+HRrN6GBsiTtZu4L1b17JJbY
cru0RqVZgDdseq//yFhAgNXDrQ99YJh0g32GZGBmRizh8hMyq8Yw0pR9VBGrHTcA
QMYQuvbfVG5gfAKeAUhh5D7enKa1/S8tTlArVBoJjoSjOgr2PzJI5XLfMrjLHc+8
G8nVdk4JjiK2DEmLj7JPm8Nc4JtzGn7xfG1RXRKwN0RxMEG9bfjhkSq+qfeNg6K1
5qGdrG3ud07ZAWaqY4RduPe0ClEV8P4X4HF5jiyjJzPyR1H7aPTD48ORAYYdkblb
MiOKzVAxA2+7sjWRveTKqgZ+0F1H/1LwFLgth4iIFwmWw9a9K1XVMgOnyBjg2LI0
zxzOL7L4AnUMhKha9kgu/yQsTHqC/9iGmW5hY/2kqYi+SkKrxf0rZYroGTzEyC2k
p+nOXknU90bOahHU1Ta5BmU/08p7iYlE4xjupia6HgJyT+JHDLj7JPgDiuRXqhHS
1WVHhJ4QfaLaNfoFNXrbzrR6ivP2Wje0+wwSC3U7D5jFKNG23VMmx3enLC8N5IJx
dATD1XYXkR6Iz1wWaLkHR/L3Otr7y9n6kfcsQAHa03I+kixXWHskAI23GtlUcQW4
meXJ1EfGDskbk7/X/OQWlZbk1rU9pa16zG7ZdJJdM5FYSqgI71rBEvYT0p1gNpI+
OWhap0VSSYxP9yR2r5OMdot6/av93Zyv/zz09qypJtxzW8ehNaHmGLsCLrt5DSQ6
473m6sSDbWVt3+qICDHIjxH5WqRKf6lvJSkb+bn2wbZPl9IvdVZwi94Kl45K1RBO
/G41slYQTBWqd22DjqPPKKS3pN9W4V2R/1EMoMzqx2tb09tBKTNuuk8WSvkHZL0r
P0VuQ7RZ156uXObwRyN+eBe0EqMWq0GX9OPPUocD4D0lfh1boGW3Gh+jrTfB/0nw
NgLu6vCcX/ZQ9PUQV6F9GXNUdEexx3OCJvzbE1SHyIe5YyTsSnqzuyIta3SaoZC0
0ClJID6Np/K+iG53W//ft2Gf5Mn09UbXj2IhTvnboh99qIjmo25fOI9S37nLc6hn
ZwrWWLZDNVm67eGVlQXMSf32EzMSkRyJoBQ60nps88Nnw6KfzINI8eN0hBp391uU
/L8QlAOF3d7c9wXW8x4m0wI6UAZFXYkE9uMQd783z6rU9y4dwvpjabrdA0vbKXRE
LF2zWfoix883C20cd4b1IXrHpRUTXCmJ+9e2+RjcqNN/Yhvb1lPACXJ4jKAIa0or
jeZk+8X2ukJgMvP+0rgoAEtjTlNgMI7wr5M51ouKWFcLzVYmEKT4aJ5YTgKfuoV5
EU+s8xMV+o6O1FDjyot33G21P+4/4uDbXCe7W6ZMe80dMsWU+POzQ0kIAcQ82ma5
9Sf9/5/Rtb7On+02kDSff1FxP0TRu1ZZeqKP18LyTqlIR0ETx3z2zDOZhmvsPMJr
Ol8AT6eC9bbrOEgsABFqn3URFqR2Yblz3jpv9vvU2ypBi+RgqziI8Fuc7W3MYqxx
StDKd0yD3nKibWTf0MQU3k38XbtB1xdjbc9amXf92sU8Bb6Pn4mhRTj3dxTKdM0t
i6EeKKMWTRxS8XZsGjzWI4lIf7qZIl8cfAnaJ1XLWmxOZyIlOmnjudCsdYIQqFAp
jfem+gc7LmFuSPM7s4xLtfYxE0moepi/7pdaPXIYQIusiNVEML1kEPUEvMfzN+Ve
9aj0q/swfoHgVimJMSSufw2tsSKhUSmBbBPbBtZJ0c6nWRPKV29+vVxhIHdyGBee
7gO0142FfZ/V0A6Z3hM2Cjo6ndPMXexB30JOwh3jiwTSFrxfkmRhIReOqST7M20T
sFPQ7RFDPAQ9KUsOcedEF677xZTmgW8muCY1ejt5+3+WEOcbwu+UfIqFQtx+9Vj5
kjWd/gFHtnlcNkcY1FffMWh08v1NBRMc1TXh3YKjN3+DHXlsWymG/31zbavKnpih
sKwtjigXrHhn+aVCLKQGvsV2G0wRb2fprlzUwbu9jf0SymeJN15e+zgmnLr6IyBl
KTNTbTQPJMxSBdS1Nq10jpAKIL4wxyH7aFiJ/2pykvvKx+wY90xhO4Yt2W1CyoR5
7VtHYk/2xwtGvu4drDObhHOo02yCFfE4fuWqjptZ+MfaLOCGir4/jMfLfrtwT+8h
9HT2XRe+5U2yOrhFN/LomQRxhhrW/uIyDPVArdnRCnmAA7WaP4fRgClcrDQ/X/ts
WcYnzUFd+n/eDs76h/iCn6zlfIwEP7LlBBfSLtBKSrlqkWAOgfmPnAnhDzg595+U
Cfah4VcOk66AhCs3ANZAHWTRHWy+fRAMG+567oWh/iwm0LPHCWpHooAyI+BKY/C+
NXkfsJo+Ofrl5Qke3IA46kMVUDBxThr/VaGvQ4BqZF2AuDBvlbfh8wIP4Gx52tNo
3pFQIQGQ5wZCC5Tx9xveOOEU35R9ITtDyERZHKzj2oZvyNiCDlD5Jp3xAGDT1Vtt
+3888BfHloZrfAAtAS9HxCg1f444VhYbcM5Pb7IJvpv9SCoiSrsGyOQ1i/DOkVAF
JfNOWwuFV/1e5tnTZw4ov8IG07OlPZC0XdbIb70mgppFphcQnaKG9vqFsJoJrLWs
WKloW13ENVZX6+e4qVwylrNiFc4IDy00/T7OaXdLgykW/FkBTwYVnp/KMzr/jozU
LtCNgNgTYN2YH5RbQahvNuiwDHV5nK2H3l/XPHk5TSVxqROSzd9VCYPf3cEqz7Yq
W5sngEFOwLIYZrEnCpOdXiBdcbKIGaVCc16koC09r55vMfjDq4MxLFq8uTpg6xTV
YjGfUDcYnJqrmEbLq8b456+M+tyHbV8dh7XK0ulx7ODQLvZKX4jbXaBhqSlADoTu
Xmxt4mP1SU2Jn9/dAY3umYL51DtVnyWKIAbMtgsFq3Wc0SmP6nGBZbLjsK/jqbKJ
EVrH/c9VrHb2KVo0hbeYVI18joxiqY6+BfBzcutGPkFaRFAf8rqyNZ3dxGlz2TJA
SeWxTg7HcQZPUxqIk6aE6Fr9ZDRhsRCc0kKQoJMSulsmzuSfy++40jky3F5DBn/B
Rw45T6CwmJMHabG9ZCg22wujxJKrPeAYNsdgl/dVNhcIM6TxBbUEKSteAGf9ctug
kzSTG5GSqrjJlKieIG8NAjFPbBLacvRlURHA+zWY5LrE648fV+phs59ElygugWAm
LMRRrOgRGRUDdu5vckxe8Q8jRjsnuMfmm7l0liZzWOdJqbv75viXcWXzt25sEM9u
gvCfH1hsuveUINEvgRN9LBu0wJkg1S4m9fPvVfKIM4TMpCuGWZWIryU4Ik2qJJmF
LMQIRGdPVLsYvwbPpXjGbi+r/v9fBlBojCf+QftVKJ6NVYQyeBMIQOMHb5A3Jt8L
f1fVGuSDLr1rzPRGRs2YR6rcwivPPmBpjoCrUajrL97VB8Cwu/9STmR8yLeUwGdN
B7BqR5RpH7jN4hx3OF6huAj2p4dMLC/IysYIvZQOjcoemlE2HxISVLQZt3Jtpk8L
ZUt/Cc4h/IQP12vWSkwHnN0AgZKuC0OH+PQtJx3mxAdpwPNRnlIGbscvx78zMp2s
aj0WXnsFShaeQWU0cy4gnlwTmAdki3QAqSjrscI8Yi4AAdcxLyQs6CPdOt4REi6U
z+8/qJTwiSCz8re8+w0Dl51mPaw+ZiPmsfcAXPQcwza9Y/YtP3dyqy2ziKfOcxc+
M5Xzon29efZDsH5rrqPGLTcAn9bzl3vKI2mgvfeJtc0hLTpwS0nJmeH+SWV/u1WA
ggKkH8zxH0TH0tIqBX2COqz7gWmhhGgGsv6ZRmMhdoIlAsXWj07A771ruhjYBFsr
durD4FNQEnJACA5OQuZb+fhSQCcfou9XzAS3vqGv6m+XwU4EYAbxV87t+Kqrmtf6
ITYhM6pfiQ+TJPTFUc6o34xOWTaQKc6wAKMvnIwWCHAtMU7kpLMqJFc03lUx18/h
QchGeRLvJPRsTjorMcJbMjWTPSCIBy3rX/E0/Dura3ovWW/vX3mkB/5AjYBtUNDS
Ux9FRoHfkEK4UDu+/GAbaB7Ut2Nrk4L7QPoSI9uRmdaPlFBHuYofp73JXDvuzku0
dseVorORiJQluKyzZTOwezgn2yzXIDG061uUyw8DFTZEZJR2LNhSJGkxshJ7L5C3
j/q1nVE//dFh0d/Kwwrele5mNRfMygB0O/uK87rNDNi9MbnPsetJV4Yr4Xrh73aK
IsCdo9GHrzRI7uQt9HbazWe/vQ7ElZWN5GqT0+TXXnnp2MVkV9Ij/jqSzpG7yTM+
R8gAyzQkjpPINB3gNXDCXcGvt5s0ivwD387J5JTfScm8C8otgeD3yCJzpGwQ/m5O
iiDGRlM/t6UBp/ItplP4g7GW1eWLoY9rtbTsCY2z7GmYfFOz0sEOk3WQi2JStlaK
qu8cyPX3YilbEhBQMBPIb6LvJ5mf5gtglaZudNpZXNhTRpYTMTvdrywO0n0NB8Mz
EroqWbjqflNIMBWFjmKO11dT0DZBYXVQ+lGLqioLivCg267F3hWOo1YoZOTs0YA8
qq2TBnUJXT3qLe+oqa7c4kVNGoNLkJ5L/CmzO9bjQTCygqKy9HzqnfY+6Iqaw3xn
04E06b3HSGG7/rHg4L6MX9hflRrbZxWP0MwxjJp13HsHfGFij2TlCu2Mz6S181UO
1cX3JpKHvu+PHobQ+WyDOqwKy1mmyY3GLuE02Ren+MpPRA5lnaRSH7KMcPciDBDd
El9X3Vg+sVGHKyx36iFMES1GjIxKeaBXPs8u9hHZOHAfzrB0vbpn3ESfGfV02wlX
2Ql0+/zFZuKT3W7+JuTcMcMNguCtn7YRuovQG2wzHFdkL3KXjH32ddyg6mfW/G9Q
QC8kelOFdgOxIq4w7P813rSclbc2N3LVjwLs1s9Bw8CEAuMh6/cQvpqf0nnPaGG9
5L6sSmv5OcHq4SRLUWCHoqshCwltrYIQ1q4VxiWH8a0ft6T09Ou2fSGyVFgdtZND
5x1XbcDaM+GndKzv6mz3lrJ6WD3ECI77sIjhJqAxD1TsENl5tRuhV5PeXIFt11md
2g+mvcH8CsGwhc6Y+1U9YyH5Q6qnHoAFZk/ttMCQugxSLYcC87y5lVr1OpmFslXU
N6xCotRPxugS5qjn9Fwv+N2G+FzjcPUJ9FZkxe/MH2ogAXlev6tl4uA6Efe+OoUd
d5puXknDdfgeX6FyOyRPEyKE/BhR82AZ9lAYxWSVcibbZloUt4KdM+nyyAZ5hxUk
Mz700YQfpXWl3IAZYvQ6Nleopz/9vH/1rnujmm+lfr8NVZpFUIMyD3S/9ZXAxaEB
AAfRU2tqfkQAiSrOSJ7NZ/L/iJl7wJjP+otFa3jQL/Yoki6QxsEWx+vCdptMER7T
Y8o9/19zGXg9OZ6ef99n3ibaPnLsh3UGukLTHdno2b25z58skN7IgnCZOsjvPhy5
nYRt8eRKmoiP0P/6AOSWkOjQ08Ys/K/LvlG6fe+MW8h/3SfEPMa0r6loxgD56Xr/
xjefAuU3LkTiI0VDnTyW7fZl3N8MMque/Arrk1F185y+c0fWa7q92OjSloV8yzqf
ZDKDJsYKFnH93wGaoK1J917k4GKNvINXftib+UYZt+xlHB2lBN3ZZ4jFNV5PpwRu
R3aeOfqqvo4fdtH1XXfBWISXVHeydt2gkVY4PzVQ/hyh8rCLBY9cGeuNS+nzDhRd
jMW/wXom1ef1/omnmuvrEziF5M6bC/guJf+s9OMxieD+32LpSOPgQqZhiBLsDqZT
D1tBrp3Tp8NnFTAhdXQNUZOVlR3vi/llb60ENF1IRnID3ronApnFQq4nTV7HwRM0
R8NSvgMYaW6gHZoUT5mZXBvpGtYBEQVO6beC3Kmmtxy6IZ5Q1oJSVE0QSGevq3px
JYHCVBs7Tpn32tADYRdWnO/UwakBsiVBJJMyl+OAIvO+hr3JIsRSKdcFp/Q+cH6k
xAIeQ3z1LTTW4Y5VwFXOw0swWVYsflnkyXsZrIGAyIgVjmTZY8ay0x7+RsteUSzF
aVYxFs1iLVCC9Ly+bl+y/f1/tFlXut4KfSMUFXU7YzjrIgpeei+SaHJS1ae4G7EL
pLeRB+2q7TM1O0UD5X+jOji/X2M42u4udJs4XHQOFqNSHG+G2YR9s4GzN/3GbYYI
2/wx9tXbdbm3aVUMt9yIGTDIOznpSYDc5GE595I9RmPtATZspJAiIuIOi9p3iSjW
lW4MKFoIoTtUg21UWaYI93OKeuoQxx+1FSE2ZYNJA7+lO29oD/kgFOKsgvK5/FGT
EFGqwp/ZkjUjI2uFsdaKLnTFWL5gDZDn/Oma810B28U3SyDPtpG+2/kV+7rEXdRI
OZHq4jb3dcI7NQvbUrqp23z6Ewbb4NDZbwVUDF47RC8G4e9ZJrz3G8j3qgD2UxbY
TGQ0LzVEUiIzftYYXeqRV1KDBFuJCJA2OGN9WBOwNrieIW9IPLA/GYEUdcB82Qv0
+XkBJ4NIjXKSjXUGWJH/25lGhgMMlTvNIFTNSgCFvjrvRViWJOzZ9z2rNi64Tp1+
JvLuLj3l/H8ejz3a5QtcIfw3gDUW3cJPNYPCL5MJNGf0eYH9TC5l+KmtzUOF8AIV
ylvIPHRDsG0gHcqKohDhJlR3vof3GKYNK+LMwX1gIVlYldXUPAznf99zGdZ0Nh8M
SlJUOz3MbPXNkDvQo3ewclL5COSfpX80hWb4EEGVG6uTJJdLN4GtR0UZETdjBXLQ
siR7UP8SabQEonJWI3dzFOKgE1l8HUoku7vtte1hkQywb+OD1OMpXu0Qxf76zYEc
bLk45D82o7deHlBj9V2pA4mZ7+2pW/O5fqqXbz4nlyg8IYBTZRWkRxpTMAm7fi1E
ryjVdvIGDMog2ix8WgxfmAtyqdBhAZB71VIjjSQb55Pd9Cdm31wrbIhDr0oN0Ggf
jzPhgAuX5U+xW9PkBTKnx5lBqWVLa9h6q/i6FR6puc5KZUTFO5leumSNWa3ITXbM
FQ6FWirLFXfkkqBUfSnyTdt0WKubRVohqNLQsAZTQG+j6Dil2KY/yzYB3JHgMqvi
pK3F34glA8cnbiAx/GZa9rfjVUT3RNhuArQE0KA7dARKeYIhfiIqEhHKALRysJVC
t1T0DG56xpAl3jQRDbGwRaw4qrAkjdwMqd0h6bwvgjC0sVDJXlB+MG6o93MaBymm
DBfYqUZallu+yDSESYX8qL24255Eg2JAsqS3LwT5EmyQX8xvvJ5i8tZC2a+ROj7u
OyoadpVNHGm3BScgel6oaLkYwD51wl5VvxhOgCAtMya+GdVjXNbn7S4+wwt/+lLc
P519gJwSPXAZ7vPRrxGO4CriNsD+Oq85iVkafZriEH9mbNjHn1B4bKfy0shjVQXw
00QLLTx7PVZn4W2Y6ku8IIvSNTMAqjEzaTEm05eoobBT452nMXFpUkZOEgEv3g5t
q6vDOZRiagEXdKAhjNOGMiR1aCg/oW87RKbqTrgZBFkIUzHWkn/r6lrl1913HvA3
S/H39eCfKzfafqtnrjpEGgHnIPq3ltl7AcyzYACjDUuf44eystmDU22b7bFSdoVb
6i/Iazxe63PMjbrN6tV6Sl5TLufV/bk5G/GnwQ/gNIkKoOlw/DO4Wdz7wPBrPwVd
hQPveDmvHeBh1y1MGyDBzG4uIHOjVWWyvFHjHgRjVwucShHcHvlcrlxXYrwl4ut3
Z1Wosv4MfY8Dngyu/8jTKcB2/ssf6FfWc03VW/ZN4FcO+dJeRhGTBrpP8WWDugyG
M0SBeCma12Fm7/NE6YCsiv+p63WSaJG2/4AxaKE7IFmkcdE/SX0h9V8wyik4ZexD
OUQg2fldGl9F5XUWl8m1xzRrAiL6a19es+SIYDj7kTtZcE3H+q7AZ+u38WEf30Ty
x2l40I/+CJ7MKlXyFsOpSiod55YOcFvB1R4agB3L7+2h2ZH1SDm10t7Kkiono6l6
xlXjCa6GkRHVplx7U7BtAEib0NpQgyhd9vgnH8dEKxQW/OjAQF5Twa5RfFR0sGui
TOV1ctHoJF93USbsDSHInkv/U8EXXzGFUKobKVPtjopogXT+5yeYxA1etnro5Vm0
D0xuaSPkG1LA2vA7ZRpkVI5FxJ4tyqiIHsi/26w/f6+mYalfJ8iUR3gfkSnPNjw1
MdtSTru7Yj3i1mbNIvR7o5SXgDWYAqu8Jg5nNK0qIOaItxiMToFoxMQ4I4XLsZVY
DuzwrIjQM5v1mijqI6a26ctQapIEBHoFd0AuRMhLIsINLtE6x48UHMJA4AKloRQu
qcckQnvGFLUfYl8EnWdvbG88WiKJY7aqY0moRqRAcKhoi6SJ6hqwKv37rAEqlPre
ODBGdCFPDw23BVHKbzUWvOLj6zY5OU2zkbi/MPSxvBvdHZDnenigFUpj0n9+Ge1x
9U89kR8f6znUiuKlHw0BIpDCBDquCI39l8qwB872RIf3tZ12OZyi0tzcMZ1P5BR5
H5Cbm81xwmQn+dVz3aYlFHfyMPYLdtckIaCHMA5YNJXIJqStIgqn7VBDUh0/sLtS
wptawTkgftlc7lYnmmD2QdKGop75n3rOkz5U7bPy4mxg1OkjhcmiXgWjEMAqTJXG
gAz52ngZ6lpZm/jddLLztWYb9EOkdFlxbjMZGR9asytFx/C0gzUY20u7Qp2/KMpr
pHfwf3nT7uk/MW3ySdS6yLQBHABUPobzSjlKf7eNj/zM9ou9Xvm+nZ8Kw0lvhJhm
jyTTtXOLfwwAPxPi9cbZx6HxVUJbFGyu+z8rglLZX52BDaWmM0dt7HYk/58ah9cj
0Q+pKQMLvsHb0/GLfbj2H0j/5nLcHEnWTzBboNZdjI6pn5IC7QHwCgWaT/CN/MNK
Xl7hqsLN5yZITTdTex4kd+Qt+kkGXkFvH3K9HVyqJKgWMlV4DQsDUrfJ5MEALznL
Zs87JJLvJ0ngReXXB4js04ih/yEXoj0hlacly5WX/hHWd2dZq8cl8YJ5Az0mgbMY
CBEGfmrjpeEhq7Ab6AN5Ay1IpERxFX4snymcQ3vCrA/KAHYDJFlZOTaqMVg4k9nm
GtEyg4ODpPWpXqLnjiDI/wAqqaurBjRZf28tQxuWqyGcvrpZMkvmJrWkr2PX+VOV
wgsjO3yDuG5u/JmcmRKJwwNPiH+7Yy/TAYj0LeKdtL31Rlh/ItNqhqVsD/2cirix
KVGJ1V8nITCYxRMpwze3/DcqEw6dOP+LSckycmhDihzD+blW/QgIdnxJlmmfw4mc
ALQJ3GPqYaX/HAOTRtybWVHmAi5vkLsf5l8JXDrhLRL3ueZ3lvAg0tHhcybaW/0a
U9Uz8d3oCNVOTnPmUUfuUXBOCn28KaRt9MynAQ/NyELB7AWaCchxKRIOXdmrUqKP
Iludwn++qt2XuqoOO/0N46NYmgiQhlcCCU5V3f8t+e2sBx9DTTsLpobe0reZg5IV
yxuU3UPQVb4g/XKmOAX2SvczN/p/wDHxcV0s8aHnFaZZnRudBz4ZqjBxwzlNUWfU
pR3afzrNPfiNOw1CGe8cbem/xcKJOKCz6vOFTfKrn4uwO0CmxsbStvCW1SompWIq
/8zHQ6oodQ/noMzq4EhvrhWIFSOVYIF74Qs8jP6IICNW7yvWu2G/v+oTIm9OVKql
hADAg8p1bD/+FIThrMk0cveGQnT3iUKpytMH98nja7We1fZp2lp+ygBKrs8c49CM
cDAo3w/cGZyKprMgty1o2SNnS4HEr9HhprgpwgFv94cx6G4DpdwWRQJm5ugg0wFj
zOWPME1WEJolfxIFdBJwGtzs0jIvQkNoMfk7S1i24Cls+HuNepCFQOZujXEQzphk
dUGsixIYZpA7/71Q1io56/kZNrMt3QTtpHmyDGF0fAH9JgsYZkM2gDpOMNzEtFOh
QdQaZek+8+tumgwfLtZBXBAM//B5LKMBrKF4NRk+xB+CBT5OZ8q/CeQRZhfp4f+6
FaNsI20x+R61J3OVVQVV5fHadgHr7kohxttjisTKha/mBqJ/zNXDiZp/dRkJmWeD
J68cJ/R+hxZTGRsRZdfcyBlukbZc9uhbG+NWU9eKIMOTtqVEK3tIyvNlHXUifQgv
8r/NNfHl6TSJRBgvRazrbVHNEFP8GrAMlDDWywm15p5rGQ8whwGnk7MvMMgBP830
VRMyZGkhF5WN9HDUBEhTt8XOHaKiCJw2dFtUKRY/L38p7IDlxp5pjN7ux4M7G+f2
2Lyk+ddCbfsxv6tqHYBalwvUKy8r7Ip99vQPBbE20CyvOhmASEQivoDAdQhKzZ2z
dgfoxCroekECp7IYhYzABHk/kDimm57mwHfX0aJ4CZcWeowKa/PZ58lu2wfFesG8
9fWC9lKghtE8mqb+hKzsSyDnKj9peZukMb6ZtxiiXTpBBlpnTLe5V2PpZnAV+/QR
24kfmzzHmbd8SHCM0xe/MAzx2WruFsZc4Ggs/QUEpdaPzpeM4Sb7GDiIg3vpURMa
/Nidzd/pUmlCNZ5A8DILTWDwayw47lyMerClVQMtXGpbusmHRmWo6BQJZR3Zfkmv
UOHd4gGW2ijNnCAl0Hst+XFztlHDCxtZJ4jFDyh8VnjvxIJqYz38FCT5rRsjW4Qa
/ENZ2DoLc5cIMoNMGgESU3I07NGwCrFMztUN0cYT5s1eanIEp013cmPdeHRMAzmq
2g/uGuwC6z6aGsrJjZwz9LqgC84zHVNTCl9emA7d1/m64twn60U25E9RPs1lUJPJ
9bj2QH3wdeG3kJrlv4RPOrzluHlThoBigYsFTvZGSn2tNNx61W+1YLp8M3QMjgIB
6PHh4uRrY34hLdmz9kdgEB8vvPSzlEj9WuW3amzDsZUSWmfg2dN225EHikyN+/II
l0kC9tKYsKsCG+ahaUG6LvpPEC8Gzkg+6SpDP4Bf4EW4wApKqRNBnGBBqJX4pkwT
P5V+FI81vZeneLnr9o6JcFBhyAT+5PPjsVU6m9R2SRgO+Q4v9+FwfolACKqaE9vZ
+E4QzHcREnZMevZsl7xrTXbwL07lHA4xnQ70LDU8kA2KUwTxnTGs3Hd9NZe9kLsB
t9M4pHRK1DtjXUjoWw2aBu/hy+uXuu1+f0Mt/jVpAzeY4KAmQmBtMNMu+yM5tNOx
340SShrwDGuMdW/l/wlE3DwIpFKfYPvzzgDEO+4MPWfkcMZ7oUkUm3oz7V9JZXYY
Q7DCk53txa7vgAPKqSBoezoNbyoBWHvjpr8O4ewa8IhJpQ/SznyTkChzlXSh3cAi
bmrv2oA5qOtGVfAtok705g9QpLhyUJas8XkyvDVZFfpFMUfviN3cOWRq87X5VRV2
1XxDUtDrgLkx8KZmdGNdkaA0Ni3sP9qkhkwP1dqDmRigIPQz3oyMDtg9fCn+lFVL
RlCQVK2/xN+V/ZIZW2XhggGtzurNTf2SRitmW2xV1Ssfgxpl8CxN/DCE3cXZ1FZL
crECVSsaXqHiPzlu8ewrrIUZ8r2iradWsBXGIcx4DpjC8Iw0Y8O8+usMOqPYnv3G
UZqM3lODjQn4r3lBNp8T2lIYnZGLoW28b90p0yR6Ifu6frnoCrNU8pvbWzNngUHa
e/1xn0lJ0XRVsa55Q4WMC7RvuxTPyTcmboa0JULUW0o4nESPjhucBdGz1WlWHbRl
MdXtgLLcKOd/0BV1g8miu5sYYu6ka1VU2oUGeBIgLhnKcUcm9wp8kTZ8Pk47hak1
vCtBgJXv9fs7AGXLja5VpR1PjOcwecMf6FXp+6PVUDRl4YpOyUUNAtSW2cT94jqH
x5lWaK+Xuph0qScqIdbVm6nwlkRmK81bJ8oCIH9d4cwMXbRr/i1Txx+HcWtGNXxZ
ThMHivg96JdfPQFLDAv/1vSjmDDTZ+bkoWOv2iOP14Dw82clRRw0vr0esdcw2QFX
bflxITTM3nR6AqGZR/tuSfesdSmktC9SSWzM4rbqpX9bP/OudLLHxP84uXnGnSow
wKZQKAkwG1OnmWpiMSTe/bVskowJJ4/wpKZ6THWOk+68zgItWWSrj9CRaEeZeuO1
EorxLAxYjKSInqsfSCAZJTk0sa1Gqj2K2dTXwx3MCzXFGyPemmUCpjlZCa+jJKTT
xXdYJkwbpcopzonpcIvHcSFjlELtOsMCl1nkPmej7hXdkTETpPc7O41OAFer0ydX
zTpsrskpuMNNTWLSR1yY/oHvYsu+/WLpki2LAFnglJQdehU5aT84UGuuS/nsGDWP
0uakA3LB23Ps0nOikSGaQYnaNhtKUFlwqN3Y+YVk2HncLVlofr80xokEVYhAVDNV
VbtO+3jTOnV/vFCsTDLJH2Axg8g3nR0Hd8nDjWgPj4rkZk6iHcsqYOOehJEgRp+X
EhSaOkqAVjK3+uEsDQKiBgxvWG5B1iQMArZbaaN6mhkel/1nkGop/MKm5PwYJiLq
qh2fkPrjrS6yxCdFqC6B5iFOP4NWQVOo6c6xeu5evLRRg1VyrEl7xElpnSt9cIUR
Wg18YBYOaCt1XttvLKvy4ACmK4BbVuAJuKGWHBASeYWY25+Hgv5FhT+XQ1YNU6io
JIfNdiTrhruERl/WrMoj3A+Csdykczw8u8zA05vzummioZi1Im1hfJnIo8ByEME+
8sx4Xvr78phnRGbkAlMMH0SEgFwV1UhuHId1TdZewDgBQXKFnzE4Obunu8dS7gpo
Nx1QvrkM80pvzt3lquyqjndfQ3HSJbfT5KbKOIfnlC3yqckOi+z6jRJkoxJg998l
no1ag7olF+qxLwbgcREYM7GqBRHbogrkhcDLXK4X/texSay36VxoXZEdCnYGrH/3
fziAQ4pINqygFQedFe5qOamJHW9s+eiX9JdKYOLK1N5MzrReDhS/VzpWoS4DQSPD
sezHlXBWu1/eN5xEo9gEq97QnDpvZbRz6Ybye0OM78keon7VDj1Ra5ilQ0pVi6de
I9Tzt8s0TaD0lkaLnTaI1B+2maFpqNmQDpmLS/TIsZ4jCBRBfT5BFfAaIpu64DVz
L2C49pkV9zJ+ex0PSF4ckzuVRCgYUZKAXD0p3OrFMZ/sOnoXdNRThSXHlDf+LupC
hXCzciuquQAYfZf/SrDEBhBzM+8dEKhbwux5oQwIUMw4Tx72APf6+6Ob8hell0Ur
DBOudHE+MvYJI5LrzPyE7F+z240DtYNN2AYS+IzYIqo5RnoviSSBz8k09tljkUQE
kq55B4rFieTPmh36Jryl9JGLPdPymwxRxaqymqHMNOsachLZPTgF4ZZtes+fQhjR
4SSQ9+X89dm+eeGJ28oY+R+v/MxoG+AhutRjgiD1s4LPqWNEdxRo4kcbe3Y7Tk0j
6KLEM8xm83ggIZ2ltQmXm6H1sJyxcGa9FbMlnRHvdlbWIAb4M2064CrgoXoG+gzc
gfr//t7Ogtjm7vwhZSoQlo5NT2P+u6RPg2pMPAdE6RFHJkEj0ak/Jlhpj2zuU6nr
og4gI6nL4irOZ0lYxw3KKgNv4jvinTwbmQfr7E10TxANbzAxkdCvS9vBxHlBgN8S
aMQFYLmTuhASmR/SpRsiYtCSZZeyxzppPUEzFLPI/0RpQ6sGnh27alp4xhKxBILv
AIpa4spjlrbbp3LIVRTtk19AXvgvzmZ48mVIR/tePjzJP5ei+rJUvpZG7H3thBgP
i/vD8AcKEObJFS9+lXvRWtU94SrpH2Hk73FGmW08XnCbbgo45UBPMjzturX1z2fa
CypDsoZt1ckn6nP8mLLHRQ/TpqaL6GqFqRN5B7P3VcEUsG2nXYJyUz+2mmEijN0z
/JmEGZEcSsZl7j7Rw+7u1/gSwGWo9GuQSJETUJJNigj7WEEHzFimgTdg8/vX/M4A
t9p5JnFQ8sEzwSGZ4X8wx2ibt6/2kMuJDNAF4hEOi7nekVGayCV/ee4plT9/fDAD
cTLdWITCkH0tSGKNdpTDeNKlwuTlxGmyNUqUQU4oGcleIX94nQl/5uQwOskaUe8u
bqVY+3RiKCo2LFOUbdHdkVHliD5iybsiwTYcNuloKqttDSFis5jD8l/aALk2dD7+
jkQ5oSuc6QM2sSBYsLRECw01Yl3BbDLxhqfdxVafPEj6ICp+AAQ7VM/A4rhQjjIy
P0Bq+JHx+ghxrOD4Xp8K2UN+Hd7rnyha8nU3CAnGrUNah+7PbY7vgIiOMXbDzWkc
nv1e6spFXDD6g40Uw9yD2p9V8O8P4nTGd+B3y5Z8RG96vXFagODOfvkqBh+O7e34
PzwT+nhT8hoa+MwMQUQhg09PdFnR+tpKNHydCEOTLPyu4+KZaFmOQjqUfkRefzF8
pytPXQH1blxm3HiilJ/oi3Gey/Ak6Dg97ujrgduX8de7eegtX1T6w2S9yt5iVJJo
1L928+3k/upA2zkJ2SzZNQrNm3onxxVv4X8H7U2lES8OhMzJCvTeuSTJV+DGvL6F
opP/TFYf6zbZH2qCDzLJSUj/BtSJqWt1IyU7A9etHQ/WEl7UnBOzPQBZ+Seq2XJJ
bmZCDA961T1DzVS7JtmV3XbvkNnCv5zSV/GHOxbRrsgd+31yQj0fNFKSVWSeYFri
ibg6tfAY0seTCKWYH/tUolxf4UMAft4KVk1K/W3aiGNIYwNpsP2F3kmjfgPgFH+5
DhKs16e5Fvy4ZdmKL9UqeEoKV8khTdHLVnn5EDU7XvoJna2feVZ34yOCjO5arguo
Llwle+ctkIJHS1b/jLm/wDj4wX6kZLjG0bAh4gh+7HzTcEv7xpScFV8VTen/KCsb
sGr4P9ELHuqJB1gTqIOrJjsgfkxuX4Pgl22WYCzv9Z9m5Y7eNXMaxYkGyagQ23Qb
W393dQtS/brXYi69FAskMOOKM8oEcrg5hxbSxJmLLclWp31beR8njYQQxOJF9MFM
GrCDd8I1d9dtGWAZMhxKbVJgmdO0yjG4YnUmn6FFUC4xK6NwmAOo3C7XaALlgeS6
XF8PCh5wPCs1um4419KKcS252d6hPZz2w3kFWrBHawOEYkMSWPMuZzfk9ZhkqJCP
SQRD2cTdHUbRxv2273jKT2vqYnUEafiP+1NpJ0ci4qBXW2Rj/H/gz657b/S7PnhI
N8ZIWDgJgwOry3fqBsLb7Lhro/DLfetMvDmzb/fn1WuXzRMSpMzZrN6MuIaHTn5M
ptpWkNTBRWSAvjgyj0d53eZU62J1SHn+46RNReyKji0/l3qB42bQe97tPwRJIXjm
4RVFAgYvy/hnoJTZssFx4Tytvol2tr03H5Nqlggnj8VJyb2TiycN5l3LN8SN8S7c
9hkNlwAUoyYYUmoFy6b0Ryry8BLHaKujtC6eFaaT7C2X1wpK+3vh/j1mKNyUOAmZ
BGhfDNsNTRdtxr3VStaOKiVu0+18RYvqB2URiwUrK37YHTiqSP7mMbUaM77pa+7I
T7Pyz64Fj4gLhe/SO7B99HSqUDW+30XSDyhVHh8M0krxYFN44yZXYKUe4YvrGgWH
otUp72NYzz+XEtpOgZrNDZdyOXAk6AW6BBu0i8fRstkFM+RZLMJnbASFGjg837ud
2449job2nVAks1GBVqd42IQ9gZnxsWL4Ne1Kk0yIUvkKSRJ2hcvQYrShmNl83OmA
C1Ffz434FgEpL2v81GqqjR9E3ikEXBaZZAs/R7DIej/45+b4RAeNvGrc2CEE8OVX
ao2EO8vTNSc+n2aYqTmy4u0mLPOooM16sFuV59+TtBylAmxxdBzzU9kRbdNBfM8P
NPzN8/guMpm0knhYAPOVN/laVeBvCJqboPYNhN7FxwnB3Scv3PKoCBTfHVXWyeQf
xvvGAfHQjtZUEogBEBZ9euEmwFk7LJVio51Wi5j+cQsenfgJ28/IaTT9i8K9qF66
haHPn9SH2831BrXKTtHHLCiZA6ZlCgAh2tuqGX/LYiK+izsWu6e/HJLJ2yCfdkML
oNbwWyXFQKwB2YyQtflMLYW3626uCfW2aTQFZLozfNtVjlp0tHxHsp1pOfEhvivM
k3APS4Gmi9YJu4xdXIYNwDeUf3vB/Dl65XHaZ8/465ePVBElQqqDWdpqvySGFdSQ
edR+tpSwjcGG/ljZvyv18WJv0EdjNoHY9zGFgmEUMs6p7BCsw6oAbJ6uBPu3B7ok
QKczNQVs4LbL/BRFFenczUpG/FFm6ePDGT+YOvDIAfdt6Wnk6T8KxfDZFQexAyoM
5k5KpHt1WitWlc4hont9WvSeqMfCsWMnoEcbmj1fwbvzwLiT3B8+0/oF+i6YDd0x
XytZ4FQ1tF98I+JT14+G7SKF4TlWp7gs9dOC665tCkXkmJ0QDVCQb9HRy5HXIscp
03jUuQB8dQSHdYrT9xqNUinjqKoCpdLBKm7+tSeE2mIbDTIbjhY54Gyc3OBpnbRk
unbSAacSzIcVgdsvIR/VPYq/MqPwY0rBScJM4tslb4XcNRTdbAskXMKixij0yB9v
AZ15rEaFkl7M4Fz2rjxwnUAS6jiXMjbaIqu2vnnakhRDjcfLhPpQZjXmZMLnPn7A
t7+WkijkKgPcbW0NzWKI5GJYkgPxgVev53Wh8gy6qZ8fYyW1ggiIeu7CtbdxPyOA
mrrl+KcsRa9x9Y4hMtJQQBcEiyQLh9gUYb4cpLgAekHjizs8qVWaOIMYo83ag5Ng
FNBa+Uyg86gQzzzBfPXtNLqyRYwh272d5OUoYhhdg3PzR2ba/xbskt/THyZSZ8aD
W1Oy8MVTVkPMB9FYvdvr8lK5y4s//IhAzHJPK8iKgDzSL0bggxAIx3xM4nvWJgR8
40mcZpq2RvcCwXfx0Wzut+mfJ3vrEA79TjGh/vUX/W+GMP/996DIjz/116ni2Tto
PE03XAwQaMjERoRdqdZMxa/fCgYRsieo8H4Z2h9vsJLU/3FQYumgomvawt9rFKrD
KISk4SbY1F3UxT3tdJDxoLYiG/Nc0w9jeoqW+ZWqlRbn9Fg2qcBPesZoVTDIRRtH
4vB9HL3AXBzzMsqszYWmlozvKIRhKYx5wuZWSy3v2EEQLvPJ0RJ+Ax+Qo7g4w9qy
7IEBrD/HU4n/EcxEn5FpZ6OBgeQ006JiQeGMzqH1H3P52t1cOKyhINWVju7etveh
8EEMLy+Q9zsiF+sDJnIKG9vVYtH6h5I2MwN2v0BnoDR60Hk7OJD9CAaKKsG40Cpv
iSqGl4xBEamX4j3XZZd4cagwP4+OZk4G0fpz9gZEjT2LJiFfcIzjhPk4JSmtm8Po
45gtmpq8bCOk3DqRcpheqNoDAzaykw8eEddHzrOBYZKRVhBkuqog5//nRd9ThlYR
vczRqdxouCPw61lMRrCnXAb93+NFuYRSVjetHMzkbaPnDpmAvcBnUM2rC0Rd8j5c
4MOU7QLJJ/7HAkMnucB7E6Oj2BukRzOt8KzzvYyM/3LjmTBAALG16xaXX51ZOEQZ
SumAsZwkOF+3FyWxMOVQ4rKnMIAfVOcaJdWz2/IK6R0BDCJJbFNPHgJKX1uCP1CQ
O7RrtfkzRHRffNd0FIZFkbYFYnDj2Cju1L9ohCTImQrIqoRKIK84bfykDtV4KPG2
4xFRhQzFJUoWtn4FOjEQtnjqdNlZpGD3QHRBgB2qr4COo9brrg3pztBN6JXTABZN
Juvwcp6zURTwn4OJXELWlFqF1sIL8nwVLcVMJpBlNh532nkszMAVxG7tkIE1Y19F
lLPcvyrtXCaXPjR8LAzBlMbQ5OH5KzrMQgVxuq79iw7h3WZZQF5N8rGXVTUq11vi
993THi5YUrHlD57vm9agpyOYPOFekAwuq11re4nbFfZtLf+D+jwawqzt/1rdgz8G
dcJ9HrXRDua0cC1dY1QUIWJa2PJsc+YCqPT5ofcc+pFLOSJTl638SQq/b0JXJyyi
THlsm7RpJ5p/6GzbvGIopW6H368PfS95CHKIpmIzYrXVI8nkst5krpVS8Blt5JhT
BkWGiMvq9sReoDUyyN/+3L6RTTE8BVa+DmW73yo6z+UXrYSqDKb3T+Wg5ftjXAIj
VQlRm4FZB2ocwjw2yc2XNJkTgYtPz0lHVIFTz1ngJRmfispIYgUQLn91f2sVvvB3
XGtPdpIElG28T1T0AXwGx0+sGLM4KKSpNrE2J5H5dg70vqnHT/jhHKKVPQY0jas/
aBitxk4q72ykC5qm6+VTnlLw2Uud1ShVhaLiUF2yEAaf3/aC/pk46rwoMdykk71M
w4QSsMh5mhAZUmibYA1V4/1ncrSd3LSXveWjYnFiW91FEroxIlDS4bCHP+jdsQX9
g+lzJLdBBQL5svkW29WoXdfGWmDnInQR3tKRq1GLdyOzUCreqlE/hewZKusEP5bK
l0NBImi0m+KCd0uyOiIPn3W1MGfWuhIznaTfmcl7XC/8r5CVmtwIArkVVzvo+VOg
/QuhhgEVul9EUvQpMlG7gnT6xEZqGUKOFcHqrYlVhADxhm68iShAXy3Oqb1bO+dB
8+0RlRsesIMppsIDAj4nEmYUmBsVogUXREYb//C7jbSp8Wsq8rix9dT5SMHh6hSs
/d+Cinf9hMy2u5AuDqysig4jeAHFytFwnXA4ODqu0abff9z75isQ2HCQUTyhoIIl
+z4BiwK2+UGQPgqpPCx3h7Y6kRDaexfUArFcJMNihywN2WU/fmqAjUgUYknSlzDC
BoraMcdBK1tWT84yQvTamFHtiPsthPyxWM0A6Kz2Y8eaRnlzPS829zzVXyi4zKaW
aUqDoj9WHXdlrjLD6g2XwcoECg/QH/+JzqgUnhxEtCXl8Xqh8pFE4+ZamDMWZE/n
Myq8AAv9ndz7J69PQjJ1ClNXniDJkmpd+5xjXhnkUOLehzuIWwVRdh2vGD3mysih
m3KV2R17FLZwZosUAMfMlfd5ofOARe1K2mupg9uNZmznKRA0JzjzUV3p7BeFfJ10
4YF5IRl3Im8veQI2MtIbIHQKodCLg41ALFwNTpNZGX9ruwQTU7LNJCgU0kIHuccN
zKgDKZNgips2RlnpnNmMk8ht8p+3yaL0Xw1JhJ6W6Ywx+JcO0+iKZb3k53muyYc6
emuYpiE8D5FvW9YPo3viuf08J/4LhBXzhjo8CxrzHmsuiXuAA7D43dBWfoiRFWxU
6bAtHmkTBCuSIgpNHmJ36WmmVO47HeLVJy9YN6L1Ds5tb3gio112zq8A5b/clDUh
y6V/zH8sxN4SMhzz6evjDbaFpczbeP/ITITuhUkhnbN/x6kGhqrtYY8lccVJNxn5
swUcawJX088zrYCz/QG61GIZh+Kc+hWqGlu0W/uyBeJ5Z7bGZPQdqu+Fcigq2Hj6
vreVYzMq6SYWesBmg0G2kcbKEsBBqAfbqK2gH6IAWKplfJpMzMuyUTm2JrO3kkUT
P8f17Mj/hVBgj5YNkvzXr5vWjvA1rc83fwxqTk/BmcVQRBkXit6whlFpf8Zrr4M4
r2tsYCLL3IA4j6qjxBxEJAsMC5XSMkAbkh+zs/WFq4fQ1QoxC3+ze2y1P7K4mGP1
NMRxB7oFGIn+puueOmPSA0T5IoKBtnY1KYMvWPDnFmUHn5XiSXZ8+j48AFhEQWUC
3rBaC5Vh/PYqd1NDl8X9Ha1HABCHgeFllHZHNcUK54/9msq2gsAqq1hoKzDtOV1b
xeqvcfTzEvC/G7/2ywTOm+/axjLrQwkLAwZ5jp931fBoj/XWuZlgiI4c5R7oSuIk
1CFacVLIAqCwKF/367CyE4y79zoJz5vxkKNwqyTePoC/e++nenHureEGgqsEfpjN
p3BxrT45Nun8CBfw5SdXikEI6KvQOn2JJWi6yejRJAYLG2mvCbRrOaSS6vlAZyZp
MMdpKWN3lp5YQ9dLhi5m92I+uW74LOanozUfXDlt4Z3mKpf6pNEv1D9fqWYRRGCN
qwhRpQytlgXF4n+uRa7MwwZI/SXCuQVmOG24L8vt98dJQk0/k3ovI69+HknONbp9
+yFM21OYkeWmDLVPuMm3NC+LWm6jufV64BzmR8ZugyQTpdOT/LWNOn7KW46bA+RG
LxOsa25BIr20a7NAqXdpxsMKMXs+iHG6GBCtE99efF2nPffaonkKB9JyHtHMcN+v
0bOYvjpUIMw8K9ZXsEGvnFuAtXi6hZWZkwrl0hRRr/TxVItC56InfOwVMNhAsCCS
nWkiy/wFvkQSKy0VJl+O2hxBcQf128en55xHwIx7Kg2NY0q709+s5rzV/7O1iN6E
oYby5kaVZWvJVj9SUv+rW5i4d+RauvRWl7pPR0M9dKFUOgbDdB0YdE9AYDPEPwZx
KUDCEhlmqPdgJCr+GWNS2eZKQqmIUE/26rFLZVFWUhZdfZAVft49fk6We60cMfhC
pXfZoih0VIdjuQfRVOgBFriaDgvRloSYxu2KBMVNop8kA06NWccYc4R5z8NV5GDA
0fZU5hYbM1Nr0MRJOou1aHV9NLekixfti78m4BTmyBN7ma8jdq5Q5Xd33Ocvz4XI
JaNZnqXZ7MNGsolVf/W3GYPZVkzkGw5w+2LEkqWffqPqFE+NJwKvUGB2qHIdaXJS
JHdw/E+Ae9//vTk2pJwQLTh/M3j2h/BP8XHCODqYVPfsJzVIi8Ai1bH+GsF6d8vZ
AqNQbyRetjhlNEcuCjxtkatSPKdrQAd4IwjKmhI+cxPk1Rr+liZDX6BQqInBnPqH
gsbmgIkiZduEnSMWB/+E2DiDLA46U3a8iT4BGk23DwTSJ3GgjiZHEBcYGqGI8pwr
UraTFU+KxXq7P1gEDdxq4AUjXqlnDR6TnC51shLXLoflgayBXMhE9KYZdqyAYOR4
qHm/Vsfz5R2fv1UajJiqIFufxI/s1Gbu1BnOvDqD1jYqmN2WnhKGiAu9eId4mm1Q
xJkWOCTZVhbkxjvjl/RgyoPIZ6vJPjNTjLhQc5RjmXS8f5sM3yW2BFvRWEKR5P2k
s+40wX4cQYUp5QyXoF3vagGs0Il7w47YgRyamYw9OQUJ2a3g9Nx994xi6DQ8W4Vj
5Q8R6CfRDubJNClkXq5is4ro86CHeH46TgDXG+y/AU2tix61rXxWpRzzHKtTDopo
q+QBJJZ935KcfMFKkf2bWxyix9jkZANT5C5EneG+ShL7OXsUk09J4WyJMSWygwp9
VYY7ntuQt8HD7sWFTZllJBOfAr7OZlkc8eGkztHK5xKTPZgypi0CSei1hUmcHS1i
M9MBKAg8oijvFmU8itQv5d52QKP0ixK22/QhIZqC5+st6UyXmtop3ROahtMd+rd8
zUXZZkPts1ndhfFL9iIFmCdfRymumbY3F2wiP87kwblDQeGpSh2JRxK0OjZeixcV
33xCzgTvzji2lKy5MHDi+pNeyN8+6S1BRK3uTRzzajp7EYUjOtlqkKQPw4TGQGzt
TofZ9mOhlcyF2FVwWNRzbGWkH68sezHziv7R3MneYP/oXFmmPDxDJ15cPS9nE9+J
0y6FYACx0ooO++97KP53kZvlYTjKV40MT12jmP7j91+u1cWd4EnXhunl8Bb/eF7f
t+gULUIZ3qS0x5PkSQOLAAO0yL5AiIdP03ePaSNEDMLy46/qfifRD9iNb0HVJG3f
OhG+fwNNDIH7wX1BmjpoD/aGR1i0htbnGYjd4hA7/+aNxXavD2pEpJ/BTAGNKDjw
ebnZBsUZYqlukIrD3BSMWrS6OIFVXPxFXWnLvsV9UHnuTzus9OuW6u4QAY/4/dLR
G3CwCXAStIyExHb8xxSlVM9mR3fhGIbuNEGhCSDbL4cb6+2iHFLaO7zfKA/LFNG9
iBIt86FIWXIBN0XhlaIwCTnmO7rIpzAnNrLU4b8oV6pRLntrmWcR2IrcUyEtlntz
I4XmUfmvz3BuBcfyzHzFo0rXDO5y/l7x7tiExuNddQbJdHZBufRbUZtv6os4AiT/
Bo/Mj/S1U/oyv7YFyo/T18zFmK761mENmO8k8m/gXEI+Rw3H5G/l9cixpfwuD9OQ
o7v7OZbXr/Z3yRs8YT/VPAomiyV6cOQFwnIbQUj/8ekRhJ0AhmaZ/ZOV7oZZNXFl
PrsrJqccna9SifyG6lBa3MxlVHPVegageDckkjxnUOCfEVpgTbuTWKBjSLMzEzJ4
voU+rDve8O9zj21cmkxaeeHSyS/tP+wI8VjxmaGzqKygR+UoJzpM/FHSwSvQlY01
XCi5QNUlgPbV8sDnb9wzVzUGB6gnEINkh8IelU1UXuOwDbpMmhoX2sF1niWoo6sJ
/RFm48Y/mEui8WniqdXt4HgE6mE1vSKpu5pe2QxuAfOc+UcLs3ZCioqyXF3cwzyl
J7XhbH4n3cr4UPa7N/Nnrc/FB33h0m8h9wmoESNShcPUWK4EVeDcXcDSr0KeWUKG
Yi0ITKd18lDNMzt8e5FtLxvu9viMYMSwCBU3ZXp9bt0Ym/BMTqTWbLJJk8zMylEm
b25xKcpEvunIWCCl93lA5ToRKywsLXAHZ5mxigskyTJXtZot++aVl19oZ923MUGD
jWBQMlyGjGsHNcHM6LW16+HacVdLrfKy7vVVyHNMrwQVGECYindbzpuFT0EXp47X
RthErTUyTw/QNJ4k0JuJtjkoVISge1g9B+48lPAwvEDRFo4kcfVdTd8WIOX2HVxF
HE2xqWEmnYHYuavqBHtqe9cq1ULKyfuUY1DfouiHHBlr+jgjG8xZGoz43VpiAsxw
/Newxi/4Cwgfq4A3q3oM36lZnJL45LZK7td9QH4fKkm71FshDcJe5JvEZ3hnnAIk
yY0+GFtvHWF+qnt57z0ZP2ybG0nCRsIXdnQLev9YwoOWaNw9BR3BBx9XLRYMDBRH
zcnwYp0glx1ibeJ2lNDgljeKGGgA9YnvTXe/0zyvaypUrGj+NOkZXSaezGA+TdQO
A+eV6Cwbgn6026YyG3pSnNd9aos+vEd27a6zcKJ9jHDKxPnkkBczD1CuDoGKNYv6
H59m2Ct7NXOpheHa9FrOItriyfLAdYaro9oO4icQ/TPJpY4kEITY5oyUlr5Xvf6f
WyqHWYRrwa+Oibvycix4BCM9oNWvd73Zkuv9qrpGLKN7wcRucxGcjtJZUorcEZsO
I60VjGSYwBZM1AmXJ6OKRLeipTnReMUsY9gg/tmqJUal54w7Lf8Fk9+oApIcQblB
pOpXrbg5UrJI/00bINuAJNKCBbrXOSGbsbhN4oBnZ1BS0FVyL1SXPZpxBYybAAFb
L/wwtTIUluNPw6FSZ0EaB5YUy90jq4fzk+OgJK1JtBwEFiaduvgHmYSdj9HCl3fl
334K/HVJFkMdw2sMZVCc8QvXFAeMNOrR0R4PTNXIOmghvPTCeXcyaEMsa+vGvRvW
WmJH68SRIfrk6JkWJRbxB908Dq+mfg1Hq0da5CHQUgg6unkTbWCY+Q6D6p4tX9k1
6+NnvoxUUGcl0wX7W3Wn0RkNcjND8Za3VqbxqJ8drzG4dSm1V5FQfeFnAeAYaxT8
WXaH3o24GTHyxbSsGknSN7S5cGbw2iWHaACxnE//PZUibpM8d14wJLmp0GL7h4ri
S7UE0GplxI1dmbMC8UwQr+P5UDukPs607RLxoCy2D+9OINkvhqP7tJphr51TAAlQ
dVuUxrj7VPaqMUU0YpqK4B4noy5pH14abboKsZPjsz/yOHrTnfGjXkQ/8ZQpvGWO
WpFc+o/HxxAegHi+43aubAjQiWGUN9d3nQl9MVlCD7Aho+lIQbtfMUy+qSBvVgzZ
/cDFej53c2HgKtc6QlLYzm6yElk2YflbyLenTzYf775go88Fs4a036xYOnhdJYQH
ZsDyNdXrC6cJDDU/nRE4Kkd158lzs13NlYoDHhAJoVKGAGd7ow800+PMmoyvDTrn
7rUFKVqDgekhbs1phnlDXHYbl4W7N96PmKaujKpdGEG7iPbf3KEaD6ym3NrB2eoi
yuHPgkrKp4ru8hg3Bhj7nn34/ot7XEaRCPcQAlrwaLdATqHw0+iVGPF/7zH42JGW
x+Mec3g1URX3qXSpGqAFYGdRhpFnkEcCU8nnnf2mhn6HzCzN9lEzZVWi2dCFrXsh
wi2bLTcT4Ca0yvaNqxFznKwspJAgW0l0GvrDABdUQS9PsJ5WbmFnSe96mt6M5OxB
i4pToFmT0rRlWPHy5GUQz1jqRRXuODXQt5hKNOHmyYUmt9GkW6hwTfYcroJ+6Kmv
LUhosHj/WfhJuX7eqprcW6EBQ6rwZouhD6h8vKkSeKtCOpnMEFxcKgODbxS2tsk2
qdbnvTvnyNqFSY4e6GJuRtWyruIOMGdBZo/YrYENFHbobLl5LMavjjlT81Eo61FP
hSg8CtzL8fgegd+rWK7AtuhWjeU1lMs6PTssgAyi4EFPmVC2QLO5cwH4hH2dJmoo
K4lhDt2L/Ntb1vgCSNt726/MK5lYSOGBntQvD/Hx5p3BHS227TeO/qbXXUFTIO/b
10/JPoARujD9j1UHJ3cI092kkU8UX+rkdNgeAqSjWDKHC0D5f7zWApQ8lPvCBh9w
VYtJPcfJZcql2+d8PDkj3ntDa6PYH+TY9tFjzJDz6wqKtyI5kNcXG0fldUTxvlel
R0HuTPgDukGbVrQVUwXgG1rL3dNDo/4hba4XRg/1EOL6g+hfindm0fovjZGCjO5c
RGlNmO5NReow/CH9tp1HtFiGoSwaqyNGEJnDN8mIpQyjXmTIBuYGfJ44gG0q9Htx
ZkmTUzU6zOdB/QPvkaHkzgy9hdHt7mi3UrJOKDIyHP9JMjp4LugLgiJW8P/0V6TX
L6VzsN+Gn9y+VNoiXh27JghvnMRDvMra3yE6/p+FOAyYle7pySK+T0FuwkS2yYtL
AppbIBCw1ZlKBsSuzxyvco690LeNoXsMp2aGWH769UfQLy956WWOlT3+moaA9ZBS
ei94K97wNwPthiZMjkkzm4BV1/p5zc319g4zUQ4VwQtSwLj5jDWZYueA9tb3h8q0
qubvPlHkJNYdKdAQXOso0WoHrQFVMEmbH96CZIX9a2Hr6urcvyquXPRwXvLU5Aai
8SZ3Yi2FrApspEYKRz5KRugh3xpVg6QXHNSEZ3X/gnzqUkKltZrxC0Wy7z+qic8a
E7zs7tMYps0FEFlwjC+icKYB+FDX/pY9EdRfkR6EaXnzVIcokEy4pr2IqioCows1
tbleaC1WYjs03zlleI+4BAq6Hnz/mOQyRpOXnMASc1U3iX58wb7m9JY5ju3tTSb6
Kt9+abUoJzZ5/Wc/cBSzgLSeZqUbu1wjbFW79nVRkDSwB0cSkT3qHvWt2AmBKzsM
ESqgPQHqKruo2Ph8hyLHCguQHX45A02HwHv7nirKCK8Lff9QLfv2lQ+HhvM/sVtu
ri2W4GrQEg3rLoE7n/Zr5zFNcd2HVjFOSjfNc8nqHoPr6Zju3ut55UeyoE2c2vS7
tIe05Pd6V2cwX6lmO61PKaQyNwvMxMwAjlAEvmEkJAGy3SuvyqoFCQqVC7iBhq9E
OFVBarkf+uonoopt4IiEXEsAKWHD81CkuDGyQZPLRTf01xxHzSppQFYrY31ToTNn
DWpg9ZJuSvUE+i5YPr64PjB8XqwtgAMm4qnlGQ5idyYNDB3l/jILs5uNULZeT8Ht
JR0gArr3hbtf9zR/CNzLZsFMcdc8i8o8of4r9OwJDAeuWQf3EduwK7lWRzrRgY7e
XjSzoylE5Yhg2L4eejM2ad/wHX1eOQM4h+l9eS3W/RgRvEvicl5lJQJDTMXMU1Bg
DgJQXRQD3qL+2efq/hkxkqqcnOhcos3fVyiG7IGG3b/E7HIDwjhan+bmB8l2i6Uv
WKbfP4geYoFKsctOOK43yEy+sZnuAnLVHpP5kyedkEr1yisNBRtYN/cPmv6IAuND
Lg7CQsC210WFrvTQ5w+htFY7m9zoblXiY0cxq5WH3zmFhz2XSu/pefaIVlo+d6Kf
YDtQZ8BLjviqMqCEGRxF512Vn3u1oRzqxt+LcaNBPd4Nh+aqpyqEQmvvAElDD1nw
6EajqFT3Owoux16/gq1dZhNl4So31ebao6YdUIAVC+j8mcBQw9Vv8vW3IK+IiJhL
aEpiTBU0SUFLCdDrKhwzrxENA1ApfuV+at8avwDnhJgH+MeaLnd0dlfuWG/2gZ/C
JK7vJnqBu1Z0OFCbDGBWcs5UC9fXrf2b4loHaKTczg9GYXsmdcxYfDKW5SDfsozK
QoilMCAC/n/8/kFWXC06YcZQdlsNoqW6nFPqDjFHLgxHwn1Sj4aOYQnm7abWG+yV
U0caAm9j+TJykX3PMPyTLOrGWnO8EvsV4VjTBe6Rt+O3TFC5S6P8SoyQyLEQ58VZ
MC5xawMZNwpkC69LRj0WOFBnSm82+G/qcOig7KtuWIoRmFdza5zGh74bM/KJVvfU
rSGQousLfo1DjQW/6t8fLWYSipNyvhAilQLvgnEUZEYAMmeuT0F8I9pusVXtc6/g
nXJpOCteu8mIeO9v7x0rnyq+Jp6aLeoP8CizfMeM2mNiABOs+v85arOqImsEfFrT
BYnTJFzPt9gZ7AnlkZjpZzI/6mfehw9FrEoJdCqZHGpij7tmknprYU4jW5aH0Q8Z
Ws+yBgIUJ/equQh64ZCSeYgG0ww2rI6GnDIVQaOB4rxLvJ5+mQ+Tzvj2vot40l/x
l60BagMoD+te/VYcUWbca9Ix59R2eX8BU+A0Hz9th9plCfZFKCoffMlHFOHY8SJW
mx88ILsYJJ0j49r45MalZ4tFyNtIsVpQnICRV8Ibzgm4YvkxMQ7Nknp+HSRqe4mV
a1+5QgQ5J5VRoOyZMWn4EJkl9RcxGfM0b7RfcGIQUApFbDNjT8AEMdVh/6x1dwWT
pH1ZEVs/sZCC2Yn7UAc/zov5Am4w6Gztx/wqDR4Ta7tN7LNxLeg+HEbmkC7zydTq
5m/9NW01zXy4+HxcCqdj9enYQ/5dkH2vGxFMetvrd/JDI6PakkzYKIaHH4unf02l
VhYMls7QVn8JNHWs7SjsFbu1lbel+swTmJrawWGJ94taTkhbQRpGbU7B30hPWQMF
lGwbjeRIn2h2jA5/sclz28w3F/mJgCHNdUSZBQ2RJ/Q2/pRgZabH/mBq57vaAp5U
oos/yhoqcpcDprmQG4SgJE7nQ9vfciSyHNco9ZSdVYbpjoiw1Z43guYWBFcYugM5
18eXVVDSDteSU01fG7pDbJITEPrSSM8yY1UlducVQEU/yYoYChTXpPAuHYYDsyIy
DqCdUEnQF6trLqe1JlX7CzNGLKGJYQHjKMCLaMIyyc0UusWePouKHtD02mRrwB4V
sQMfbgJ1rFzmQa/PYNJzeZwAIasThIT8vVjkkMoVVvjAiU9w3h64LmC2QeRw5LzV
NLl/fFoMMnJwTPZJJrMJIYSDS17PpTXpjN+6mwzaznGQUAP61Hula/kOT8ajv4wz
vq3PmBQ49WsDUi5Dog5fckdv1aGrSqm0uBG15Vcsrpno3nrQ9O3CcNQlsR1eLvVn
iOnSq84DGwqSQqDxLzBBA494sH4bPHzfqyPW1zRHUomp8Jd3utikvvsd9LLdlvS8
iryILKkT3HY/T886b8MWBB9ADiWs1qRr2x5I1KCTax1uNA+UygoM++v/H26ePvij
cxwu/3CN9qm1huD4+H1p+JfdM8vWsLTWj3wqZX5IidhP3UWOITUbbjxSv45HVLgB
VNClvBoHNjHPpvTHWa0VUGsaR2AzUGQ6uQW0MVPO1Y/5+IDG2Y9StK6HszLSOb+Z
IxNZgps2gBVW4EKDiPSQHZeRGxd/s5naVHlH2j9U5SDvRG8gwcUCiWiBzpLgjOfE
3cMy6p0K+tQD8InotopxI1a+8mju1togReJpAvter0nLilxBP7NPYUI8/Ir0ZPXJ
vMUEIpqq8P8hhtueX+mDEt/SoloEZt9YjQ0Y51JcAw9vg4L5cFSotMOsr8O9uRUS
D/LPvNzslZ+v6iw3yd9q6amk6Di05MXCZFq6Dgo5bG/+HbU/CZYlTeJ8Mv4wZoPt
mgplEaFwtCLrdvNglCnQBoU6Ixi5XieldR/KnUyRnTaJZlQXKdSK34WIb5sr/ZvV
sdyr0S5ILZHwfrLqZp3M0gXitDjmfxv0vQAS0bruETi5RqVt4pdaF+mZLQl34IOt
2NxeH8eLEU3+ulWDrJaAah436kyF5IBE4TQvhXwIOQMupresr+rDjwgPj4Ld1ggv
tukr1a9sTMLBCIt3/3qB9ssVIPGz5xIBfa6581uOHWTQTroE7t/0v4KnpkQK2d42
NvsGv+1XiojlkEDvvdWBL7xJa0rEUm5y+OJUIoZiZmVnyqNjKi6V1fy1nGJD9/ta
ft5R2kRHbABM4O1D1LPgJwRtUUnOdCpDU94iI5ewvdgudAWf0v2vjGdoXUFrMTAj
fldAtTZu3heVFtyyn83xV4TY3mk+i7u+HDhCgJ6TrOuSwvIumLHIP74SZmcx9uCR
W0dSQfYjQOSs/GqXvG/E10Abm2ZBgK8iPiscjZcSLR3rg4qeL0VrNi9oehQHbvSE
jCHu8Wt2TGo/cZ1VWS0D9HSmYLwfSR3nXpnyv/xQut4Jz4WG3zTPCkKeyfo8X4Lr
89wCyCvhPDTDB4Sq6pC9zn5kd5aXa8WtrkZVq2e/kdUWxgZWzVsuGrXMmv0GJQKm
YTT9Po2qBa+wsyRsCYJDm2vFMz4nzThWU7QPqRAO5wwpThCG4fTJj/4oJSrjETvP
BHpE+ZXpF57hb7JFdES7nn4x/Hi1gQchCEjTRg+dvxFVgCsEBMI2uJpPMS9gppJ8
YccuhxyZHIkDBb3m/0+iy7K6Mze03PX0dqKDBv4a8wPfBGmMpCHb4I5dKwx46h8U
RaUgB+9jQGIQ6RtQJ/Z3m780YrqK7DiIw4LWn8dCkqFlzm78di3dM05TRb6IWDTa
RWz3I01bvERXtG1sdt8momO5b7345w37gVk5kCaIb4Dn6ntRGGKTuOAraBhh5C3t
tYtZ80CF95ORsqQebgYK4kEVRsHMSzEoV87E3Oa53XAGzCHdV3MPGfmjtYKUYYw8
IqcAOOtMSH4VTRat6/poGFCgU+qHFZ0ykmcqqPoXrjk6XvtDEicGlc/p+bs22oOo
CoNmkBRStiHQJ1B+5O0CASVuCqQ4o9QrKtjMnJlvDhbJ9+AXrMnjdC7Sik0CEF+/
qkUzzcsQObCLQ6GGxrPdu/HbNDwE4515tY7WEuIFnSh9VTl/U936zOM+4puvjX0Z
FwzHpHKeM+ahlxQAkqajLrh3sau7CyMIdVuV6cIv7grkZvgt7WWL+vyCjeiyP16b
7igyb8FGq0wzbzKGvAlyMrTh2lTLB8cMWtL1KpNwuzm+xjGb2xUjWRieMTgJouvQ
tQO04GGwi42bae4ZWvL1chYPnNWsQDBk2EzoIq1AUwA2LDlsBWbV4jOWWYj9H1sV
kNwr1M075nen7z8vV8tO4PWTzN880dLTH5ejwJQ+vFcaykJKYBVIxVBB24v9TVHQ
Q0v7Z6HYqcxyiqFAv5JhuaU1msyG00sblkwYRFXLnpiw9qo+DZ+lfULxjPmACT9K
Avh0qVRzQklXiPDQ72Bk/8ZCBJHy9nsI0MSPS8w8wI8OGYcIAU9C1dB9PtjMYHN4
lbp4seHeVrlwrLFPyL6ad/9WjDhbeHes7wZDb3JQcdnoi33uvK509kVuZYZiaKcG
Ia0GqiQ7m5hwVKyRzdlNCvUH3mKGowFtOKlPgGNDU7s7c5CjSB3H8TbSE9IxBtrF
Qhzs534xpVX9BSZaimCovUqx4TPTCbabquYrpUw1yGJKyU6YA/B+5plqPqh3YPLC
U1VkqsySlQWgT4vkn2oONjJ1UE2qliCPQscgrNOSg13Yy3h4nvWq0vqh3wvLgNye
EPrZSUDxC9jpyN03aqzNE69F4hjAtmvoP+WaDRl9E/C9nrmWrnxFfG553B2H7cDu
WvaaE7PwjZ1eqe7N5MxQk4rJRVEWqv67Tg1nMXq7nBmzi9pIbvYYpksX0PzRUjFK
Ndqlr1hr9B8NF8LODLD9BbwWpJzxLOD7L0woS9YRYzP3GBVHApBcJ1sRxR8MZmRj
CtrTuGSQkZS0iHlOBlNQpX7pSAeuk9XUgDeqH14zovCl2vTMlEtyCQtKYBP+CsGm
NTqJry/dMC1vjK92BUGw7pUZHs5IDIfDB+hwgOvXda2Sgl1VQhkPoSSXL7rEbMaF
tPlx9Yc4apVSKDXKiu7GJsMOyqeVUAPo/JEFBMn0+7rJ7ELjR0pOTAy4GPJpFQnY
dUzsgSnsEbkjf7SSzV0uUlDxwzem+jfXCZA1q+fWQNxWAosem/CDkNoX3So7qqw8
NFOjG7KhDRVnCbhHbFuHi1UINdGisk/IQMey7+Fqhk6gctCgKB0cWO18I2T+onYf
MNh04Z38H7oLFwVvSNLyVfDG1Jggu6uHzLexVwptfhlW3uBcmGe3ckv2+3wvaozb
Xadj98LYjHlcVK3EsiiCemT5vZILFiBGcMzkDXTK/Dk13TOnL/uv+8TLSBUBXbla
aWOxBkm/5D6iJac/nVA8JePFKyVFgtRdc1Z2g7UMRgT1016SMLFGnQclNPKP3vFe
r5Xy6jWMhiVlJw0Ydw5c4UDvy3NqKTMcAELLPGxPq854IvryNGl9NVgU4BF86n2K
0HP5onf3uv/3L7na6tH2DOCIHxQkTWKQzdwVy8hAnYu0x4A8Lqh9SgaUhSkV2r3Y
oJfVLAliK/x0qpF3yFbm7EmDGUSsFOEc9Dly2SwmV+COApGh2EABt9lu9dUO0QAB
aPF4QHb1C5gWzgz8nWFRv3qXxVi1DKY2uxZbU9yI3+MXSBdw/5A1gunjEytMhD1v
1+X6dD84ilVNnzlEjcsoJmhwH3dkZAXj5a001elAnz4Mcz1HEJ62aWMDC/8X8Vi9
2JQdEn6u0NL1/QbGv210mQ6rtrTKWYkVpOtafQZr8TuxQK8Fdj6SI78bJgNLD/zA
t98U3JMsKGprd7pYQseBPkIX5sIdlBgz4zbAN8ZhZ4p7hArxpplosvIc+S1Mzl3w
5IsVKldgk1DQ1J7ccsNBIeQ9ltygjnwT2IpEGc8G6ZloEXZ92axPsEHj0APThV1u
lDMhLlFvJPh+j/A3G9zNY4o3DxGKc7thghmbsSBozu9Nahcgz+yssLQP8bcLjdsy
V9acU3UdO8/Fa1cMLlEDqYNWK1GBTB4qWjg1oETajFvpR+RODCvlFsZbRVwF1XfQ
NImWs6eCBVCMxkmNm7z5NOGs8x746eC6bKoUFjoTXLouyxG7XZHG5ZJaTpJXKdo3
HtW5LtuoTBGS+AVeit3veEvDrdhCpxdFInCkuiNFXzO1HeLz/OaLPUE6o3ZFnIn6
FnDpJa4lmA46baeu1yMYMxY80ebV+S7UePYMhEWSQwU5QOJb8A/35WxZwbNPC389
lrvFNNtQ/b6ONHD+fyvzP3mkcwK85pwA8vH5CRhQsIagUTQAgoxrWqmtlbX/QzoJ
JGrrVsNnfknuvG+Gvea4+0cZt7wP+N/vrkof3+HlGcwEArOA0aPUs7hhdiGWKgr2
wJDzPhS3AHtZCKenynN6I6LmwgQGa9EsKh4IrZ1DIKXcLhkrv6zO57y+SWAQ9FML
WTypxR6tHO9d9JbpX/x7rBe5bZaLIhb34cLPJoupaglk5T3FhWaZlCLIghuIFnau
+g4tBTUsxX0W2E/jJ5exsbzay6cvBkGg3oCJRbolqqeUzs6sxjGnKjPfgjAP8YlU
OinjcgJiRwV9gHsEsVbgd0Y0AaldQL+hkwSxsppsOdmcnnW55fMNNlhSmJ6vuIQl
KIx2sIJhByrnC5L4BCHU6XJyPAum+za6zVuPEI7ydxmQSCOx2OZ1FWb4XVi5/GBO
KiK4R4XNht/NO/VO+iVDaZSZFi4xXoV0Sy7VPmFj+O4Pn4XUcQ+mU8wHwkK9cc2R
JpKUlsrhA9wBQy3b2qBiBCdbN76sb4f8V6pYbWgsrNYXdhZCd0VqvxpaiMi/7Snh
SJQdP3VqWSSpeFi3FPy8atxUJex138+OIDQLHeEbPpA6Zz6asIGNAsv7PzEN1cL9
sPJrvACy+UMAUYBUK9Jctn2fPHsetYGU9nsqsTvjNiAjg5D/MrKXllgVs8ZZ/n7P
s3QSjg8pRjpLyI+8TgU9ywjkEqIO+wIKsSrCCerdr4qnt4M4Z86hBBoT8XfihxXx
6INRepGKQbpbuUrgH4SuKpbmh17ClWwKqbtcOKPyw+kGNeG2dK0u7/457mdeVW9S
+ZiE8FfIuQtScFqonlrrqRTAymb2/GjPpHHG820HGowgS1enT0KwQwxE6d/UVncm
GrPBbG/dtaVBOce4GoDPXmbs6agbbAXY9Gk4cSk8y8jOMvtkAG5obpZ2eLuTqLDi
cc+1dOTOcbKQ9AbH3dAz+IGZimPNoo+WCgxk6BnkRmHqKDbxiX8bl5SmoPIeZXwU
GXJB5jMQRR4wFQl11nexutRWhqbd1LVAf5fFKMa43HcRyZ3TlCDgwG6a73ttJyD1
i0En/QZeXG9AYHKxy+XtQzvBcQsamw4WrvH6Go26MycQeBtpmGlA+4wBcRYbYRYU
axv//lLEhoHHb5nB/kEcsyA1uZxibruiObdLepwMxKpHE5p+Qu9KYS3cnKd7iRYT
+n6QsEhd2sTY11RwKavoxmjwvVrOWxqkYbEdfBAsIzLoeBQ3nuMRzzLzzfeU73n0
96Kd1hHNkj3hrY0RIAjh2EE6K6Hbhar603jdAhQDOPxO9nk/h4yrvSTXWtQWg5VS
ufrZaaeqG6Nsh6tVxNJ7ML3qhde/3tHwWugAikRwUsDWzHIGP65ZaPISVzvkhohH
q74xF3CRqoPQC8/xUDldwWLhSx3JiNlqPnAl0wKrXm92x7BYPE4jdeZgCUSn3peW
w8eq59JjVU6y3nj2Lw46HPNN3Vn89UMS5g17Y0ziGUDJMitSh6Q4m/Op+4KLHKcU
6Btl4v1My52Hyeh38r9yUpp/e9qWp9SlfB6rBlMBah7lil6iUBlR5jEwxdfNoz5a
Vf5dInUKBwbtAia0QsLB9WrAeiqEYNnPcjpYAYYo0iCNFYvFGKh+ZRzGK3A2ixyr
KcnOZgq3VPUpeWqjjpxTHV9Atzx9mEz/eIO2frSt/zX3/uc1mdlQyGxjseWTYSgX
1DDHcUrurQXPF2bMXWp/R0LCe6Mu0RhzVO/Zy4vJWqW1dTsEY0ioj8QzQvx9r1AN
sfYGQp5m9px2x5kPsemT2uz+hu+LiEgINMH1nkg+XcfRhuUagp14DxwBm5XGie1N
dWXuli1IiBWFl2hOPj5m1tRBD3CWtol7qGxW8aY/QyHg4vTVpGZe5dyFCzMG42kY
TKYr0WZh5ihp2aMW0hpTHx6cuTgxksfBoYJSGHFXCLYS+bDY18VkYXzAqpIKUrlx
G70/EPt55L2hLqH8e7Ed8BMd4XNWpKq4ivHEavBs33LiHCY2uaR2Uit/I7y7DnPY
B3m1Z3n8EiNSi+HBB5O9NsDEyM+VzQbnzf4hTGlRxO1OIaIxBy7OnirP6hlVBwV2
z6l9DNG4wGTTgqgf+fK2/n33JEzJ4kumbYM/B773E34k4AbxnNNcuA2QfW0oZtFh
1umiUaH5ErI5ao/6urBXapwQ8lY67evSsmNfMARfve67n+9jegf5m2y1NynS4bmV
1fbwiSDfQSqbsxKBWtPoI41928Hj3k/MNJOYA6WZ83GMO/s6AyqdsTLPmV1JZj0H
wG/yEyeUbHl2+04D9PzAej4Znmj5bSUnatf+t8aNrVhYDW9Ex3ckKeEETXOWPr1H
3HCIH32g76uFCyHYNAJ7uf75VF3/R+Obx456qGe7vpFHXSF0YGbyyUpJxS5fAEnD
HTmjnVj5v32JyrpSj5BTbmVfpwXp5PY/4sSnDkZMMRis8kaxgoVPYpq7fP68HHZ7
nPytcnVqnNk0kMk4tMVo7eXMqBTAkeG8UACiZygmDD61r3bTRAjtUWnILlV5szOm
vabQ1WjeC74foCyvzpFvivu6TshwtfTVJ7vRNqIbwCWMUVznDAIwGbI669cSPcyH
+dNSMBmoW6PE/wAoitoCcQ6JaM0zEwJqv+0wvksGQb7GVB9mMPsQmDFyswHt+tZU
EIvhc+Zw58LbCrbpl1odrGqhRBIiFuEcnJczGPIytjZe7OR4JmEak3gGSKux4DTe
29CihElLWSo4jOUMFTO7c/uG0tmvmuItZwNBERm2c7vQs7fiOOmj+rKoTNIdy5u+
N7MtzAMgsceQJtOpMff7Ro3dGJmei9RScpm+GgpsO2cXIf2HGZ3sh89/46FEuJ4o
zUvdOI6tGnAY4ywMXkoSWLPtZ8y7zWJwla3XeWlcePXwgSliVq3fq5btkSwtVVvC
eha0O8QGLUIUtVdotttfvsBtq7vZGZI8xK4FdwiCUTT4kEoylCM39lq7qz2Y5XD6
xKCxlH/GqXRNAvMQy/gnGuBBFjz2PS916bh1kB1oNTA0VxwOz9c5YenY+pBVdT6h
GVPU4xeaUQZfRz3jTlPYRh2EPw5skY+CSizJS0VIunXS186cKpwpnkMh4OpJH7zf
bhEQaRf2/XXRY/wuwx/UDBaQEbK9AYYH9vY6CsdsUYPQGx0C63jJGSTmKiIj3to1
B3fWZrYMSa+jTNCnBoec1TvqTXOU0ZFdqeu/P41yX13ZUe6FU2TOS1eu0Wiz9ZHv
0DhP82gAbLpbDXutBufp6BFh4pJTKfwgjxrC/iuuTLgRfTG8OWOjJ3jYuRknjNdN
IrQLNFQr8fp8r+QEYEpVfbcn12ut1cHSQV93Fd6pg7ZnTLHgALjOdHOi6Rq9Ra5V
zxyKWzZuMR4g7u2afIWKxwgpVmGBEVz9o2w8+r7SG7YEf/VNRqhp4HkDiL+dxN+y
7GiDfctI8nGEQbpc6IQP5hf4mD+OkpZGhVnBhLpmTL+Q0d7R/r2DVWBomQscDMKz
NPzXJe+Z3T3DdWQ6pBBOo3tZPUHCgREv6rmhzQ2N5WZAmkGIVX9qO1oLyS3QU5zP
gwzRFN7Lcg61jGwqzluMpT2roqyxvd04wtooxPTJ8p2ovZx1LevD2Lxz/nzdN8OI
3lqlIyc/oCuv12DsDe+/R8n3a0j/TVRxhhAnKAOaIpxxDpnRYwH43rDA/2EVuAj4
zxSgIRkB4VTuuabfwGLKdcGsbitJRplUbGzn3YDA9OxBEbjJAyrXQAzpxRsjfVpu
O8p1TMv+P+l1BYH8sTxOkAGgy73SO1i16ytXiJuEbnhGrQGwSxMf/Xt0FjV/WtoA
T6jNBdBEIDDSgr4JDcm3SCOnGvlOLiMABP8JTXm3GyAKEu5YNFkdr8TFOcIszt9W
4SaeBAh1GvrT/Rv5OTsLR7HrE8iAnqpMnZxdTwFFwvRmt4n7CyrELONnMVYUlk+k
NUnw8tR1Y24G0/cJXYo2hMOjzjkCSGFBL5Z7chR5U1zz64M+XMhUJ4PNHm2DASaw
VSzALoMoWZdGJXO86+6+9k2t8m1zoPbB2B2dv4maJo+fRWCwB/+lbf1fydZXRxqd
9R5NAEdTbuyVBoxVypN2Fb1xOQ6GH4BdAXsDCW5mTVygp8Nm5K73T7SKaxA8038U
xEDZMWuWFmvdR4o5VJYptj7WXJ9hiNaJjxu1/beL6hsL5Cm5UbjU+/Q11ZW4A3tF
VJ/x7tQlhj3xtMO/Ml1NrVfgKzdheSGHvMZG1pQg0yrU40MfwQzaIOlPfva69yg9
FahgGYlitLRUsux+cOtsF2ZPDJct69ah8INlUevIAKm3vyoA7gdbJl/vQb5plRmr
by8N1FxqcdPyGvG478E7FgxYQV6cK25Y/jKXUc/RosVLgZVBCyVtS5iVXkC80led
32Zuv4WBqoFHQlU8cbccdJGJXjU1LKFVEI/7tKBScOWLovqt+vapUB9s4JJTmBZg
uVNHpc8ELSYsC//xgXjfhiAOs0NMGOzKTEujTwkw2Qtriw7M9TwKrANx+xlv9so9
PxfmPBrEE/GmEAWZ+IpvHBM8bdqoJgNOG2pGy1mIjeQOQ5XoxIbm2vm3X6WSLk8a
Bu/k3fBxjrfvrXyuAre/uTSCrRRG2+vUO5zo/QCwN2xsLP4NVOsBfpFRe1+YIDbI
VJ3jkT0+59qVxUQe/lbppqM92Z9I36jeAHOnUp2HpadWq2hH89PKK8QKttblDT6P
+Zb6vWT8qrf3gtzx6Fu9JFiu4NHq4e9wVqprp8LPF1Y4cvhW5dXKeKzVfuWgOPvk
WkTXWUooK1agoAz2EGcNgTruQChNYvXKbOooZbAaEhTL7y2SrhUirmO+yd09y3i7
Ku0csyO+OZzxz5HIfx9x2fkHk6ef/6vt9iB1UaPdCJo5fwvyifuLKqLFq5GvT45R
dOX97qCj55GhPDhS7K/jq9bOLJNEcDB8G7N5TJnS+kp3Qmzh4Hn8Ule+ncyU1qXT
0hpCVPs20hjR0SesWB3twX21hQS8dl8bDTtw7g30826Y9bWruu3/UiJyxdrlU4Rz
T+yGIP/rjspo3KPMcQUukUGeGoM51bQMoeZUe1wHzJ6WYuDDythWTBxHD2IGvTnB
58FPAWzq6M1JPO2i9O1avH0YXoHkIBv8/hs7ipTbulrbRTKQTKC6UVFqyOxjpnqo
TKyduKJL2nUGAhQTClbFI6t0WvEzly+vp/9bXoZ/fyF+6SczW28vFf1mXv+a4D+z
B/a6mflZxZ+rN+rcChyxElpcuVLPqnQOKUQIJthRQvSNg8h3s6dXNMlhN0OjMzJR
GkkgxcXvjdS8kYN5xTI7DaEZRBPX7Afg7i/QYzQlAS5f+dbun4Iw4SHjm85hjHW4
v5UeTQq54nKn/+EIlC16gtPZXmGDvJnuXV45eU7bz+09Twfi7KwdV+iT6MJPSz7b
8vLuu5tJjsnxJ/8ofxcxXTSrct8jZmHBpAU4IiQYY1wvY7N/TuxQinP33wE/5hV3
eWqi4drAdThTglgGFnzcYotyyk/6XIyXPGaanQ6BicprkxYwMHWik288DyXSCAjE
B2phSp3a3JW/5MZueVDx5WSHQjGDZ77zrCtKKGKGffUl7RHJ5vLetcOB6aVLYqqF
1h2nAMIFB8YOwNckA5WGPjXWYVr4mo6GCLXrkMCPRXwxhOeV8nTg+XJNKvneXBQe
y9Vllr3zbvYHOPitw8tBNd/shLX2Bb0+kRUPVeEMai2yRjoD7xVaHVDW2ekTczQX
u3IDB0cZluromiL2d96iI5tYCtea2/GpsV+f9xLDzdiTHSK+oxumJIQ2w6sJsjjm
TU2BOCYpvwFH6mtM7+asBg6DzrXoNEr79fQWb6BQVCVBhLU833VOXVqEvr0qSLlZ
PQGuCspevE8/YDhawXe2TS40gh1DZricLyyIjf4M6Xpahq0vKq/qjMxe4rciW4BV
41mEvVAISG1YnSldb6U4oeHpKOrxAYuIQZpy6rJoysdmwEJmewrJH9pUKWJg4sNa
3D8XATQEzSa5CbBpy23SduFu1OOJE6iioifQvf1LFF7D1VvWoZAKbsmKg1kIv25v
xoZ2pxuK5uQYtKZGfsVYavoygOkF3385ckDSelx6K5ShX/BxPTL+U8rrYq+hQP8M
TcY+jJwBwzs17DQTFryhF0h9cJVf3QSK0F+pdV2JgOXNnZnbrptDQcrJoSSTh9n4
Qvpi8nDsi+WJJo4ur9a2bDRnmD6vxQEDnfnZT8rNPlV8POF+5Yp/DiAZNRe722Ej
Hjfompzm0hka0o9BNbCRavnAFwhuL8Elsp6W5folURZi2dXOph3WSn4bUa+m1yI6
QLlMVJGIjffo7lnbwosc0MhHGu/+jf0NuMt8DeuqF6H8sWYEPBi1Zxh3lpmn2QTe
gzllmBitwksHxULmuyEEAkPn5/sZTbaLJSaCNSGWWC6gwNzseKiB74SOHB+HaUUi
9Ic8xKR161MD/N0jZJ8cKiGqMm5TbGCo44xioT0Xf4Oiesjuvkdjbit3VenYAdHA
r23dAjjtzplwzqkN7EjuDzyQQSdO45+aWvH1mEq/q9ctVtBWJQHbYjn5wk3wUFdu
+Vyla2qXpY25ZMaoRDyoZwdCyr/MjONiJhqwGzSjmKJlhZI8oZq4NM1a6Yr4b+wT
brsAscCUoHt1p6LDeAKyzuRixD/lvm8eV6F4jeLnRWJhTjUSWFZKOiPRTQzlVq+A
uWEY3kF6mFdeHYtuP3ogJRKaO4dwfzPZK78J/wbd9C3wW+tbn5ImYKkrI8fbPIPf
FpFc9NgHYAMGLeoVDUbNBT1piyxA/Zq8+Tw/XFVIOWI8DMlqx0OPjtCGDll1fbRI
64sOsXUhv5zrDZSEhfVOYjyjnMNjS0VqfcDKKuciNUvwDx+94xp8HVYwpWWSodyU
ahCR6ctwke8mljgB5Q0OEg0XHTpceO+qRGPS+bn5DqNG56oCbUwCV4S5nH5OTP5a
8NGoDoGN+7gAjVsdpaznqr/sD1sbwd14cxkXtsOQxYncRVW6L8OGKmU0sLsqX90R
vqlg6hD6hgYP7/+ERtgKJsPO6kv8Fbkln5jDVLzCs0cVSBux45IzmtJt/S7Tpiy8
UjI/AY5OsGH/AnKqCJmQ7545Yu7BH2Zj1IwVNadcCDddamuhz62nsooJSeVwh0zK
SiEYlnOAUe/SYFX2D9QsiYQpYE0gUX04cC6pxiPBOEbm3UIY13cdI7WOarDtoSid
hgupOn4X6BcGxC7ajAv1TcPX/2FgVnwofE7ZUUQrTUDb8lFBlpPKr3kDAZj/4jLc
ITOTkgZDF1gpNggQ0+li3OtEVwN9bApk2n6KE2t558LBG+E6lYEgnGkdptTVWPJX
ZdT1MaNt2+7fY6ltYeuZZwvXakmC2o/4th+kzPwFFeX3FTP4ecDpczTnROerWxNY
E8Ru8kZffuGt5XOcfLc59UTTnVdFE/Nx/c9+DOhBebdpMIe47fi+txEjGQCYkOyd
1xkSaywfaZ6nhyaS/nDBMY8hT0Goqlsb8MrcOujYTaWFvOuzfDHncdpY7YcbTwBy
Xn5TULn5Oj0XwYdVEyicnFa5kSVzYyZvV+Qbkw23GAMsAHAs20/j8tRQO9A34f9A
4+bFIukXpoOrX+JLGlbQNaXa9JH+oNktgO8hSKMkUkTMAmLqhBudvbNif9459ti5
C92IOIAakalpnuNkL7HlU2ZwJCvBO5k4hU4xgITWzsyTMoZXdcNvdmM5xuLtq5eL
NWOSp+FCX7tB1hz3Lan0hoqiC8lqcI8J0XJ9ThjMrzQe3TU/Ujd7ij/Ooqzkcxwj
rSoExgEzNBgSIDf4hGBImT1JpORrZjUPZB4l2ZL0URuJ/s7jekp8ItiPCW72wCQF
TOAjgLwRZZGpEmuyMAiGZAsO/SUKF88MtmbG44ZYueFj5lVVyyfxrP/MkMDkNJuQ
xSkt9OPdgeQIOdCBn3jQ9xUG9Cf40johajxa4n/h7Ge1O1F+XGP7B9aCthkcCnNy
eXNN1nHAX5eSf9ygXyZ9NZiUXdGT4SaeVygCwb3zgmxDDdIRfXC5vFMa/5QzZP3O
dd8A6OPfqrX+/nxUPFo8KilGlXIVZJQ/uH2/PI4/43OzYzYNDG47l1dQOZQ1BBsV
yJwj96w+th7E/JRrHPj5RnOaMKW8nnJAw0csuqIkYL2VqTRkY+7jkI89lUo07sSj
8nhbA9Dv839BrTiv4YvqSCX/HfYJbAqG9RxO69tv1OuublkJplp+9spX6j7W+pYg
Z1PQfnPki6k9JicnuizDLSY+1MrRwMUizD2YvL3BxOo/7wNOAfDy+ukibKnJc4ws
PX8/p1OSCLlpZqtdzmITTbVV+HGmEH7+0HllnMjTZdEmV9F32UqW5GCtPLik3mrS
IHMGVpIYfznzzu8DEnxfKuPIdBPVTx37FAS5E1SgSkcIXnDhjh5wZY88PPmXkZDK
S8y14twh1XfkAR1nSvoXEm+RBNnSCJRoBmPNbv2SC/1ozT5EZ6Ltp1UMMF/TVOaZ
fxc+jEw+kOV6aSs72cOcT5SsZdR83cQRlv1dbsobZu2yTF6P28pkytwBtFLHOqbV
yPSQzkoVGuup/YygyMLZ0esDWKCFVv8MkK7nBena64ux6BLPwM6RE7Y8OM1aVSgu
Jy/bWtv/SaeoyEqRSrRRdD6DOJjIB4Pb2/v2l/Xwho6QVuaSAh2CDbaPhENawmh5
R5iq+GF8xXoabV5pjtRU8EcUO5MGAU7nyMVRuCLU36uE4/J+2M1JD7BJnrm6i3w/
hnRyC3PUltKbDBLVmiYiZtPuYFb0QGm5zkkl8Au+5CLYPgrNNuJICjdvV0igduk5
oFkGoVU5n8o4T74fMob40XKLZx4hysitgWZY80zd/KaSU6iVMwlT4gnnwgj73H+5
JJkZWHgSawpnv4ketFV4MYLOOOCDCKAdPluRL4WFwxhk4N1VjZO4L4qkamJblqqA
WlvTNh8nmodlmxfc3M48zeX9GaPW3nx+LJ6POFkWW9V3oH8pPBm88nozcBjfF422
elU9rzzjGaCzbmSxNxFN/10EtgTNijrTDSSu9ohMH8MDJMyoiezJQ9S7bQuVwpsJ
1h0jdqi2X2RuLCvtWAG2csIUqcNjkcNhWZR2ukXh29rOUZODTtPY5ieirgi/KK1j
RGmDBGd3Ne7VZnW3ykaOaflym00kvWycS8BQmMIS8ifo2aic4CImGUDDou2Zbp+i
xB9+SdceozTwLsAGKjS1pN7oUDAotW0kAmJ0ei0GtzK1eTJZ2xMloWCwttSFz2/1
y849Al0Vre6zvj+xnKFQTKeE9apMBuJhM3HyVIRhj0sN+IUszXAMCXHWo1CQQjUO
qBoLYSR8TlDhsOoszvCRd2WeyxlG/oEb463uWN1vitNC9yKG/F1WmzzJyZIzMIX7
THhwvQR15bof5U2/iuwbUzBub6hyFh4HxQBkVV4uDPbEp52WF3nCdbRYHQBfs40/
GILbVeEvUsdBX+JbtWa8QeNJ8dPovMdseFNZ+HgiCrUqcmZhpLAEFF4LOvYo0wMK
vCcEUaNYpJJylSiq4FQKqireP51TvJgOYc8pQ0c8cx+MeC7ZbNTHD9AEKmqcCDKu
/RQxZigBJSVCByzlILQHw9Xr3tB+WJh2+E7x9pMsW56QhwSFXpoQVq5mvtYjjr4m
oQikuwaEQMJ9+/syK8PnekhqrD+QkXeg7dDBjYh12sXLH/xBO09nuAjrv7ta05VS
Op7z58UduPP3JDYWtOrcsSLB8HhIHoWLsEZZxYPDpCs9OiHvPk3zOMSHcy1cL4Fq
VktV8GtthbPfQp+NLn1EPq9F7eLASMdKPrV+KvsZiPiFhgmlg/HvrgA9QbPIhl0h
YzRG/XF23uvv4xfXMk00283mZDX4B6JkcPbdK9pBHbwaChbqATxLlk1ITfBXlQ9o
1FW8QEXP51vw9uW/JEqolJWANUBTejb2CurEjZoVDkRC4VivUZO932AAyIPgVWfb
qVFeBdy4SmkzC7Xdl4FpBz3OCQMo4K0NO+GW4qKl7RvJFSvoPfgQoNDR/URB8qbz
/br+Hz6eYEpD4InMUDhtYPsjlBd7Z4qGGYYp2unJZjhfAUl9PEHjRNB0aceItf1z
BviTGeTwEuFbrBM3ZjnAqfALDWr7heG0n1FqOE6WiCtbJ9xQOXvVMG3+DrJDK2+9
oUsK1Dlu1CGj87W4e+Ne9hiOPIhhQR981PbKtWx/mkspwvangfXMROOu8IWU6ytM
WEey3dx3AcRsDP1J6flLKAUc07YzywsgtaQocnUupdyEIWNKMJB9EGKQ2HwA9UoD
aqDlr96MXC9kYOIyvQ9m+otgvbOXvgmOfRQpRgMVz/p+meANncm7ZFaCTFskwb2F
j2XkK5G9nLYBTRqssL4Fysh/hQiEU3MIRJO3+4c4mRo6Sq+/XcO654qpx/weO4xb
EL1JqYFKnrcfHCmBE8Mo+bzFLOZ+H0btuIvu5WcYcmxL6tGNVZkIqRUrgzy26OZR
yymsDFiyUo77J39cJGHx2eb3kYl2enh3UxiBNBtuOSioBL48EPPBH6aw50x81Vvp
SVZi2vn3ynHLGmXqBCGusU/d7ghmQ40VtC58SrlaLooluyOuoH8tHA+PpBFMNgFL
gEZl+kTJ6iyB2LTCDnxwfZgrYgqsWYDUm/09tcyx8BhMMarH16Nbs4LKbvgRq/9y
NFWsTJSknlAMmmqav+heLjZ7G1tNJBeH6Oa1lS8+SMw1O3ovYsVjQeq1spwYveeU
pHMGun+IAqNVAM2iplmv1fGBBJPKs1YYunzyAt7dP0JOS+LuVZp53wQvo6XLXdcS
IOW7H5HqziD2xpl9bUcAO/dnFVe64VEE6Hc/NHo6kWLoZ4xKlbMxC98++CS0Sc5I
evTbkPsLr3Q+eUumPxDs25q7cdbe7pKTRWv4RbgpkCpIHjNuUq7IPU+rXp8co5rN
MkPBbPz+h7pYyUTtImDZK+NYpdIQeQnvh4MByuzP6r9kQjiR39qvaEMMB99D+oJZ
z9mSrna9ugIkVM5aVJYS0YhULE8jPCzCaEiKfYAoH80Von4WYnk9ZPRWlaSLxS1w
KuenklVKipfaPJM9cncN9Yh1qA/ACejzqsoW3YddWJh2YJrldlxWd8QE5MTemdzj
BOPFUHixSL/5crguRQOeMcuTuGEB+sem+z0wDW1Zva2YVQy/NDnQbeJctmfFrViZ
+22R5nZdS3nXN4KXMUgaRIn0ooc04MXc5ynSttGLdysX03OZgYEE/6UVpzj4wInu
3XxuCpEffw9dlZbcLl4RgzspKcsaWtr0ae1brUF6T5p14VGpa1BmfI2Dbaw8WhH4
Glk9sgZZ63xPmR3ZPaM7AA3o8VVzEVzACVGt/ge798TJlFK6TbwUaIEsW08FyZu3
eTCiM2Zx7AmG3T9wCniYgRTTLAx5YlHST5H+5g8n59ZqefQZGmsUx4RLxoRURDE8
yzccsR9vf+bo1m7QrdcBw4wdQrXTiExQ5pgEZtaWCe+kmcT+e+2W4i4FYS7WvQCI
3eO7v1fiiT9GqPLWAA8K+mQpRkcZmP+o4lGigaTXn4I7CJZM5sQG/q1gUjbfiJ4r
iG5beTY3KeKcQmYS19sh+zaJiO05QU7CnBT5tcEL2enR7YFR2YAW/KFm+d+HM1iq
kMlHDLSb9Sesp+oUUTJz2UmCtwqR4bWKUB7Ub0+4XB8oaXoo9L1kTBGutoVRQ09p
mKYFVFbifax1w9mSXiAhiVrCCVOC/2WuhDy8sM/AppBzQwwLf+jaCGlxX1JZ//+Q
q1kW8it/NUEkL3QzmO6Vv2hsoPYKfa1U1im2/cGOFLGITjUHULzkRZJa98G5VuEs
ObjiVskkrgf1GBli8KjUz/EyCkOyl5gxOjakwca3NC1tBRjeQjjiya6a5GCkF2jP
1j+m7eGCQY7/2x9RZWyu0G9GH5kiMC+/L8RWQehVEazW8A5ygof/g5mQ+43SmqXd
rrqJ7gBnNCu2DeqM6VgM2adZWEmgRr0G8/iqsKOHiNhZU62OdC44NYB6yCH0KO7I
drnT+zROeCy1TtSyTf4EjKe2+YwEDHjCUqhaaEhdyLEgxQOGyvksgEL0ThtaVdg+
rCdnILxgn4FwPkUcazoqVXdTyJya/4iVtDvf6+h7WhsFB9Sp1c2GYw558fyLJhsv
yNmlffeb37SNUPFww329hy6sWgrKcmxLG7u5tHFvSXFUPR1Kb0j0LsvCJKgDwNbI
fjICogX6rF5b//cOCDqbt8w6Y2Mpq9tmvXAukHKXoAEvhxxGcmzdJ+zPFwDVEJb7
UU3h3eJSHxq8vv9GO/vd67ZigjeihIh68xLr6HX2TMUszag28E3LhcmqRfJubKDk
x+/4hFVGXcxIdGCCxuU7fFbJDw+2JjjCS24DH8W+XRAy6e24X+RTqfBbGj8tA3n+
mTT9Yny3z/cwVprhir/oAQkexEtc49RZAJNkWnUxGWndFE5IFi2Aru/08r5PWjEJ
wz3JIld64o3QYb5qBcOASnH6qRHuDw6EPcvAUSBMXSOoiFtI8UXj7FltT1JiDL9A
19OfNfpYld8mSDyb3dL47VtXV5rhEIzEzub4Inj7J9eagsz3VJVGRIDWR67h8zws
Dl0iRQL/F8/MjLlVk0yy3JGbI3i8KKVgAGxm8xXA+U5Yhc42AbAteD7LLXCdU+EF
jIb5ODdBpfT1b2wrz9NAiwo6SHca39mzjQ0OWSqZ5X/z7luYCtdf+W9+RYk14wa4
t0ndLRqP1w21S1FmjuFi7Z+OPxr2302PRmSTL2yBwhkY2bupSaWWDyibnzhQW/Rj
Dj8ryI7pOu+VLZ86Cn2dukSfheiplkXlDXkc88nOReclMmilmmeg8RT5HwC9jbrr
7RW3klgqzBlzTG7bRlvRTJQ9P4NAJLM3E1JOj9rB5hoBi07xuwOJ3l493oKr37b1
a1edqbJPtekZSHKYLacXFhFGDvqb0SW+XPjI9Ezkjo7SlqK6Qjwso6Mzs59LOWF5
Sle9gGs6n2P4Y0LVI3zYQ4w3S+P1BeUJY6BcGR5+MUmToGnWeoxy2aVaotzfR046
gaSxKpzNMBTNCnpLTel+PCvzNJ5R/NupbMSgsNRoFYugdarbJ4WP669NEQx+aSLp
/9AyKccWqs+mxub75jmXLP/vvKIlWP8XkxKqmqugTeqcs5tHxmgoVZqGs5j4VaYm
WMo4jSj+QesyFgRCaLkSEtO+FoEuisWXBYpD/dAp+VUom8S0YP/xhB0OSkbzw79U
YP2g63WaIyzvWrhusvsHTMtubgi2tNSQJrFQsXzwt2sBZ90pLJgqOo0YFRv2ONFY
hqo06PmWsk9hquq5nbNCR3R8LXV0tn7fI4N9bBUZuYxWi82oytFwI3D4uILXemyd
LcFyCMFoUbaZru07OeYl+Kcc+WvRqVAEKabT5Ujc6wuYwSxXHJxq2BdDdnsAGZXK
5ShbHvt3iJfYzbqoocahnMPU/Q4qQHTLnJaXdtr0bXSA4ZOBf5WrZjKNDvJhNXjB
3kudVziWy4DezyUvGkmIX9ZQvBLfz5ezZSG/pyD7iSjvzYB0qqLBGKkNCo2OZIeM
ye9Yj9A2ZPENg7vFz2xO1uJd7YiRH4POZzbmIdu2hO4whZpB43nZ5cEjFEzYv410
82umW2PAr7VRznGK6WyBkGbsEG285CS/pdhbtYnjXr971wi0GWgAicC7frGLqK/x
i/FPadXvflnIwx7VSs5nPOxMAmXDC/GQAS4916CQKWSmJ4vHKZEdN8RAUYWMafPM
EDpjLWUupfME+a1TZjWSe8Gigy4UBrbp+LKU4BoDGOgAP572d1S+Qaq4mwH9jj7o
jaLSdComvitX6gNFEFq8X+yD2ESLoUyxrj5nEGkAuDPOo6SNibveV/STvlNLI90g
ZEJ8Ba0CTBe9qocNBBaxhy+OtbtRTjig8ID4R0Af7gVogkr0a16saj+N3DNYJc0P
jPRC12psVIXLedNmmPeGHo1unbGIzz/12IF6ZDVX0PaOsBld2FWTe6YvybFvqwHw
DyfmPtAPO1Vqx1pJaP7yx88nhI3acCz7CAbcwJWOePZE3LZIGnU6Ee+Iw+cHzRSC
oOFsaLqBLPGri2RKxMeSF9F8IIa9jBuOugWdfiwzRFiO9IrCMa78cG5lOw19pzPS
1Pxi7g8mVEv8mqjd7VQOAkL20aiax39klxDVze/AGRkOTLsaDJImFajz6W05uSG7
ktJkpag1zql/O0oszwtWR6G9VrshRd1TqnqS5k9j/ZRlrjYTWXGvNl3LtSReRWom
7vUitooniTsBuF48mY949A36n84NR39fDvWvOLv9tpJ/8EnvzLlSd/pNWjk+akwt
CyZFg9eYmApoQCKqxMTDCb2WzQFHkrZv6kcyNpNg7469eYhC2YkPP+hvdySz53YB
ahagEMnuhuMT7dl/xm3whpsmHv0w/4m9N8TblJUE9jzCH5xNGeEqr5jDXolJrxcK
mmebteftyJScj/frlKSC4W8LwsFfEWYJz2hCHPPJABwKuPbS72+M1qAggQ8gM8xH
W2cxmpZWAKYZRg35jF3HjkOKO0R7o5bpoVbiR6942N7fm/JwOX+yGoWWilPz3eZE
8c9cGB7gi/uEIWekrR8EfSE8GCIJ8pz0relhITKCbPppXGyfx6ufQ2IY8CMHYnwT
8gYxn/Hbl6QnG1hqHZxu5lBtpT3yWEyR6Ql+NBtjTVmlgpJRno1lbt/7iondUszK
oo8uSaMrxCKmRAmjf6bGvU9RvGZm/5uRudlUxrDDWmdhpgMr+ibwEtDo4NvA1d9g
TYxRYYlcTZxlkvOmuIzI10A/xlIveK10iAonZ55tRYoFE5OD0QADf+Rs3k792Olz
lm5WfQigyBS3iHfvGTFrtMyni9xivywrEx++lBLLoRedDZS2u1of2XBmORR/YHr1
1UxJR3horHqFd6+C+IFeina47OW4WUAXNHB82n6N62p3sspBXuuyQm6GTGQKDNuH
Ye/d1sYLD6GEwkvJRxY4oF086vLpacqCufBRKcmWcfLiqfEoZU0jZ65aqdDDR9HK
ymXjUioEpGkXVrzcb3vSK/8Ssedg+tkVi/HIaxCC1/uMMcbqu1uv7ez3ez5nxIZA
oKD60/7+AcUl0EdSNL9CJyHIsS0ETNQ/7TuuCcEEpP8pVi0BwNBPAMN+mWzj98md
H3gcQCL4Shq/0gartq6LaUw+nb4SlgH484PqX2kRPC8xaBSZdfP4G8zl5nj3GvlH
as2GRnxN0oWZ8nLzmZ7S0ob+Fe6S8MUUyiPnTQfhUlGMFqXJRGLRcgsr10Xph+1C
ui4nkm7xunc74CIm9nYeQya1HIr7eZ9RO06Hu4Eb4WotraV6oYF2xnSXZW36zmg7
XFf9Hi8Pwv0470gNnko9Nh80/mxgTOUjEhV5iVRCliacioUXP7JrelzrmAvrqBSE
Ak7HazfKXe7MLKNWFnn+mr2X4XgY+MVyLc0+d8k5OfKtsM7AQDxJnOmBXi3JoFBx
UIYP8yHyG1u61cbRVJDqXOloOh4F9vXowE3yNCCzJiNi8dwSInPyz2NvVLwha0Iq
spo4i01/FJtX/vifRE4tZq1z1x5VWUoJsfrn3uKjINLO9e2j+jKhzAfO+ebaht1z
beuwwkJCCWSW3nZQ6rYyh5FgT2q2/M/G51GJGTnOhp1ZakVr6p2wrU7JYXWouSbj
pPRxEhZ8nkgJo9Z2IOl4BSCEqg/o36NzsNvIH9Rp0VnRMUHCZQKDg0FqClsaRS12
vllD0qXzGu5tW9zDgpRBePvFRkoIwuFjI0nMU4lJO6iS1BgEd+yERCFFEgskR8gA
PHh1HoTIy9N0eSDlxFACspkqM34ZssjUlcnMj+Vg3ylQZ6KQ8U+jHzihREX3/qyZ
T0LdkTFv7JXLlkj34KS85NEIbXJuK2l/RT6ka4CwdCbgsGsADybe8qAHQGBlCOcI
YGb8QdV+StuDvA41JvYtHVNj0ZUciyuzVvLbd15shVQsDtUyjI9f63906SQR8R1d
VAC3cx90fbypdQgG2lgvk6WFag7S+Zuw4jNxEjTD/DT8byCyCZ//NnXE5/b3r82Q
LXKlzZexbwYuGznRLM1eyDpl1Kw3q5f+MKcY02dJ2/SnkY2JNCuLy/WSCqEyGGb0
7BnFijBicLD+QXmbeyWL205eHZ5Elr6svqHgKaShIOxMfHDh2mnraS2F1DMBF/ZT
VNe8GEG4WqUClPo4uCtPw4CPmDjqHQubB+RvT9WN+PNlkY/mI4JuDYrYTVF/uaZg
UrxXD5qMQ4Uxnzlfzn4pUvUXSxxtAfiq+7YyCBr3jpf+kJcDe4fH11xIVJFxUcCN
dFyAhsElAkcBWo5KvB0EQY8Cxr9iePbwybB1AXU+OLxXz9hL7VojPMpdxjdeleAO
yUlzgIAt0z3pxzVgA1MNw9BPU1L2UNAjt6dY3haSKY29ahctZSp+cwpx2VFg6/+L
9JJbhrFM3b1ba7dro9oPVuiFw6kdvbcjldcCCtyQhKwKEmCz0QAxkEYO/D2Dfbm1
KbhBxPfGJxAreKZc9dleXRMNljVMv0pShbBMdFU3ScV36qBHKhuue0mV1lU6vDED
BLNNyxqH5bfr15PQgljUKThJLPR+H5GNDu7XzAvDxCBZt4U1dZ8WkhbdQvS4pBjU
pDYWD1laTz9XR4clZmPlJOsiJBWAY4Vtr1MNMD/OsXZWXzYoo5+Go4uOvz9CoN9k
fa6rkItfbeNU2YKYbBnMLXCBGiS+bxrV5+rVXeq9hXnYb3+d2mQsC5c7AlKV1eoz
JQ9rCoJ2K7OQO+zNx1eUwpYrhspVfMYFcfTDgTxK9Dujj+g/UcZn1PvjRSjVTTC6
7MNKi2881zCXdiuVard+uuNbX7Zw5zqwcLgTuoJIggRwA7/QREWN+IImen1+V7wO
WLd1KT65lMADPMilmbEyEXeh7BmAguW9bRaiC8kzBQgV6twodqKUR23lMegPmGpY
Wyek74U0Xhz2Wk5e2v+Bo3Qn/Y3GkpY94kCWJWkF7pljwe/ZdzMFbiMLofTPwrep
58oL+JxJYYf8GPHX8ovQ6entYgxldiLDXqdDjL5I0Y2AYYdD4yhgOKmTZlcEEaSl
kQBzPwIQex+9GsLpfcDXwcmpfuFQV6qAbAuqUi2wBh+9EXeu5VcJqHjUP0K8M+t7
+W7GUF6rZiXHLzAzpKsW8e1RJQjw011Gp43m3OC1GxuW43ELACa/bwg1UgWSeHAv
H+kluiZRRPaQofzxQ/d/tt9NvHBbtUrzJHRIVBxFhygj2SBRL0OtBA38O1NAPF/j
ZXQi7TxvDe7YNch5zRjjt2PvGVOZU0rtSWxuE3ZoA96s1vuaQkAvGpEyoBogNAQN
WyYTvWzhLND7YW3w2C4ltXX2j8pjuFAu8IAx1zsBABXnyY8Sru/tKftZSIwVPH6S
Y0drXgEfA9sVjPg+LoS127DLOnKi6Rrv4kZZuTQcSHh3e0VX03rhGQyJsFfgOwrn
whUr0LjQHTVJ67H1p0hvZxv82JEJVxOftyBOzCvAZaHa/p+Wwkp2viWEE5ngVsFV
NDuzXRnLiD6IWI8zeNjmuEJlngl7jSELRFXCiH5ZmR84NytiwQZxvWiQNcHDJjCb
rYyQP/lj/xZ+Avoiy7DRxo178CiVl8sjl9NN1MZY9ZVx4BoE88RZueqh1JjlYOit
TWn7mnWAF5FkAtbEQMBZdlVo1D9Ar7cFcLyg21MR+OfzWd/3y/jyUowD3lzv2xCx
a23LgLaW4cmDsF53A58Z3MYgqNrSFkw3JyXb2PGFwTy1SraQ2fbvDStec/u+bTSI
zMwfN50LgGssiOjMTDn3rpMK4oK8rfbJmBjWAMGuo/Xjse26xCNIPf0+sRmKKmp2
p7LS8ev5x7sUuJLz7Rv+YWqtn3Vn6Dt0RMpm6fuUDMmc0yLxkQy6r6mR3dZJ3eO8
c32t8dlCUoBv0a4Z0r8ytWvxO+zWO/zhSLbcE5gNQpRmcXZFbzEBGR/sVQgHvcgg
b27Wn39ehFZl558tDH4Q8cFW2pa8J6+03ep9E7b6Xau+zRPOcK5lBcbmG5O0/FwF
bHC11HStkE3BJ0DHwoOSnlnGx0p7IdrA9SW2pFzyFi6HuuQutUItZ+ssQ4G/egdA
1fZmV/qIL96y1WbWda2HR2O8m37hD8caG6ub5wVFpWx8GfvivIE13XttLXCj4LJq
hoS8nnlQ2MGl8A7nGgxj2TsTSSI1UJVNRyrLFXaeX9s/+iUWuU8ffU57Tg6mkAWk
RnmgOUOZqIL3rNacwAVihIZTEBiVa9rATrkDrrAFvVTTWf9y7ocpzK7ChAbeCC8q
wj+D6G9Iw63zB58HnFIxKdEfhalzbF+ZwY2lz+KakswjS5rosCTjtICVT44zFbsD
Tsw7Baa3Dsk1k5Mo53oC4t53WidqqQbIYWJ01RpLOAgkyCu/xHvThq76Myq7Zm8T
i8ytNjia60ssJQXH2rw9fC6QWThdoXKIYqNmuTR5et+0nrK+l/floISnwRCqGZJ8
DkRNNc2/+dQXMzArDOYTqMeRB2PVKnI4IwmUMwGl8pH4KMk29VXuje7SllSkmPUF
YO7CIPlp+1GARYmX9LT5MDMlT4m8BQykF6f9Kyv0zlSMsaieehzgpFYDGJXoaDFC
QsvJh05ZVy0QZFGiGIqc5DTnsVJZpaJwUEQRxBRfS0HIK5M2Fsu1LSoT5tpN+7S3
OR0L+L657lrpBa7LfPI4R5cxkbvCh1OOBMvmbP+ODjxwVCCns7uFQSIocWpLMb+b
cLqHein/qEb07LvvRDBfMDg6ELJoJp2fMm3PivujTjV8y6hJNMFmJIbQ2XOvahot
TDJLFiKv1xWWwVIgIy4QQYU0eFwbTqGA2LiLc5BGlIe6fH2tc1d7ELXkWn96E4SQ
4Tid93snUANHGtJvZShzfgIGs0qv8WTBASMR1kFdbE4EvKLdHg1SgZ+6Br32FVyO
5g/Begwj/YVCU87J9h/8pKtvx97CkDqlmc6Hq173B5m+v6apyICH/DNddgr0UEkr
i2mLsecoz6P3SZR2XiAkvRkKEWbwCJXgmCrMU4FSgJSBaewNcPrrCP2yx+SY8wpp
DzSYvlC/DqXM0Mbbrf7CEdqKvAhWGEyrqh7q35pZbWwuwE9jS3+YYoGBmJysw7J1
7/r1C9o9jNJc1d3jG3JBI4XaBWhczEsxHS2DvRyDxnORbSpsQBBirgynouL+N6b6
gEJt/+AAW8dS6+aZqcygNQbB8cv3Eh/lG47bnlhZVV5QpGtCgnaSRjB8l3MPE3xN
L2tkmWMiVHDK2Scr424FTaRN/7xyLAwFX1FVyS/CMZmDTRzIOc2lMQCLnHhYdZnT
ItohMmBBL1nhgUUlewjtC+pQnVcfnh74HkaQQbt6EaF1yFjJC2ogTxRmWigeKoSW
vKewS+gt6Y+C6UZ3FsDA+8wAb0FpLBRrBIF+N5Ez35z/z99xwx0gW/As63El9+Z0
3JoBomIjgy3rQoqgDW7O7Z2HP0EmpumiMhbppMLmBIp0Z8bnZx3ZJFzfT0kgdGpf
hBLt9tt9ZYAj8H4YJ/JF+k899OC7EMpn1AANaskd4wfXB/gO/JJma8bZyLVyJTw6
ErJFg5TqwZKFu30RvRgXUGbEcIOVZb0SDSdLu0byJKHFScRgUnK/MZJUq3eApO5Q
pT6GdATcBsfh5QHn/7SLaVOTmcPZb+8fgtfV6ZN3zDjT9tL5QqO6eIFPKa3YF1gj
nNR8ax/MS3c4xTUEJJ3JPz5Z3Z8TqyEWNrkyQo8cIJdbvaFjiyuY4grq7C5JLFOo
1fyiRtOKO3H+0O1j5Q6nxcBSt2BS+UJRkXCExNbmbxRxi46mIzcQmylioyP34hje
/LvL01p6Sl+8Ygo8BZ10hIPtCBnYHyiBR7ZEhqy1Dc3H7FaV7bpPWTth6IgD9v5S
58z3w9gmKFnACrg9h4RrN8l2krfaN98OzCJ9WCM+yfr6namVYK9n3qE3YNPtN9k2
ZNyrt8K6VUuZ4rcRFyuCmQQ8MSmBdC65a8KLDV35exzv2r4GAeHswXZ5fx3KC4Mg
bzkOC1sJzWKXiOdSL+mgxSRBc8LrD4A7Jc0Al6rTTWjw36E2VbNNghN/+1PSGRTn
a0wbe4O0mkiKc7iuQjfmJ7Gdt46PIfyBLV3aPhaozlzQ7fVvtsR8KgRdupyvlcKv
kpgIpu3oyPjVUJlEABzI9SR15SKHN2cyG6/f/E+WsU8U1VQFLuAFvIf/y8oPnzWq
ifnAwFrGqew2NiMPIn310sHKQQTs1Hcx/U5LqOEjy9UILwEzqF05OTrH0NCBgK+w
4n0gvcwfM3JfBueZxYiF6sY+XgoRDnjvHSPsDiakTW4DYo264DR/fiRGALylDF5+
1xPpQajKpFrAiddZaOgIqf5ahAhN+nJhJz8cVydUOVIQ120smBrns51fygccoGGg
zEbUuYAN7o8n7CtnxLC86CGZAnBPjBJOol0/Htl9z+rCY19bcx1uDFL0aDZimSSF
022MYfphPSmUpk8CLCEvhRp9mHkMPt2ndKaQwx8IKiYHwyVbVkDtXhVOhelJg8su
JZVrEqfDs62r2C5Ktg8u6F/eBQGQxu9IZrnGkAwa2Q+MowM+LV6uZLaPUMuc9L3M
6KLaXDXZm7xqiKqCXlkXnWWS6IPA+011eBpHXbEPrNm4wFNZ/9BWQJdqBTXgI4FU
JR46kd+kC2MIdTOvAqvAAwYWFyTZ5CvqDuHoQo94gjX+qPZ/q+bNzVV018KLbI5O
QPfBysi3aVdMuZtQsf0tfeoHZO7MLs/kYw7xMokP6s/w8jg97O6gHFJgxbJ79szc
0t/AptYpWarKKjtrW7L7GHLRgFCLDGEJ4/vHe5xcbyfc7THfxR+rvyLMBoDQmEom
NmxrSHoM+TeBMx1YLWEhsfekRsjzIOF11rXL5YzZ64Npr5iynhXmCRU+xoJE8hLq
3fZS6ydm6HNdF+EhWE/dGN3wwd9h+gzlfrgg2tVQ76/NCCB6ndw8SH83WuT6P06L
sdyopazd05y5w0C9CnLs2d/lOmB38F1K+fy0oiTH55MAnME86nFKWWX8FOoiXwHH
tOsOaNFjLhTEDQ7gpcjg4kNbCx3DGCHjaRCHVlQPHDt0mX3aBcTU9IT6KyVww1H1
v/hoY5wFBUly3PDQB1YbWFDmKPoayYDi+stEdw4+naMagK9+LR/a178H1Si396yU
IeIYSE07zUSq+VQC7vm6T9DvGyuXLeu4Nn3v1TNq/zArAVb9Y6JCK3pho6MVlym3
JPGSO+hrGYYRD41/xHzji72p72GCgOfOFJP8fs4oG+VL5PfPdxaQkZ1TqP4+vELt
HFpf0pF4y0Z0vAE3GWbi571BriU2trCTY0gSt6GUOgAQcluOPTvxn0gQU4JGOp3L
L+PpmIou7kJbI1c2OBAppmSNOtwXnrRl+0JCfzvgzhu1kK2ut/Tc7LtDHPCg5UyE
VoT82vtlGsDO/FiqmPcxEni2Rpo4jzKRfALyFFOpELVqZws6NE8U/hMzulDSuGaC
iT+ZrI1V2wYunciinSiKjRjJr3QOymdVLSd93foLoDzTGsKIXHKsYW+SXALgpFJ0
aiIpqlGW6Fnv0eyDLuUiQS2BJ+monsMBP4tzkxyDW0G/Ao+4D73hzwX38ItKdUsW
E4wSnWIu5ON7FXuw8aFloOPSVc9m2iqXvZxFfsEEOLoT6Dojur1fmmPT5QkBEGbn
GZH9qQYCC4Xbx4qnxs7IewrQTEK4qzlU6y+05uMFtIH4Yhn8XGDCv2vFYUJ988da
jDdHSmURD68b9YNF9fU9joN3xKpwHwW4BxMQyTQ73j22eWaJW8UffA58Nj+FZG6r
WL+eWPTD2gbKBNHdt97Od/xJycJimBvJVzUX2sLEosANDrpnqQumNonUv5In2hEN
xnntLhfplEZ9A9jyi8A5Q+F6lBP47anZk8PhZ9O+Os1+DHoouElkK84EBAkY+3Kr
g4Ofif2umye0B1reHcRSsV1pOAUayt56Yj8jqf/Ag6fPSq63HjaYB6aG8GzY6Esw
SygjxxUTQm6NhJHg1BrHcKIxdf6TaHcVBfr93escKaYnWIDK5XWsGpXkoMXNudin
7ahPSkxfdwkbWmr6SW7KCdtRn/LeFfSXju/6Cy8JwKj/RYD+uzElK+SuvYIo/4gu
7RDukU8jJCG4ocCdq3PDFEJcEjJH1A584v1JTckztJb91J++nvTeV0MEiSWCAtHm
CBJhbOnzxoONtOv6vaNVvt46O/VyE1RD9Abx76vbKiz9IFyfLgBj5Fd6rPq940Qi
Yx6JzMhZwaH15SKyekILjfGVOBG5Pa5QNUAzbqXYceqZOMTtoPJusa9S89dRQTHU
NWHumSqSqaUnNOfBztSaaQtn+OUt+CTRuXEErHrhkffFxR2mChagYkdtKqaJzU6U
dhbuc56HCC4dY74FI4+HvemaZV0Ial5T8EDhj2YUO8wHIC0jvJ3UEam7/ekGhgnF
XMeodG1QDR3+ds4sMnDW1ESV2zaSrnOClDPfnrpezTiq6WPAUABcxN2tX4GAJrov
AQVUC9cqmVHy43UkRnaOT3BBLJMDmKvo4Yy1dJbd/uEgNdGt3GatTjWC1D6oF0kw
ByxNYQbu4T8zgkDiaE7LeQYw8HBBz+qkSqLSdwLk/YWK7e+xE4d/OtUjiJvkj1gb
Hx12C9OPhUgPJZPGORYTEPlqlawhm0GZ5i8pYyJJT6yDur9mez7hHpDgcav4cWZb
YEcwLBjNIJv1aO/AjALhwp2k2CuihsD0W/IR69wfNkdsTGilAoz7LtdSZdrducRQ
RxQTyoAt3JOu3zkB+PXIVWNjkQG2nRg6NJbeYg+VVj9ln4V+r7qdSI9Ijpkne8pz
aI15LwXI+aQH5boJ3Gdi0YXMCRXfT0rdT3KRMNEtYUb/ZvQMQc81YrRscSR4d8Md
zYkhXQa8ooDy3UvyPKaCYa8TdHsJAwfTj1RgyPM1Ub4KD5Otf7pCCSES8CK2wqVE
LH9UrVrNYg3Z/xQNxluqYk/9Jn5Db7i5quiVuatDGdsYzliNTkkYVEdnsdlpezrS
Upk4Q4PwQ3Rk042bC3/Y4TY2YSG8OfTA54mhfu50FpdzYCjZXwnEP4KpEIdNNPjX
wiCzyg4g8We27NWDWHDmdGaWY/GBN9O5FZ0LlXLZ09GmzxVmgSADItYu7Hjnmd95
+OVm1G5YeYZHR/ZfupTg/V26IgWu30mV8hznEcoZTD9RWMietGwNcOB39KopaB5I
G4py27Ttdbt1+GZCuQMP9h27xrWB0lM3lO5yTXa7tWafMtf/f/niqO4OyUkfZeUv
hJZmjooz18QhSyJKzkVGzECxI3C0IrzPK8sN6oUIlEdC+r5I5wvYpbnA+S13FTaI
mDCWAEWFVAPgqYI/CzqYkeCvYasdQXaeHUHHH3WQp2jToje1vKIQ7Of5u6N8S2XJ
1hRDFwJrskplV29hGx5dv8/dKblNhrMjntrXRkMybEn8I9MxfaQaCqU2PzzhUXHn
KPM5Bmyr3mHWzpKkLS9uH1Le+sGP70vyMkrmPAzLkTfIQEuI99ca/PCsHKO6P56J
YLcSV3lM279YV7uJZtmXyFyQ9JsKTbqCv4IHr5C2ReqYZ7LBhl8h86NHAn1RZ/1Q
y/ALQ7JbWIIO37Bsf4Q5lF96BsmuSNlkkJHo6lOr98SdQA7d/Zo92MCD0ZSksPnK
3tNcdwwmaD6OLd93aZT5rf+eJR7JaRmG82FbqA4j9Y0dmF/ozwraDlI22n4prY8d
G/aDr2V7hE2gSRfZSTEMbvpgFndY0qu121sPFtOhpGAwTNXnR1xOOhkccyDHiD1Q
oaapSNYgUr6J2DGTxf+QAbULKXe9peWZ57i1UcusXNEtW5GYmS52WHB0AlKOnLbG
2TsLw6wFVyk7y3j0ND5Pjs8BJMK5kpbtegYyczZFPpX7oqyoo/op4hfRHwzMRHwO
qiGM2tSFpte0QGENu1HFjN8AI/7MkhOA+zTsbnvnFccjv/ULsVqMr1wMr0/bG+FQ
HXunSB8xNY9+1o4bImc3tGxddJheYJq2LlS+deFsBN6hF7wBmcsmG6k7X3czXuN8
KiFVeLuJpj1aOy0keienL27qc2m2digl1uLSu24KV3mb/97uPTLhxieNkml2HWlR
oGi0Arg3XWyLk4fQY35RHzlU31QEDyenjwdheF+Q1SX17mzecEf8yOA7q+YqQhZB
uDyih832HnXoIgGAsurVhW07aJk9I35oKpqCN31csmTtOSsSCc6lHJzHIPhb5ZY7
wEwm+xAazzqKf7Gc1Z+r7k0+Nd6gp4M9fZgje5tJThx4d6DJDDjtIloYNWVA4U5B
sA7wNQl8vTvMXC29/FISuK1LXnvq7VFk8dJm8cOpbew/rHqHZ8IMmInwrzqwfKj4
Sp3LftN+OHAuqjl49Y2hEf8XbTpx7BD+m/j7xeuCsXl7IiCEUuBAWrwdfaFwlRHc
ogN//u9Xvpjxw+vnC8ac1kdbkqFOspegBkuaqyxV+wnjThZWwn6Letc5JpPzzerf
m924rob8SyoLSJdEKr0MZYTRHdI3mEeS4+Gxu2izmwl6q6QqBytD4tLTJakxC5xU
dHn0bkQYZbLHRlo3SoS4SEQXTZFSA0e3sAEA6DVLIHTP74b9E6kkKsT2fFL7iUmk
rrw/gvik9Ry6hFTJ5+lQu7WvSKINaLdPPS3ZTzsZ/4RC/mqgs1B3rwj7/DGo5uIy
GL9JsC+FnXppd7Bg8TX1ehSnyngyYOOszBIh4cqGumkd9W0wGAeQXKL3s5FuU3kt
gOyZUFlsUq/Nt9nf1aDy9uUQF/iT+Pb3/wB/0x42rqZrM6d+TKceFEVbA73TTtVX
kKG76lVt3CULspx/zNffNd5N5P3w/a5WnBc+3aJheT//tOWf/1J9/6K+lNqk7N1y
8rZGFqNHM+R+Ug8CJtyUqF40xwgE0ZV19nIMJSbMJXsNqwgw+LVtwJt5JKSHZqUx
b0hGw/s0YPiWXULtP/gEr2FR1BvJnxqs91Tde3A5EkoyHkFJY2hMSG/eH3hwEP36
5X5FsSMMmNc0aJ8W9KGQOhvz7bRmH9gQTdqkHgXdsDjEiTZYJQUqGKmGxVERPAOg
1wWQJ2fS/U6CL7RU8CWpH+1tda9Qupq9bM8M9ts9ETXv5vU3bA5x18Z7gEi2PKql
N6yLQ/I+9czE/kuMSm/azOShe9Fs+cVtLflXMstHIe0uLk5Hlf7ydZzLKoMrDyz6
ishjy9qomRgZvrx0EXfA3JEa/9uSiFxRpbccDqcMAWYX6w69NJOnU2i7qGY9P0JD
FuEmohMtiVydSr6kXYyAB5p2dEPiizpwWVjPxU4NHPzDvmkoHgd9ZUDJgkhCysZ9
jgKPTMfa7kPxhvQHw6HnFLby26vjYUozIH02ESvJUNbwYfVQGa3sG7OTf8TYYqhs
QPRh4Oc9XvICh+wtuJysZTnz9vX9nNLE3CjZzd46Y3+fR2Iv77NEEBXrNGHSQJg2
NVguYY7wt9PGPEFMCfh0Si6Xt3H/ZhrznMGlSjv0y6aZKWFuQDE6/6EyhsBeT4d4
VOMtJOPUjwSAYwcJ3X/oc/oESQk2cnd5UaIkoxdm2qvCj9XasKwVgxl8j97I58rP
gnmtumqHXCJqu6qnGaRNY9AWVA9fHkSpYQq//rik0k5HWaZk64+/yKk7PE8w2R8B
NdkSgBPI+op69C8jv+zIDIjNfSDqwqQ+9Lbry2iIFZ7cllV4o3HG3sEQ849ZmW+S
L/uaDzsGyp0kXp9KsVbfLCIxXeDtPnRW2pUgYPj3Jz1TNFs6IwG+KvD+eAjoEDJF
B7E6XLJHrYBj4+fc0YlDs4QD3jHl3s9X0x35zD9DeUD3wBFAeAEOFlSACdfRXguR
uNSZOrbxKwnug/a1h9bEG5vK9OGH1Nb7TN4SXAllNSXcqJglxvhYnvU9uPtRBuzL
8Ha1vEGmA2XD3o+M9c0Q5kj8eVyUIwusBS2ROb538RQoF8V+nksMb9IK+i4keQ7X
yAtQvvFj7qKf44oz7YScwz4XBcQAP2ajLg8LxeF2xdeZXbcSS7I3fehB5nYCRsg0
zBaikSmsIQRr1hxdmUiwqIQaJb1fP7R+BQyj+UiLj4nVY9kDZ3WLVUEP7H8S5V46
9pAp+tUVJgkkqbmTSBUw8di7EiHeMgLgKhd39SCIQjvyA++KahHC2mFC+ufYnYy0
QE3NrZSuTOtnfD8vYLnLhq5MjC3p0epvpIsWPfi6F0gwXp3NphdcKox0zsAK+XEv
DYm0Sh6WHuUaFi+DxPamaaUqMQ4rF2r8SVPnzmfu5p4xfnYlZmR2nhSf2jp8TZzC
IzRuc0d5EROKu1xMyB80y9ub2140EuXYVD4Yl3mrikJ6GBiJSNzXIdiGxp7g6jPG
x0rL/oYNc23j1xzxIT5v2LC/1N7/vCVo5hcFIKRx7/42vXvLTovAk007q9boeZAB
AXP9d+lD6DpdGqpeeSkw75LtM0w1QUbeQCBaKgH5z17clP7ELqs2+qUpvSYGcHaj
Pe92kE0oxXcAs6kaYNQoNXAan5S0yw6xSdnpnMOCCO9EqQ8Ii+tkmuLssqIFsiXB
166DzY/wM3mVrz/JrBYPMgx/jwIwY8HH4PzrfGW9OwZtjZIj6bm/N/bSKdf8vjPM
ruTMyxCTY3N+ob7iNLMASI6Vzcmm4NTRqlrqkOKgQME1nfxlKaE6TVXl81kEDcPo
Nvdm+y42GbfvqTGkFIse3gKfY2RGgj0VCq4Haovy9v3bVDuHddi5E5x52cUclrVh
jLsHFLRQEEHN1uoEDZFUx8nfxIxPJGulGc1NaLourEext31BxzqXQPR08REnu7zh
MmX3WiaumhNzdgbls7IzLOKpkcJ+/csDdtLv6mLTsIsocTtoPccUt9BGQAbT9ivL
5e3TJ9fv0uZMiPo3kyH4lQbDfrPK4lobaL3AMRsZVJeSp86f641Gr5YI5CHw5pyI
qKZrO2vONxENhD/zTHhIaK92jln+Wo77JfXL+axmuM17aX7a+hmneYOvvGWu6eIe
nkuIbgPpTlqBo7eDQd2JrB6IPJYcfymHxXo/JAS1x3ZtlkMWBhRqgt88D3zjsN9O
TvczOsKvSK8B/M+gl9fehfBuVzZoT29ANfPGEx3NWAb6pUVOBSjefbMX9FawTdr+
AAAzr/WoGp6Ihid2IeWF5xvgymJxKktTjHqnxDdUWbjegtjvsf746HVnf/SUVH3W
VNn/kZTwvBDm4gLhddcyv6VRjzi8pD9FwVpVB8YYwZTKQ4Pmo1PmVUkvAzHIoOB/
n61RC80GUlM5gBJbE4VXruExZF8Yzbom/EX4EjucUyUzrlEYkPURzPZjbPeEMJse
OLBSsDR+JOX227Dri+RknTtxgxE46Vhx2Hl9z0oTSkXiXAIm3PqAtWFzjwxdAAFZ
l1RhAXIGvBk1ZcBMDFvvJM/QPGzbziViSr1TK4FSr7bmz00+0B8VBNrY227huFLl
6LnaXk5e+ddeBKlKz/ainUsYeBnT6p5EQhvmdX3xdFqIlI/Shx8yctQ73WjST6lK
ONhB94qvTNWH0hY3Fuv9Uz6JoJWW1t8qzsqN7w9oNlreitqW0Xhj9EcLrfR3AuV2
8pgJNa9vEN9Mz2e3gt8HernHhoOiPSHn2fKn1HtSuJBAc50eE2zQIdMczzbUmVg+
7PyvKIfiaw2tAB1+W8jeU/vBF/2rWH1r3YyCKFM9b6sNgkBaSsYCTWwnh6Kfq7Ca
xhPK4l42WNqf28PkonW9WIkyhJ9YUhxnl+mFt4zVt3yJH+JbDXEcaSsuT6b4MTcL
WK3h17R+WirbEJSOTDif7W8w3Y0kXcVJ4xy/l/57fg6+zXYkZpoBWtnojipebVEl
R36KejF+RAYxnAYVQDaPgW82SkG6VwA5lQS4MZ2RMp1N38qUidC4+37k7Pfgd+59
bPU/dFJKXYp6NtBb2E1d4HGDfEtOWE10Nru8tZKDqSxMiUKy8VxCWlqfejoPUqJS
syq6NXERRMLz6zt37ZFNYALxOc/RJHBadxKGpwCH69ych47fXnPxkOGBjblYKCJ5
VEflZwB1/V8J34age95fnQexjnDwTu2Cn1ORbs8shAaS4Bz43AdfrVQhU5O+kFCO
jjYzbnY6dw45yGohgK3lYLkqQRiUQK40lwT0/SwfoLT8e0Z/6w0sE7MMg1pWcjVy
Ky7lsTsuBGCvoQ+JKcD8dt9YSwYoJRkHz5BVhZ7DYespo99E0xcherizNNJHi7vO
CPpbU1WcYG6yOo8x8RlRY+iFdHYF3ILZtR8NzgXQNp4ZWwS/m7Otlu9uYpvSUCOb
OO+A/3F3XjXp6hppl4ePtqrE7ijMuUDJNNF9+Tw5XqeO5O6txBi+hyMwG3MRiZiE
oVwxigh4kUvnHhs4x1ACqYv+UbXaxyr92hOMmfvgdbK/L9HoXuYrb/aS1pCR21XY
H/PuJf6GwsLe9RiRFC6ycqi1KkHT2Hkht1j9SMjSDWxJEiV9F6IMpmJ8Gy7qJteM
d1BzeraByc4MnuGoJOhpZvTLkoocNyok0NVjGRqYWkLkPdrJ6RRSwFCcmzXadug+
KBZxtb3BrUtG9xAG4GzEzGVH+O2iIjcOERCj/UgVqk2DMrAyTSXXIagjDQ7XOZMn
7cgDfUhFIFKh30gs+Th1JBzIIy4pgq94COsQ+DZwwwWKSQf4VeIQCFmrC5weFZ5e
VP0xbmVtoXODTxooRxHhLqePKztGD4zp7lkN4W7lu5ZpgRmQxoLuoZPRUVEETOL2
sfLgfqT1Q0rbVOgPmfmEv9fB0/nDWgY45UDdAOWaVqKVqFvPab8XObmsF931smWv
DWaZtlbVAoB9VjdG7xrbB9LYocnKDHQS3Cx/5VBGPwIqtJXrqlXFZJvyqXtKUxoW
64VnOqjsSjshzocQInR/II0YW5Rf+2oe7WfUsPXOjMcePv+Ef7RVZs/E1DAt7ZNg
iGX6b0Nm2uJuJ6K7ue90ittRj/lf25VNfmC7WjrbqitDBBCcxWzk70HRouNjIrjc
dCl3aa3bUZHqz7WR4abWXZMtK+JN+g+xcQ2qIXsxjHblgnQ7y+6T+nCpHf6uCIII
NP+ppqwDu/NKltc94YvR64x+hBvDOGBB2OKOPlGydW9QX72LJe6kMLFsBhuye1k2
d8IUMvxvdiByrGMqLZTnynRsxr2yTq5TNu8Dr3Haj4hbTKt50zT+izTZfZCvkMMJ
5JGP0gyhUZoFmoNcZaJif7lVP7+RxV6oQr8Ip111jBT+DnuU4vD94xk+0LbbdKDR
OBMlL9s0XSvEQbFKxJQYgbAj8n1vwB4IvwgudHpC6V2CMXxGbnd95G+/N1nr+4m6
jjJ0WsnpsYx46+wrhpsxxgbDi7JfvCgfBjJ0KjEF7MP9wPcN7UdNe5sK/vqGSU5E
FE7bwRikayNlzIYwmNKiPAboKbPn7rG63sKsxAcWFfIZoR4jKPcjaCWpKy1F7W1f
hQ8PkiW/w52QxMK/xrv4U6NuD4JmoAhykazNcIK+rzU+UzPhmAA9BbPfVdOlvb+r
yRj1A9oJEoGfyBC0qjUjvC/kYC2wrvZJrOQfqxOw8XkRWKSXD5ZLcwL7bHjF9NL5
89bo0Ogk0rzEYp1YtPvrgexkE8bTpotGGsNPuYKo4kEiVEJJBTyVAaMDI5xUnsUI
7/oOKNrLDrpLKCyQgfxIBbmIe+wmiltP9oyan/idp3QuihASTvX/rt9cIXTIdRHi
pnnstnfBTTRTb+o6LAqF/JkcM0R9D+YqEGO6Iyegr82pkMnvp9u1+gN/G1YN6jx5
81MU2y5oQ/gk60J/kyLC4Iht1OmoiVgaAhxI4j6hjHkY3UmrDTCf+ZSpg7X8+grk
hoA2Ff0S1BveC86+p+TUGBPKJCFBbkWor3QNWFMwfuZPK0AtOrjTmPqeNpMYDygI
G+Td4qNAhcttKYjmNcnme1G7Ci+FNYwb4r5/pbHnEgs/ThDUvss4mSxpdlWAw7Pa
DMd02o8bIMHQ4lqVHqajSGwq4XKkIRoSwQR/yWJof/XzAWMBbfK4/G2nEStYhNsm
Xq3idlDR4qA0KcwjM0l63dpSVxYeaa4SPrPrvRafKFL8I0ij+wJPyO0jfZWb+3Jf
oUibawxWY2X7Y0wSNXb7+FEjfeNVP8HI2ptmpoqazThsuY5I59xVPf5jjyNaTQqA
WlUHRZUW2Zj73OiXpLEqL93d0DZXxfpvasy3FouVDkByE02uIP6BENGoABv6wy7e
CcKLAuiNuPmwpmRpgrp2fcMr47j3qI2PDB1ZKEwwuEVY47G5AQkQWMmBZbANIkEK
XCiQKGeTEGjYL5HoFuMqAfsUODChZ1OmxmOxSw5CbJl/6PqedJ+0ZIHHvfaXhDP+
ltswvxa+GUDAg0lPp8b6BL+1vO9vzCOvW8fP2bElNf7p/NYzOTLxIquziXX86WMw
0HbcExfFZEe2Rr8X2h27+oLPrWN4cRG35sKqTkZiH5tC33HXTHZ3MssbjPErpF5j
xljXPJsQ6kxaSRR8v4g6sQVnZnt6cXjNsC21fxgFzlujScITimOzpft7ymyzZ5g2
oyV99UeNJG8iUe8On7bF/l9kJNM0UBeeyrEo4U2UOUTdwLoLlpmuPEi21w5whFgs
JvXY3w9dAEm/IuE6DkrLlEfHKvvzcujLsh5JnVFqw6O29MwU5TVEg9lt3MbuICGG
N7yKzYxp58nLp+3i4iiDCSOHw2j/oApokd4WWvreCb+LI4K/C5zx2d7tDcVLW3rW
mY21BttgYaQ7dGlFPY6yYU9FxejV9dmC468agMc2bHqhh2g5PzACs5Cd6xv0DX1x
JRcTQCXrxl4CxT0u6Lyez+YGuZCikQNENlITtgvZioCxxNUwZmscSQJJq6Y54ZVW
Ltt9nF9/35VnM+ZpIWUBKN3Fb8VN9Y40FCWgxvwNsijGoeLlds+UtQep4R2O8k3y
SnpboVvlPGVTk/UNtBdn6khWVtBvz2+t3qX72sByLeD2QhozCAyEKkqm70e7A6Nd
q1gg6045MVrhOz5UvbV7P00dng/RUHTGRWQ1AFbc+qXvN9zOZNSWISI1je4Vfn5q
qyYsNGMsj4y2BZMtD2PCZjly8nWDjlXd70DEJaaGC13t3wOQ97YUpEAqk52P+bKW
d+Xtpkp17a8PGTXV7gp7strpJiKBsupIaAxCrs7l4ZcHqzOGtF8evKL4E8VHdI/O
mAsKSTCkG10adBVVDdSaQvl0QoMNOGiEt9PmqWzTMrMQI9QLTBcaskrtZm0+0mW/
LRrXT/VYHUbBixgJIKyDDyFqlMiWrnM1VzotoP+Qo72ndl9hWnLe2Efox+iRnAzA
aUX+Gd9AgAmN7/nPkQHuoWmmnJPW7SxYDcgu4l6qfYYYWRVS3OTWhQxy9fsjUsEi
vKLlBDI/IkJ7W901mxXx9y7f4ZUXnxM6sALbHg2H4nvfVOnlonzwwQKcYF9pzQZJ
ZlCZVMQ4TQdUThzgbS2S7Yyw1UZRhLYNewRrSC2lT8O08dgHZwDpTMHuyEEyA78U
XMD+8fMN7HK11VPv31uh6D5jSf1qdVXTU/61LkoGlakIzalpujRMqB+1sFgD+hFv
bEj3Ao1uamAejiBHI/ShUVPETK9zFYTwuCI32lC76mcawAdlkXXQSZw2L1Zz1/AB
XCRXOHIw90EX4m5bTlCVPMVC5plGGVj+p+aJwUFA+lecHT1YjNsbW889SQUqXGOX
M15hODV5n8myTGmPSiRF3Vnri48qW/UNnkUXc9qKCyDUqRKrxWPaU2bkTLe/TcaY
S6VMSwANddpX5jll+QKRhBDZd1qRD5gSjZ+lPxWgHRkjKUUzQtfGReLRul71gyBf
Lu1gKJ2R91wWA37SI3w7dPsnT/JkXfhWdhhl9ycaM+czha/Q1qtpcBjW+m8ecIMU
GWaM2k8Fbt4naZx+lM+zPodskjKI8xQ5by5/p638fFXvnGommPQD9u4XiEOg9z9P
2+VMvOPcbNI1ZkxI72OqRGtzqWYTGrZcKjb+99uVbGuW+pQsfVuGKe4R7LsKy2UZ
Loh7K+pO7Ebk20ZZ17+ueLpqPFCNTZVKdfMWtggIQaiA+qBiFBvwAHwIHV0uuPdv
ebaXkxTPijbh2SXZCRCxRBUk316r5cd7O4obDOnw+11ygGliaUFnpdl8Dzd6ZIRJ
pv8k9PGl6hpYLRbLl2JMANAAyHM4+PEPFZqolokUbiYj99V/vdGqHDACpac8aSAh
lPSgzhtHv9awbyiONYzDn5dsGxFj7zqxr263wp9q/kD4tUodob7SeaIeEl/MDsKd
juR5T4LslvedbfhZOIwfEciSZaatYbwTqHvQm9mVQMYY0lp0kNQ10Q8W71RL1YKx
byp45fmLpNgyOOezIqRyDxqXPmX6fyiwWeTMnvMfKdMdxnGreDZvyi8QO6YMYLON
LN0IAWMI68wZSz80FjqX1GD6b/EGNIa4/7zwfmw3bO1P96AwOHsmkuPh1U7jXCt1
g0CfLotgyeR0D5b8E4FenMgjVz5bJKcFwH7YBu+81kDKroTJaPHgTnhNaDPRdIv/
M5Q9E4sxuTyMoXv00vXA8LZleruSYcCkkGM6NwxbxeNrbKO8NURmRd6S791E9tDa
k222sD5uf87+PSZVmV/73LkEdVDUH9Hq1JyPLAXgmXSQC83LO9N+oQ1TmyQ9q9dZ
Pa27obMRlqxyqZaLL6sOTlaQAZ/0y5O0lrsv7BIkzWribxJxAhISfQ3GbrMwulGz
n4h5dT2l72JBq/Iogn72Y8du3dDCZ1Ds7UhrdG1GlAwcmXwaEAZFk46Tqmb0+hkU
MqUl0rJgUzO5eCXa1ABTEkpd9oeSK5olzWPSImSmFIDHO/8H8kBK3Lg3QxmZLB/L
iqyVpXBnT4F2ob76QmEOeloHr6RHWq7aHPNQe1EGjYzimys5tWaQBQM9Sdd3+K3U
THMGOeF2otz0bitVQaNrmk51VMJuQkif2ReQ5FGRxaN+ybr6DMyotDt8iuMALYSb
NP4EaopWqZkiEvq+Q8WtnPUxJeuBy0mBeJ2UjSdNBrIfCAQDFDxZi+rj5eJnplpM
Wuf3pH81e1j0cIxKkgaU/pe4p333qhegQyIaBmUJfYla/OwoUNh36+202LLX6zCt
aMe9fmMb7hawwEX5InNAz4RioIuQz1PfszK4ruiF/C3lPJZxFnvAxvtW73gg2+9q
VMaapPMjidqrEI17KITGyNsvViqGr5zzrF5xXEAD5ugJVu/BcHvZ7fGL643U1KAq
nGlHcp4e3sIyP+YVqXgW38xurMq5oqZGubECLnhnQQ60i7CluCiTlp4ZeslFQEpm
NEgfBNm2XD4XW1Tu/dYb0NIasaLSSwCG8hQssyM7ZgrnOFWrqtB1CCI2vAsyvx8N
FVieM/VORrVh/xYXdtIYu2mH1JLrrVfuRkm2YCqCEMM9+w+NfkaUAlqC8w3c1rtB
zia4ePLhbd3XL2pKiZhLH1rKz2TRcw9pttAAqGcQKsHg/0KQJaq1YDpdwrviNDl+
vw0oeDA9xWOaxlY7tQGDrjnUEOz+qdXfBlo140n2zleKAe2L8kh5mmxw9Lm3YzGu
ANAQBmV5z1h4Nq8H0x+RukMCL4/TpLnp96C8bb7lP5cDDAgi99bCC8MTBsvIFW91
n+nSP/6qE6bj7PpwkfGtujhFkoAZRGlwmSwONma8Y647a8ML6kXYgmNpsVpmHsAP
xpFmwIctWra+YYP4XcFXpdvnzTM5h7Iprztg6kkfN+H9nR/9APLw1wOEIytzP8w/
jtNVOODzWaQfHQb0IJOsGQwaQkIgje9Zmv5/P5vPlrBK78RbfbxDR+pjBjz2xSU1
uMjsMvmdvQlfl4VR6lp3KbAStLUMK5KGqtsvPu+t+CUehLCY195Bc+cJO2AxAV/X
Z/JRAcEukzCGITHMBFghcHJOEUxKJ6YBOasvgrz2vI8BhfpQS9yzObJVvXlB8z5z
im1Ur/6764vA5fUizCFLdtEAgPcV+kwwSTt+VfWbi7Xv1GxAfTNt9SLIuRqo3iQf
jm1QUq3p6VQDIMTg1+FKsNZXD0MYF+5QVH9MzOMxd+SWqIMHbIiiI/IN4ba8GwBi
iex/S4JqG62QV+sAPtesyC+CMGcuawuLBbwJZghffklUuXfSxFxBASUpLOUISOr8
RawUIh1IqkUSzZOe2jOrOUyws/0ab0vNM9oZu7oT5G4fZxk9u70Xoq24W5BtQ8as
kfrTAXbqfpIrIB41A0GisxEmQjaSNPvKKh4NHc578vmU0lVAlSTj+PoWNtInE00s
w4830oCDlVJE8A+GRAUGiM9sUc92N+y3wlMUgnVHmCV7DHIbsgE62vUq9pBgwczs
ExLHKq/Y+f4zNUimdGwA3XQzLneusHTnMGihm87+WSH7dUs8wGeDRxUxf9m0ubcA
f4QY9LhyYBzzUwlvl3yjlWdSnqt4kCUCOlYg9iM/PqjtLkW/tlGyVH1SxHV+zeR5
hKx8rHWwrAwXQvyba8X0Pz0niZFFPldP/da1PdCIsq2PqeuDrQaDz9O9NOS8YzdO
7MCq6e5dGVTmsACSoBS0UNwSXIIZJdHuKTv7Oed+lCgglAEsTIXrY1M3XswAujYx
vMJVWKdU5cqUclkR0yKiFVx9KKu8HVB2ErDQJLhtcGb4Yi85q1yPTGwwCWyWeNCE
8KtJZJL6USaSJTlPd1oPWmydu281JHWdN6nnuSH8uaEPr1r7d3SOGKHG6WE8Y+9Q
KIjjeQ/Gn+PAXbCA5tUTpSEMy4m/SOc/5cjJeQOJMLKmr3OUsCb8uLUNaq9TIgOj
pmGvTwnTCpknQxdnyQjvDUrx1yIBJ7j/UsCXKVJutEvn1wv0geliRBgZjOKcTKW/
tWbpANrUsMT+hcYWrx4ACHdTHTBlj0AYmr4JCaJUDCyvBFK6W5ogfFh+7aGQQpi5
t3mpQ8rOR8y4gNg03sTuL1Z2rCihb6gfKzP15G2xOwvbe5uPtUpJvBGDCmoHnQpx
S+bwqlbKt/loFTIOHLc6GHP/J3vTDEvOL0+OYMmAnrneghqPtFibvQmSNd4QHWCT
tZsQGxqAzVg+LMWgA1YZSedbukyzjwoMaBWjdtfPujPVrW5jp6EqnJttUF4YHOgH
T0x48o0fJoIiNCf6FxKN2CmkojZa4bMZ/tEIV8iW/2sYMTCuv4b+BogGWBqFboIV
Gh6Nh+hE/jBdy0TskeEP9E71Locp01xiVgtg45zztib8HgsblGq6BDpCMJGJ4KMW
Y9wP2tJNDPPN7McuSqo57/TPw/hF0GpiUgcBUFZnvCtps/sNwxGOYZpFWrg7MHos
XNSPsPvNQs1ZnTybZeQ5TxEsR8iqfKsosalB+FBLAbzdYUxV3dMyzW+DIFPZL26j
814pkpMyYo4Yo11hDPU8lIBp9f9i12QFgp7+NS2zpORJ9vZyDMzXzp9trSxRFxNd
0bb5vIXVBwpdiTAOZqccX1JB8rTuDC8PeQGIcWH/Wkd8p9Qojg7/CLRw19ZZpiBA
FjPpUCMbQIgM/q6USaKX9/AKY5R2MQiYUvAYo9kjr2KYlyKLkutmqjHx7RDkjzo1
4GR7RNZuCbd2HPJzoCAVmt1KdEbdbRkVbLcoR6zelTy4J460D2zupGTTaxLpVVNF
DcGHOaU1hyFriYCOXw+PNSzO1BBCjoXMIyjoasZjbrEkkrB+/h7LWTZcjG0xg87z
GbztjJW4meB4CbmS83mtRAT9hGZdiSycwsl4FBy48EagFizPMmQUz/EFnov8qltd
tVFKGZud2VLIxb7R1FsSyxM/6aeMAvn92pXuqjBsj6dhmQeSl6FmFUJ/nq4ETm59
WtRN602oEsZSl2DiaoWtw2WPcEbNGW8TqnpWcLkmZwc+u5junXDnSO1b3bFuaoWI
D+2fK5bneZRZ7KGHusrOfINPySj9yK6rMZlo0Nzl/jC+I9Z1CyvcRcJOUWtiqoj3
yPdJG7I9s8Bqi7COpJs0HxIdzOeylL11F/HpsPLxg8LOkO+ISU6aBa3wsxABny4s
mSYdhORHQCiV00mqFDRGf3pwvN3uiEDT3G5tzWVnpcrzhIMcUsDfu4XFzA3Ix8lP
7Xg72IJ3bZOXMylCf9fq+pNvlDjPNCCrhlu3dM8m5oLnXXb/+W6GZ7sHNSHYoKxm
fvxCCcGQnjnyvDIKXpyuqcCMKGu4ruQ+epu5yLVFNUvLaWAqiVOMdm7Gm5Re1vEy
0nl10/+ULQ8Md5RrowtlC31LAU8zriJjrzhq1TibcdM+IfAm6W06L44ImPKi+zd2
fptGvXpkSBVtwndT0A+EC3IJ+E9il54SLekraSdIsqMyNEFnAsMyaQdZ5lohOhwi
+CaNgZVJmGiqwtMASn7IO40Ffczg4sOqfeDcK8Wwwp7chaQh/G6vAPLK/a3eCfKU
5KHMy0BzcVtgwOv+fwORDllMCbevo1xhdZm4OuunAlvPGNnNlJJqHETaYZfB0s6b
YF42ZdnOqi2lRxSCVAUNd8519uBg/xyMJs4xu8L80V1pQZGLxl+RoFa71/04DcHv
kc2TPQlQ9MLUihbl3iPplhRQID8Z7INuNDnmmQbJBNUNHu1UST4Ucnq+spTgsmt2
UTYinlaCiuWvQJReVWfv5zAexSkTD56SnOpz/qHLgB627vTBnLkyNOpLBpqFqTA5
XwZOXO8hLLDd8DW7oM/2jGe6emudR5Sza4IKMH3UcAPgUmVETvl946roWd6dfglh
Un12r3BBZ9/7jhyr8OFaHn9VmJrud+xw3paTqoV1TBrY3Kmm+NksUPMI6g1vBylM
eyZ/xQOhQ0Pw18Pil713hcfASL+lHdMirA1oBRhWKzZCDr1qxpNJ9PkfinHbO7mT
cQnnEPd9J21OR7IzYmCxFSZ2LP+dWVKazpag2DSA1E2MHCYeJbt6ANPJj8WO1gVm
TS4cVlgLi55XIj+UotEpaDzJzmj+8AmRRwItFuzHS9miPchkvKUVjSyduPEkSEuf
CwTQnaUBmE+R19a/vbgbYbygpO9r1uZPEqtWvXfKyFbDTvcKW3OL1NmYVyuQ9pWk
+4XO/OxTXZ7Ks7ZyINu/+i5/gnYUePgBxAFKSwckiIncN2K8yzj9jBk4oX9mMRe3
dkC0ZcijGGoWFoe+jk2usM+tDPgFLA6u56iu6bL5gDUZ/CwUpq1ukSuxb1aw3aWV
BJal30/6zw4hQ3+1Bl1jz8IgAtYBuAcD40DBLgNsJIWX6WuoiKQOosCMAa1dwxxU
onn9HHFlwNoib55AIAAcH+CBu1fHnjJmNx/oST8AMIS/qPL8ZuN2MHqpLKjFOICG
f0i7JSt2lQWb7xdg2O2tfVx9440hquuyJZOwS+4k7YlMxWhiGPsCiAEwD4581gym
T89Hl+RYL9LO6vKxCN3vIETCQjTFi99PledT47dD/a3uJq24tHpiYwL6higxkJ0c
5/MlUhOsyQ6XzqUXQbl8LYVtNw1WOUa2Lj4S3BUvYVIlyagkivar2AQ/0i9Gxua2
OCpx828aSmSPFJoOeS/q9Dr9QjJl1OFkWfx6RvKSgZCXlJnB+EApeEbfTH7ZO6Y4
3PM7HNv1j5DAZU5ir32N/QvCwyIt9wZvpiUqXtiPi5bGZOaNjtjHoj61SiqBt0Bj
yKSh6EDp2r42hyyIRMKAB27VDlj8cPBLAiuZgin8CkP50+59kb9BSRatKZ7I5hOF
NCBJctyyHMMOHo3rmxErUA49sDnkJPZed83eoFSMYieaqe5niSR9p6HAtefagxvr
arL82Z8sJ2/4IgixdWnzbAhYEgHugjzBGlUdFKOe0moBYtur9dDkja8A6P96mfHY
NqTU9Uz/nFkpKPN6mTAYiYlF9+3H+dixBXvOsFZ2J7cwG2oKqa7Pk6ezdcv18+Cx
e1+dmC/Q4w3wukWOkJI0I7JGC01M2ZtWQesOVcYL9M+AqQOe7H5Df+rBAJIW5Kkf
ggnBVg9Vmic2mG8zLBWDZOYhZZpcoSUgOwppLFlwYWQsMTE3FPD5T/YZjqY8MD0A
bO3egTuQEwGevmMcI/pY/yJ95UwMiW7w6Mf8MudK12c11+t6MXo+/vioxIBbzjMU
E98HonZfNhZq7UISFjbhlBxo4a/5TehB34FZeM4TfjR1s07jko+14j+XCD0h4BVP
3POAl0asektNZo3QU3TL6R8c68oBpnzi2jAHj7HwG9YWSKjebe71yRWhUaMTqwQr
icj/nF6T+w1dM+9EuT+bOcCsCekZPxE8qhpXYpzJifjtQ07CUSenCPcz5thvEfKL
Lj56VZb6m9kH7yhdLmyk8uaqYoqaZNXx7PPuoWpsaMdEbdJLj7yvqiHsikmZ3BSA
yR0EM5YRk/9VtT09Q6hMf8sm/+m9MK6dDrtUo4vumH2y33HMBTDjLl3bFbhW+boI
sK1yzsbDx7FKmc7L5FVaX/8zZlcJWBiPnHOCcPVoCibS9x7Up1BuWUqs7dJtRyxB
SZorMC3e+RLHb0e+Kd2MWwP2djb9gYsG2LMj4nvcKM2EuPHrW6VBXgcWHBUPKmBl
GDsE/rUZ28urQUPx/NdA/eJd33Irq8HdYvEfJw/C75zaNB0WGCWzaXdt/sgh1/D8
1hCO2r0hSWpP+f3L1RILwv40GR61pn8EmYZ5vXyFCxS51VF0Zr9zgSD2R9viz7rD
GApL+oehs8osGX9wJcn4yKEua+ohj2xd4m43vrXO94EZapo55zNolq3kGHZqi+sY
6j5ke3VXK33uSZrDkPLMuW2RhKgVllhGQJZljoJObPiWzKL6mSRpFfm13cZQ1b3z
0KTFK7kpXnyJx3BNW9HE+S86Cpdp/t6jIFyTjHK0NGxoT7Neb60bxwDZZuU3FA6N
yvO/sivvwD7TuAm44KgONjBRb5orbc6D6sYRdQxuab7lFXthjP8foIYSlkMIcmyT
f9P8R1k4xt3IvQcfrteIcQxU5timEg1KYcY/uVK8sU6bQnO0275r6h5l74znJ59a
5vGZzlfmoNcV2EXKB7MHO+jmglf63ww/8lB9k1wRxcUkRD0V+AE93Ljoxi4TORrt
cx97rTCxFTwkyTmdwj3XvkSh0LAmXQeiZkYsFsNW+oXUfpVPwMK8isX7UZnXVKMo
uiHrp3T8Wzli/eAsHOOnu9773dlHG7nBcCjOiOWWhDBeLz7Cu+6LMc6z+yTj3bK4
aJnWSICnasAPCcatPk9NEpAf4FV3c7LP5QleilgtTo2UfnDB6fEumtwafnbdk8w+
JadCEXJ77kX702QN9N2bJ2G1Ql5SWnz6QxpNitvN35ub1V+9ThWc/ySFboXZc5sI
/7eiVyoYJMs1mf58OU7ZXPpd8spBYJlHYoWtec6qZHCP89zYkyrcr7nx6HeG8Wkm
v4mUz7vf3rNEb7J48LqrMFKt5gYDLpWV+cGTdd9K4Kva8eZLQpkGHHZChhqseUjb
P79gtVRks0V2ALYs8mh+bF/f91vmeR+JVDpZZnGvt6nlvJyISay6SWWzOQHSuagt
Pyw3oyWh3hsT0NFopoyubqmoKBpPCexuP80RuKPp4vmiAQMfRJtmFN3M/yKHuhpI
MT7ctW3s+AQppxIdOzle9lRIIbm/IzuVjVVpE4aO5fDaSODkHzuofxkKKRGoXbDt
ad4l9N5iusCQFgVDdElv9ZqOqO3XtVL3lKDYIEYujLq7i4k2BLpYmrCr6KQd/z50
YBggb/adJQZ5Gnnng0PDuF1Snuy3ZwbVEsV+ZMBWVRZdwtaMLxlwobOy30QVKupp
HTkNcuT/cpkHjN5lSJfnA8yYMRWdJmhjMLtn0R1kbgOoCI7dz8NuX6CESM1dk54s
ZxFMIzBwRG6IK4XHwUfkVRQDPlWawtOHZCuEUgLNfw9x3Nz7qNNYmWgl0gSJy8Ig
88YB0cGSkUB70++wx5nDr7/ZNajoLu/N2qyneAu4Zjw5We6fv03Ykw/F7XPngUGp
A4ohRob0aXdl4BSc5Uihdkpfy/FL5X1TQy0Exxq9caCltSZte0nQv+bvJLzHnWHX
9WHV7fJvo+A0gf+7ci0yExeLdaS4b6GOx00HSWiQi7uz3ZvpivmRuF4BdXSSAplF
yIpkM7POxe8zGDsPDgFp0cIg7LQvi34VyJocCPgDDr06oZ11mQj7t2UX7yMRli7q
O2Ya13bUbXyX/xizgteQ+/gCTZi5WP0a5PqiUDqSkU3iJIfwf0j9vcjj4rn5oih+
Y6C2CMAcd6T1RdJ9qIVfSttJEtdFwNXoz6ySu1kZSaRIlc2bBj1CXxxQqGBGIJBg
IB32wMw/YhZRe2S1lA5o/9ytPEAflfH90pdexob0L2osRyWDq2//HVzsHsQyWsPF
3NqQaWQ5TYZwBeq2unVL7uYzaG+HBHLmYaCMAEFiJRct1yskWFtGSHii1PQOL2D3
KAl/wCmo55wtn0BPwHKUpRkXdyUlhDw4FxMXexbFXbBkTiQhIkY2qIBpCcesLJOI
3MaVRw4hEOT2HihDLdIMheGZ9dzZWfzILr+u7mjtDriWUk+A+dzmZfEir2d5F9xX
/0IaNXdE6M//dIVlarr6s8Gxn4bDefUCG2Li5jXmGDEYfTl8x+VNnvSqopc7q/QU
gQI+26BsC7cQKzwz5sM20cKijry5qcn+yDTyY/CacUs63lSgf0L1BfuBndVRv8Tl
MF3LjqcoWTP1AFwllbHhUMrxW+1FcCgZS59JzU2Z10MBUWAp7Nuh5aMIX/UvekNm
5yVIBdVuWbUcgtRaUKKNfxXArSTnkEg2xLfjI3GuxUOsNDrOnCrNTv/RLJoHVHU3
IZmYEPcQzda8AfoMl3KLONHh5cKcayu2tkXwspMH3bgpJUDtzACUrH0UQ85Hu5TA
fhtLNIrzfUx0nujjCCkEQCSXsHexsmZSu9jGMS/Rq7SBWs0jb6FK4ktCfkc0sGS6
i6swu7lEoHwqdE0pDDOLPOppUvIjp7KPyWvwqi5vuV4HAM+1rqLFviAf6Ly9LJkM
qIU20MaPlC4mmeU7NqKZsB9kBPZdZG5AoHXXM05jtRgeaca8s1qo0LevHKTOq+Fz
U6HP7D5QSVksQXnf0+oLPEez7YPuxIx7iPPwh9u8ZPKYOTdYt0rBfYEjn/6ED2Ja
Y4aq1zJiS1H0Go3BLNqJiiji/DXnOdooSldkPDdd9m7MnZWIdc71IiW0NSB2w/tI
0NXT+PZUuvvXcrxlDIYd9mSNEzxo7P9Njrvq8b0cckJPoiv6+Msu4JTnWhmbtfYU
W98AWclaUruVkXupE9ahSobeGpoOGBTYHOmlGiH8qoZ//flmVtQ8BZZFVPJC5VCU
Tacudnniewj1ByOw4vCpMWTChdFj424xiivKZG70N4NTtJkHyGiJRCZCZM82vwkM
r6Ue8r5Z5Ic36jFtyVuWyH2LqAvkT+qZE/5VH6+bNz9LT1LE4sYDb1ZQcFz9hpQ3
hX48fyxKEfl/IggsUByhNw51Cz5GOkKj6XiYOJmvUJVGmQho4Z3LXMvsH6KwSXDn
7rMOlvv2Ek3Yqldf9eGQPa/8JYvOgMgSRJx+MHYt5bjY0xxUbWx5YEs8CEbt9HTd
XzX+QZN3Wfe0zhrSqDSIRwcy0qrW7ZGuUqwbIFkig70xF0THKDD0ADmOhapTknCf
p0w350vTMz4y09jGiVa7Jrf/AHF6Yq/66p5CNWtQK17n4+nrZWuTt7QVbU9q6e6k
SjdJFCQeEPIKbZIPkDvyZ18a0kt8rsuPpjrJwLZbAtzFowEMPOZ2JS+WYtQ80hDc
5L3V8JHxq63tH1GlJ02ka2QEYi42mMessMkQPlfR4Ne72nD9Zq7m/x9JWGif+QZh
k+iQm2a1+ipkd2gn6D1a3uW8jl0Tzj2Qoa6DuFDxB4iegtOfE+/ehVrH0fT7R3Qa
Ect/LmLR2XPZgHXvY/QhPQBHD5vrf6At8KjNAUtOFlVcMTxZBXxEIeVkRJMhfzmg
bkdVnbsnLKuVi5VnhfHAoswAXjw2WQCnRkyyVT1sPHJ0UD5JlKovGcJH9ElR3OHM
tQifaAO2sg/Z0gAF6Zyz7FIWsP7dlxkD8uM3sujdoYfPTie79LD4C6p7yKtEP6wY
DA7BW3QL/3uIUpl6M5DYQ+fjcumxi+PJ4GevVo2tw1id1bPshfQYIKArALVzdSX4
UnINKaMSsriqY/FWwUupHDEsVNmOhqBn84meAJBhTNKKbOLTCpoUvPW9V5l9fYjf
5zK1pImHgSIyH6gj/AdPugavX3ayDyDssI/baHAgRpZTrSHhTafpmV0zNU/0JYX9
m3Z+KtSzKJ3khCJrD+OqO1mtATll3g/lC9KYSgxyAM+seFS2O/xHPza1Cc6ZNJef
SfEzyCYy9ErfxsIVKa+OojMbzwzpI4d0bzEJpFNCDBdzSQwFYORIz78QivR8I/nx
8m4+mMGMhSrT7tZnp0S0HXmDRY/BpMDAt9HW/3xXD0TIFCrX8AcdTLOSQS49vRkR
HzN9Q518oP3zpy4DpAPX2ihvqNZxKusoHtvW3DBONxH7A2bHstbOrzE9Gpdxt7BO
Nz1f7FJfClVVNwfvggTq1ITbL+DL/txNNgTQqIXFrOq5LyGLEPj4tb3f0Dby/Pvn
Qfi6x/Htnqv6c7l1+avrSxiRtXl6zkOWSbAucligC/mPb47ZWjzmg9fokZX9KQx2
DG3ldPk3W3K+N+XV68sQLv6wUqK0m3uAjRyNHO4Lp5XwQ20wpimjhCnPp45w7M1N
S3MdISZ/VpozcsqzCI9JGfVwpqzddATII4ru1fnA7BzmhF38BxrkFSv/5q2CSu9x
PaZJhAefi8Nap+y5/8BWQsgfMRSLA1QNUtRHDyvbiqiF5ocEYhkm3QENez95K8Di
suBhZXL+anp7R9gD5j3j4AlKfT3/rAK16asD+d+3cg826H1Pe8vJbJazWEpT4aHd
jTjis+MiQGahZpUUP+pzyHnBiYR+wZCSGrfnLM9YP0pn05TLqyuHNycfLikv0Vh4
evsQm1YCoGDbY91y5J8WD/9/UQ9tPsvQc2t3iZsArP6URkUkbqy4zRJzOiJSlhAV
c+8g86zXGLby31ueS48cxrpmIeSeGBM7E9QvT6/zxpnOaIG/Q+o5c2n2dCWJfzdg
TNMeZRWGK3KpIh1ZX6s+hFIflslRsz4CgAKOoEFRRqgIgFE2WKbbQUqNZw0//Xsx
dv5U+G/mihfdkDSGM0HLqqcIu5xoGIEZeE9CIkMjOIvZ/7rDKvb8O75zW1A+/1Og
p/hlxGGaq6lxKs4pBZwiygALubFAXCr8lIC5SaEkoCmufNhn7U0E5EZSlMEnQ50J
tOMhSy2De1Zvbz1Zsv1Nabpb6C1aFcY2GlgF0f1X0I9Mj6CeT7D80R1NkL6p4qCP
UzMCrxyLyXA7lIihziN0Zaxm9GdeO2BCQpBDc06oD4sCgjWoQDaDk0qTPBsSLA3j
2x4dlGqlCi0AOzB+LS19pRSJRykUps4PWdruZ7g6Rx6fi/CUqEVvBoMgIzO/w0Ub
RIE6OrWx7Z8RZkA//9okTltf4ujuj5UdjcQSmBFEXGyp+p2Km4kpSY64WKWG3AFy
yNHFKA9zsUnETjIWzikPzsREYpBJ7mihdg32vDRQP1pYmRl3gjNTKRV3untBcMfd
nInYPSfpKm6YUREOLQZjchywdnZMJn/ZpOMSk4Hm8oWmA2xMbHH/HFm8W84ieiRL
1Z0/og1ZTJkmG6kwYklX6/cyMR95qc9W1bymAJKE2QIEOE7TC7pC+gjEmR8SeGo0
BlPBH8NYDNDPwWemuzZaEjBVKNwnEQEFc9gbcekYfZ+xARkjWzZLphveaMLfVHWG
f6CVd/Xy/w4uAL2P0GEqlE9gsBYyeg/EVSJAUHzY3vZP5f5Minth6YA9bpsNicnk
JWCrRoYZpN8U71TdVQSEUkdjOWTeVWdZ9t8KbaTvKjGA1nkXTC0Kawwin3dNICVF
R8Kz1NMt5SlP9rdywNDjaBR5jhsoyuboeRqnorgdbjM04CQ+QH9uB2/Q/5lOVdRX
35FiUZgD6qZScgRnFaU5fImXrVIGkHnN66/XK78PcnTUETWCeAe5I/97hgFAvVjM
nuUhdq+c+itNaGDAkuYQflsNAeiaFqmOBP5taTQZij0ut63/yVvj6VC5WvqMoqfO
ZPoaZUM23hhV+J/XSBTbRJl37x/sHNb9CN75BG2ZVHBm7cRzfiCeBq3pQ9PCeeaF
oOsnLWFaLqYsBKZpD98+jMDD2KgQYFslNzF18RilaZX9hjINddQo7kxzwrysw0+4
hZfYMDAMcntuRYMdI1hjltAyog4UfzsmBVrGUQuWEApVqyj4qnHM99CrGc4TCOve
4LYWSGuo46M9fyZcANdEay+88zGJ6IBEOwjisDPG+ZRlVivksVOLqKiAqIbARLPW
dfZ/SK/Xul/XrxL0Ax43r6/R4izVJJOMDBfMxOQC3o8JKH2qc42gDXB8zeOrfPBJ
`pragma protect end_protected
