// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
E0Fj/Vd28I5eFcfSYIGE1xuOO2HpBHVb6IoCGIWPpzFsKKnYmmb6xTqwOqiy4g8ac6Of1SoRFv9U
4ANM/pLRV4kS8xEbEBeoyUjKBH6gpsUcAZh0ZB8XUBrKhSQmSdbYesDgzliU8FBbHeL5QcBemitx
PKtO1USjHwWLxml/AaKmFhe2bAsPTjGiPwLCkifbUVJM53LyW7K0OP8TC78lWk7mdu//Dpl6ktyG
FNLBlbklrkADqL0rHm+KX+g4xWaQ+j3pFTdSvg1wQg++cgmc2QQCjA3COFQqar7czZUDs9E4bSI1
gSaQ/4+DsugHCVgwyC209WueuPdI0NWHCHMawg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
nE4porPgi3SoQhhyyoP2wb1rgQE5lhonBc2dfrYvWLFV2Tb5K5ZXz4BWGi7lj519zj1j8FACPAgp
H0yA9t+jqvsy3uw4oP0tb9aY8WzNaQJFVBqKaQAMW/voFusvoKJ8knJnZFhW6m+YlxGU8V0+UqbP
J624U619Y1w5Sx7ogCCIM6otLkL4ffVqi4Pbj/2trj8XBBNpcvtnuaoH8xd9szTlUrbtVwpaRq1v
Z8dMSaLv0jsuh2Bx3I783y6a/6L4XOOXFwg53ZxK5OjI13XrjOAJZ/3FlB2NBnTQDJ/fWuLy2i3o
J3MH2s5Bd9TgqPqQxk0cw2HN5XV2d1T4uB5q0g7SSs1YHCgXs5khU/Qo8dQQrNoELcPN+sdDxU9V
NQ1ZDAF+egMJs9JLeluEPircgRcGtjTtCtka3/vlpPhRy74R83vmUyw+dh9k7WfvgzUiYof5Hktr
X4op6Hr85oudVZs5MKaiYAMboUiism67lJ3MVs8WvZ+4qUCQBDzqGTHaClzlsDtklrjARSePerUH
USF5TjqUuBKJkEsrsfO1s7kiYH9mjcWqxNC1YnLz3wEIeR/FHO1ZmjRgh6cMzX/012Uvp/3lbnLl
i+36zPI0RSxsfleipI+Aw1xSn7SUOdBXQAlgvfu3up/9SZBxX1pj5dmLE5bKJDHZEK/okq/9aGwQ
l2NG9YoQqB1lrExoAHUb0voXjBhlPEglpA0m++Si0kV4lGGMxySbegiUTghtM94damv7ozz+AzSf
DqODUpHFo7dFrgCpe4RQowh5+xv2l8flqEpKzkzuSrvK5HhadmmkYEx7fbxj+Bb0r4qJaNyTp9hJ
RQygNr9TLyhVJj9Sg9MKOiT0/I95+6dZzMXPFgQi2JOrPoe1PBCveARz6lK7GmCSgkEpFrFLju54
Fx+sKCKeWigyjsZP4bWjeUD9kbjo5keUdsS2bTGRYXbDQBa1HGX+4HNe0Z+ORyOCchgAPZRNUOS9
ziddrSP4Y/vWtmiLas1CH5yi3yHnJ/lcCmX3V/o6d5GjBeJNm0HJl1jSnL+dR5FXjiVYtnWJ7DQr
/ANZ08f7tuIf8pRdJeUMgEHgvtK4PGTJ+Vk1cMkIHdFxwlgeUKU8KRA0aPQlk/Q126LwvCbXIabR
O9ucXvjEIdeSjLgFXZLQQNFd2fHqD5jmfuwslPhv3TypWYuOgU7QImhDnBNrXV+YeQpFo+I9q52G
AmLW5lGyA2WiAO0YzOZOlAOT86pWY4osoejvgDR+RWv1VDmY1u5J4UihcKHntPZ2jtALjeCf4NuC
ioqizZjaJLdR5rPUsz+Ao/8C0a0cPZERCvpySxcALegT48+MybQpojTLFztsOhbiIIKb0aHX/Qh2
jJ9SrjqUJsMUSAjYUIjoj1CE7Wad4gD6Ofx45zlCDKPijzuzVJTNlZYIhjgG4nq3VFLw1KzPeJqc
u4/TJvyo5e5nhZ4ZJPfMzjjIXluaylB/Ix6CVtoXLH+r/2NpupIi54k9hb1tEI63JrBM5Xi0g7zE
5zkiUqlDD4y6DKS6/25jEV0U15TgeZe52hl2Ifuz/F2kTr20163RvhtXG06/c6dhhILSsrnTtIiA
j65aLIKOx1rZSO+r+J9u8uMhealpjfH6zClVuvcVoQ+8266nAGQAG1Dt0sP6YpDtgUycMtej4zME
IDFyapfOiWKY9ZXd0LEiccC1q4TT3EMk4lacFFfxUb4udfdYT39L2FKLT6/sg1fMWqnn5BGVRW0L
HuN6AmmgjbN1lZtSqGfcoafJe9eA7t2Ex5hb1l7V3bAgCHsupadarLMcYAZkb7mm5OhbU37isRps
iN4ADliav4ahtgZj3DtnstUzjepbgSiiuPQa6nn4K44fKJgzuyjkW7mnizEJzZKdW4PJWq4RshWS
glI9ENPtBH+6jOzMlnCAPXPBHeZYV6o5ucyUHwsYXzLDdJbGxhet5nCzVu4BOsgKGa14U3Lqqbs7
Mlg7+ILYw9LOisclnH/FBOHfdzXqKk4g/dRapqvp1YOygVWqlGSBDwBiCpr8WJxQhhPgQmeJDXH+
zB5INjdW3q5lEPAuEPRSuQ+f2K257Mr9drIqWR1cVC+9WI9PICjbKKd3dVj5G5SnrJczGpXpVjAS
SxTaBDgA9ItsCO94eq7n+obsjJ2AvGs/B4mKPPIrG2LqUZGbMiZW0ESaKHsylzrPq7VOJY0Au4Fv
uAUESnyaoMRi1fdf9SqvGLBgpOpYSjUOJFlUYV6FooNh7Jq2BurM6mgvjzFi1Y+JTPilX7dXfaB3
18oai9b1kIKSpb/beoYQ4XWbglMzeUPWCaGYvxdl6kGK5DBymoDQLZUbRCwKkPy8m3khMS0W3oRZ
jq6zX5e8Fuzw8UuqtkI6uNZKZfE0SwAroYpa3djYnWSwiL4GyHKG6CMbqhYNTpPk49UpvRRflyTf
XEUDDQAbhYbCPaxTlAbyFwlfEpfTBKj5KxqmenkBghWNACtwRnhcncE1TGYLifesqRic6VZBcrg/
n4ifXWA7FXmiqlxKYwkWK7H0kdAiTuHjMpGOxCeodVbKuJwENk+PC81ThVMKo86BMwguhmlqhHVY
A4JqxFTkHvheZlxCsy58oZ+9ip0lCyyTkAr6bPKEbYIZBYDmuy8b8jw8ok0TrCdTp9HlkNk44T/9
10W8mlwuYfpNb93xfHk8DBWD3teuKD9PnR41vRgAxVYXv9iKfFLdR7dfzMceYJNjzIgy55fgDBlh
XGTugszkrKhwj+z8IBDZ2qLsl8xr63dMogRIQGuAgnAicmSVoxsVoA9bOKXfGroIF4MKOE1h2ibe
ORBSbay8QDidJjB7yr31+ErvYbxiXe7I+wAYSmYPw7VziiUkAgQ9DgtF28Cu9MRSxw3JNu4KSNiY
hPjnjaNCPI5MaL+4CINGA1xBzHHiiNTeMpV3bfqqvXIDaiEZGBnGghci/1SncO4wwcySGThUJ2C1
arRM9DI76XYlanrRzV0xy6opXEplE1v6aO8Nv0wm0HkGnq6DFHBsMxdy3No5Oi+WWLeGIPzgkM9G
7lUgdwKOKVBTSyWn2aH85Qy/dpNpDyocEiSP5Rh9pGo/tynF0KaA0irI0NagwP+xiuGvwPBkAT2l
9nj/Y5XSWzqHvQNssi3kQNNwQiRKyV4qISPawdQ3QDFXZs75l6o6Fh1oPebIV5STSl6nmKESNnYP
NhPkEma2Qwji5MfMsB66RI43vZWKI2Mgs/ZTsoj0pF90p896Qggy0I3zWNSVXK30vwbbGfuWpiTy
reUgAx1sUlzrcZLzu8mcsI2ZW3aIN+RViju5vaIaBTyggKk7tgEtn2R0iMSJTh7nPB/huTxBFRxR
La0rxEFfqtZld7XS09UiYdGcOhlmjCOwmCUTAFlE8s9YZhQG8bRvGrF0pRmqQOi88nMu8EBPzVe+
DbXppfATEOHqtqDsh4+gBrYoHxN10TomMmU+0JU0yuXyC9JfrSJ5ShiDrWZc9GyBBGkhoeLi732N
kdTqpmVIHUZt5ZZsQh4OWvc4OhdOZQP9HY6UBW4Mwl6s53fKJRoSU2GMdlqAd1eaMb+/KkPq9s/+
U01iKj/9tBc4IwHEb6Xye6OEsePWoDo0y2Hv0zd0NcAcD/VhsEcWceQbX95HRkf6538iUB/DiPR8
qteneR07qJkuj2+mMbZwG2SJ23+PhAfBYufwSaSf5N1wEqDDTL9fVKF7CgsPGL5F/vRzej6a5qfl
1JbD5veZfxH7iLW6bN1zABzJUXXZXPA4jfV1ynImty0zdaYzGxTQwZagzbO+bKhAJEsIDgR8KD7x
zqXHcjS57AyPmUMYIAeD9BnCSqt0fVTEpdoqsD8m0kxYzkqNpaZlesRmPvGqBmYCvaERo2sf7MW9
+KVN4vDip3xR3AqMKLMXBykupkNNsQM2LD+HjNNInh0rcAtpCIH4kjGakc1zZ/RjNCRRRl0925KT
sJAaRqh6L3BpuPS9aDJjU06ZxBJ/1MAjQpfY3JxPVM2c6YzxLXDvXNuPRN51iiq0kyzMEBB3ViF5
R/m3Ybz0IbR/xE1mHM8mFS9l2M6MfPq1FN/h7RSH0PeyYJLOW16vF5tPZ06vfPSCw5fZYCAWjbH6
IrN6o2ZkLPWPY1vALKm9fn6slbZ/9lpiW6lE1Sikj9jrKKasAEjsWFoIR2ovQ5FAq9Znfc6OR5jR
05/tljamDU8vvWHe7tn+Onaa3LH7k8JWwzTTlT05LRnvMrplpdb0x/4n0tuT7D0Mpfr+Rb0S0d4x
Nbsh/8m9FEGbSq/cJntGLtguOVccR0oclE+u0Ka5lqzPMeQf7IuIvVW/MFiLfDg96lfe3UOhLC0F
hUD54S7DJQPqYb0CsRrqkeI788Je67+08FXW0DQjScq5UZfNDtFqVKYCRcoXjlFhOJGSgjCt+N+U
o10E5BiFUScYf3rNTB2SuIsQ7oyz3xA0tenbo8LPOpX66atH3p9qdtRCUZp0jomKWKlqw6l29/tu
6v8yiyPhTWok96pGQRAfwLe23bdIk6nZ7XDokU/ZaeZs0IFNUNy1YWmeoTOt8MOFbEncQ5LTrG3e
icr2bln9uTYvrcYBhoRmur+nRQhZR/hh8+sjzSF6GSWCCO7+LAvJLjVTpJwotpTBVc8T3A6p+1th
7izIuufhxSnT3pN1+JFdEEwVFcPIc8zvxZaI4DtayVoRuiReJOoCEQDjWEbafbmVECWAwGju3x/3
o5/Tpw1QUb9f0L0w995bIGYIYcXDHTtIlqd/GYNIwwmN4o5RV3SJBMVGcMHNOVO516hHNgAnNgXt
ZSSnl4FuQrxBdRm7hllaHJG7G6C4kvWb7GUPEYFBvr01wLBM9nSqBTt/slqDL07Px3BhCTGOqbD4
myjr0wAwS0q/aOKzDgKvED/pp+BBUQGQ9Wpe55uso52ZB1ToAgnyj4gKgEhdJS+7xeklZ0WEKJs4
Q/c/JHf96uZnaHcuOYysGff1S5ECXb6K+bHGRpfxSOIVNzXWNmBVU66xZ/dSnm1saCHgWzRPLT9u
x8DMwqhlXb+m9DVBM2/QL2xUmM9+70+x1i0/EGbJPFjSGXae4/jPMQfwV6t5afxSnnREdfgTGuS9
qrmlvLxd5oaraTOxhVOWZ6eo0HC4wdhlstcOQ+/wJtSSzxCjsACLW/lEySt+NROLjuVz3e3vpEvk
vRF7jSplvBxCrh4ymPjtWnLG47jJx0OXOrLuayxJQVXyY0CK9qWxc4lY5oFiK42h4QZ7zUw/2rDt
MMwPdTo+w1HBr5/UubP+fEe2vtutsz9Rkcy6B1MEmW4zCwJgxmv8sq8SVVx9Uu0cPylB+DOAuYV2
YYsRSALBKX9ahj+ypUR3/z0hUfxABArhy35S3ku0ydgbx19w+RWVVru18gH9OgGoVCBLz3mAdD60
Lnn/ABEUAQ9U7FwsPhdjMbqDKkL/AvFOgClz8LLWgoT7rC/dXrsHnNuecU8WpuNkJLZf15NY8sEc
IoQkpuIVm5sncYmLlG07CKFKJWwwa0B4Qe42joOce6/3zvIm0iGxe3Gq85UrlV/T14R0Qu9102xv
eCiuTUmC3dYgvJQDWQJGwq+iAmcldBqHXLGR9TgdjdT4PLJgjtHqQkLczn/Egt/8mixG+H8qXC5W
AqF99A5RO0rt4IUfnGL7tFXjyK/ot2TZGPpmQ5veNDIdPQQU4ZTETduydkiC0iu/VJ99d+ESKIss
b54gPaukHzgOHRxtwHUT+WplefLTEePPHqtbFNKIQoQsgDubGYVrDJPov6f32ZNRnJ3Kn+5lFlHR
k0PGWCF5L6a1Q+NPSsx8knVrF8YbZakS6GvY/sIG1zOYJbc2pxDH+J5o9nZaahy/yB6fhMw2SSMN
pk4LWr3iQVpWFDjORFKjkrdYTo1CWFSpLjAemqBmTW2c55DMqh5EOaTLK8b6/GSAUKppHblm6Vvh
UUtpN4m1qNszLFNuX+A5FOp4+nUdOftqOR84KaCKdwjzxGLQy5378zbwEhykAHog+sYx+spqSSog
6DeKfNvb/Dv1U65eaGom4+4FS5KX5MG+/xyZZpI8QrIDlridewNyHk0E9femL4bh56oWcWSnQ18e
nJ3k3uR6+MvHos3nH7JTknMoqeZJqnFaPzFyXz+js7cIjg5FrUzUvUA7m0y0s5FjA6IofhYZo9Vm
umDLpkyRQiVGnbhvvgrpH3BAzwtH4HOxg8vTO7f7UsbeR3nwGx6g/GveIHJJ/jCbHKDSkKxmXvok
qK5WKRc5vxRiQBrP6UF4rETeyDDVEIXgcXIe0N02/vGZWO2HglDd2QGJ1CqAsRLpN3bD3vgJpf5o
UJ3HHWWP7VbN3hv3LaUX38dic/kpq0qdGnV1DSnWqF22o6dqV5ibY0H3nVv8JL99ybbYWXYS7DFt
OaGzQaB3KCMcPsbY7frPBPc9EBMWevmbtgokYxzus3geCivKTNH8X2de6yQRSQAbAkdflHPBBOBG
2XXvu7RhLBwXLey0phmORPqB+2vyoXruod1UifWrt1dH0tUTO1jwBL/9ju1ESCwZtwxVgUyYTd8V
bG0Dlq2NDoB7cDkFoVYWtcClfjytwHeAYCyFaqc+tVuUbKkXlERFnQO7EtJAgrLA4Q9odya1fmqQ
S0u+uCm4YlLwAw9hCjbo4a0Soq9VuoqXQPl93Yat8/EJplfW8FpCJ0S/4/l1UQcBscGclEXDJ3M6
ZImiwrZRDGMv4xEuqZNp92dtxPjmaYeqV/IYSl8GHaDlrkoBngPmx2H73QmwQ6Q2EJE2K+tCn5lp
02qHscFhhjZF4Nk7X9Z+qdDeA1uQCrdvKRcVuqoJKgpmOfPQlSYaNqWF9P00cKj16vimIOtCvmyo
fij6lAiVW1Q3l+JLOeKEl3EaxMdeBVfGJjMacNKzm+/A1Y6fStisrOj97+3nucF01+sRzhfcClUm
978oFrT7aIbPe3aCgUluVPLyhQUY31+qmE5weFip9buZACNZE8GYvOqLOt7/aPU6T12Nd4S4WCsi
rQk0Dngw3SwtmwmVEUH3IqSAX86owdQIt5ObJoAINtrZNXSQEiALHrw+S8Tqzz3QRFTSurc8akO3
ZmBSqUCZsc9Xl+tX6fQbZmlxZx8HS8MD2UggX6jjaNl1LU+c5U7T/xnDYKNTYwMRECZfszz1EBDC
4KcOd0oA0GQanzSMLlvPGsQ3KwyKzSjxIbzPaPW0Tb3OJJ2c1cVudjMRAetDfcgILvW5M/y87xQ6
wgktH1j+d3PQ8UUvhRSha3g5BbDtJdRhAsEluT1P6lvPdLNAz69rGn3K9F40c3i1RwL5GQsFfKko
A0elA2L5oA2sKM+FMk5rXIfk6hudwQ+1xulemE05v/vBLLi+H+3HjMVqcADRkY5bcJ2HeCbZih+R
0EoT9TzVV69PXlZK7RNRE8fmiOOTzrcDxsxePXR9Ap4AIeYiXpiurui1JLxADcAR2vmVp4VFar//
EX04HzpFvGTwWDm2gtXEZIIj6tz69p/9LkP7V4BclrhC6KQvSxGsxtzXtFOxEEX4eQNzbaLpSFZ5
aBU0l4lYfih7q3R+4TdyW91sDFT9LwGcN5AmzFKt6ZsdmNNfUZzqrUebriQ0Ci8Lz/z9oE1VC4PM
9s1/eP1iXiQROL49UgIh1c3WlnC1+D1bkpiBsUU+JBs5llchiZh0q92b8890nRbzggr3jdN3XKIW
c7HAaRuEmSiWFVFfWc/BhQ/Ds8Q5/7znAddTuRyj70mEcUCixsV7KMgNOTn0f7KK9n58vrD4TKcl
ykaCOSYuy8v5oTGjUj20AEkANsHeN0JW5a9PaUckRDXCOL0Tqce2Ry740cpx4X/wEoEBwZxO8elA
UpN+aMQP+hIKLz5pSTEY5BBjTGq4Gb31DDar2cSPksGPmoV7lVLWYPz8/d5MUynJFonezGIwmAiQ
B1yh7UlIskabpuoa+WHvT2NUEcc4zvtmAOWZILMaZIRRtEs3DVwKstr6Ebs5Sfx0luAQe9JX81CJ
9xGuO7pZurtnML5Aajyff9SqtsrHR0F6a0lYsu836IPDwUcbv74MNOwIQGZQgQDR3hp6PfJ4Qde+
ylRfObdpGbJvTR0JIBS0jUmkS2e4jjz5jglyUAVDK4lv8Rzm3y5qkP3licCmrOfGU/EzstSGm/uz
Y2NNY9RqGkaNDNUuNaO/HPUmtqpUgqXLdH2q1RfymtKqNa/esypR3SmxzJmIDyzQSTwWhTceLEzN
5jtFnAi8pc7OhUarX/30B+qN03UNvdagN3MSkAdmISw4qarxvet6eWRCIxg6hHpjQ0Xap0RAxE3J
l13KFTE957+oDad8tt3TzBhUCVQdUoIQYqvd89jGg1Rk5GLvonrdHLILPHEJPb6JeMPFU+tGl/R8
1DfIy1+pUGZ4kowA2IYzbiRJygN+P1iFNRq6cQJ4+3J1/D62XCHp7/an6m2CaYxWAlpg+SeBG6r8
W7JJ0atqnz3NorDWIddxa5bXj3f4/c4ZY9g7vz7rS1s9LniiuKc2WDyHVicphxuJ59WCxOSCi9QP
YxAn+BheeJOVcvoJ/j2i5PMdArS+KH1oZoNh1xB9gp2hyCyaIE0mgzoDG9gdTPYm+r45Y7KA8Sd/
WLmPSEvKF7vMuWXS6L1uczcRVghlEfs/00YrFsQ8QqWiQU7Rzwh1eyc/Rdz4AdqfOJftVyt0Q2xY
ruFF4U1hKMDAXdwPnGEsnDY5HIXhMZHJeinGuf9DjXU2JvC9e2X6FWy8YKklhcChKIeL5yX2gYzr
+FtzhfeDfzp/Jx3zRcVQmXoGCWz/1ipn8IVIEMkZwL9SrXdteMYQtPyV/koFV8UCoJjqFExFfpVW
fPS/96awtEhsdZFpe3hCIynfUinAUNOrQZgosyPj3JfeyaKjHUQ7Wpn+3fBhYQbmL/BiRzHNxJBC
e6fbD+dcCj98LWJHDEyJBAFMOSV41RyldQW5+iEGq1MPLd90hzwtStd726i5XGifDZhotaH5rgNL
gCMffGNceknQ+Rc/yK04qeSs7IIq6qLFQO+jFAfn2pXS2eOlmeJpJ5UhhFciu+gOAF6qN8uZUd+H
7aon1t7qNlkEGoENUzvpynTowUNf0hjbmDOxfnACCBFcm7T6CvnBhQ8KX4XDy53AISZyNxKsShZ0
8HrQ6YIy+6oLfrUyltnqwPk21/lPgR/gVhP5IKoGxV6zXBfhdc3Fm8IGoIJuGu5PyKXb+Cp55G1h
rTgVsl9GghX0tvxXMxjBfqcgEHXa97S606WNY/2xvI1o9iZel3Q/3Gf3eQDgFAxI1pMurfwFmfWI
rk03hpgkI+qqxwWXheslrQuDW5s2l0jTuOt7UpQHOkOO2DLFPBWNoSgO4Yr7F5WdQ9i4u9V5Ly9w
bYWTnSRPof6W9u3r4WzpF/+4CMYYoLeRT4lekUosfa8wB0DeOKRC+c4Xf9y5e/O6QIhSMV92973X
StrrGIDSECssAljlm+9TqefB/coBueGDPMriCSeJA29Mh901q8oHEP7gtH8AYp0IBO7i8Mygg+iA
vXYawMaZN2ynFuwG2pyEogRGB+zvBgtxZwWS+dT4axgiBOJgWhPIAhuVq8Tfru7KnuYcd2gxsT8o
lXQeD0Cu3w8JksEe0M4HJKyhfich/nmcfSTLC6LXEmmv9wl38W11Cf9o4j8pH6voGDkIhMTolbnr
I+ybzW+OmdjYiyKfvl+Oi0SJu/yNnklcqRVKsA3Fdlsj7y2pDf78qluzpy3jwBAzw1EwptB+6W0P
QCl/02TTnQs4GWZJNFQnkMpRqP7nMYJ6VBvgQ/I/lD03SkTPuBJle8qNE3hgqbir8xyJRe4pUYhv
ZKsv9Cqapy5rYnn9zph1JBfnJOEy9v2sSEP0zHv7iEVKV3Itr4ZLKY4VI/nQzeUKroIeau1bfGPB
tsjOGChCwDLRNFux9ivhFdvxW6Vm6wnxtWOY0gVRYIg4wyVYZ+yLpKqf++/QTAx5AU9KRCv5p6Si
halBxiqqp9M8WJX3U6xXbPbHbS0M0+i4c5DysUbP+ZDro2xPWvhZeUt56DuQHOCWeMskJAmJRzff
EsTLWMzU0ICnPlHxYNbTmvmC/RndPqXkJBlPw4Tp8MvpKkhh25LshUxO5SOIGdoNNIjQUqmg6QF5
sbc0Yv7vAufmOKtKuvppoJ+G6HLmOWfKUsuGwHHgbggSLbtoOA0Jz0DRDLhU6wZjEGE4hD56gQk6
TmUMk1JDo6qNM3rRtsMGiHkvEMZVzt8UosW/pZDF7iZIypSNQO/u7z5HVBAxYUc5gl40MZXZnzWj
D7lZ/F+iHD9xNS6RfB+6ndGH93G+7ZiZ5RzrcUppkCfG6rEkB7YpjHiE+c3v4TAHjQYlF05o8JEa
3Dkb19qSBLmMkFdXwWpv21Too9XGSYe1Kfciz6wiCS1tUZkyxxiUyWA+7DFC0259qApInrt2VZVg
WPPFZx/1vwcV5VhnMtG7gOL/Mrj7UFaPLp4LwwOcDJzR4zod+OZ7umEMqq6mN86kV8XKoykzDYCB
q+PbdeSaBbUIl5ACjkizSDv1+olA5UZEOYwfhI7KQY797k++aagavTuOYBF2yxEz9MRXV7HAh9On
5V+LB83RRXMC7TPfvRKLUwWI638ArxXoRraRpv9YMSHCrKB+IIe9GEEPGvcMciVgAIlIzIlBrSsD
5lbzLpTFB9C4v0Y5rm2RyDYBP1ejyLI6aEcqQBr8TWaqpubL9KzRa+kdYGB56QLk0RbzEKfygBaQ
aXxBjuxEkD7sDprZLjfLjmveMmtW8I3ghEy7wXFnNAA7/9AzdzpgK7of7JLBvGpvRXXnfgG5fsws
vbNTZ5HOMnBExCEW6s8LWeQljW5kCdbzHaGkffpoAAa1nsZJdrceuIcKyxLXEF4zSw0Ut2IUlHsu
FrLtcHwBdIrDm81sGLe01AjwY9YRta0WSVsYUUJacHuzRFk1IDdOEJFJeGb+dlzyXsnHSgx1y8CQ
6tDV3aiFzVl2ze/pq9hD9l9wT/QPj+4zhhI1pqVHEl5yHbKMPM7H2MABdUWaaeElzwIBViRXboC+
iROSzbC4DxEcWChsAgGBfRfhYlwU9GoYZGht1nExvxjXprN3VuVOg2UyIzCEnQoDVIxrvC5VAJtv
PcOE4FtEYqyLgUW3VT62jjY1wKRHcYLhwfHunfyHRwMcVL7qCjsS8ZEF62JOOgUae1FaW16iQ2wN
/OFInZuUg0QK2Tjxor7DCIuSymTCfVbgMoSPt1jrgQCBC0C6h+qoIQSHR5PR1zizSfGPfMoIyJ3d
CH7pZIhHgAzdetiC9q65I9sYKAShM6D31bvPmUCyhQzdOHxptRCYMQr+lPnFoCFN4kijY4y1IxK5
uBZiIbR6AUrrDAphihn9Bj9KK3Z/GyS/aw1JinSUeceUc6G5Xs08FBAMqFz3kbizswjD0PQLzF6Y
s0aOg6LghGa4B6gmfYVGpRKXPCh+EpDNx8mb/TSEDfgPavGZ6f4DFfAQ+v30jmqbWx6q2JzWgYAC
QqbqGggyX+Atu9YiyilKt2Jvj+/TKXM7dzeyQCY8ORQxQRVRO0FycDc/vgERql6MJzAy8T7cNkUW
RsdWOPPQUJbpQHSeOp00dMvxiHBdvn6Ky8ITs5fBV13CREHJ5+pSLeuDxoyr2zuuvcZTXCMInkFL
esvg2hgw5Ur3IO7gwPziOePb0lzZ1nbsMhTd7Cc5Ys9WxXnqdPEoTADFXfGEcTJBW/DONPpATYsU
/XYHDhZD99V/nR+BwuyFDq+VGZlQgfmPztPQcXQVX46WihLStJs6ZNRm8R59N67FXLeI3bWS7+dg
wfyuTIN/hJlrOXCfVHQxY0BOMS1Qi+D5PdWx718Za9ftC3pvyX5hnPds95gmfQ8SP32QQJHCyU0P
8SpAtFkH8ZzMLpl7kxrrANYhXkhIsQ88gB/EVlIY3NPsmZtXjAVAgkAZmeKOUOUgqi8v0MCrOAwd
zWRoCF6qLT9F1d07BvI21DRQjfT0GUlY9Hy4u95d1SS6uHXlOEr8zo7a2Imx+HECpL1U9ppTh9sd
PvL0ZpGgFsS+IHzwMctOkE9MjhEUns4GX2TZGuwmLiLcC3E5QNVqqcq/UL1JLgvWRqV4PO1M6K6g
XLX/mcx0MCkvSgAFZn16f/2lhlLEgbYwBlS7GZLUotkVO1WRE0xXWFC/8HkRTaLxHaJl2E1XOiFF
T2KA08IRoNSHxpOEZDuSfa21RViVfnBDgLaJmJh/JY9cc2f42qlfI9+1sdQfD+z7MfIyu9S4Hnbp
b63NbReSnvJ8Fpinw5Asz9KQpEFzb3meFWUdZCZN7cf+MXe5VDh1qZmwru/DuD1GOexLVstbXFi6
RNbh4/h26TdfsBdQDO4Pap3PqeVYOpa/5EdJAofmohbzF6TWLRuJyiKdnYP1P64gM3CA2pYBYJB3
e9MpOQAgtV4LSW5Q2Jy+3we5t5SF0NfUDIdw74zXoGIU9ededgoC4vAG/dVGXPHGIFaXOkbcTtgw
Uan3UrIizdUZjQdPCdtJZcrSXk6KQx2rS6oiPJEdQJopOz/lqY9cRf0B9OWNRnG08qpDAaqF7eH3
vQSIPsP/Y0bcN/Bb3AT/hx+2QJLKRjhI4FGioa2n6SWC33HpRp2eg1MUAfZbnyee20FWgigfKhgQ
WtdPzJ4apVZSzLUM5Oe8YtmiG+YZUR8qSnk1HwhlfCly0Bi9FDh0A+7Qr3kO87fIgSAgL431Qfto
XjLEA/vRnoUWCzVHLJ9uFg/p3OKqD8HN4wrCWe+AWOBahXk7Sa0XW4iexAZ0DXuKUWWB/chRljF1
Yzc/8PvvlO/NxAtRz+FgIEec1B1RzzGjW/On9+8qIapGccO+HNmnZyLMHy4OT53i7SkvSH/N9X8E
8CMkN2tx0EnmA3Fym5/pn7fxGuSkrzAK7n4v/gg8nqvlpwnlBbL5+S4f89g5JD/vJF8eg0Ob9ZEq
rxOMRqVMrHfc9VKzkGlvOhZhAe5nxR3LEYjPCiaLzQ80tg2Y5fq5V7jCCEd2AF9Unbvj5RHQg9EY
wEfeKkSzPUpiYgzxwtZf1BG02/XtBgoaHTdY2nn3IcdW9nmSUSQxrRQNptEdE1ru0GHC2y+1x64R
avx98B5KTMOz7W+EGrI8BsoF6XObgMJoWzsXjtB1PS7HRFjnHXztQG2x9ht+tYYUrY4++KN0mz7L
gicgYlnHp1uFIwwAKKlA/fcOB5Y/mJtHr/Xph0+9pleEBz4t2GCXFus+2KaqVdM6oMK0kovh4sQV
xWUr7GDd5VAr+u6/35KW/0nPz+xy7+D+xWg7CtFmYUxQ9GwVAO8sxVV5uCzvdsDrb52lOnXLcakL
RJxHQlVekpr9nWQ58n6v3G5RgS1b5ZKCGcakjrqrvlwIT/1LS72rdsxewVeimNfzQ7TC4qveg0TI
fHl0AwvJwQeRG7aygBnwC6qg5V31O91PvPA5kAXRPaL3/I193ldwmyermcGvVRJ1LKHw4Akq3MDJ
AW8cKxUtzt5l9/rm+4rWFMBc2AJy/rfjl8jSC1Os8mLXM9874tLPIOqXpFthtqL29MH/p67jIdWT
1hn4ZD548ZbxGpceZHtRJ1I26C49CPE8RI/VCx1whJtJq0T62mk4cre/yC10VPKdQY3SGqYIujlE
khe6Qkg9Vxv7zcJSZI4uxA/zkdjpnvKXfE6ul/Gub1lH0gGkJjNxsobNJLQsO5jigl6r0pdN8kH9
tFRyPrGFIY+GxYnrB6PXa0M/V62eJrzi8aroGz7nwZzuDXklZJegFDeJ0GF7LUIWC6ERFa9+K+YB
N53Q8M4VuD6MGK090+YvyT35k49IjBasv1jbpKjtq6ngk/jh2WOsRDQGL5Dq/sdXaRU2CJmV7AJS
BZ5TvgW7fSFEVbhbvgQUT42CQ4vrHz4bWvhSzIfuU6Aph5/+1MnjqaFDnzNCHrgZktEWT5jOqwep
sCj0aPG2kiJ+AfucO05aHT2JRXUBgErHwxHjdJ2pyGRnoM8zXUmux2lHWExsgu0nzcSp/4ILDzx8
oeurr7++WD3Me4oTQAFpc48bbAqncSKh8XbWZs8/TPbJ2LtPNh4lICLjcWqXy9P60Iv2Z2D41y5p
CHE7BvuSD018cesvaxeYDQjGq3tYfW4ylBGX2xFBh6r3phoieSOZxxdRf4+pkpHzL0GWNE5bFTQ/
bFpKrYQ7068ohXTD7jXIXMl+LCwDnXIWeY54EjspoXBjSepuOmExLfKPasnSQpMMNMsbWhLeTYHZ
p6vGp2Vr/QtpNVRtP6eNj9/7iMXbz+uzs3+GTTXrs5+wD6b1tFnA51LHiYbXpKDDdKgPMdK/r27L
HF0HpQmfLPLrt8K4WgDLp+ERY6ScRlFy57pOnE1B0JR0AUXVXMDC/BPjdfqnzLXF7UcADwbUy0Q8
BGxi8V0+XlzNhTkE+EV/pMNvTnmfpI0I3kWt9T+tTQv1mvqyMEhY6u83/u+F991Ds/iF91jTVU/B
iJ+V8mr+UU5B7DjDYGZN0gZ6Zg6Ce3S78Ix1yQbu/noITqBF09c1tzKe5jlROANnIFkRCnC9QsQw
fqYmCl+5oWj6QCJAGOrXofBnwoxQPBe3j0Q/qB4lElIVb+0UybriptvRHMCDX6pFsjfRKolBenKv
i4z8wDdO3+hOzC6z/VCdI4D8WAifNFuats1FFv5C/JjJAoc5GqyQMx9d5TXq/Zn21IfYO2HrDmsI
+2ghaZYuQKETHL73UUK0DMB4rM6Iy4PBKVQBquYIAEVwUKcDMXvnk+vAzV73K7nAhb2gYiXUxERn
G0lB7h7CSd2TXOenEv4nISDN42S7Kw9SuUogpqLv3MRorv9+47Na/0KnPOnyBTh0kWnDlDRbYDGa
aBw4UJJASZZKI7IZyiQRy9VQmAMy0+Z8FYuYK7GRr6rhPm8qkyz6JBkUce820yRnXfbxNC7xupib
0BuimV3boGEFvfx/ZaYTSqxpVrY1XAB5BhjEYzkWfmcBMVDff0Um3FBiGfDDvw/aaiinNo3ZZVK4
C2C8AUBuc/9tc5EM6nY8PQ7iRazJC2k1Gta11PI3I5fgu8T1Cdx8OXAcaxY49mwCYCRe/31WI+eF
Z+B+Q5aFp2EUWxKdbSUxKuWElQTFrC7KT0xq/C08Z8BfjlYoVpA7v86zXGjTuZVyzkzqdoIzC66F
TVD9WSeQJnPxfyexZZxdolRpz86ID4V9+SUDXucE4UMTYnOYYT2HMqUVpFi84+ZYgp2PbPjlDKov
IjVcjSRwOW38PVJhN3fZlFDR2vrhCWFlvND20xiuxsqkh6kRJbx+kjhIvponZxWEmZvPIPGWAN9q
pmF+MeZ9iUEDJ3P44TDIiy4D3ipzm6NWl2x3fNJuOvPZt5+vzNBrv9DDoNkobnsX9n3sJn/OlsTd
gq+4iYqVhYqQs2a2oW8rYlKVEkYcQOyvK4GWI9KnjEYT8w/1X3aXnMf+Avx3Nq8sdz5dYMZvpeyq
R02VyIihuT1p0Gbogbzi6NmMWrmd+JDYJjKHo5cXveuE/iauFkLLFc4BwK5NJG6vxntaaHEEeUDF
ulMtR83vDhQiCNF4b7IAL59888PppHyxFiFRg8oHsS7gC+AxtkGDXoowtTM3nfAHv8Yb6BbSTdlM
zAaffJR34n7GFlWtu3UZpVd7A9FGg5BjlrbtzEvGAwLdZTaJiF+iUe4+B38a8bb3NRrmdpM4S1SW
KDSy7XiYJSkzp8xP8qkiDJDyGDFu7VYdlJ7u5VpSNhece9COcQyaEHsn+U8iXBtrrQKGUALI8886
kEw3EzZ7T4G52c8QprEYOC44SE7lTKO4vGXwdWMwmV09LVWAw7A8Qq4LOMRHpOjli3nlfRSIQTGK
sl4lowqCODivegx0fZGc80c5boiJ23y+FV8TjAum9twGidB6h1BuQwqachg8BgpSr8pW4YZdzvc8
GaLb++cw1RbO7y7Zyl7Bik1SEm1eZS6b1JyNZQpGsyzKWTGROvWT6BSrfriLs+iueWw8r3NocE1R
yMpnxHluDgrWUiHhAfXgFTpkZdVmV6rZMs6yht/CQvRqxvh+CaEwY9emIxow1Ww3pkoXRnwHYAvn
tLQbnmMJIIry2dVxc+LBitRzKJ4sbkVMUU39TCZhAZngjDdnPw4EoupJdQMOpk+XPf1qT9gR9kf0
FCc9h2MZORptQ85YLF9YaZTmC7ya2mrMYHHodAMVh5NP3QspcPZjvLUcbeb5h8dpQWJVOuEWGLR6
nG4NspZYtapNnZy6RknIXqwbmxnQdM6IN/e9hv90uemXs0mI6IX1ZMqnsU4b3eHjuP3JwmbbGYQD
5J4PD/L49zZyryqFOsLi+eEkP9wcgLshMJYmiG+CCjaILFjzYr78AICflicQvwjNWDcFuSdSp3st
V27ccHZJotuKPe2/0pE4HtnSw8nlArkpdcxYlmoNeteBi6aXQO8LPPQHB9EDsqN+CUbgxhrgoHiu
KXsFtrixygruliVDjzyOKbi7SGpXqIi302t0t7UjICaG6r2bjZKblDjIO2bGFx8Sofj7ToxEprNF
ZGgi+eiZl8v3GFEKHaScd8unNJK9l0RmfJChctN9ypjPVzMacuJWhNP/+k2CKqqPvt1h90lwgI1j
+rFSKe55+N+IFy7sSJKifdiN5dlq5c5Lh6zft1Q/jH4Bf34XEoVTr2zVDgcqIMeCeMmcHnRHl+uC
RqfWSm+VgzZv23mqvBQkf4B//oTeCNymkYfrLNOSOzdn8xNBj4b/VSm64LSCnay/Cc+3rH8WUZI7
btl+10saxH2TQ2HsEQ/3F8c/z6GxIAcq8DiAwvhhvWfTcl7HidaKHXpoAVM+P0Jx7uxQUD6Kk3zy
jfabnM+lJc+ct5SNF3T3P6oQvgz8I3a/ypLXsZVw8dfttZ0EnpPAXISArofvN3pljlpwpa0p94l7
lWH4we9AsSzKEagMNl8eeRvbOkcIgAQvN1iK12iD+SHXFPkQs6Cnie3qq5BpxXv0LFA9SftgYIks
Hl+Vg0CI+PeNZR+ENNdNvydLaVl8kLgqhA6AEoqUjg+nxRYEOAVylbCWf2G/z0IWC7xe0iK08aB4
eEgvKsXoQpiUHdqakgcZHrrym60AMFzYN9kaMg9VeCQwFeUpboMXsgQS0EJ5pcGb3jQB2wl99YQA
0QiegJISiv4J0GGfJo+6aBGzbt/jP9DxQCCpqp5blPX8ThfBLkOsC+oP0iG/VT74RK+Ul4pshiV9
QQiNHirBtHnvCmuYgDrCA2Ymf88XMrWnY85lUJdhwx2AZGfuBrnzQyAO9lH+W3bwX6bUV9476gt/
GpP8hSTgkYc0J6XF5NTuQi4gO+8g4MYxxDS8WqOOx5/IF5PbJ4o8D+V5cmvrYEomHJb3b+APuSHO
+VX7suSvcA6uu6E2EpXq1T6oY3PyLEkfBZjQiZjyuYgYXyCLTlQn86Wp8Kfn6VVmtGabXQrSuaVQ
9OIwFV95uxdHlF76fZVmTrq9GnAe325LACLoKk57vtK5bqRnhD7hpWfdXgcmSG3QRDbdmFR80cDz
mBaVqxTwzVp3lWZunnEFDCSvdmsyPWrCZpAHzpPcCEdrK3VDPunkWo4QDujIFHG0jkL7iRcnogRm
R8Zjhab8Ki9AnPaGCmvvW5hQ/CBNSqsMN24ZlBOZ7MaFCkf9W6Rz3OvKPMjuXWeY5iP6S3wwv+08
292T5V1GPDW8ajk8JG08DsWXcHhXJ/BseXH1TyISERnIIaqsHCautdQOR1IIsuHWEpZrb6CQP/te
06r0l1OwoN6yrJOvVRyzG/6krbjLws51TmYOtvLccZLwPGLagqe6VEaEGdoD4++5RQncffyjXvUu
cLE4SME5iMP5TRSZ8KKWNN/Rtdi9CKMxMNgMTPj79epa95Ask/N728tX5XhPOmg9K33AkDIC8Zvr
lbjKw0i8XQuHbHuJEnByt15QdqHP7fHmdlq8KRG6UAOhkCK4hyVI47oAAeYvmFL9xgf+wTz5PzGD
il9/FWuGozwzCHQkDaOPZ8L1A43ch1stIaHCloyv3WW8V63VT22alC7hunS5Dg9aTf+bE392tiU6
U2/wR8sqVjy9hMucbqPgyTOaZ5+58BkFZ/sg6kaakBsJVwNFKEeflRenNR24SOzhnK4ZLklfzzjK
Bz7oji9yUMInqljABeNppKPlWr/o3D4AlLXqFyAQ1MtXHg2uPFMrnktGwyJQ2kEqHPoYfmMQ8NUQ
Wkh5IRouQqnVBwebZDi26/mNGCM/5GUKMkhDrUbC2+i8r8BqsnUvvzeYNUDHMJ9rLPSyml56SQhP
kyB0hDSaPft0FCnXnwrypR5MwSCOmHChnX9kRGXLuLcKwYVovsm+xCCMDzsiECP0t0RFVoaAPgQQ
5LxgpmvlvHLyLnDJ/ixrN4YC58XnHJtNA/BrqKD1qTph9KyHSFGDKtUAMJz7c1FcKuZskpq7J7IY
KKpZJhS6pj1GnpxOzxqyh6PJ9sDme9KxeVTpz3li2xvbE/iNSslmabggIAKsHDTSfifp3cGiITaP
Ifeg2G1b0GV6IiQ5bgz6eCk6Ek2e7ZQCUbfCqvoKXZK95OLPUaRkE77A4pFVNcPPTfISiBzBW8Nh
IG5WRf2oYiaAyFsM1UEFi42x1aDowSPM/T7XEn3qabYoqSHtbFNvi+BgJI9rw3TnpJecEj3WysNt
OQKEFL6xOWVAYteHYGjFWlf/aarB4RqC/ozIgokDlDz5Nh3kW2GdFu4QQtkFxXCl6fhEfmBR0dQl
bHi0ULhvrp4/ixQcUSOK4dv2cJ9qvBkt6dUQGbtzfSNMIAq1Pqo/yCDiDa6MMLSoAheogG+1RyI1
33M9jmIgVq2eoUULI2g3IVUwI9kOfD1ZjqgtRW9vNWiGi/ph3LQORJa/Pfi0Z+RCmaaT5yAenAP0
Yvw12cYyVuZp/kBvFl2Se2I0a5iRIGYbrDw5lASlggrrVAYgWrhoGtKEXmu19nLOsrxIc4RcM7y4
/v5F2YPKYcrIWZeWROSWG717+w0n9xqR3WSFKaTti2ImENhoQPzqCUiMkJkT1mk1z8oYkXVE/g2A
J2GrhVuD1oMudUwF0/avrFhhwiaVq0Iy4AfOQm3R0WIKKkZpHoGfewMD+Vl58x3GZ8ll4RC2hCSr
DXXX55GHyecGho9OZYCp8adnGF98S3RSROt8bLZca+9S7E3YDw+8Tl/LxcdklOXYx4+d8dl44p2f
DnhOVUOOuaOuuITZHn8mSKJ8dTtLf55sqEaNQDyD9yKTHl6Uj9vWLjy4yDKJjV0eaheEZm91puAB
rpMq5UjbaSd22IOSM7sFRuM106G0RDofYAcoHQrY02CLjBG9p3fQLCJ4Soy0in/Re03tUDrinZko
g46jn5RTYpd6KZg4VgPTMV9u1nnBmIem/9G/mAxaqixVPsq41WyxBYKI7bS2VHv67rbMUEVfXzAj
kBOCb+KO5pCSMRFKuo/pODYIxzyvSGVYU9/YHaK0BEWz2Teb7Gcdpt35gMJ48T+v7J3ohx0T1QWJ
Y66m8XsOrFCUebFg7+RCrmGVUiTgEt7aDOEwpG0cINKOLvLB0W6eSxuv99qXMEy3yuDI5VcYzofC
EhrhY/2/xlrIsVUU04VkhFtzbfe4PJexowOtkN92RUAQ6/nOstkKNKDL21DJBEC0ePgAda7E/uDj
ClZile5IlEF35aDxU6paLfFkuATYndwI0H9vXwcb0pAa/8SrvI4Tg+d4QNdGJaMQe8YQmvow8pUm
U7JyHF63fFiFTwOYZSiJPg2qcdr7Xetaw995Oxodm3x9jI3AMTL0tU7YtHw5czyY/2hZOnwwn9GV
w00aw2HQIzkaGZskZOiBFg93VsQu7DyH69iXTpJ1zDq68tgX5GzRacSQNsj61fWpMp0J/czZP04p
0yYpZd+3cvNan51vB7HrTHkAKshQ0cs6z7Bd6Sg7WJcbkyis3t0Vpv0T61CYiOdlH5t9oSyRw+cM
4BM3e/RybQ9h7bnUM3W+vPj8FBSuRz/ms0AcmStSVpb3hpDMq/CtLkzKLCgbuzEHtRanoHkn5s5c
+1tYyesq3U2GYLhfqHeOD3w9QMQSNfB+u4bKVyEQ4pwrntUbCgPgfkV3HMJv8gcjtZMHsgd/Pdxd
HjGhQkATH2SGWfFv2zvvINxilWJrkPjjbQw+Zj374DDXRQgkX/qSZelkeIqPBqu/hxFAWIHRjWtx
6mWASoLu4Ocaj38TeE5aVJxvqxG6alK0WqorSpVa712AwnUf5X+2Mt57GkiYhEQGKBFRBpCbop7c
poS1oIalUgJTRvHSHa9FihLMq2/+Mppt7iHE8+WT0hPAnKCSs0FRsmTdMUQWm9FQwWFJ1rTqAsPU
momk47U8jXQ1cV7p22NKOkKxCibH3dRGUvqwk8yomppddBrLeMGui+WUew0rdA6msTccgciDr/gt
2QXS6VM34gWCCkzJQSJPGbnl4Uwi5vmVZQ+YcXZYhro0jz9sWP6f7NfkuMbDDfN/IAykmYwuurfv
8wIn5OZoSH935ZZ4BGasMplGCqk47bxIkhYc/6SGx13TfTPY6bPxw/P1CR545IiOCgqjw103U/Kv
exmD0zvVOTpegeIcNbMJszutuGrs90zH/H1VmntJmDV9pytvNeVASIy2bHkR/hr6YzxK31VVxPMJ
qD4Mq6ro0wFukMGa6PEl7nf6CXVc6eyVsw0e4d5cG3bIdq2e4zqYbvjDlslnnq9ESv6IU2WTBdP+
lJl10q1aTt9acFV0S+N7Ccl/BOSSMjJpZ5KdOyEpTlhLu9el5Wn47md5PKqCzDxeGfKuicX4QVXo
nw+DV+ciM2vq240jcWmh2VHmZSDhIdZYhnckVrDDyeg2EZBgps+N9AOwvA1k/WoymKVHMacEgPLr
JtsDNXZ31KxsuRFzyDv5K3HXKN1c/ZsrG3ukjah7u12kwPzjyLLuEuKCn+JITgqgQLcTCn4CX3Y8
tWMHV7JdkFJzOvE3Ae7AK2gUJBosdGuUV7fc2gBvXmC4Xh0jZj+WOtVP7Acp2+Twpw+mYVcMjthO
KmI39e7E4UZZw48IYxHNW5xznA09Im7DBUlXFNXGrwiNxQSo+GCr25gVYf6kqiPTDOLmbeB7s5qH
CQOkRuJfsWtlWfdXlFfMlo50UCZgjW2V8JiRd8JvZZFNlXy3WqdS4dSmlBlPBkkGZP1C+MFHQ7L1
0T6TiYYUgxYG+Sf7a6zx9HV+Ct09t/czDj55F183g4860v3WkhdNkuyAOODngsUciYL9AbCMXEiD
WKJRZlLwe75w1DIfN5+eUAr6to7JWBEbCDNI69WIQhP34I1ki2dUooFwmCITXvv7tvjyyY2f6JEm
vCJKmZ8KIi3ZL4PvR4eAPCEpd4G9goPnBFG61fUNY4Hk26ZCCRibBL7qu6o+uU0+UkaSgMq8ZXib
+aHD4yDUexzaA44Vx0QcK4V2iKkAM+eTM1dbcNAgQ7Oj0Bn/okxRjuR2yZsw9JP1yMFQ0p1lRpVe
sCigKQ+wkIm+ReQ2pyQXJ2IfiWtZNiUJpu7l66OtDP8CGo91UXLfQBN0An86AeRMAiw6Dry5SoZu
hok4cCpW24+flZXk+rMPD0Nw0IU6ygpDSbpTYfRxiZ0DF+7dS9ZbyqRaod1c0Q9xhyxW3/6Bh3Ey
6M6wI1hQIzelshSRTpq7HIzcRFxjvXDoOZsLPqnWA4YENulUMl9lxZf2FrAGI3AEDKEXgIxcvmOx
L7/mF2bh1EL76ngs10rkqalVb/o5XHbv1eNl4XVA29Z1kKQcp8meSw2PkxIFLHKPedVeqnQKYhNj
CoUjJF7sWkkQBGl+Q6mN/qVmnTTswAflyAWrevQYh4ACehxkmaiBg26sBuFrTz+J6dZaCfvvcsGm
vsy/iUU/HfVXJNhBksVVlSTIoNrmQHUSLuDtjwKo9ybt7rgegIuRHcIvljCfE26sYs5AGKVMZFgV
TA3bTLv/gHug3L1EZRYG1fQ8eXX3gmPw/kh0ciXIh6V7IQe+ZkTm2E06ohAlGdUE2jB4m8BpylBl
FkMwHIm/mdzDC7vYTco5WIRbkkxVFyA77lyBhzCr/0K5oJo6cbAolEn0L1ldPCMbkS1kZcYq/kGU
uLfac58vmfIidXHJskLKbPNkpBzOa9/+yzJo3BAiYRONNry0gtgB4N7HbQRWw295CaE/5u/2FsOg
CiZcGYk2iDFqNr2MBDSgesjVMilF+BvP39YHDiPVHmyKCnA0h689srcAZkqUD1RxXXHfoxoHyM8T
xldTOoOcPd7d3Ci5m9ntAiS/7BspNIz3wBdurRhOEu9J78uv5eRulTmnVcB4c2vJYc97VYWXgoew
zJZIjk/or0QAsmPM0egjE1hUXneu/u1POkHKbJphmUD1MKWnARCu8LY4uFUkhI2VcZ9UqNPn0vzP
l3fUYuyUY7zefg5MN2cJUgfdV1pjyrIe0b7KWHyStz8FHOedQGfLXZugoKRFokLhbei+GElDbcyx
hF7KspHOxMqVZU0FpCf1XgtMRfPVPtzjGXQQMUF9LS0vWGnMXQqzz3LKO+/5WT6svaMW66ZfRCfX
hjflJjAvDOlXOJnBlswCanyGfQdUUpgdL99XJTZGhcxlNpG7HlYqm8THkkRt+3D6emNn6XSs1yvk
GQfIN5HNgTWOzTTfX+s609wf/VUt/vlcaiCyBVO4c26ZJSadxc2wo+G3dZd83Xqyo3c/BW3pm/77
f1spifaLwnbdBpQlnuVe1iYjVhEgcNnV8GaKqBC3hy04Dxe4sCJgijqpXRaIc+j0chngAv7ZedHy
ii6Ltlbf6z0yum2jkZd7YzjOMG/OfWbo37bHevmGtNpDRX+0DdGIbVXSfTJVG50k7JnNjD2GUhOL
dfUxJ2KkYIGAJn8nxZMx/ijQg1nDUL5z4yIduQEdrRpYrIOVqCfRiZ8KhrZjeROquU7N9OEmVv6d
5Ag/Z4mS8VgNjNagZuzWq/3JGiGl6lHTh4U5zahP7IUnTM5x/CZ7MVyExRHjR58+v497jq7k0+u5
e+REnL0GGs8/MNiCuDNXrjQrIlkK6XLR11kboJltklellJoIidb28SLxIKkTVTou2nXeFZrAc667
Y9zgWNLsxgqV6Hrx9Ev/zMMMBycf18BfsEY5Hvdp3yRPW9lu21ZPewufR+ZrwBji0ytXlTZGq66K
UWHORd1xeOlJlptDXh4eEbm6VoswisyF1pVN/SSujnof3Ycwfa+GsDxSbMhB8u45/p7atP9Wb8PT
lS959rSXl2xTzS+qyqwYmgFAIfN8Q0W6zE5MlZTLt32rH48JyyaB0W1L4PzIrMejYgAMCfuMT3Lb
V46ilRMV+UHj3z5Bo8k74uzDK72NPdQy50pukU3pZEhMcJf0LWQPPpu5zPw08PknB7GewHgoaNdr
rAwjCTxat2wdphou4DWXYNp9LgdQQQviog6HiVd5bVavZ0/8uc312G4JdxgurS81ft1OT1W9cPzm
vJy+x2yd5bLCiUMgpASaqmgvy02bw2oAYd7DRL9D1qwi2InJCTDuqAy2TheQnZeC4MMUaFQJdqnv
kGEhUV81IgMt5tWxVfUYHwgnIqNjbz+f7EXsYh8puIjggRo2PT4kb2pTiEP+VV138ik9JdvOuiWP
KxxRHhFfRN/Ln3KWNB0NuNG2exODjo0qA/RB5gaBjyHjJgcY/qKkHZe2xQZDW5mAVH7Pk5hwJA3M
xgX2jlk0oS1k4oaBy4hGONZGu3OXm73yYtiDmUtItxpkttnt1Hawx5IpIpvC35uxhkjoLDdEaxnX
H3T8AzqEh0X0DAxV1vAmTP4a48SnwtkCuAuwI1etrxhZmNhe0O1r/fMC+HkQuU7z30UzHn8Aaghs
7lWHgNJy/SfuERpvo19r2TIg7wbLUV2zxmXE4wkOAdjlbykb2Not2DmJnImQLaK/6O+wvKuIZgV6
sF6G0TdVgUIqIpP3LodtO9GTl6iMPgrCVc+28A4qWKSUH5eoIw6zOhLjtCpOumuXi1HYw0ILDBXb
WHpIGkmE5AVbKazKaVDpM6soUeGPClX95XHVlPzzd1/eKCbGTDpJpiv2WLX5S4afhJHzrlwkJLey
1h0bWnrZN8MYePSlwLueVZGSRhAHh3cfE4abxALc8Y4tvfvRNcE5E0PIFRzuQZwVmFgMQbgP86fc
4WHCZscsBRht2xI1zfYDvLajVY4LlxLZrvAFBX7J6Ryq8qJUFRF0WMo44jMXN42OW3Tes9Q/KBuL
X6ScjZuUkciUBgkjhpYGXwTvbsY5QEUrcS7tDRSzJ+8iaJNjCqz7l1bnLasBntng1tPqvGFbY/BT
mHylRTKOg8b29FMoPBSs7Hn12J9Vt+wxeObl2huTCv67OHEAoEwpTjaZp81SezII0z2XLIFjdq/z
wveKHeoUASRg/zwaoq4VVC9cGo2RWqmugtqZlL+JK5t51AODvgBJq6ArPduro260J/3Kbezn84CQ
PoHOeU6zm3BDPPp1Psuc4gy4jUBbJa2rZyYt6EJNt2SiXSzFXpbCmN2X+9j6L/bqmtQ2N057KlVa
OOFi/zO2Wrl9EwGDLjwD0d23u+21sUtoOmd86vKLdTwbkjBWnqpx6gBcCBh1YxtfS4i2IaDjTDxd
qMRzQQuXMvS1mfXZu70SNkBQPyOi2DPFqg80BNKWk3nAXig/ScqheNFA6RCLDfmORhKJMefWyjhl
m1K1Ezt7+l6gvz2R+RNgIsnx/q67E5YhCA59nYKIEwCMSHgmsdKD+imWxMYiDSN/qTHg80Sb8TmO
JUFgAtj5EbhuXPL7TtYAjNeiSh1VIYsBbI/0b4OCitoJkS0Qg6NjE8zR43saACLI3/XnygJaoSnk
i+YREoT+0dXEkvhYuGVPC/aMTLc5zWirfSYxj6pZ4UmF+20qC+Kk8TZ7HH/MiDze2W3B70qHHzbB
64w+3O/hoohb6GF6Bc16Vq9OmBfRsuBPiIMr+u8S2ns1qDtaKFZTrUBeWIIxVzYAIFNNafyd3I/0
XFuIaKywuYEnYMjJwkLWJfmVBPrLZSlLjfRIH2uZTQb6BKS1jx5AHkAucm8kElbMjhJZ5VV13GAh
u8rJe5hvEqyFGTgZUhTbpu9TxS8kOnClvLieQIgemi3b63oZXMBBoyboSVGj81UxMFJFbK6w/rZa
954Fkz6MrYte1Oc+nzLA3uTM3f+6NiMLG3IcYnnpWLfdYI/JrReYgRudeSDNSRQJzWkFLsRCfZCs
zqFcNd4/DelkXnuaPl3usMtMGHrTZWbbGaGP3bXPRA7c6H0zUhDaNtnTian61qKyl/locfh3JmEm
EKrB7qL2qp97MPHSN+ZU82xnThoL0WXUdZ5o0aOAe940vu+Ke73iJ9BuI833Lo3oDUj/B+K4fG/M
Z6JPcxJM4zk5NuPI7pVnPM9DjN/EkAfer6JNE9S0ncVK14QAT0a2R2VI3c/1ITmKUUbpQgohsFYN
Lq+jeJVNTtrNscocj1ea6Yka0pt/nxp6I4xxd8ZW0CmDjIOK3r3vPA3xiRidwpkFAdpvCda1DRsi
xSNz9jwUyriN1q5N3MN2Nz90elJ9lnrH618DEIgdxiUoevD/XMed8cU4IxnxgwSl/rvnG1X763hf
IZFzl8zThHLn2F9HaGv/Hgi8Df2UaVYmV+CmcAzvoIONKAvkrBAlRuMwfpkUN1X29N4TDcDWm/ev
+JeIl1uKO0/tbS1AQrdZZIG8gozzq2bntB+UQQW1KPAVBN/le7nR1TAtOl4j7jKwbzAmcicf4Tt/
mEMOC4nInpeZvrzVPnO3sRo+poPyTx3sG71GXH61/tkAj6bzrice4MzV+4PETEUb71FuzJ+yXDSo
VM6yyBaRrAODixPngpoyZ82DbgPTUTN+hxo375qgipeDRs9ELXhiIEbHLD90C8i8kWtMFrIxXaZF
MqBbwAeg1TY3IjgKrMcpWZWnERatIqbGOB+nxrTKY1Mz3szggQAqZi5hic8kYZe36yvmyguLP/ev
GILNWdxZOxSWwujkfYBZ0QTfH812t85u2izH2HjCwG4tjXmnxRYQzR5zM9oyWMjxm8TPzGR8uwyS
EM2mNSqANSyDOiRbL9TZFFsLViYcRZGSlVWSLCuFqDDzhmHmkVfS9rJx8qFc7jhaRukjsb40oB2y
qc/KsWKBhfEM1jsTMjHUB7VLY00OIRFm+Onzn1QoFormNKCL2mKm28/b3bCNq9ywBv9lihnHQLPa
5V1Ogw5+ag8pH9ekHUSh/qHy4TYSSWu6EqpNSqht8aLnPoC/xbGrYGVzZX7SH4gJQNX7wM5eWdN/
AhtW6z+vpymtwE+zVDW5oLUBeA2dKhlMfLoWvWeh8s4GLPnaHR8j2fopWu4yJRSuhgxVF9stwxqW
XEns6No+qKWFnwfR0vBn60TvYQI02ShbhRCGy/phPFIEqA49966+HLYLpAYUVXJkS3R4fciVFxZd
T8wOyvaVBh3yJYmCOGd7+JdJqyah71tMHanrA5vzeObE0ZgQ98tcSxBe0K3w6m3QdejXZv9WAmaS
YgiOLhso2ERK4PV6D0WL4xoQlnGb7oeGT+xjx9XMovRReN5FcC2UjTROoswSNsJKzjI60JA71Q32
7C7dQskEePGSrvALCuBHNUgDMa0oG/4no4+q1q49PBk0XO0ITYBxxmhBXzJYdrM+YJi+NB/JNSc+
vyEVSrBp9MbhpIbaXZC36j/TuGLXB3skYnQp9ST9w0f00VuY88zNLpx048mnOyGzcQnOq1jUV6Gc
qtq13G2JP8gkemJsUhVwl+B1DvRejp/ebf45WIn14frwhoqg8lQTvmbRqLhhDw857mzAaZRAY/9S
EGGRpMx/bTBG60RLPUJFQ5Tvnh7rzHaBOU2fQS4wbxx8iW3nA0R8ry7zVGnWSBgD9MD71Y3sdAsN
JI7ljgxUMDyoSq9iMexCtuyEtVrgKMjunhXxtaIW7CrVii9AY7JokurR/BEHbF5VrXNxJ4dfloIu
Ww4Ho3UdQa56n18WXbLQeoeWvxhXnvUG3aUcEzC4aRvwDEQ50u1M0nLmR+drQ2H78FZCHTaCy5Wq
OHLvy4gGELd0VtL/Syjx40fcTSHkJCnP5RsJ9zLwQwBjS8tObGm/QHnsEZ+okTg5KLbPRaStfqbb
YmSh1vZWgDQpc52pudPbJIEuLAIC4G4mx+EysvSg8ZXgpSAa3Qs72vlI2Np0E+WV7IBXxyXEuSiO
uxoeSTuNJBMEdRLgp2hCD+aEeObXZFpA1C7GBqxzlxHeQG8LxyKn9lrcVLvvl3XPTa1kxgXMY8h9
ip7dDIrlvKL9NC9qfrQsqxnE/uUFMr3dTuZPZEw0xOn+DqFNwXDT6cnL45H+tUZu7HdAkcTsY2Qb
5cWeuhWRNc7Jbu6RmAURprHY9h0n/sKToPTwqyVMjMGxVwiAkR+TuDWfjKnEAsiPgSwJdR4QyKOC
/ZZzmZidcOmbmMX6lxbw41DT5HRhpMytzY11fk3DIpM+CXcz23IYcSqvsvbXk9sL4oz9HMxhgMQd
ZVBAwOgsd4OHKVV3olB1cOP/fyCCOp9VT7+y8N3t+o0j3TpGCFagGt+qwG58XVmR3pvVXalGJb1d
3bGRSzDuBWJfVPZR/44C7DIdBOr2CWPP7eoYzNkGV+2I03UMfYN1vmv0Yg54yG46c1IY/kYPGb2b
QkH/cA2ArSUrYJDNsYFLOfwKORZ4dXHyX+qPt83JAR/th+PRQcs+zdp7xukwiWcLMCULYE9TD20x
1fVmDgqGoDXxH/ibkXSiBa2xdeU51XQcSznywwnb9fAzmdTaKF7CIC0PHHiC6gbt4ZCRiFi+f8Mj
HxGmSsbPmSCde+zvISD62/l2KEmYNYxiBcGlhEle5hyG0OXf3Bop+a6YREsPObYm0JAN5/n7p9M0
9niCyYAmoPfXCNNm6y5EF5/9VU7wVBdPvDYEh3Ltlf6Bk3BDoqoEbj/if/MDadV6Vr0wt6eg2rPB
sNAfjWhIrS83oz2oF64+3q4KcszadwULetbckkil5egTXDPtuKbMvjtpwAlCHgvuErMwsZoGHyoQ
UvddJyCEjucC2JBlF52Ma6ICIWh56dgb47OADksJO8621AzK7Ibw4QefRhT1Dt1AF1AYSPGXqqmY
5PDkdle4kwc1Hl91mwA+nALIZCjCe0iep4CBm637iu/kApAPhqbuMJfJH4uSUT3P+qd69DFBikwg
HlvWGknQmS2KpsPkr1SoEYZ0dSxxaPS59JhwqtAKxCC/zq1rYwPEWR60aqRZU94woySDqoWhi7Bx
ChZ/RphffzrQkWFe1whtu9a9RLvILuWsBXdRtq2j3wy6aAIt744z+hy/scDSv3vFYcZxwWjbpZL/
TvsynmlyFlpS1/iqAD14UbvCJtmGs3at+IxwDcxthLvxlkZM8ie+CCQrjfrlW5HMUe4u7z7kWq+W
VzHn6fDQDnQAMAL7yqHtMCjdMCXPN2EkiVKSVxGLPQj4p13QvdTRwt8uw6zuKDWNwWKC9vpS8Zc7
gxXpoS6Q3hKLSSxU7ozVOz2JQMfyGBwM/yzPjLU4I5hU3e2ks9iNFYKVN191kfP4QinXVyufwbj0
9EqWelBa5f80xUdocQzEUB3Ho49g2whio31cBXweD2A+xbytvgxW0G0H3IjW/hrRn4CGe+rv+0sK
jKX4lRCL3SxbbbxlF1Nq99qPhEaWoW8d3qKUzclpEaiEOqs7GfnNfhGaoMOtrw0ZUapv1rnRGxti
h3M3qHaMAB2uEd+5aS24QhyHQF1GXk1AJOBUVW42GGBUOYFTr2GGUlk8EshyZ/ef5iC7MmpbLEJK
CvnNf6h2xq+tKYW/5XpEZsWA9THzk+WTJLeCKoJAGa3F8MhnGbSq36KisI70wH0liZ4i/dbpR9gZ
fO+jrhI8UX2uNz/vU9TY3+Q8RTNlgdWN6u7KqwM6FZhfP0rRcSPLplqBVoVDRYzp4H+cHyBv+R5v
TdFkqCKfRFT8t8yAdwE4DatJwOcnL2Wf/58xbWUHTApq7sOBVCt8wl92LVZQ6ePC31D8YlVwat2k
9g26kfEXE0VCM/Uk3y31sNNj+/r46mHsIDRd27/prsVv5ayZ/eeu1bnf7P08qo8+Io3L6+TVxDqQ
tmDSGZpCk/k5H9CGuxOzg//ezh6oGkUZ5DjK3RSOEuxhndyAeuf1ClCRnwLtxcwfAjg5VU0s0HZd
TLipl0U+bdXx/khon4KpqWFjYZ9uhG649HAQAmXCtxCmMEmEPqWglJVoo3SLjk8BsPzxYIJCvujr
B2jm0oQgNpzLANCjP7wl+7BNPleOaHphLLSvJaamu4Bgilgj4d4Bb8e8Bcl6w1svnIR2ntWn5HgW
cVm2tTBFjDIOzJRJMVSVrqjRW+2HX0cHLKcDChcStKO2q4DhcbYnnErbzaogJKev+KkqpD/RfsxK
WZ5JnE2nywRTdMXBoO9c5Ht9lbnI77pydmWfLgM1QX0zUZgjm5etteXQOaMwn/dxv5/HL8FzefJy
finxSIGS5Z0/51E4vvdd/Uel6Ki+TfzEkOv5PN5SIdJu+vcXPK6vDu+os3Iyn7AXU7/Cj7GRyGRa
BmmfgOLls6W3JCirmZZPoREl0WKnf7sNhCC/w8FSzwfz4wlBX0m+SXiVos4OAQTj/PKeGi9i0yXR
v7+5V1/cSdePyJZdlUPCXgywbw/pjB2Y0C9pW9yB9Ua7O6kPUBlWaYLCpo/5bPF3Yyfj33EiLHgr
XC2lJQn2aaGtp+YyrBQDzVYxNPaJ9seOTSoRQKyEUN5yyjoX5CpE9BoIuwJScfZdA/srLPyXauRb
ODwvoGTxzoOhlGY6tN9RCYzFTr0zteUh2KglH9zmWGm8EjkXT87a6BOhrAx4A5I3LuXHQtCyqskb
0+kvyg7RXOduiAtoJeKvSRTsssHuVN74SA3jHadDKouOsUDQ8O2k5qI3WF/8j81RZ+7gslSQTenw
I+kk9apf8rlJNkKDvnP5GCCiokYOZVnKnavXKEaNWfbDakt6ZL8JtGGtTomX5aRzVcPfCZbAw5V4
ZON82FlN7jWnkivnpch7zKGZ70JTh4t0tOPTxC586l0EKCxjmW2wAimP9XGyLMwQ0dTyRPcCMRao
u9qd2tlxCwA3GVd0/L4QZyUxIl+BZV35ZIfpBnh2COQlHXGEdtWgnyL8Cwc2PQq+yIsDXFYqorfR
L+ZgJqVMfxf0M98h7DtSLAicK1A90UlLzyslIZiaQIbwfzlzanm32DxwwEohOCV5qZBThbkal5Ab
5UoI5iqiZkBFAE09Meizb9CRSUAKGd2sacVuH700LYFTnE+reWWQr5UB38F8M5xbWNxiLUCKiPSA
6Fv20ZLJfEhSye5DsLJf8xhZaTQSuGbFsdIXYzATwiIz84P5zsekm4dNCimHkJtZxokE5gW2jHVZ
BQRus3zCzz30CBaq59cMbHoGYEC3vZFsAlNyIwQBX/0XIPRIaPIIlupgUeFbfGVeiTC60ouCQ305
b4x+sufJczJsZFEvcrOn0x9UAAO7tqOcBSQJsDmqArbNhSvux7YK+USYNY7AVC3VUnGbmDhgiaQf
0x5TqfvmcytI43HzCgxD6XTMAfvQ3D1Kx363ajVyn1NCw7X1dqFIZDWGgn+t4OO5WTP5bbsoXuSk
P3UBksS14teljY8OTJ82jZtnsWTCVdZ+95U5DJ2Hk63hbjIJkjqvfL2NAzEAEU03JHWYd29B0+q5
uNbLalozxcN7JZND3i687SaT1yhbgXbX+6PsuMrrf3PcI/uEwFILN3xAQGv0rwTNiuGPHvlT6L13
nVs87Ib6dAsmCqhKBCC6qYXsdlpqJzzgPpABHuIM3YozVuhmpuK094425Yj49/cu9Zx8yF62bJPs
7wIkJI2I+geIQ2m1w/x1R3+kNU2iQkq/TmDDGh+CQyBwJHh780bSAyiyqObclE3yWBifETwlU6R5
wRRRl6xNzpifXuks0FgMpSv5hgGUob3EE4nhAE48O2oMrrpKVnABhw8VykiurO88e9WC/Blxg6Fc
ybqxaijsZwrqy9b8JgHUh68LQD89GNQTZbZw3vk2EsWW0RfQapENv8NNdr8r7KF/VYX/rLhAD5v4
nrLtukkXiksITCstRNegdWb9T3/4lP39rFygWtebUHnXUdLuO6vhZDHqSwnXj+Xrqga2InBNCEM4
NJ0UXyNxETojDr5IudU633031wr32NAXMiMBuY9NxsP9OAcoqj2M1umXDXX0vF+XuEoYuWgaNEr0
MTGBU/ZAxV0dqIuDLcdi8lxjTzZrc9zWskk+L8K7QK68nUT6yUAsuW155Je4uKwS3FBkm266FneN
/TghSSlli5eZekG1Z1fbInzTS4Ur4rJ1RDFzlNHcMC6+tdEZ0BdKcnKs6PQZMsC6O9K0qAyEKypn
2EgH0akds4UuPb0u9yXr7LnVNoTPOkFDcWM74EDqMs461hivRKvUBInHc8ar2Tt8oLY+6DSEkgUJ
DN7lPbDX4DQ7At4MvExOCi5W1wTykrLjgcOyRufcBNZO4J/mCrwlOBFttzKroH6fWxcd626v1dPm
1FWat9vTfTbpvs8obszVv56TssKw7ynZVjT4UZCWxHP8zDMfRNrGemO9WnXAP/3vgAC/nMVR7yuj
rjN7eo0x4W59AlVeW2e8fWqfIXM1T8JZUb2wqrOYYVZF4OsFL59Uw7GbE2UfXAotdThzQykSS8nU
DlAILfJ3AYiqMAyo4rorOWi5XdOsBVbNzBRtDRBNzjUZpkaFo+oLnVDTr8Z0d689DdaYOzTpkBQN
CzPooSxRkLKGZqj62SIoSQ2FtRq7xQHFh7xCO96yT4sGuQXl4w41152XZ8F10ya+Uv34cuyEhJYw
PxM0Yw1MAmjS0jr9zwTcVH7No1zWiidb9kAd3QjJdGWwzOTYeUNSWjNpkBRV/Twz3c5eE5lHOCaN
L31pITk2xDG78At01gF9VKtpw3hZ2CdfH9AqsA9vJJ0Xe5ZN9K7Ufx6bMB0mvfZfvST1DbYIAi/S
HfUloXxs5sCiIWWsFVtHfqxdaVMmIkICVI/Tg1SXGHjSm5xi6Dplrh8TB6CxB/8hjqaTUtezNmZO
TyNsx/rjztLDRjyxSL5edLacaCxhgVGI/0c3SVHTTUkgi6+YW7ZQUS4m0Z8wQQI7+YpIQb9b0jZr
ARRj/P66VQ5NzE7AeBmT8DjBns5s185PDBBNlOCGQglZPjk3QKSpBXduB4foYSyDotV3TnZgNXU/
agwHyjJugdYMTHT1k5jYtWaNbqFdloNcaAN0KjMmXvvtL6f90u7D0PlCxc32yC24vYsjONhiybyf
PR6/Vz8U0PM8th8qSJMOz6m3ikNmp2qhMgk3S2qqqF4g3gvyDtELUbma7PoxaAvFyrk/FXs35F4y
2A+8C2ig8LvMAkl8NYvmRqhTkrnvNnTGniKGLVPqfDFLIiT5AkEHnIPxDoMMaLDcHB5xi1mHiOUt
+WeoEeOeyDr1XuFs6bPlTm1wTZ8fX+Qm7gaYCIkhvJUiJ53wCDhU7a6By4kOrax+lcP2DtucrDq/
LZseun1qfacfzMfVGCRerMPy96uySzrhbFfZS29TkkOT4O3xmv7woqVqsETmsqUJ82sE7uazUgUO
b36LZoWl1vw0BwpMxDgN88PL3V7dDiZ8ix3Wk7bIDF494M1+7L8QvIpINGwgbmDLyrzAvHFzzDXx
Y3FYaupMxdOYxUCveFas5C/vjAe6NQp/bm76xY6/NC4hzvfeED4yTxivngdrF2oJi8HqJzXjGQwL
7FXs/iRvDCTHtn1H0BIYWmYaTIx4ClhOcNqMvkjcfFyXMTkZkqOzIbWtL8ZWmKX7ucuhDuMBDwmA
7oo5NeNowFTJabmGs548HMO0LZCka8p7yc6gxFpQyZqppVw0SGVfhO+ZfVVZieaI50Q2pzcelQdB
RNXSC3oKGVkSw9MwwcikPc8GWvz07+Xcxvoae5WevAZIRdqrZ2Yf7812ORXnaETF5zwVqyw0Wadr
JpPcyzGtUkWyBSCrdSQITcT9Z2xOLAiXivjZGb92k9Dta0zTzhz8JpftTqoSzg800Sf+FyBjS0EG
NvhykYB9E+jcf5od1en2kRizBpe0OfI2pqGVgPMFiINBzIleuIMJGjwoAzBGpawH77LjjOsCAv50
pe0+tWHGGw6a02GalKGi9ICobzHWpO2FDAFlD/CpXHV2rtRL903aOo8/NWZ1xTz1nEU94m+IIAtY
IYIJPbmWVuLlhNPT/DbYyGhal7hTguCz8hHKOalnZ+VdHQw7ZcAYZxEHikbn4HPegjGijvB9/eO/
Rt93bnOZmgpQBnIwaqsqZTxowpD6ir+vbsD1FfftwHEr7E/PfoADyrQfbPmeSpUwF55LkwLngNy4
SjTlsMZcsjPK8zzEzGzwKVgk7cYQBJpBP3tgUEtnX6qmuE71wfXNDv/WxS7SNGO4s7nNlwAcSGrY
H8XJnBCpm8hL5K+G75St4txwjoTbmVNps/X6x+ez3ZAFwukYpudXHVvSHJA2fqRTVyNv1TvPhgrl
h/brJy97ITXDGt6rMeBo1EUpUH2cShx0CGxF7NcOefZ8k8mGEXSoeZngYxMXwOKOA3Py+H6yEsPU
SMx92US62ImpOwmz58w0GI5xfEvtfhKXuayS0fXKgiULC0/HlMSZKQg5UnEvcBTGp8K9RM2LCe2v
zUSpNiRTZ3ks6ca58bxRrtrbnnl6+y1a5RzGmS+vU6o5tjxcZsxQEfJxeuKUwyAwy5stDKlskLqY
U4qLl/mw7LDTDRrlm2neksynnkgdNOLQ8wWZRsdVZWJpKlZ+GW6VRGnSpory9jjOudDCxcJX9JjK
ctqfJHsCHUZcaKp6hc1r3lVfkmUt2TBfPofF/H7rgptqkIL8hfvbz+kRTFiQ+KCFyiI4EHkuktc9
EIVlWg0UHMFgQAwJyLmvQ+DuPjUZqG7qm08P06WpQa/UMHRtvQLpElVD8xYuLKnmdJd7rpmTErrj
eJm+iGE9kjLsGgLraIKxqIxCGrYjQeWUBkCOGFmQWZmrdEyQoPNIhAZYJwL/dUNCX2Q5LGE8EO5L
Cp12EeG9hnBsYEXa4dXSDe+BgzweYNgpjRbBHQ071aIo8vTQ7LmrXcXd6VpwbD/5EU4faJVbv/mE
/jBvRCAMNT+JnD4MUEdopOVPNYFo4mjfs7RKghFTgT3WJklIsjf0Tc0CM8K06ch+qrVf3Jg6DMzO
CCOQc2Z9XKX6GrFYVEI50K2eGmHHZGgebPg0tOmKX9Ctvr38M+UoRhPwKIVp+3EoowrpbpO/P+M8
pvhzoOUhnhE95Yk2/ABd+8+X8Z6jR138bM0KflU6oZo9ES7o3VjxnxtRqnlf/CJUObail3WUqmLd
14qwgJkROksEcSesPzyRDs36IecbEg0qMobVSCcOB1BthxMBadoQgr7UQDprkHXvJJdZ5egAbQ0n
Iq8bTlpFfHLQe34G5ndpZUFh32mHz56wxvyfhh6qxIuYZA5HCjwdYti5gw1cOIB3fx/oh8bseNOQ
1LK0wY6dQ59wNu5ISOPoh2FvdWXLd9pWIiXjSVV9FdnASPv18XN2meyos9RFNtxqeDN1ImvCvDu4
jX+1bvA5//SAlssmUK/tXuzvRnZ4w4ocTaLsn5bHVHWxnocCqpJryQKuanES07TV+nT65mL+mji1
pcSKt7cdE0e8tnZcS7H9u7YujFF1AM2c2SYk9RigH4aXZWMtD4HVqDhbRY5KDFvBzNKw4YNkYi4Q
z0LukabXMRFNw7pjuW1psc4Dp46cUdNpAqSb5lDaUIYqq4BjSrqH8QaOgAn5qANw1hh/obxQBmxL
lS4a+YJTfUkPXEVFn9Nq4W6PEerw14ox9sBkNpKKLpGNe5tMzS0aRU9nsnnPdhvz+OLvtuUtfydk
LszatOMAZscBzXauWvl/9nprQ/3YxtKKQ7pq83bbYolCcHPysuw0Edxl+SE7rnRAeBfuhWWJiSEm
j9GBZqsStBbT9WkAxE70jwl4UmDvpLrphQ/d3sGtx5udotYpdTNknDZSbqCpivm0l4eOiu7CXB/O
4cX7rf1AdPuoK28IuX1ZU9iUvyZ57JhvLqEaYql9Sct0K3rjC9gKx6f0SGmTYmUHMD5tqSroVvXx
DaaIOq3j/nrUDGD6zL3dmg94kL8RUyEqM8wSULOWwi9cQvUOi+nkbVu3znz8zhAD5BxS2VgN1W/Q
LR0s9K6NsXKSReqwavY4RekvQUAOuABU7WXggqQhX3VK14LbpZ7OqcJsZ2tE9iZKD7Rppi4b5wLK
zMPaXhTIcJdMwRNI9n4ESqUkwQnhobiKjGrPwLxSeTrUxqXJCNY7HPXHwAwD0mIojiU5gmAVRuA1
dpoFlYsPShwQWDKCPooUBRLriiwl5iC/5KxKNYGr49AKFrxlzBwd52Z2Jo/v2OpeweqRxVK+bYjK
kQxS+bEMwX90YVw/sqtA1jsDTyZeFUtTcLmlhcBzkMVikoesyl5e5528R5VIyzZkatQt4BKUf2Ru
3l89RraV/iUO97EhP1UCmajEFz9utYO9uh8QNlf1Xc8UOlIgnc61OH90JNWXTQl9kZNomaOoOaHV
Ud/Sgc9pfOu6ocUelXitwdppgiHBqTcNLZFxXDkB6AkDbVDSQgCqsaQsi+VEdLpM3zOIqtJxkGQP
axnanlwOf2EPFo02UCeStvsoggaF7g2wH/oFu8Hul0bvyktF91kmT4kbLEkHZ2TsJPTHOvRgC+Kz
psBOYhoam5aPUbuzv+2QwjUa7gzCVYBtAAOaND9kVmrNTkOE8zOgKIEs2rxo89UJVZ9NKkK5nnyN
5idLjrtIC8HS+bYKeoxiWNm68d1IN+/l9aMB0+3JD+ADUJ76UtO69E5XhceRUPywQZlnLLQELQBt
nfXmvJ5kMJh08oy+DbQ2m7s2nHinUECTlYryRqaaCKk+kFId4Ku4C9sHSa4Qngz0GBUgA+RYSu+B
pwWIspzJlMncEgmsixX7G5PaR1WSncGxwNpOMC9S5/8yp0nW21XVNeGt88btpW7FI0xQEkpG1pjv
GCkE5b8o6k+igD0p5L78RY6wV/yqLkGMKdsSxaeADnueEsr6lpmJ5A2J5p34GIPerae8HouEoH+K
8gDuVtJahJJO2SPjO5qntTsrSw+hGw30/M0C8M4HjH07rjC5YibBjAeyJfxnvZeKfZmsiSv7H4Kz
WbO8iZa5p+R7/7fPFtVtyUzYX24oPLgihnI4FByVpVHmOfriL4eEhphNif8yF2lzk55sRxf8MU//
LNn6UG7vLRfOPFqwmmDa0Fql4X+xf+VRDDtv0ZF2k/F13KgB35sNU8bL/gnwtne1PJGHKhvlo63d
ijQOJeskneYlUowu90axuYQZVFLstD4/FwS7FwHw3fD7S5FKcMs1y2oBX+jC+EL3Lg/J+JT07//Z
yrKcDIhxK+kiYoVkwbf/GFSwQjUN6gb3g2iqVIaF1SZ1pRiVie+0CWqhlairAhcgsTJodXrYLJPL
vAVqywRbTnVwOttI3DepBLmM2DMXlV41wJTycCfTpX326xxP2kV3iEyhvTk1asPrN4VcjAWcX/JZ
EJnz2jJ2k3oc2bWLwGOuyB6XYSUKkCaB6FksISMmf3v4gQxgCC/C1nzL6WJSYPEMAA6CykTVITve
rZ0O0r0pxnicgTgJlTvmVjysMfRPqIm/q9SI8usK7fHYAX+YNmWdHTB2j660DSPeYOeLHOOGRgDd
T+CQ8MZ8C+57zWzodNpbovUbR+6G4HAfJNpbuWf1L1wyLjw2g2Yy1epMmtl8a1LBALwd+LldiKah
csCnRVXXtQwKjStuMDuKhosjARVMeAPvP0+1OJVNMYyDMdqwPX0+07ULLTOyGWy/Qli94EisTZs5
vQO5PpgQc4M2NJ732IKaS4dmj9QOE9++9MUbYNPf1qJ6jPXMGjsRj+DIoFPmP5S+1DTJA/+YF90H
9VbtgUN9VY92mTYwxR0KBniMo0E+P6iHerdq4JE7ZnuK1d7+wfJoxU32G2wdy7GKrP3OmBJ+1VEN
0v4k22TI/1NxP3Frsda37R6opiPRTQJaiD65U6FSprDKRZJLenL/mbcg7lnAe3TX+sqiKgkaSEYV
blGro0Trx8vSGhtisvBjDHYwKnKXEGzO1pefy2oSY0btJacMkRScXhj6VhYCVjvtmUZLjFBrYaL1
ra6RUfo1BHzep9kKQo6q1/cgZbO3GsVwt8gif+qjVhJ/7lN2onni/h2IaDNrU1qWwvkpxPXvav4H
LrihPoou3Iovz5eS49T6eSfzax1X6hRLq+4hReXaQCjWJoQEfGDnL0uqbKT8McFs6fAvG7vvuV10
j6tuVxBr8Gk6h1jWeVAiy6XUwmmyU4Q2k0A26sNveE85L8JAC7zE+08fv8mAaVA3W6lB1Ww4pp3n
x6uswgaMWkQjYPC7IMt63WBgiwFY8toZpEnhU01MgszUJo34kq0ZT850TWIFy3wYo0JrdA4CujoM
JnnYkt44+fLHugIoV9/XW+l7oGJiGbqQsk/9EwVP2Z/mBNrOGAay4RiA452TzwsjVrzFm5GlYuzA
xX6NzaBtclea0Mnw9sqhHNUM/dOBEnKTQdK4hVHF05OQtfweKtWB6nU2MFtCMkCmBBGBPIwnMJRG
u2NHszXa2PyqsK5zHfZ7BHCnoK/mItXWrV6GYXZK0SCCGxQnxq2LLZMCQVfXA08NkQmEa4cqv3CP
KLe68J6XSm2b+lKCR3tv3NTSUggBqHy003f5xvJYcVrGgiJfr5aLBtMGRO5OwTbDg4k6GrUVK36f
VEeW+jkAruo10LveXohQdFHzmngXHFj6KnGw/BvX54K5N3HBbOdEobskXWhAPfzqyKsfDXpRwWHq
IVYPB+8s4y13yMXs1F/I2xSjLYcKB5KZL9Eudg43XleVPnaqOIPl6kU0ka2AoEChPBmxIZs5BGjr
2r0g0kMGmry6kMeIY0HPJfCeu8tZPHRse2Q0RM64PL2a0wC2P978dqVQLMwTidGnsCWwov+E1Ddf
6zPHv71XYaT2jSJJo81WLdKihoPEjPKFGKvB0nTTIAnU0Z8Q2tD8zQy/SSPua5WtIyAXYkNWlWs7
ePsiQZGbRYvvFnCqyda793KpXDH1VVfHGq8SXVl8La1XAcY3hOZjD788lvkfLO87xugHkDgeCqnJ
bAB2z4jIWfw6eQ7pVJ7tt57f7t2nmvOQH98/jjuQMBqpOweoBdVwZyFpoFZVHNnuIDOxjdBBWRr9
kQIcQBrMGtwk/YAeb02G1MbDQwWVm55Haw9hWOxtVPunjyOEFpX6s3KqEL98PGoBqlqEMkT7vhmR
nP6XKF9I71PVA5tJwYbkWVUEVBsoMrg2ntDJzq5DwUppAbyNZ7eZxTbL4mcDn3LwMYA7UCETnBrE
GkzH8zNvIt3xzblR97URb2RsA0Se5UcTw0QMBAK0MtPSHQ4ISrYBEzMOW+c0URChGW/TvXca78xe
c9F5+3Dwv7jx1uoE3in5KD7xEvctu8uZU9QLPXQOgH7qyKpuTWaEXK9oucQr5hc+JX39V5V6K3P1
uxrHNky43QGqJu+bg2oX1rtPSyGvxk1LFKmfzddEoQ8C1uDoMhJtmzb1jeo5yhxITaco6Wl/AcjJ
gAQ27YvumOGDhkngn4Al6P7fwVaMM1wSQtBb2FomQqRFiTDTsBc6NWvtCSB5ZwmfYj9VjAaW4EJZ
iN6IvWDCnq0pQkV4OBfTQ3ADnJr+Cr3iIu41ojVJXfagiQtrHGdfQ70ncy5mqkHGp/x2ZOdw6H06
OHMlbw7LgXR6PRgfz2rMcot8x93m46dicZjDKp55yQ7vd2C1mfxyF3bNy2cVxI2VlrcxYNYG31ix
AFcoCbSszwHH3OF4q5L//AT7kOwKVZLaxgYlPlrulsJJmKmIdb0ktK45FISXhbhb9qoUc9uiNIb/
GDQejWJB+LY2O7qRi1kjt58RwfuovlZLWycu1A+/Rhefy4d7I2no9yZn8Yh+g5sjBVu82nL8dLRm
EZR7n0ISo82UXQA6DbSgOZ9Sxvod7+5YYKC6QiUpzrtNjfz8Dbj2l6u8sZpwciDFecPAmqDeBgMH
IJcVpLIKuzhKoJcgtpq0MeAzUCfa3yF881+IOBt35YayiSYPQ/akDTpXfObMKdk9t3vBj3R23K3P
AyuTb+zXz75NLrfi8kkzkm6vJz+vE0wUMK9jMcmPYbm6EQBuunI8r4UcyOKHiJRjUPCVLLP+evVd
kqVYHGQGMp5xwo67FTiY3azJ0giQYPD6WSN057A2XLrU8wgz9XDIptgZA+Gu02/Q1GXXRvAX0agB
iQl6VqSSx3PgZ4Fij6X5qXsqDuSurJN5cUk5o6wkzjaVqUEyepOmZi2Lq33Y2slJ1wgCcoAYCdHN
CAx2MtjNySmtWuugpnVKr8j6cZFriUtaHt0YdzWs0ssz9GgAKGHpY5c+DhF2s2ZZwWEc1Ic6CPWz
fBlgN6Ks7uPTaGa1JWsdVxVPPCbSkHAehGM4ablxZCntp/RHmUHawjYg+R5aMf050J4IfvTYgMsX
/ypMW+/0kyccfjurYzKiOq+04PNmpRTlfxwnwRet5wPMpJIXAeT6lRIc/8Jil1E4aeAYOgaiDMPT
8/21SeRFpruv9lt37w0pWQp13gcfhdpJctke3HXPGWtpVpNpydfvOe3LothrwJC+ph6/KrFlJxYd
ADgTfW/mTg0/r/fni3qMZFtpPzqtbQwdjXY2s+GAwMJZE7mIN/qJ4lY2Bv05hjlW7JiLV2zrntlb
aUcmeMsxdZqwOaUBbA3ifL/n6we4HtDa/uml0Ox7SV5Spu3yRBgzuXTiD2PjrAy5dKIqcoZ838Db
x8e8Qjs5b3Vs2gk2byqX5PqioaILPbb/SCVI8nNkevCOmAMq4CT6Uoq+zJpA/RBQRp5U69P8ffzg
vW37yn1BfPlw6kUsSW+iC//nfHw5Jnn6jKzbBVnoiKVly5IsDFQ0pDwgX2DgTC4HTh9w0iEKUAZs
jDoXsaDINoSfjUU6YZJrx18MygiubvJSdP+Qn8qynt8ocKEXsEjznBwT0lQ+IgHGjPrfleT5qQHC
vgymOd3qQheceR4suADNjic6zVl2NEBgaY6HH03DTs2MnlvtkPZHAbZLiZ2AE4Zpw+B7PmeMyO0f
fYwuGgkzezHvAAcMqnDWM0QaTOe7W3PSz/doHKvod7zhKw8gdYZyNlbcl8kXpCUC6zIO54yw04Uh
ky7edB91qxjuUP3oLMCfnfOvTRhcgt5VD/ggbSMzkTDzAfAuNa86ASs1SCKn4dL75MXHNW5MO76W
iypXXdAOhsWrnh5hq0IqF7+tNc2hSVG9ExxZSzzWSQGw8/NwH/u3PwofEXkU2wFB2DJBkjSW+r6E
7/pu5JSiqPlbPyGcQG0dtOU7bEh9fhbvx+fhGP8o5GepkmEVAoWP7Hou+VuaHI2PSlMwKMFr8Otx
1V/SFYaIp9KlowqjVUhpAyxVb+Aukh+T68guK33PVMa0OMrPkDlRwve2xHVXxdiIqmoP5C3ULvhH
yoAg9aEJFGdMvn52wUhZu5yJinJfG7iLLjMMh3KkBXc2enbCnqcatI/No4uuPkxWruZZxASP9Pw+
nZIbzNcqX3eUAkopxoUXwdOvyqQWX7d1dYQCk9MJ1Ix/1ojBx3C0w+lQxFmxAt3YmPVlnMFS/ihz
aEXTaLosnEIHN+911podQ3NTpO0aBq+ulJqvzCUx0toKsCc5/PYWJVik08sWZO7hrTSq0Zs33jce
XjP22nvIJYvlt7Jo9slauF0BMyJuYI2htOiaxFL7uU6wMHVWJsbKuUWi8hwWaBIfIRh8ymQsdHNc
oZx41aLr7iZ2jg876z/cTHZpVRZb49xVRiSJHNf8Uwy8tws0ue3C15lU4utUxWO2dyiY0nGHibhU
b1JH62YsvHtlteHABG+T/lB6v87hGZrSMZ/QN5w58kfarwtZmw5DqBeMEv9WPXSfWdmqdwC6bpZ6
ZJ66BUTIFX21Op2I6B8lqC67ChdrSTLX5QGNJ2a9fSuwQqTIYyzsIr5wujHeccA9F0+NjoFBvlUk
A9ngnibio85F4/IDTdUoa7pe6jHulBzBVcNpHupvMw0UPnRy3EgDsMP7tGmomUx06vaFsjM5qqcy
xvvd+mmUWvxU17lGJKZgXy4HPTeYsTfXc6+e/ZFp1f6/PdBdEbPVyoKYSicQMes9ZOgsVk0SfrOJ
YbeRhcZYeiMElvWXdqgRObvyvtIuSBoygom2e1FJjiR7F9Uyjr/nljg4frqfIyJojT7Xse/j2dL9
Rqq5E1uiPJYfXIqgToaLimD2GxvNaFAIZR3Z5bJHD6KmNwV0G+1WEy/jaFfU4vTCPH3jx4VBoUUf
jRpqijI32H3gsktwtO0dGBgv0wzRlXIZ1UxNJccZq82RSgcP5fAzjDkx5N4zKDiyK0JxVY/sUAxm
mTefV48TamxqFbyoi+ej00+/9o/L8lef026NZS1BXiuD5bgLUK+qwPSDIK1bpS+NhjDE7H0Q3s+0
Fzw+q3CLU4MyOq0G3ilL/8pbRt7SMlvpryW4EI5i1uql3z9fPLRpdmOGQiZtHl1pLQ86MamJd0L2
EOQbHfDAcE1c2Hn9Xul3MYOFm1z1ZSaQDsBdJ0wDtg0UizhpXeVxgSfVoXQf238lClZL5He7xhK2
Lkb8WqefDU24yjWio1TiMDwxV3sPQOMXAZ5lRf0Z1GeyHaWgGhMlmYr8uM4nffqYhRTRIfDiAWxJ
qG7qZYsoY3ZRsLPwfjpuU2FmAOuKOBjpE9FINN8XRa/dB8QVYjsOTVEu7Yz59WgHgd7FKbuGgY2e
0nPz1WnfOAiNkOeGyj2sMa93gzFvg8Q/DoWDpTMnMh040O2Uq6hR59qxpGO69tF0ft1gvEhAYFEX
iZ2sVzu9iuSoi08aE7mFyhveK25NB8S+MlmBV1r6i9ik6Xb10W7aCdC2jqIUSe2WSj7dh7AIsvrn
VnitgkGekW1ZlcvubTC/A0nhDcO7l65A7TxjGQArGm4q2AG2LOsSSYAee32vssnQAz0ApguoLi59
AxqPsKw3YZPKtmPLCiX6QxstGqB2xpW1E6aTmRhl3RxEYzOur2jouRrG7Ij8ygyuC/XdthTBCqYS
X+pbr+bgMC4uO+spNNuuwJXO+88uF3FxmMmCV5FyrgW3sb08/j+Vbp9J48DWUlQZtDwFN9k/CFPE
q7CYJAFRtH4oiiwsdpnIIMP/j9f1EJwBUJFLTB+2eC2/VIhtiPWmZgEkzFFBszy3vDkz4xJhnsCo
5qIM9QaAeEYIkSwC/QXno/YANYre2Injm9uEXb6S39pznzOil+VPR33Ff7pWU+d5lg4swxjAYaWV
2ogX3zTGLP2Ci3XU0gQKwxfPVik9c0G4JG2LxCuxVE63ak50rAjC2/e1l4E5sqi58TSvETsmHa0Y
TgD1hDvcudkxkh0s0j5TtCcUas4AH1nyufIjvI7irdobyjSAcSASKxPwulK48k1NEaYGMcRMAFR1
Nh8KJsdsLdfxihr+NLh9QoXaJ5/mwedU6C/rEZTI02MCGwxscZalim00b2kJlV68aWy8jQkO7fvS
/ltpGRPbIvC748Z+kmWhcKGjRC/tANMb7pQlnYSyLAPDTbCZJNXmGHIOQeTi1m0icr9Whs8/UzoS
DcMWDy0Rm8RfwrEWHgAF25TRKhuxkzZMvy6fCqEn0HCLrvJeHQGmcoSUMxct6uqtMkkgIj9ox4rR
Le3uB2Mfgo0aFdX+tkPSPHkhxGlJiisxKtkei8XCw5bM8kW1YLOT/S8pDLddDXRqadxDSoFQa15X
OsIzt/rPZMJirP4ONVJYRPn6ErpzluTnMGqFRQu99gnbsKARwfzPsBb1iYTv3EhlpdfhQkSCxbr/
D1LWGL/Fv5ZJ4kICDsmuucZnXTNA3TCPLnhikxb0Qnd/9ObUsDSLbCgXu4mFrCZkYy/nTOXJ9uef
TibWLRNyRal1AWApO8+u6uzbhp1W56silKddpuuWZSP/j/g2UrThDkKkBjXQ3V08ziB/jUAT00/f
zvTyn+Sa+6pSYpqVDWNSUChF+gmL71SJgX8QjuoUmSnIpKuFgdNOqI2Y3UZN0icEcCP7/iXvs0Lb
9QQEb7Pe6dS0DZsoUHDXHp37Adu9bqDmuOvqPJQJBsLSj5HtOAdd3Pm4YWyTrFdQYV2EG4/a6DQt
xAGIo5ZkvcgRHJBGk2fzknyJWW18BIkTLxvbsbslPuGfPB1E2szQNbbky3Oy3TUqISkA92tSYdu9
k1IQLrqirvkhWJtB96Mq2yQAnYxmEwPI51GCVyhVZ6V2J/2E+FqotVhb5JMPfvMbMfA/CcHprDIm
hqjp68Lh8+7uHj72gij5JUx4ynnsA8BLonstidorcpzvO32IcoDRL/3b1SZrfYgvCK1whD2lJxq5
oVrTM/eqyGLo1lqlQLR80FejWOaBGQuHJ69Z824t49WmFDqXsRkGEPIvyKnUIrx2lHnmQiZJ50Qk
95CQNohMI7XVNdqZ1HBGgtQgtiyyCkf2rKCsYgyIls2Dn9ODpVCmfJV1i0fnbar8yn97DbCALNSZ
nEQhBQINeHmlzMzFMZ4v9LuVbb+yfwq3DXCfseskB+JrpST4xqY5WMk3zgsRA73gsfqlLXs4r/aW
vqAn9JIj5t7lZmP46nlhkSw0CxkRiQaUX6CTWgvxjdIIYWSotYqs57D4gfFm3a5MJVPYgooWgW25
rC5e/z3Kw+t86r83qnmQIiuO8r5ZbxX8VAe+/oUObtm/ZcV7o36u+JPw4HjKV30yQWAuZyZnjZrI
yaSUNrvtuOnriJvkFJ8EIeMLNhNdApdZs5X7kkdVgViZnKuWtZebYM3mDtkIzNa1Tfcva63Nz8QP
cO5850henZCDzTw8987/CQzcIALV/jROwVc4xwmXK5bO0TGx5sNK5SsZ+nnSCu4hkgWS4vCA3wBp
1Jf+2FC5j6dQe6dOcqYABm97uKB+mV52bts4d71TQeN6NI5ZHAf54mZznbX7ZP+WkOFukv/uLcsQ
ila//wF1B7GFsf3sJOPQwidVbdf3DiNt2Tbgx9RqzAG7f4WkiNEDo1Eqp8W0RkPWr15BoDMZla58
mbPBG0dF+lvMcOws00WGCRulhDgDeH+3EG3EbTLrgh6psDQKKvqbI+gbKQhuil3FitvouHuZgxzY
kdemRVa0NPdI4CP0pMtBtiu4Enhw8e9q6dgeS4vO2jG5DeQ7/dZVq4PncuLvQ1KZUxkq754WXsxa
I/xEDjCSeW1l+YGZxw8R2y/oL22qtQ/5sMgZ/aMq77UPcq4Onp+6d5FkwEtQhJYUQj7FsCurR9Fo
Vu+y7PT/W2cRDc+0hbZUErVwOCh/fIGadLwKXRjwhmDe8lheW8w4t/wTynQ+VoDgzVupNvD7k6qV
6H6XJbBtnGVSLCXyA0zivUhjlKzKSa8pcGNspkJNXITxlofGnZmB08LLeXyIo1qUUsfGTm8ZO4Bw
63Eh9MtWG0lZWzn3fS2thAIGIv2enUwpRZF242ztUr1Rdp5sPWHSjSGjolzbIkOSN93yVJCZQY4C
tXJs2czQ08tGn1dwQQU0hijFWk53+aN1F01e2nyqMCtRXtupc8+qxfdZPR2umVfzuAaYbskpP/dU
TPZnIykr6SPXYTDdSLtndu2pOffdPGotz5B4ws8yZKKdsUxoxIRoqIfEV97d3nf8xNn5zkfmNaiV
WKAXq2nRl9HZ21tSjSIJD34bo81EsUCryApA25cZXY+nZ8B30lxCva9z4HG4/UBpPSLWbvU17Emc
JPx043FvWioaQ6cX7bZHqHEwq3OJbHzF7nak0YhqY5nhYkd9aK9PV3K0a/UCC3YkvesTBvDnXbgS
jzi9ynHLcNWf2IlNtB/PwfNjlS5ybJNJzl3IyqVISTmBFzStZZDh30no2MUul1QYHTh+Qi0/VLld
bFSDAvo8xeK2ymdp8KyTIn74pl0EgB60509co7YRhLERpC1ter9J5QqREbZICCe6R9IMUlIT7Cr7
FrPyngyJiOoj3Tp8ElpvV3D+OZDgy+HQOTjLzJmXz42bko5+SsQEVQ147zc1FwpP/aoA9c9Y0fJn
WmPZ11Xm6dh1oD19IRiXvfeJHYaExH+QAZQKK1bUMD2+pDe/U9ygrZszsP3zwtKPgUHIV2rMo5x4
WYYSzGlo8u4GBBujpX67oyMcfdzS+Vhs+56mo2Rs5XCPV4fUYmg24hiQIwdJpTWRMx1a/pYUhoOt
6AIH4uEMH2Zo9o8HD5fy+5CoVfII6x5+vNXENTvlfBAVPJX7g46wi+++zD+4g0yQTKyss+PK7f6z
Im0HSEVIY6UqGq++RwEwMJyR4oks7Ld73xvLs0zQIsbdbJSQ7vg1blP6KHK3HWAy9CGKwt3Ib95Z
2Pkh4scG+U/SRrWuIpE2j3iKPDrUAq5PgVrLKOMnLL+Q9D9HaSX2HxCNex9nVKJDDd0tl8eM0VZG
TmTShVq3MEVqPeMsefsEXjKl6V4jugQzSEoyRUpazy3kgp22ls5uLQOlk+Gt0mzxrhlnQnaY7MQb
oYqmGssJr54pDFRqSMxc+d8Xql7eA0a06GvCg3mrcRHNP91c7EzunQx/gsF3tQDuyUmaTqMAu6zN
NKVmm9sj44B2BVXANyUtFK4aXbvzGayXfbQO//unc1uWfMHOsDwrE9LJyF73xr17k3Mi82998qF9
reSC+RJQjQ4nb44bxNNLlXfiS/tj0SDlqhJoznpMwUMuRkQL7mwxCM634dawIRkTWlLGOO3aT2s+
diRjJJRHU8jE9rKF4hnKHhUSgKZQ+nYe4naEneufJW8vXr/SSDCDjk8hYYMo3g0JZvp3RN6YwNXf
rHyKhlo4Qe1PbaPUiraW11Fj/JwRfX7t2jNuR/jHw706o2mtLmUGuKDwaEAiPcQGJdXd2TVRqrWa
AmTYl1Y+0o7dEoyMYop8aAMauKb5IlGNz12nz6gXINHxPCv0dGbEPB6NWutmu2i4mG9iJvk/p6Mc
FGuxjcrYt/52Ol8eKmtdGAnIM1+xSc8QHFyO1eOtCQGs8RJz9hHSb5N9MlOqDmhcAs7Rh1szdEoh
5LdEMolxSV2MPjHzIBPXGXCjwRO+n1D95znHJDk5QiiQw9yS9NoTVhm+5JkvGm4DuV/OENcRojWw
1smysxT7i9S/1YVfBorVD7t24PX0ny8WniXT9ESGFJkibWSHX/qHGfLGc+AcvU5u8xG58ykfklDo
AX/D0UbV6QPqnHYkz8c791MUwkkdO9wuOpBffklyJf6jJ7g+E5MJ8AQx4H4Yu0xEs75UemvYB3S5
4F475W33Tg1yTG/F29FFus/jo746sQg4VH+63owTaiyYi8timWCSjBMCWioPEEYFSU8FdHgczC1z
LkCPZtlsc6Pf2lcwtFrM1NV+lL0QqpLKiBg7lIkNqplWjVQ6oKnce6cyCMKJI86W6V9KGGK+DjEe
+nRKj2fm4q3ClxdHxbC9O8W2nOQc36wkusm9PqiI0zmULpZ8U3vgV+j7P0xs2UDSCxOr4gxzCNo3
dayrMl6o0bUOrjkuPItQuDlyAwZbH8KmbUSmjr65BIRL4ASprViwgMkRsouMxvpCZs/yZu6JXCo4
GWs6MSwG9nHzd0OykmjRDqCzSyJguvwDKaw5zWNa1lKNiSylCzP/ccaZRhhcoX10lK8vJ3bd1mxs
EduT9v6x5KFPTGxnhB4ySBxTyrZb2I+LxgD8hnYEWnEYFFN1XUjFhAmI6DwKcpuQYyz6tZBaad6g
IRHNxUWKAQ0wCGrhJQDGSO5OWOa/mjfCBGUaTrw+3Z274vZOJHbkZ02Eif/DYuWKjq/A4/NvrJS8
VvMMmibRQApXz5KwytR/t56yyUNTEnI4f3cKxwI2QS7MchypDA99pzVt1YN6QBllFs7i5LRWYtXK
bkQzVka8hOehwYfcJRfzFtydGvF1+eyNYHpO3ubJiJXs0ShWMEAjR1xnbKoOV3wYsg+OumXySzLA
ynyaah+livCsjhC4dD28sY6D24sPgWEnzIt++PICKxt6ivX4gtWqjobg8rHOI0/XSre8wj8LDj3L
hNJ1Pjp1Hz8EKG2vc8mn/T9TjcaHPv9JPvFaMa5ZoIJOhSwuFL7IYPnyGOWTpP5HEYG5zs5sR8Gg
DXCqUGSP19fliVNEIRpbJE6SmPOFKZZ5PAYK1C/OqcXhqP5HVFz5vStoDZmqTm3IOMQai6wmcd5m
jz93AakacjZv2HyhwmWsxERvmSQyz49NQr4Vsep36bp4M93PQc66JIbbRJFw2x+dhH+SS5yYGQeA
uTysi2mYH8VEn7qd1p7OkFBzoewSVQz5d9AVFPkjYobGqoFxeC4Qjwuwe4pAAzZvn3rMy2XFviYb
JasSj6BkrCKoaYuxZyf7gRDsJSaexjGHxEATF/T4uIBY7hY/FXiNaluEXWp3/dVp3YH52rSDVNvD
gDPlfAw1kHz/fupJAoWNzMqXgUjXEr2Eru915xX8GIpp9TvQZIYQ805c6OKPNSXPdh7GIFDT7caQ
kaRvjqpipdMJsX4HPabE6Brljawc9TeulKdEx091WvQVSvKTy31mLfPP6RtN9JvDlIYcqB1e8Vlp
dsQLxph/2Ge/Dj6TkpWJqTmwSHDrVvgsGIaavxuCp5IFAtx/Z5oBhJmRTFmLqnmHSHEdZ0oVDyUM
t3ISugDXjVGBSrUAzAf85MixnpB6CLwRBj99o4p/dD9FyMlEPbXStBR08U64sKhBlBHuDafpzHPK
Uc0Z1vbG9FG2N6DOFUqSI8vEBZHuxNOndEa3vGce8Tr9BrtL0I8Emsah/pCQcqVPg8rRYs1gK1Xu
JNXoDF5MO6xYASWyNck5M43OJFY/3DiW4P9WNtgMx4ibjYnLlg5mL6myD6YtVJMyt4WNFO3u0syh
VHvfuSZbJpBir22REgsOzXIEJi5NnEruvAXj9NKc4UqsEcBoubu0Lk5JnZIMCh1fGn+LCeUb3Qbo
1i+QKKijNPdNPADZPYxSpEnbDZpGVAEfQMbQvkO3tG/sViZ/+bwttL8lFc7LMvKgAOnanq3c7g0o
xQENg5UbuwToWULIhvwNzvMOZsKgIBtbZDBPTypxU4dSiyaEovATF2koW7HUaS+u3fREyeriuHB3
Zrr+t55KwIu1KL1B/flB48XSWdL6BJtZDv7oHex5qEsh+e+bqT6W/A79UosZsTueWt39Y8m7vqk3
e/caVhGAZd5EX/flXLKI4V1ZIMOi7KMwFwS3zMkUcDZ5Vl4Ryy4m68ZaI1uIanwEpxqd5J/L0iIg
ocqgpjdwMmMAqVK3HLut6mRLtP/uYerRExYGLiwezo7K++OH3ANJOw4Hw8kp7LCMCk1y/ti2r434
Gb3R/htl3IFmaheSwi55TlJdwHN++ZIeBO3VEtdc4Foy1gAsLwRpMzp4BmSRq9vK9vP2RIw/hluv
zvCebhVfgj6JhPDSJw8vnyfIYL3N/lXJTMFifCkzSovcScuGWQXb7Mq/lr2CsFcoxiEMyzQWTIfh
sYHOLKXGcObZtSnK4LSjLomulBma1rlmFjJeLuHysbK89cUltnqNoMCniABUc9hSPRX0wIBNjeRf
GF+xY9PyLDGa5u0VSc2tPoxyXs23h8zUorg/6FoiYJzDYeUarR64KwE1P/OAQgnrDljJx6wEDrSS
201aZzwGIRZrH59oxzW2wf6qpkaTlVgc8WPJtXQcEahfnI7pL8s2B1EbXldKglfqfnedjlEc1FX3
IZ1He9m6bTNw/9t5OioclaTW0JF5y5+W9khZCS4qeg36/0fqnJnlIMwDozORfD34C99ffqEMcMQR
mpenAiO9abVj4apn4ZZVS/2xKj7D5kEdVXgElVcgqBeCSqTo9GuCGQX18ylTBpPPkH5QK+U1xLFu
5bdT8tU60+PpW4NLUjRzr4APomrU0InYmQ2Ms29AqCZoA++1nRMXx5V5PzdGj5yipw3SoQiYSYbR
SZ7qlDgOgmK7AhukZXBhrHQORWt7+kher66AK4bvVk1z5vKoAC0Erp8pZETdaTNJLIE9SN9Wb/uv
yFAe7m2lUsjUZxoeKHuw2d5IRmidz4pyJSpDSW/s1ShcXOhNzEhhaSx3UoSAgEd9RzfR2HrSqEC9
wWzHjWwrkrw77+yzFgmVaiExwTO6lSVDH/1Tx4a0vaaV9Qg0rQe4SYknelkoQZjbpVnHotJRU/VY
jX8AUC/educqxBONWC0qMK+hjb5fKk/gXFX5MNT4ATy0TCxj126N7AzMoSQDXh8llH3k0XeK0iE1
0e0pFnlhGRCDCgox5iiePkm8iM+F1QmZ4AzZnHmUWY+XL59FegIx/VXZGtwJRhbP+CHIG8/RW4pK
jQH25RvsHTHAV/SV1tDvv9p1shyWqPYBc6ylJlPP8YtXwsTbso7nHzt2y9+qW1ZDaPL5joZiVT9p
Z4knsHBEKLuRs5CLmy1i2ajgMADolClawDewu/qZi5McA3+azhn9hAeuVOnYBh1ClSpwGjwerGBm
X9DFxCxjaSAC71bdh+rop+MR0JlVrQyKWwwFK230fENKfydwRzaCHbHwdgV7UkJFpjva6X3rkro8
HqtZNC8h/qHswymq2c74OzrinecOVswgi7uvEha8lqzr0E5lgx+R1EOIrx8ZWQqWM3TJyYr7OGwT
Fr1X9p9OlLoi6fX2b0d8vQroWY2e6n6wj8fPYejsUTHurCyYAZmZl+8DdMuGRoIRst22oesX1G4b
Sc6OJ/25K64aaBZkr5pIQ/8GwLNaso+KUKq0HAklozgT5Om+GpynGUcbWeHxHzTfbYxrReJBJhrx
QqTIFpVBpv9CcjYdrd0so3q0aWUY0VBm+TpmhIhFOUXvCW+mRWRCmiFrw9M+vk/aWScJDVXOg/Uc
3n9ypdRiPg5UEFGAbCmgCYDVr3lce0OtdJ2TIDPZcJxF8jtpB7Su3vLPzB/aD9fUhd12O8AmfdJW
wdYeQLHIEiHGVH4pABTfFxjxnKATgVgrXrkNqBFvyhTWjO+/ywyQx2sBYNuEyUKfM4NV+Ou7Zn0B
j0o4WoOl3D+iY6IXszXSbc90IgidH25lwnb8YddlJ421fesppMARHXX7JfjJnW8u9PUFn5NJSLN5
iFXzDgphL93/WODPn6FVVgTTErsSYK/W2yru7L1Unep2qqreCV7zCJfA78/KpHnzUqvepSqQR0st
aeWrwrINsXk0fIVj4Lfa6oyZfanhyotWzplnLecFsKsomQ96YjusKWcdtwQb9VmX6vbXXogusPob
erfkmiCG9aadhC8bUvTKuE1G/nWkz9RwxO4c6DX2KS0nN8TyA1zKXtg/UA5GeNn6qr5a9QERf7GF
LJWAwgCWpP2LhkKfxvHee/RFl+ZMZ85PeuDcpGa5bTvtwAxvXH+Iig+oJBzSoQwGJ9f6/K7GdPfm
FOysHqb9PSg6J67IV9Ys1b0PgytivxiKKE2Qsc5tYNoVJYRN2yJ0KLBpL349mddVmyPiijWSrBjf
mCXf5u6MW+tYqtYG5a0FybYppZOFwSJThGumEXfFlkWojGyCkjPbHJjhZi82mXlfJzSp97iRjiiS
opHym3QJzcWQdAs13F3brRq3215rUcZ5S6+K+n2dgfnXfUsmd37rogL9+Cc2GctF/xt8azJ9NsID
u4Qi4XTHizwFouhJnTzx42PxUsZzlPajksiYvh2zrmCwxAHWNfsHABHeeJlHfegbifj+TaKtHy5c
L1TTIRJKp6kSA1MYldV0FUCRA43gKFaQYhZuYvcyVGP6vBOjSRepDRuUloNFDySwq/fudJIXKatx
VZ0YMbYjKjUuo/QmMXAmlQRUWt4Mp8KtNkoXxu5qtgPJBmpa5EVlsUQks3gkxCdNdSIEfnj7rdK+
zzOpiBi/abFh6HoqeFZkYUlAAR6Nl1ancrI6MGO7BRm9PYI7XsAmNy3jwoL1FMBX4bKrpg8XHbJz
/NHb6Xy9sismguG4rlfFBmITfjhKUiDFamFxu6IO9iNbItjvB/Mt4EVJJ99rdmEqYrzFdidDA1LB
KON/sCnUKw3D/C6rFuGYky93xX0wEHIgkQ37p6ZTuXqhgrfIwN6zURs9ZQhzwzezmxXCjmLByodq
zUW4YUVdxezLPvCcLJ9a1zjbIGLowXO/Pzsofpu7aRnJGhFmeDrbW3llAhAJwmtn2gsLwsMRSbLd
YIgdMc1jefcxKW5fKUte/3wFG4FuupoDi0xi9in8VEHJoBt67n8xZpHRM7ilsP+pqyfoZQv2Q1Px
1uZZjtxE3fwskLbRO8sSizTHTuDaQb5YPVu/lXK8SLngz0mJje4r1Zra3t+YAuiXmRnNxTsCGXW/
ABnaWiFONRI0J3SUN8k/gXWiTVkKm03pymuP4qKeJWx1OOyykpgiArwZZnrA5sORW5Fa/PEm+DQN
U7+an03/HYXphqus8t1dKtYu+v91OmtNi9n8raIZoqmWkY+gtRpO7F5ky3f0N8iJ0yU79tLaW4Ex
Un1GqHy273la44HKYCVhNXziMTIwlcYYbg6nHED/LfieqUSwqXAPztXWzG8Jd0QvjCuhD8eJgvdI
bCja49dae5oMnoFjxas9k6tpOfuXOksH42zccoFA/PmoR0XnRHexWBN0NKioOF1JA+KLZLKc6z6A
bvppaKIir0Gk7x5grTW0W8kURgGnqvJYcqP1MkaYl9qKCylZgC9VTazbsjkWHJjJewhCplAw/57P
WWn9qdA9IxmtBNJUNdax/YmdbjFwPoxTGEHpxmJhX0RvpMe0Mg+bH9/a88GgBdu69iYOAowiTitV
7KW+VI+Diu9LT6mSnhafErWeVY7LqTTflqnsw2VrlJNZJNhFXmhq5l5dzo2Jz+Y9ZGkb7S4DwyWz
FAv33kae6oBrDq2Ap1onRNqMIT+IM+TUr7qY6tftw0ZcHUogdbbOrUFnHXlj43ZydvGPsZrgWF48
07jKqBcSS1EHtR8fdyNOqoxlto31pxg8PXtBvhAEGl8zt3hKRdJ3LtY0+Pa/z0VHoY/rKt3bftGF
za/VxvCAoDnlFgW86vQ6tvCuVKk2zlSwB7Rijqbv+6KwZ/onK2ehIxyIfKRFaIMsjppLx0Dqa4wX
7WAxmD8Olq0RtKnfcMrQboj2tQ09CntJm0qI3HwdszePlgCwzjKLSY4cxrbo5QefQlrFGcXpIFa2
xeJ8lrCy8bkF/ca1Nj8qeio4os07BjYnudBo8Snk3yKiY/8cwlnYEkkKHMlWqsYbPnOeI5YTatV4
lXEpYMaGjoKOWiTDTFUjJ168svJQfZQ1+gbaasdZebBuToPYcnrvSlrvhsdL35JGk9fYcfZWl7WU
bmOAIroBIz2W4t6laLozUwmYpKYmlVxsoIkh1M5DNXzamijCvYEhxXqUh1V4gle+QvAVSln+ODpf
Mj7Flno08T9s+Era3Dvb/1gwZZjp7Km++Ej+oxyzD1k7fT0uq0oEobTo/k9feOQNtvCEZUWec8iM
/jlWKIQSt9hIkjvV3EibKWx7lLNUZLbh6Ohc775cCpv8SL5CBPMrpCqZFwF4lAr7GhHuvm2/MgEQ
HJyK8h0tpos/FcELQAcXTfcazVlrHIOVYrs8kBR0oKjCB+BDA+xG7iys4YYh5DQN32GgKzSEoSrF
iUDy+ypXRRVL5t+dpxFHBkSXRYjcAUYDFQ3xEJdh7iFbaMIcu3g0zhb0SUSeD5v0rOCrrhhaPkFR
Nsgm7J1CGed9LDbxsa95/DwCP6ZraU2SOiksQD+rtpLJD+pCYF60oy1HXGfxIDvr8CpN82jxGaFF
GBGoGn1x7i8BsKex2SkZt6Byh7GSv1hnbxax5mJDm7XYSSM55EQM+NIClgiV1o3+14ZMR/qrpsnc
NBTgGHw5F7AdLru5f1YmWUg4e9o7DNqc2ZsMHVbgxXT7fIQB3qFoNZkSsb2S+ZSBBTr0FuXeJF9b
sv9cqPPeOzyyjXVvfNGnCndL6w00Obh8YmIrSQMEQZoR+vcb0Snax2J2t9LQxCGi6rm9O5ohCUtE
ef8q0R8Do90KaUKFjvU51uSULw3m+/Er19yuFh8kSSHb9ptkeadu86mkUSS7ARDJr+/oGTowAFSD
lWLYat1rQNdSHGCJJHFB18xwC1S0THcKTOGdmNAG3Ya0VLTllanS4fNgAlxbYYa8JPrXXrybuJ0W
sodpfVlE7sU6gabOZYIosF6uxVPe8wqD3tUfRsFMC4SdgmSw65X0YalprpdL0ZqAA30sEqhS06vR
RZRCIGcQQhk8ZZEIGo/yJc5DpvQ21YiSqHHaPsBORbGm0QCrsulCPoObsQhJRePs5myQ5E4vMAGA
YrCntBEC4/Juu/CwVijIWjn6l2teusr5v1XaTWOL/cnZg/coPE8XObydm/2BQRBAI2591Dj+B1Cu
oFpdp0qlTWjaKF0XkfncBO2BCK/OTON6FHVHesVLU9M08dU/cBbqn+ucKXfBFqBlpYdA1j0j1LJ9
cMgv1fSD455PIyHmAo1ODDTo8bKIU6VA2YbTbyPRoisuJHpunxjTSWWpkcypjA6bk35pWxptSiQr
9JOMpKZjp77EW3hNcSZhgxYa9TsTPV1FR8na4pkVN+Cfl6EuadFLa50MEY/od6ucZZTcLpMUzSaG
GKTezfTMD2n6iYE3d3I2nzDTz64vYjAFEcEY2CTkZeu/n80ATxksvoMGWMrDkt8q0D5eDxhYI2KN
6BhevCVVAEbvoFgH1y4eeZMVUu/3qgrOaIA7/2UqOq7cuWqnkJOa7UoVgbjWx0gldOlsKXpuxB+y
bKXx2Tm2zCVJ4Y2fxIigzLQfoeHFtcY2foNoJPlijxl/lrs+dkdArjsvlwPVDaiQCx/a9aNWuvsJ
iFQ9T42Nmy79nTTNaFIPr+eSHW+UZ2E+UqTSIaBct+6PIpCJjahV3oOGB3bYbH668NA9KOPqCv5K
/SYRg7pQd+5guvFFJL6TuFE8vh8xO6/P6vEbZ1yv8iM3Jpf1wQMy7kDz2i8aMrx76h006AA2gL00
sY19tVBxob4ubZdcRTw1kuSC88pz1yoL1vnSJ5zy402tm1O+leiygWCmJ9Gy0Uz6TGizFBMb5BaD
M9HDQwBHLLauXZaBEXtQnAqiVkxfPFaodn4ZI0Xu9TV1AlnMz2OotC6zIMS0jz1BHKKvI0m19hlb
RYv8ldRIopFm5ik+L2Zv9ViqewMltG67ahTwCOfyTomBbuW9Rlk0Is0CSH5fMMlnbtlfiXkUzTik
CcT5Dcu21p9Hk6RlO+nNif40kYs4HmYIu9qZvyKVRx5w1s0ja82h+rusCriyYTmmTxge7k3Wkgix
2NaSPaODJyFC2ylsHpr3nngKrS+aPtQCePVWu9P32ZfGzZJstuOi4xmrClGg4cEKQ1SQP+z6oAVI
L8r9zy33twNXDy9emZGM948afyKiaptiP8pyRE37PcFA9YbOMHRmlxHUqrHvCFM/j3niCKtlAtB8
/pQ7JyuQaI8a71kW0OKX+ztE8HtBv0nWOSEcpilOEWQMmXVYunJILOXwt8E8hEEByv5Qvf363G1x
+XWZqsjWIX21UGAfe59LPjCNk8j5ue8F6e4KFDrIpSnJJ08XVkTq5ORtQxK/hJ2MdTYk/0n+h4ea
dxVAfz8VoqM8+ouhUSYJn63nltdBqxFlED/ackEznH0S2dqQzT4gwvVajIacDB8LS3M+6HV2pPrk
IDmSPfXKpE4Nxuo0gdvFVfiiRhVE7qUM7fDV0kjze/3m/3K+oPWTNi/Mhpp4BT9ZEvuo9X6mAsN3
7TEnkBCobKIUVWVBuRmUJkZ5L5wR1rGXpYR1loeCGEDKN6f+NzUvtIhPf2SB6Ok9yJrnUEvZnsVy
SUe0baqT70AV7MZfMMjJWvoX/MdXNaMhyVXDlWI42343TITVX2B3En2OijdzIGKRGZPZgefWFmdC
RraomMm8f2PRUIc7shG1zvz0YIs0oqEn4TB2yLPbOKkunfhXfh9SyTXCRqZhUOlOmNb42JfXygl+
p1dbS53JKBc/499qrKiEPdVR8ggeDyE5bxSVxRrTMQWMxR3A9EIp39HH8mb03IYmohYayKnGDyWd
doKtTqlvxQ6cGgpcE9yAqVksrRDSmhh+eDHSln9zhR26j4yrSGD/qipCdEbOSipffbOX+aKAdI3T
fzzJ0Yg6jeYgsTWFKYNSBbxnzyIQcMgwyjGF0Y/H39FsKp8SZvDGiyv/2Oz/RCWz9aSCW33u7tNL
6Q8dDWRQ3MJoc91pxtLZJ9hzUfUn7vLClgTR6MNTCBpu1NoDJXAciYVQOaW4x/BoDBGWOJuNjU1R
IgrIHFbTf298yvymu5B0qnFEes1jyJIxHBhFDdY0DPael3Iuray9IusgKDq9MsRu6UK/Cq9Noxe1
nFy1Hcgoh44HhX7T3oKcDBUakhkYmDuxypTR+lvphICdSxV23HpkWLwqzGFSZaRiWXGhFpyIOr5f
66tbaSb8gqYv/cdKEhN7eVxe16Zo9lgTvZwZEM5yOfnJe2PDW53eE1tE0on4RuMuGfKdfnOQ3Xoy
ui1L4OK6BbRUWQgHiYiPh5o/CCzu9UhbtrodN2kyOGC+Hp7KqTwjLhWoo9MUNaxQbMBcRdcJ4vsM
yG8cpNLF5/8eUxlH9XfFXKNv/db7niHX6MbYoGwzmmcZlDUmAQwV9Uk4uthu7+TWZn7KuvREQjNF
iYLI+BUSTj+GxPmv35BowM2Pxhybf3xjOJIdbrtsQUgCsjVHcq4VcRIOE1irPZUrkJZ9aMm8tZGU
BTPGOPbnjP5afyEOlteMXASWEmLyUE49CPyRI7HJvtWB6C4/PokHPboh++tFkUyvUN2D2opIxI/d
44jUhQ1hjjgNL0mK+D3RZT1Mg800/jh7/0iKOQFfE01pHfZAkwjwU57/jRfGWFihEHjb/NKmIdmm
oUzK8gmhJfOkjQ8jrSvwFij8i3NaEbpOlvcEiGVp01+IfRv0tfa4ivWOU+SEDp11fHcTxrGTKf8p
tMtfs3WNiuVQC4BPZ2PKT1t90oerj298+YKVgUYOX45WwvFPji3rl7aZl8XyO0D4OUj5cVg1twmG
dKJwYDBXJ01sSFzc/+MnD7docyP7aRvOoSIAsrBaXwxRaOEzLOI7S/Jwnz4MXntvS5cRkTB9Hv8G
Me1PxzYVxWMvIWhkssW4D8D6z0FxMAH+7OV5XQjJ7GQFQUVJczmNYYH1NvcZ/zzFd/pNFVWKCGp8
1URjIr1BzfSoJgPtTrNEcJ0UqaiK2x31a5maeF9IyD3wWZkykKc5byUNGOWKphS+lU4TF8l+M22n
L/1eO00nAlF1XcOkKu2wdm6iQZwCErB1rMgdKh7BTODtC8308KBeBobyydwFSlLdorDkSObUvcYh
05L9AWhQqFALtjkOSHcPbxhLGlQkSYjGLfLcs7p+vhalwC+DxO+kVY+6RM7V83tUbhlLA8sixdg9
IoZdv4Mp0ag870xAWZA7SwpgFwIzHdOsub5YIf8j5YihhN+RIRxWRQSADffj5GEmkf4WuytALxoc
tnlLNhOcWQT/VyC/o0FcsbZJ3afNCnqso95PNYtxAMspQGnPQftfs/8LQ+aH4DdDefNFCnoHZnK+
S0Yhc1NWTfqKu2gJ5BU4BuuiFAz/oJ3wSG6/aJPF8zgoShfWNfhFG+GB7jRIJreglIaB/1xhhOOZ
/nKZqulTfxat5mryR+lQjfuZXvHfNsGRurCldFDA+ZGmaG4bDf1pO/sJMiGrcIIc84IuoFfeZ3Z1
wM6+9lLoz8LlJkbMe9j59t/dfNI0hmpiTD6+bhCLRZks+g49u1xs6vl4FuJYndd7d2pe5+F41R/z
ZetASYpxNQWX2LMJvVPa8yMiPiW6g/gPpfBxyYfr6Bw++Stjy2hb6gyZuF2xQd5Mpyoioto5Zr/F
gRig1KrUtrLg4MmHGX/61iLjZMZxCwKr46x6p3XU2Slj+hLSeR3TE5X1n2KsfkVs737OL/SaVlTS
k1tiGQDp+cyH90gZLjXLyE4lx2euy6zSPpEFUi2jqGGuXO223UiMilDNFGSObx9ZtZyJR1+k8zl2
HJNusma4Hwzp/zot2jcSCrXvkImNWbv0tSkxPuYUkFsuLVP/GV4DC6VRT5ZcejW1xCyQ6+1C1Wd7
/lURULFKJxKdrr50jc86csutuS/t+yrvbBde6B8O+Ka5xPjzZR7lUqqh2f0X4nDncZwxmkpAS8WL
yYjbwrtqY+tMbSk32MEWvBkDhmv/SsZmvkII0tCJqv+Ijel294EkhvwYgaFam+fURMC4ZE8/TKM+
FH6YZAaU9y00TnvmHvNWpORMOVh+UzUa7Pcg2t0ej628N/Gd6YRk0Er1cNbJqziDSlL1Z21YkoZb
m/lOSnEW7oz56hI7M8U0v6JhleBAwOpK63jU1dy4CSi1qqAV3LHzpmS560IQLQ16tpluics7MsAP
nka54DogYbMuKh5afe3fgvbuova1TXjVsAtg/1fVNYG2EfpuNubPJFxGCLJ9RRZXIyuwbJ9UmLu6
seCnzrL4t7JJt9mh0tSI1Tl5hB073dVYxsc23Wyx6xnwyV4smTWUVQC+72NfriFxYqZvM9cmINej
JMVO90an9SrKWwIUyRTcEA6IGp1v9ohfcBt8qVqYedhMc8/HnvyOiLEbNvJVUVtHMfjPs5R6xv2S
D3vZOeq7gKSDKybCLJeVbg8t04y090Nmd0vQcEIvzzKnXDLhfWpneW6dpVPuCiPXKdAqZczKXsTB
3oZ/cEZt8Ry/3GDXFvaQHd+2wuPOWPaf91+vvkw5SlZTRNH335uaJSueOxxeNdA96yorFJ8Al/AD
Se+Pfg8LA+eq6iBkHoCWboVmPzw0R3Fw18Lzx55ocoxkrDQeRg9TFQO+topHlGfxe4JtniS1QgnZ
9UbwYgSZLl7AqWbhnCavQef4LlAFl65PhQvLjf1nqLvhctyhSIEkRDGuBCjsf2SIeYLj25qs6r4t
b8r31jloGRGJK0Qw4mjJBOkHFfudkcKHqhwnVd4I8SYVSMbNWMtRoRaWyyhIbC1hHguE7na7Hiog
UrU5S/vQ+rZOD5izfLJPsCERdd0Aj2yNeY+DL/iYV+TVNvCb4OT0mHWucUaDQjfhC+ffdLqjhxZA
spXgFGBaMmCfMVjcScso2Gk0bCXrolpTdVkx2+v3mnNbUEqQcH75ZX3sQvY1EPgfUh4F8TA0k9PB
98OPgMKxQgOKjL/IbeQJR44wfucyqEM1vR70cMMCSIoFy53DqsxbCkXjRxas687ayGDOWsSc86R4
B3TVJ7iwJW3NA4BthwJPYNLpANrRf/0uDrKGTHaz5AqKILVsdquNIHBmpXfzVroC/mYdFx3G5QMA
LL6KOcUte0r8kd0VK0l9+4J/t5uZM+1WafRtT4BxE6LyR2LNYdjiGNNk4jDr3QNjarFsQXwX1fYE
T7I/PfpYXXPNG4+Ai6iU0gtfS9dHWOGhslpUdDJZf4/+VHEG2aKCW2Oj1FLTRcaeFLrS61YCAttu
PAdIP8kQygleS11iObNX1h1OauGQguv0jy+NNs1PaZsy64mCdR5BsIQjx3uIDQUruishwqUsc7QF
0zAFtXptu5pYSrmf4riXY5Aj5edGZfw8vA2WPG0H3hOCeKoiSvgHQ6x6eAsck6q8OzIv2Cw0Webp
ZEEpT+w0/aprmZRDqhekdf0PDTKhJGcZ4p/A7YvDMupGSbQOa+hiKggeSomXTA2rsbfwxght968y
eg31+aUzVchwtjCP4p0FM28MsXGZtbeJpHkptGpK4tP1QaKyQo5E95fJqTMnAVYcsGME9ed4/iQj
G38XZ/SMIY22bSIQ/o+wbFQLhsMNU37LWZP5SyIjTXdR/T+PH6R1AqLFqsf6V6Ew//70KgldklEt
yN6p/8TaVEpblQWxAVXFL9WmBfM7c2o9w2K31d00P95wSed0/zQ3Qei1v8VyXbb33jGfGtseHBUe
cNIkcuXgeVme+V0fRDuTf9x/69JfPK1yOj1IYbvZKtODjeaMUaKe7eg1vZf65Of2pDK2cHYd39zW
xThNcyvIYTpGmNJ9qlR9mqRHzjJGNs65SoXoN3EdlSd0jfggQCWxfLOTTTnBpXQHcXPJDyD6kkqc
1yavpZBk2HCXkWUcmJ05lbsloaf0vXNcQKmP0Bi3the2rZyNVAll8TpQycGOJNkArIi34LljuFRC
bii++vc1yn1sqRneaBFJ0L/bY9S8hVIYbcG3F2uuowhOtZmF/fB5KXZlF5XlAeNKyXZhaQPHKaVW
QiT0pjyBEg8lPW2yd/kF3Yg4fTBqQUBnbE188BnCPKQ+WHNNKA7/DC5Y8VNqlf1bD+F151JFtEgI
rFfWGQtNJSLKY4/+3E+xjXNkf4uSLH6Oj0BqnZPBk0jd4PmI0LxUP/xwTXa/16EpTX8U6Wlv/2hR
Fg0e8ljZMHCK0XZOxCDbjVHBe1noTPXZwhLRCy+X/PO2t5nNCDMcxuz8WV4bGBbsqoJ+gCRoxXQG
4uG/uxPi2ybkLZ2kBaVdRbKub4YhrYiYVKbORTTsYxiP2dJzCOl75D/BVOeHtGt8PIGzL0f+KEPn
Zf400jAES3hna1XD6tSeVcZUw2+iicz3UoAs1ESJATa1NAa3TWJJdoU5BPaJVZKSsCDsvgad/vnQ
Md+9sLJR6XKSQFLpeGW/mnz9byBtFMRPA8XgLQUghtqlO1n5EhaK5foqbvyW2p/OQDImfInUivre
VWoB49nJcxkNOydfqfwyELECNN2jxD33ADqwMmauppyGwkcPFIbfU1Nztd1vONhAMQLp8kEPNcvU
igAC3Toz4d2RU9XixXRSCH83XLYNwxWRhLMRmrSKgRaq8QX0ltcYeOSwqP9PHJ5zOriEhRmveMVy
q0Wc2TwDswgCXi4nOt6TxWo88M3zv/skwu/ZZlF8391sHs32CbjsfSFip5TAAXhGFuutgOIc6cq7
yiBvKLHDH0Hu76pVrEaPpa9a29ePuU5rsIdiGHVYZPTJ6TpLcBm3iHBNE31eMdmDIszRfywBr97P
/lIvLVrX2+4jONoWdU+m4/CS7nZe6o6W1RvdEqfXipnhAWWM3HsTCTaFQvArNRC3g0lXjVrURd9O
gJSdCrsHW5hmRVNB6XfRUf8vjShsv62sxOUc+/rENNq0eslsW8swFB/UYClQFd1yioI+6ca1mqRn
oy9VT+xUHiE4HeQbWiMJZ4lhsg6W8pl77vKmKBbIc0ArC6ieQkl1lKMYyJYnmbPa/TgrGoZCsoYD
LLyRE2mjvhXdiazQ6mzkTt0W9ZCvaqOirIOTYkuVa9yhlAB1QX5UN9piV7QDR1iiwfc2ISUr2+KA
rzpYVAx/HM/dYm+Tx6MTfJlpEoTMoyVKooXg0nnWn0ugyeXPDkpyQ6hZ29bIilFrdFRBFWj3p+la
HYFjizfx2htrP3v6PM988tXGMMRWaur2kApKwUvj+5LQkakLbsC+bc/E8/ScYi7Uq4AkbZNL47Ft
4s4rqQnZqYqmHGTlslEstMjqZy9qMIe3zF1YlGSnqip254R47OcOiXUpZij5o4dODk425WdOIFIQ
w83It8qGGZaLEZAZrWYeim2pViV3T1JB71G00BqOzAJz9QMAWuwL2IZsoEv6sEsWmyaXOxZy70iB
O4SpEYckXPAJ9SfYCielrnJF2q2079JCS3vq5GO7sHj4XdsSDgLTxsO4UrRvmah6Na/xBdoT3OgT
FRmNLedRv3s6VsTpjY50kxHNrFazJCL+BCfkt6ndIMZmiExo7cgaKb9U5fULOCTnbTxkNM91yJFU
FesxjhBUMY9nYP7Lh4j+m2qwUzDdtCpkukUN/yLGJp+No3NUVeJvGydkol/CtQhgp9ozIZkP7IqM
50O/RQ2lzW6fyKgp9HD2bzNVGYJMLskFANE3iKTznne5qCvlEdYsL5+eJ/M37r0B+dftf985oAx9
YouXyLa5FEPvlPTNAYUVAvPweWJlAuWkPaS1KCBlUS46uJ3z6f9hBdbdbXFQst5pZznp7Ptxz9Ww
Wj8dbUvch6avS3+DGF/Y86Zx1D3oHsa/Txw+RWsMk5VTr45SR8sLlcY4k0bHSxqHK1s0qsbNEyuP
96pMvvEz0+jBOCGCX4yGEseMkoig57JMdTsZApJJTiBh4/yhVnr1Yed8gDs1TNLRrKyXrg8gUwKq
kzsishBI/HylF9o+jXawUPxR3d4nyIHUYqoimc5nGrCD8g6J0+BwyPMhqgtRdrwo66DI9lZFwPxZ
RL/Z6Tfm8MF6FILijbcgz5ofdA6WPLapl27yScioJb7vXOgAkipO4gHeQ0DiXktex+ubsfcipUqO
klJIqeC2F/oIUn9YlnZSbq5sYmTR3BZU0q5CNf40A3V80tv6KScQe4c6KKWYNz3Kn6Y8GWC4DwGW
rvr8h5T71CxtZEHo9nZ/XT9FavFZnh4HvjTVxULEQqUbLNNCKMFBfxE0/fLmlvwucQJzHbYHy7Xb
weXTR/JH1ZBoBlIXsEDFpDCLt+rQMHWoYB78jk6ShWm6+Pcck4d7NUE1orcx1t3/1yte3RN4A68F
/UwaQDb+HIQ1V+oMdoP+LvTDUcqDQcC4EhpYAxLoRTNF6yApBKCNEkTGpGYrBkOm9nX/VjedGy3x
mQtEofiP1XnKFKsEcOJ0BbR/Rms9eGsTV2kLtX/E+cag8D7AV5yQr8TkcXXQDQVGwImd3o1MbCgh
+3VWVwUHFI90CgOxJdyAoni5MRuBTxM4fAEvcSn+XVOnl7YkyfEkX1ph+JzznIs8Shdwkq+XoyGB
BNfiXeKasIqNBunz+5nvoMYX7alvh/fJIvretgl77kTsw7Gx3qZ+naN6kaOeRIviM9xZcpkMkNjk
Oe0md5ZvIDmo65SyecjY3a5zn3rMPjtBNLpVVqrrezLQ4s7mB5V9D/nXtJrH+Z6w7ocsLx24dbZk
gS3ROu2PhsmKahi2S03Pkmm0PzIEMjBJK8ptlZ5bR2gg5PTMgCie0QbqundODmD+JvsY7AjOHi0s
+a8+U9uNfDvZt2IzN6FIdzPOrDbV4ac0G2FVylMdD5tMqV2Ka5XKvqshD7qa02yABthKZ63yWc7n
z5Dsg8RifVBC63mk4ixU4bBZFR7p1NG6cC2FNvejTq9sI2LwW0AA+VSjWNeDRKeK00f8dskTAf00
MOYxUFrfkU0gv5LXM7ashIeg/miAyVBoDsX8Rnb+6+QIwkf/T2CsyIwUclfhotNIcPMBycT5UGH6
JbsJcKNcCEwKd6ekBtxy746pceClkYXB2wyHVCxADQ98HctVViTdI4mn0BEjvBAj8kSEbtfCgZBM
NSFwLOs8K09NKo1A170e3iJYwkcXMCfzeMxOrzwi+nB8AnaHbQKxr4vfeGRu0lPg37F0tFn8vim0
ysvRnFeQVWO0JEWIBKzSZhXE+fMmAI0sup+P8ge+zu7KMZfsz8Q1Lz7FDnbTAlx2CtrbYG1D3T4A
UClDGxMjo1AtvpeV/T4F5Sald6FlVkdUJPkBK4Tzk5Fq4f52JRVBjyPJw4+S3FFS3rZY88N5uvEj
db2UFocOFIxNdRnDPJu4bhtJ0GiL499OQWT/8dY2UtRkRCgXWzv0jJ1vNAoDIMjji2xnyslZ5I4I
XRpMn2AHE5i2YIAtOBIpL8wJSDh9QMS9HyKdaW3kZSUI4peJEviXeuU78kZvTWlMRK6eBA/pQIfL
0yyBISZX2JwZgMgyT4cVcvoAPu6yXqiWeDskV+PJiL9OQBAtHxkz95OlIQ6Qr9hagY92AmqU0Ruf
9AYQ1ZUynPFpnlMWk30xooDqetf14f2cC0DW9xw8NlqW2ZC4GrcJ0Y/eRLHWSoxDJGCwS0cO5ebO
ATXZ2f/ZnoW+N1s4hLasmSM5W00UyVJXINTuqtVpfjUO/c24oC5z0VGYfvhgNobnQenyxMnkMmaa
AriSb9GoaiTwpUfbxiZPdtsxlwuCoM77pO2qHWLduiVNreWSzw2I91vKv9KzovNp7DR0tAjhwriY
DDdeTaaPfLbTYjProXIypajukngP1IrJu2yDh35fXFtroFP4jNSm9h5DarLS7a3eGbL4SW1kbFc+
VB5ya4Qg1xB8wj0Pzc2LV/RUjkCO49EX/6ta+8tRca4nZnwBoUwCS+it7fU43iBpyoCliDpUxI/s
P1HB+5M1OaAYrVvEp2+My6622tjQo+joEDsWJ/gVhU7OLLVeeAApSQWFhTegI/mcdZLHA/f8bdig
d5Qsh+BDjH43VY2NjRZmtRQZlugt9chAqqw3hcVs/PNRI1pvbqBJC58Asx/5ONRwdvjKfxZHANyT
2A0VqUewXam5dbNgtRSYquKnM17Rjro5+B2BFgQ/paz44lET1n1FdqVq7yOxYiIKzmf7J6Gkc/vT
9e+OjXzrUMOVS4T1rfZ8dd5XU/Gd1F9nhwQoHbgokqEOBjfi0VQMfmsXZuIyb35USk9y0pFUXEiC
RxdYd/C4k5FFo9wWVY1vWBj7Uvvg9ZWglasjPWVOBzL2EFPjR59fIE/uwwRoAV0h9XXTvvfhnf5+
Gvl9q7T2VVJzZXOo+IOQPTUQcyuiY7xTu/TYRSoTCYGNLVAGYVSMa9FdxQfX1KcyikaHAbZ6woWD
je13ODaE7tMaxjfl18c818e0liHx5iZDY7cva1IqiXHZOvXjVKryJlXJPZ52dyJfUYe1nyH1b9Ox
p06b5/VXJCbzEZB5E/IoO5A/ynC8nIoUegPRt6KAVJSsW8b2UOlwvSTUCX0d7sxP0W9+oG0hqc9V
ai7ecO9poc6S+FAFKcrwo4+OyTC29PotPk6Zi8RCJO7CUtGTf9tZ7VIAJ3yUIt7Bz0+Sr1gisAZE
nm5bVTqzylh3Im3KcsGv+BASZLrfz9z7zwu5WxC0FS8QmtlAjwRZ5nS6LNXDyLrq4LTf2vaeDkvZ
7+0hhDs4HFvV9WxuwzQRm4QNQedEs9HwboAQ4tPT4IFNOdr7A0Tls6Vzy7BW96S0JYqForYKQwuq
XGK1itNx+SbJhmY3ibJgdRPjo7FafSLcHxlImJ+xYKz4tqubanlAkg8YsVybo0cDdySqyvPjEyqS
aPJHEFyFBvGiM5tWyhkCKPxTKv4xl8fUnzxHjFydowWTy7CzkMk9GZWkETkO33Fwk0F5C+1KbUqX
04QbRCZhsNGWu4Sk2vXcDm1Pf2QWIi1pOpy6SVNqZ442f+zshlmZGw1fOwVL13vi4w7y79x0QDbl
J4xcAO8VYID3npyOfRjLET+MDj/2cMf/9AhPHgRgn8tKKoPOUfIzixKP+oQQ8CxGSubib21VXDy6
VnmKXT37CVnKufzCQ9b82ZdY65Lqc0tp+IceHP4GReteoFpMAT5Euer1qqW/FL7JTVUulmobWWJl
ZIHSXPjkDiN0jhPJK1KL9EqDmRZZXzIAz1NDgx9Q2zDaHLxgVwvVSChrD5h3r00MFdxLVBb0JZAz
klhPEz69ZdFgHf0+OtUM2eInrsU0pauSgsRqWhFlia5se0giLfg1LA6ysB3L1Z6+1qWcFU+MBg6p
cdHTybOXwVoNvovnWyDZWi0O1O38PJ4nHOJXmOREqF/Z83h9VtIvEn/0hXKiTByyzsElauiTv05V
9gS82bGqWs/fnfru0Eo1hURTaBR2FnOqIfEencmjd3VdUzRXriqSnzWboOoncHB2NY9wXJyYYVMQ
Ji1uhd12JoseCOvF/VIzrijOTFYKqXEDcdPG+6UrTvq4zzzQwWbcPagi691DqogFHkEio+KDJYLm
8a/3cmBk7XKxqOWG6orzhOd74qvszYAQrNDF5x76Y6Eq5Q+f9WSVQi/wuBDOqjxz6XQuxVmfjcW8
+IZ9eTI94dldhoG3ZFzoIHZxHAfVIvr/K2uKL+hlxq8daHoURUAvdVL0WCVlkhcOn6d4BjQtv/9V
Y90Mmzt+vUtWyTER6vXTohb0R8iaDLQ6tQfL4ttV5E5ijKGH6z/st5sYRwkW7dHcLahVCSI/1yvr
IA5U4kLAkinqVpn+GWu/tXkGU9sbaETpFLmnNcXemBNar72kOJmjJ1IKtSz9+I4DcuuRrEfD8fCr
8gntTEL9pGD+Wz7nM9jMcmrnoIs7HX6D0B46PPX7CVTkWKIZ2t5wHbtOkfG8p8PqD6AyHSs2kQjY
h2ISIOkCnLuymwr4cCxS1EIt7W1nec8aexTKCrPKM1JF2qbZ+lyaA/9vkafWg+Zvaag/HDAww7h4
gk2xdRLvYyBHyrlZYT7NAoFBhZY23AQU0hY7ACBcqe5xnRreCI7l70v/QL24PPV84WNN7lAMa0q3
J4ilMFhqpzMM0gEud3nFJtD5GMTKE4/Kv76FwEd58nZXiJKGKoDnrM4SwSeolrQZmtD2LqxRIiEK
Xy723PJi8bfZayMPlTh9bff6LvIuWmK2bITHrtnTi5LZxwEB9O1J3zsvFCh4xu83iz2nY8pduQ3b
Q00d9dSqx8pQ8D/DcbUmK30OErefhpmBGuzxySgbv+FXUBMG6y5VJAu+TpyxdpGT7Sf8q+NxQct4
cNE6ZxgQf+jnP+BIA9wF61po07Pa58Oc+28suzT1hrCUqgRHBd8tHPWXA5nWO6uVxxLo0KbHmebn
2m67j7ASfIeO4pR4280GC0iNlerq0K1F5iheBqlHR339/wo1t3Hx3pLucskZGlM08ZuRx7hWrlVC
t10FlbV3ofcV4lVfUYC1AqN+qT0Q0oMyhpoO+ZRde69Wkmmj7rnBJu7acoAbZboSHQ09m/W1UYOx
rTxbMr7/R96mPMH2rHKydD52OqwKoedq4D7fd7s/4J/aS7mOj1Sm5o15HrzmmnghFrzhGYVmoGcI
hgZBfNtq6G+ynaPFY/tP4LXvJD5aPQYk9kACLxv1oxDYQclUFZLlFUNadBkbV/8TthZQFu5fv/aw
/yBSUSuNM2K0nNmxqYMn2RebBJIa3nc0T/lOFhph8JG9QxVX6JtmJDX3ARnNkkxeSl/+5NCa0sfK
mdBBarbw02ovGHpKCwVGqVxv3tR4mczjtqPOSr5993rRIbX8rAju8Jede6JXDOzHvW6QVDUOAQQS
1H+ZUH3TgFKbH9hQDe3GhOK2JM0E6+Qg4cLi0mtf4y9BSNz9zXfwUW7dOTone9GmhS5UTRKdfvIS
PX4Ctq6hQGrQcVc3Yjkca60Irl7T+eHMXk2ys7ZvTqJh16Kcfz1CQyS5hQLJwxvEcHBxaRHcx3rJ
0uiVQZiPELtCbDkoFxEQC3Gbeij3+Ll16rziirfgUFlmj/aiwzp32kX+XVAb3CUEz98wlp8SNEeO
rCeW6RFhYwzBf30oxetmF37xzXCOwr30ZMwFLN6md0MR6SC4xMLum8ilgdVSjD4kRQDIpkJf0nvq
k77W3HhMXS4GhVaQFhE4Ymnpf1T8MWYx1ct0m/zamMArKSQ4GBC5B5AeWmyU+WJfT2ACmIFE+oxm
t9okba5d5aRwPs18LsxZcv2JtB687mH0Du24Q9N+HmAvm55qmgw+QRqBjlWqZZhe0VCnZI2hTg7Z
0Q185Iv2tzk0pN7cJTwoW1Q8dlhuvD0ADp5rd/T0vZt/nWeD3SdOMdDsQkUmEaoWtygXuDwHbAbO
5yZJ3/l+lHRMhYH5DcPQhf6sGCl291A+3epS3mh26nnZJ4K/Zbng6UeuFnuzQ8Bs+4WQGEUjBrZ9
oC3mYUYsaNlH79fwcL7gc5d+zjr0Q9v0N3/VOxrSrR86Byv6KQIukg/3A172Hf7APLfp6WFOIs3S
OLPS2balzQynMe4yLi0oTgsy7PEjT2DIr/LdnJ9CqWh2FnSi/qfGEzf2eEGWoG2A9wQTmzjv1jCv
SgK2iKewoh0TyDkCQAGODNud7snR8bMZN9VpR1CJX4H5c5KG59oXZ8GpldFIOhayNZNAq8jrS87Y
icmiWhLXIgpujf2V73qej18dMvHjHQ7TypXYYcnbHQaN8ZXorwDHexI/q2CxrAZ5uPhxZpwq9bPh
haCJjvNNoddOxTeX87WAC7bXc4vFtJXNcDru2AfWtkrdmhCGdRiHFUX1CzM/kxjCjwC2QCBRgx0P
EQZ+J/Wik+b+m3rp0I+tRSy7RsbgT8NpzPQy0Y7jLxdgoS+xJkI7ZZoJSCjVZgzZcsI3ALIGgoF8
FVYR/kwb6Bqg4ggs2uDYnnMXmz451H33woAb0gdlZ8YuhmUc0mhxeHsj7R11jD6Kg8KB0PrzZLvl
QlXbEkzuhUqCBnFQ0pxJ6oWrbVcHcEe1u2nHzd+d9loL96lbweConUveg0gfsSWciitdIbWgUaeW
2puuoSidymKshXTKSBT9lWtH/0j7PkuV93/rXmOPdXkWFGHPyMnGi0iJs8+dJNpY5A5Ku68ceA2F
w2q3QhMzSMpofbT6qpJdv/TpDdHjxHB4o2b8oho25KYRhNoFVEsAtBNPafQZaEk79UyHwysyMHmi
jV4IdBBEOtNL+tEWFBrRDb5x3/glCmCb7P8HGtLPi6jlv5h0o0F7SC+HvZEacq4nYRRb+nIw4hAy
L2k0DA4IQ4wnLtx3bNxdznahuZxTWu7m6fQ3ZZqCjDNi1RWgFBJTM2dGc87n8k5tU+YPsCwaZRlp
UrFItGmQpseqkFPNCYnN0AYDlHgueEwKqyYnT1rTwG0v3yv9SR7a1KfgtEsWQ6jvryel+2zWIEUD
UymrTe9BTn+ZtkurraUsqOy23eStK0A7Hr8rkEYGqRRwn5WeMA/25jEIpg1a0eXcxLSe8FGra8P6
82urI0A5b1wtysbpkKLD4qSxlv47BDg12l1PYUJwzWwNaiKcpB/SShp5BAFqT9HN8Nnfj0mk8r9f
+3EpHGgvYFOpsm2/En5C1+t5InizsY9wjSJIMPCqjA7QC4QipDJB+qyUh5h/rfOB2k/3tTa+ZHOy
q1P9g8CGzQugvLBTXQukYp9K8WaU+tp1TMGYZb4pDhCSTOf1LzTtj54fhhOFxbO2ResUg4DB6VHv
IY4q14QYfL92sY1EfN0NMs2//TzJNmjA8Qx9ASwLtpDYNY/VV58j7Lj6iLtEYkkSXFtt+FOBy88c
HqCHoCud+Szpz44vDnK/ebd59btvWAKN639sn9a+xol4zjms9eJrbBJwzNNo21YrTlScQ3p0Es2I
t7xFXUKq4YxtKDuddYL9FPIvoSuG9Qax1XX6bgStsbmOofc2FGQcxw0dr92euRCVDByN+Wy6fxnC
wYvNWKmAnq8JH7gNsUGGDGINSa82eC47LxrsPpZNOOGVyblFZpKU+ywmTGscsxZqqYea3vVv6LBw
C7ui+59sdOfXiGvDM7IeAL1oeQaWMkp7zQq+r4zW8uScIXqe7jReJfclrBRurXtQ4j+aTUDGL3+d
yYWFNyZtG2DX5i0SyI77U2p+dq8EDEyzCIp7DhjLUxlkQSotzHTuEJ8iQ0XYgQViMH9UdNvH01el
kR72sz8ZgCJ0SpBuEfDynErfwY0g4QwsEhN7VJWGVq35Q7QJg10cn+qfeJB8xY36ouNLd/iYv0pn
HKlIGp/ePW3mL8/R7cGjagL32vOelBX3aYQo13kItEiJhXaarlpTg4svl1OSOjEzxfvSiAyQaExt
aE4K9D+yA3JOmvBVlb+BH9+s+UOjphxKbfITN06hy9Qs7DdpgkoMBLYk0r7I6ibI14h5tiSrYkg1
SBFD/VnXcMElaxAIR8GEVf4hLXuUl0ZxzERqXhmakZ5EsP+JGOGOJNK5rdG2oshfu13CeIxXgOvf
BJCAmFooUMEOxX6hFoz9CNGOmYKC487ozQrhJw8BZytYVgeIMJzX2Q+n2CSgcBXM+u8hbFuy0LXg
vyODWX63RpJedOraj1dkCAkCl/nceOo2gxPsByg7ZYdgdzZs+2XjiX+AZmKtOdzB3+bD5aSC18hP
oCwZKHfv7Ff8MTQNNgGvS2Zx4brcABUSVPnAYpgH6kyuuueRx8VFhCAib5cBHwn/dIBhr0nnjEyN
URZ77FQbh/r24L3OcTJTvVZYMbLovgMeXt50ynPqxBiHF9HpbynJOUo1rLoTZDWydt4tvY6QazW9
JafmWtaNi72GAyrAWrxBrY9XTIkmxXR6T2GaK0W3mi7XwZw5WbVEfsZhp9yp6Q2L4vQ21N7z0ZN8
NQiMLITppnxOZjusCE69rOj9W2rDvvsGgMKQFj02lVUoRZBSD4GSJtY1NV4wvHX/whzzxYK/BNX1
feTS6v0EN6q2p1eQXlrAksdyx0M66Y2Go52K344pRitW4otGqNHIBXHRJNfnziNO2gxJd0jrVmQi
HRQ6upJ88QveAKpOsjw13vDqrV7RDaqvTPrnJIAff+13NqCDgoVGoYa65FqiZiMddtFRX83LQ3cS
ojzifdNKLN1p1WBCtnDYMBQ5khdxQ6SQ7vzXeScuM5fPW2b3O2CLq3QgeXnQTowqfbXONXNUSrXE
ag9g0x4L347uMluqDLfZtqokv5gpT2jcj/3Ug4P0L4XNmSOh1RSEg+K9BFvH46lvZAmSf39R9dty
01mfVx3GaN+YTIwMGkKEPiemYkN1EjCCCKWDbMYkZIKQy3flbupeoZy1n9czRe28wsyKt+nHuBYb
HzX8sXfyJx9r5Cf/bG/TYYy837eTOCfjXl3HY9M3ehgzvAtUzFTa1pnk+ubvRwwzw1r72NfJVkRZ
9zC5+jW0vSjmI/xFezxb/98jSgY6lz6bOzYC9cLKviHbTxnRzAM59q8SZ6Hc/qFfBOW72YG3XQxB
AyjjvWQ65NmONn2ClcG2qQAIi1kxUtEomYUTUJBYKK7U29/yO7vH3gNWojxAZ3t0lm385ADOqB9+
yNQnnxJdQ3EJgKAbEBHsVQ0eXk4QLxtmhzzYn53z5ILyvSHhRwCuLPlFji6Ar4NgXhEm0z6YQ3xW
i18E3E69K08RprfF2rKe0jobmzf4GmCi0Mme87Z4mh+6AeiVQyOLjvNUFyNdvXJvXX6USJKqpCN8
y4C/UiuUom/GcKbxlUs7Zq9wRyfZVWQfrrHd339CoumwwbbOJXZ/iZGsKv/EdYgipVvgjY0v0IzY
K9K1WpNGBeCdZVhvY9YFkhomgtRm0GrUI7fi0iCKiA7rXggLygtHoghx5sr2E5sAuJDFcyDWQYP7
+gSHfo9rHCp4X3ZyWkJPa9zKdzFQFZDEl6iC0ru2ERJ6jsGu5baGTn2yzKl6MVtpkn6te/iUBBTO
Vvlu+VP1HTQloH4zrecXfuclXcX5B93wVbtjO7LA1Fm34tikzoGCOaHsSvTph5m0UfHU4JEH5EYb
+i2wAvGgx7gUnjR2QdrT+cb53bb5/YSGxg50oiqlWrJvMNWKlH+MR+msTdt+nq+gB0JBtj0qXjqh
rgemmZvw6DHsO+GyOXvrRITD/stgRDiDnsazNU83PS42005T2+wRWGErvLKPdLx+jI3k8kE5PWkw
KdMDkHdieq2z+blswULqVATHZX54vFqVkAugOHjZFp/dHxbwv7Z3Bw4KWzp3r+1xEMlyN4hafibD
+CToSQVyAbkzG32wBWMa0UXR3+lIfiW6H6CEjfoLOMsCBIhnUhSMwQMFuBZLU/dH9qQOCfF17kHX
KJ550CLNVJJoiHqQq6XghTyLXg7WEaktWwLmbp+Mpk/m5/74xoxc9VFzyJ2nhjsEvEhXrzbqLaaH
bGVUi97gJHOPl1Z2t1C9aw0Wwh0LyxrDh2dpXq8Bk/L9a3dAayQ+tzGWKiFL9jztK/4rHYvpCBsp
UXb2fnPQZ5qdYUlLEoMn/wddqAsbO+TtkeZMo7kyVUBM1zbVpPOaTKkw37KI6ZVe8YgaSaua4u6E
3VZLo1lVsKfgkObaJwY+QdYtRe3qqbmzY4bIs+1DjbelZbRwa3OT6rUQgTqsVc+uNQ3K/pWziyi2
k8f+fQKBPNhBKdnxm5iO1d5oS6wcH6ug0o4ij1F0ROjct/c664lqU8RUHq3Pr7meENkdElQf9XDY
vui1tFv95wBdTH3hR0V99Fys/CFGiHD5/BKh53wPEhmE94j4fMOvtUJtpc4je1xA4GAbjju3iK27
aOVsG9wKZ0OWil2vy66gt6T7QbPNEDG0yTemznFoKw+aFiTj6U4hSFJMuVUWwulBBYKVj9jSnst6
tv2cm74JkGl9reWK8UKtU9dl4a9yzm748sxAo/kw1Ukxezs65Ly+mfV9t3CqVNhdo0dq67fb5jQD
/gpOatfg5eqg4B65qxoQBcICTX2d+x35AjAAcXITQ2BQRSW/ogdrcXacSIbIWu6+SCT/r9dVwTnC
oDema3aI8Wx8IQ293jE9Cp7MkdIGBNduz+xKlof1YS2sL8kKN/xRq32iv5iyCJroUPb2dJxd2pb+
ZfA1VSwC+y3ZQsM6iceyZY9SunEilymimBsq0z7lNDliDw8omhN6Y8A7M8xxSgl+bVQigMzR5gTw
bggt5jyFUyQQ+kYH4exbjLBkwmIUPAducGx6aQHCIkXKCxlyq/lJ6y5Jy7SUiIBELgB56u5Qr6wU
YOUC0dhHW+1Co3wWpHfObNA8hMh3td5QmrQcnZvJ0FEJqbKTjc3Xpsq0xUg0XSkJRqHyocpnqmm1
m3e+4L2iDUDGdSptFpkYjYUnI6460j4qAxsmVpregB8/kgBUHM91+92rRc6TR38EwqirKsDvavNL
+bwhH6BT7rrKQdF22zBgDWHaoUdydfNFd2b4x5xW/Bfe7ZHIAp7dYwy0tFzSNU6jTv/pnLb5e2u6
ZLLB266yg4WvhRwkiwPjDIZQAQuQZyKUhIYjxvVOg4r1QEn+lAa3Dx+xKz0m7q2QIj/uEKXUxZoY
9ildeHUbs3OxSB6Q24YV28FrQZCNHQH5/eI5esMbYEYrS4GmaPN7KRqJMk60bXKsPm+ZzwJXn/9p
f87R0xT6LlJ7AqE+4pgJrHLBTlQtYw5AdlxjwrYiKnEDr/AuWtuPYGNs3MVDLJI9Lt+G0525kUWF
B1jVx8JQA2gJzUy70VJsPqU/9l6V6dGvTM5JOAyaySx+wuHJvxryHUgKXa6SBX4j1Fdko8BdSm7P
mIiTiQmzRo1U//WUV62yn3i8Y9pM22TI/KvzKk0spgqUsQofU6gIp4r7FHGA5CLGzZGvUhlJ4Mg7
m85PeCevfBA7NdX2BEzu/BHYSrU3WWCZ9B8ByQXYM20nrRwZWit613KWEYp0W5T+Dq2wfe5ohssa
A066GlTMYsZBiPIY0XFFAAsMRSVIimbNgPJ3f4VUw95akO5vua6SeIS+R1I2n2VzQ9gu1+5w+Agx
dAjhU+oj7F1pm+Wbwr7g1kipOqY0fJOecW2wqvS8HGbwgZwPXq7rUiCeYZe5E7EDftrGkSapxlRB
9Lpu/qc1izDIinlMqNrGyRauSyfvTTimdSCYc0HbMk0WggnN3mek4t3I3svpVMD+HP7Tb+Ea23Fo
iPHwQXRZxfK0jA0LVX1Zdn/r0weuIB5f8qFbwRd4A+tbaYMN3ThImg3sKFePU+qY9IAn9dPFoIOH
KXjtg5NqalRTPd4cOwpMTb4jilE3DgWbM+lJhDFoDKDIhmR2a4HrTkX0ou5qnt+ZELfi4m3poMbf
G5IlcmjlY3nYXZ1K7RShnOaP0WEGMFgCP6o8xgoYL+XtJHGyRW9r/VHlyJu2K12NZCv2QImBOqNK
6YGgyWyKYIM7C/AHjspTykai8W3jcRq5HkU9eqZIJaZIsqb2mu1MNTWUMMXEwgF2apvYDf3nKUtf
UC2gcRQow8IwuyR6GpCfQ07gQsE/Tr8YAI5Qxd4UyxlDFCnW/jU0E7HtwqTJjF2LwyCoB/As9HK5
TrREFIe0b140P0TCQTiu3cuVNgssHXevg2H4cAAf+XLozAO9buKD3vWBnOiR+iBYMDduePQiTFJI
a2Tc4xaP1b96qcyvdI3xCeCF0Kcm0a1bV1ZMdg41ezFxrtH1UloZ81sasLwRes+Pmx4z9EanR4pu
XIKTU4izgc0NyYZYENj4SKdjZfqeOp2ucm5wi+FtDy2N8z8mkeL5C5pfSNt5EP7BBw9Kvp3Hs+da
/W7AxuAVkwO1o/L3JOUdsPgPNbmvdOuwv3okQV6Ny36pbaoHuRCbFOmmwfHuYzQlYW7KWIOah8dO
tnrtFEmvFGL6J+LVPHMcwO6gQ+8Tpron56fi8X7xJiY6PtEtg93b1/5aX9wZn7e3Z9N4Y6MX8w4g
a3tkewZfyztPO0/AtqLTfcrnKbPWBrW0x/AFf0SctHJoevRAMzOEL9QHTSflnJySsV/E0LhTwSSS
+3QBZ28C+inLu3KjqJJmF9DSnjpIs8TOw3wWCcuY0jdeU+5T0pjvcUsldYWf4FYhVVEvz3eFKHM0
HpDq0Qz8rU38uNu5rQJUu6pQqYTcJ1AnfIuENxf9dEsKSLFEpF8tsflXzAQsBHdFRBb7VTDqVHJG
hXrM1mtIHdTVh9TBKDVs3t/lYFzdku4123x5iAPS8ugxjKJZe8W4+XiG5M+Fuir0FrbaBYbgRiR0
onYbYykadIIKpqRVtP39yVPvwnCEn8crWacxwMfL2efbFLyyFdxofAFiuKqSB+YO5OTAwy7Acmqi
O93wWq7bEM1ppzbyCQeA9KIwXJW1rD1/jkFSmP3yLDhbasjR0Rfkd7913CFf4zi/bq83XY7HnoT5
R9SDMn3gzdqxlze/XETuNTLhPvK2OmqDd82XC34dzh6NuzO8IKePPekwU3rDvITaT00tpzGEva2g
jAS6VhYNIS5M1y4hKS/pKxNqqIForPWEUFCpgsEAaB3SnUx6KzuA28Y1ohfigbb5CPoDN0wP7w30
D+wIz8q54n3YlficO2Bgvh8Xfr+jV4v26m6st4IWW3O6JB79XSys4zCL4Meo9EyD5wuFZA0zHl25
tLisllyCN7U4b6aGa2mI4skQjIzsIU+9geFGEasJYB868fw8TRp8cAV4ob4Gakif6Sq6mLGNGTF9
I0Ers6CALEn7bOB3trvbLCChcSXgV0X5sHZ2SLTNgcOp8UAriWOW9Abp18lDNrsiedIGb0Vrl2bn
4XorWK+jB3H/nS6krMw+iClMJV+oE2LJXWOg7H/hI31o5G8W5yKJPD6CV2uXL+fr2R0v+ujnGuxy
XrG9Wks5WfXTAoWkR+PtPqPc+nAdKKl3Rc4Aa5VsytN4Uovh6bWiksSY0Wo6tC7sFiUTnLbA7G8D
XYFXIq9j/AyEpuv70IICiZ6kjuKwTZqqOIhEptR8cXrKNWIbYtQRjCYZk3KKm9QrcAMcNaZ3lkAw
k5wrSyK9ZN3yI7BVXtr37WE4+Kc9FjrxZlJX6GeNdapvv1tuBpQbOAXM1cQKX2AuQY2OndWbjA0Q
RaroYdpByi5Aqdn34mMRtslxzd7vnlXs1QKeTCaxAWHpuXao+qVuc8aWFsW923axov2lrwwpeMnI
m7K4KhhSKQh5r/VjILawovi0WnZ13jAR7Sl9vhLHUxlV5GCtkeNT92sfHl/6l/8oVNGX6NZ6CDIC
c/egMMQxA9PB5zjoccZtZ7eDfr8Onu1b1HBSbwxyRzz6QbpoZgQnVXh55/DNlY1Oe4f1x6ipuiS9
7yXoBXkd8TWuQ7vuejCaNiRQ28cy0D2arV/+T84Vg2Oh0EOirl3kCWh3TmBEUdx3mDXNMYgiaU/G
zN0UBtwM5dBUgPPpALn5X7v1G5YmwXptHRhDFur/kjL5FxvKrBB71/lwFl2F0S1Czc9rC4T62LGb
BWAbfwWy2ufkhAwZK42H8V8dMHd6JWJLfY8mH0hMGpndLr9GuX6gT8V/9kWwyFD0yZUhB74nuX2N
93s6Y9aOeK5AMg0MWQkcTKQTJq6zuPKiofGagHtAYnjI/IXOJJpTbOxIhMMGVMJXnz2sU0gzcz+V
y2RiTRD3W9u9t01UNCqw123P781xHeiw+sQKjVXd/WH9vQ/3MrCQojfEHbveI+xwtsEGNjfATPkt
f11uX0F1j+62XMrUYXlPSnH2QnuNlMdqnVI/X+eR4ekwaGCHSU9jWXS2AfMbtHqUyxAcrIg0aIMO
jHkdrcfl3m7knVvWXL+jQHcjV+OPrlIOsSq9gcDiojKfPxYtQJZlsIYO8KHTMlp0eikcXn96PIn/
FpEjZZDdzibDoF8z7np7q58JS3W5wkRBr1S1N3NiwKQviBORWRtvbouWSsgPfnNK3y0URxEK+ru+
1Pfq69bSr4mHOQn7u4aH+OC+e9TD4WiE6wjC16MBfk6BMvRBPHIpQ7mAUmcG0HSWB+GVCIkFBjXt
DUDroJe7BR9mALOzEF0k93Cqg3m1iUsghIxNzYxQiVYO1XURHvA1DVJWPKnBJbJ7v7sgJdCckF92
jm89sIBESsdV8Hd2audW5XzdcMNILzxhd60bqxYmAxdFb3LHZXZVrJpy7pRe1L4eUO1LHSHq5G/y
3VBFEwkU1OBVt6jN5Wv5nT0HJ747XwZZo3Se2fQTxO8MNdeF7neqAKStEd18451tfTm6KKsfstNL
7tkNQJUOnmsg2sMvrMiCjgdki2D3YL8FuQz7zG4g7nBWvmH9U/A4vgDInasIw6x4YjzulueL5fHw
wg7MsgnbWUfHxlcl8VuO06O8jZjNKXyb1ilaYvkQGCg4dytJ/ikXgd9q+ZZ/Ukyyit/kPsrBSiaT
GTuUmoZrcWVtLl9OoqiwOdAMaFVtTgEO96IeLASFJC4OP9jNJ9/51y9mnNNtIUwHDvoqxgFyiWR2
tXeZriqnoMwrrXqimyGF88Q9PPb+JokXrHouw39m/2s00oJuU6vW0R8MoHDZ1LZ+NrQen0Teb+8Q
bPN8l9F2+ipaKkSHnbOz1TqyhWRgewQ6b+QmF3OpkIZ7s7+ZWRUDbBmtd4DqDAMQY5ZGbF+ip+/6
T8oxftCRY++ioHW+lH3bPrDwQQ4265hDxbMnIk2f1GrEtNaVPrjZb2YrqJFX9zhJ5/r8yPw71ogJ
p/sgX6eSqF3PSs9PPkMapeDR2qE30KLfQXaqqvO2UxSFc6MuD694Sfdi13PHr5Ytv2EFN4OOH6+y
1xhHMdX/icGIxhS86HXT3+pdQWO+RuCDmUiu0GRq8C+7ET7N/nS4r1Gn4kBEGVpkIxXrmo+CSLGR
MSoo5XsfARiCKbSiE2KvS+JTcXhpeIjAC5u/zmz/nQ0PjHI43QyMFVK8Ska6en/F8uDuPhXIMZb7
t9Fr+wG8fdLBske1sBaZsf0sM9C9PI9GqZnig8e9wWEIJi/0S0L3fajuEH5B27EDNceNX1RnwY1J
QjwzrhfIcmGxFCl9nHs2yMlop1VI/h60u9Ph1+hfT21y4TCXMkxh6qGZVCysf/h+PyrehqLZF3Jw
tPBeKBAHcFJbj4NQvKLdWg0xgw6HrwD4ZEyE3qz0CUMMFH+9yh5ocpNKgDtDYueKXL5wkFyw86oA
+vq97ei5Ti/Opf1W7wTNKtd1j0wDGRVxnaaShXP30ta7lkKiF4VLBK33j43yhh0r76N5cKgy3geI
9O1VJwcj1Vehx+jufwq9iwfpjmAFBCLLNkiJ/a8Ow/fIF1/95teLH2Fbe953DsGcscrHbfcw2DQc
pvpWW0bZqovdwV+M/M/4eherwq5b91rZbEajLGh9+c1mqmT/T+Szt92smVos0TZCheHiYpU98u0q
n/dw0FysjK5Xdq68y2bR1+jh+TpO0p/ivqpIE3Gtkwv/eXrhyOpyNmlKS0Ac35wgJ5acxAQUpTHk
qffMFPbQ+H8pubhKX+5H+W2ldLRYbSKUwI0dBcem1u/8TeHfn8UNX260k/ysCp8IqL7ItrgKpXEm
dfT0tbKAsONa/NmBNG+jumkJMAqYDRaDV0D78zAmYDUCjGT5PJ11ksaNDJ02k34FT7Hk4LATWVA0
GUUvO7UmbG4vGCxkuyf5RABU4dPP4l9mjuqGOmx1HSNBDrNAS3b+ukfK6iPT3pT6RJSa+IRQN2V7
fxLIg5qrwOi01p1F02L0odfVJQWdpY6YvdHsSi44fGd0X6npW8EzetSMTWXQSKc0LOFilfFLWJ78
kCM0CZmGmbQv1pqOLtPr075IhZqpmkzbxdcPM1R2rg7QI2lhI/rCqqm1x+PQz2JuGOjRjrIZ5fju
CTsFMkaygC3vXQq5x0UY/P90RhLuRDABrA6jaJydjDO82cLmublIW3Tp/j2SmShyOuB+lE/NQTXo
8byuhxdP0ZgTY0nJDDprASEW4UTq99mt/CJEDTC2OiAPaxqmxe/9PkduVfyBBH3mbiAiVvluQH9+
LqZKIhGBk6F6M+fUfZAavLzeg6tjo5x2w44RgjWjYpTTLUWFwMTU4M2G7rEpXf6lRTheLuHzbX3R
LuydDfkL+1GSbJ7JA6YhtUMsD3vfCdcXUxib1lsxOAMgZ+hk0LyDV3EpmjXY2kitpNpbenmM+uC9
P6kWQeqGhybGn+5PLy7UfeyCxQbBQ6Hvp/f9aOc52AJNG3v94mKDVCVEl9vClA3awla01BJcKZl5
jnPNoELvaywzyVlrxjsROika5VukG98O5qGob3SkXwfx0mMD85WfATXGERV/DluLeLQ6Sbu1/BeF
KraBUBgV4jBzT6B/JrOLC8PO2e6f4df7PlSFQ2bx+WqVG/wYhhV9R0uAU5rNPxiG+zPIEoLTBlS2
oorJQPMI8EFQWG0ak1EGA9WnmT5O833esj/9DEo38aLCXle62Bjs2g6oJGEuxcU4iKiBkl5lgqRm
tCXSZdalxYPDGPf9j+yrn4aoBCpZbhOpn8TMBLEbTkG3Klo72iwkn4Pwjk0pKkPimPmoqfhqrmah
NA0QPmc2AUfGF6D1P/98cMDGq6m07ulbSOfCR0hUePJgWBSTF/FtjvLUsg2pHslz9qY/Pxe0LWrP
jsf1CqSic8Em2/XrNfSxQd/FOFRh2V4G5PHGMJ0SWtA7cz9bbbtpxF1zxFX5QVngS+atEvdUI+B7
blh9OSvdfvBx9O8ONz8IH9Z9f+QzTB/ru/zqjbXYmKi+RsaROYV96OJxo34+tgwUF4JOOOx4O5wC
NO3uo5+xETiIUFVQ4Emzn8ezFuS5n324LA==
`pragma protect end_protected
