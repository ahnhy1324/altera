// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
P+N5JhDzuRUVitXhyynWvZWaCUUJJd0vzABTwnfAvYtuEY6T/Zj1ff9j0x4jSqpq
/sPPw8RKkPb98OQEZhY+pfOaeONv1FVc8CM/P0qfxHf7ivt7qsL59D8dVJr3RACt
XNgnzj/RRzdLy9eWToqxiYwiRxp+op4E+nECH+zJoLQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 42768)
028FwGWDBDBjA6N9821gmVeqZLLAw3NuOdD27bcFUOwdgwUGQOvl1ZKKZev8/KYu
g62RN8Q2YddddBHLjqfTSQR4eMH3dWNrnvQzGG9L3O5PUzigBrl+RfDh8qP1DKAX
8VYhO6XW5wi6YfnvD2V66X2ZcW8/895UtC79FpyucHUxudchLemJYxpKWbGZohUH
MaW9OlTWRopp7sjqscnAF6BOoXoUltAWNOTOJu3fFgyopnQJZt5z1nep2sz8WX1S
QQHOlsc+IILIPLOGsqd153kfpelWNDW+RLMOMKLLlDb0cf2iFPL6dPSABKQAW25S
/ZlEfJdyjdwbvES2TetyI6CT0uR62i1dYEsHdGbEObTuPkl/ohlg0DCW+smOpuHz
6V+R+StMzYmD2L2dkuxRaHzFgiViWmPYEQWUI6VrZ8wtBrYyOE6+ElV+sI/+0PRK
h2mXASiC2OhWDVuKEbT+CBm3gPHDGb+xkX1i4/c47W/ZHqbsqIM8nMnO5y3cQEws
kwmtgKo5uuOryoQPmBs1bkQR2Vdx1yL/FQO3xJCHGB6ajztf7bUxF0Wm6zJJUFTG
nOQaFMnzJilaMiqtwS+p+g4mTlJOxccQgQ4fw1X5bzgBDHIfzw1D4Ogx2tOTEtZe
HJ6PQNELssbTkXezprSPYyoEr5/jIj8ZmTUHBUYQFUqs8B4dce8Hq5vqczdvLzy3
69IIwYuP08GOHzBuFxmliLIwLLjfJwa26eC5+pcm0AjZsCoSvJDHQ9QXxEPgPwHZ
FDrZYebpZ4ncJ12dp1J5qXSVOMyOD6RUExmHCxZWyoECTfgoK4kJUVsMXarVUslv
mYbBq4vGw4oc/4RvRGTRINCEHtACEsBiUfkxkk4bcBWF1abVxDE+JXR+2tC6lClo
GCK0fE2L84XGuGPPmpNpMEYK/dVo8FQF0JmDyUPOOcjPqr+mx3Ue4JJTc7vF01v6
oQOyxv/jFU524lIpLHNwrJ4pxBAoI6btD7dwzi1GmFtDu/rwzkC4iGj1gvBtAJxW
+LThIyiKUfm8zq6lrtXKUM2Q8eT/JCxY3KWcWv8oeCX3qNhXz6moaCFdHGSYZ0nc
13sFBfnT5eXwmRNP6lbfhfNL42v1fZks6vaRnHhyWfzw31gRqSONMW+HpycKXl3N
wR25QVIrfK78yZXI/yZ+rqgw/2KAJPckPTOg/pn5wp75mvuckqtpOoQkN2c1/hw/
Va/2tgt98VheF4ifFJkAXvWKvSDU3I093sVj3QbvTkJ1kTiYXH1u8WJ0xcQ/oSfN
hgt0DUyWoVVY37QpK/dqvzUayvPeQPkiPcqzk6805dwP2/7/4UTwwUT1U11BYxdO
Cnam9AHTuacPX4C/G/U6LTeW8JmaPV4YRf3qslVHKCaPJwWE5IGOsi/VleZ+o/Dz
WYvXkxLZ8ieKK3urJTgVf2peEHtrosDITcsC2eni4KN8dzPtef4d5iWkcVamrXgD
+u+Le6+aIJRlA7yjVVg7w6OFVr/YwZTwZgfG3qnNvPSYtTniPNUNR3k3bfkBWyX/
qfmTufV/SHp2bhfAjIxREJXfaZjGiYsvtnmKERAksGJNbV5BNmJta0Lo6oWfvyBa
WIXvXj5TbX3Kc/vp2S1uNnT+OTOgoFsLzQ3M4Mb92jB3sTij/XJKLE8vebjx9uMy
HGzaV6DRwXy39P0GancbATzklthFxtZahqOPg6qeGw56XpKzSC7i4nizTO5MEfv/
IYVisVP6QADKh8dx9wx2S+82CdEWQNMvZsMdHYd2XbYkZeufr2FmUm2qPBFLokvg
jXbYexDYa9HCi0Zp4uanGyB+jkByEYyJX79tMC07LqnVzAODLkYHO2mWuW3jYL6R
PJVcdqzK1+IfWhV5+DxW9Xh82/Kkj/X4/ZaObiFg71lKrilzYRYYqitorjRWkr0E
U96uXrhEgabJTE6XNddQH6jfIiGGlb9LLPxUt+4qi/lnIDobmuBxlm2jLh5JcP3v
hhe0cDfyop8ci98u7fjtzAkMor6z8A4kD7PZWnvAa95Hn1GPEbLxdFZg6VlrDjH2
HLp+dJ4JIt6XL6b9zPPVBqseYqXOBjCcG3182x2zgCwnPFRBTA5+EIcVRjx4lg90
ivxWyaM9SK/mWEA1D/AVHrLbbIy4klNHB62jNWJHxOfHC2J8RANh7y/aPjYqPaj5
u/XTtAPcF/lYyc80GRddZ6Bj+w8d8t1qCdEexrU1COM9n0/SHC0rbKKomIC+svX6
eiQD+g8J4TzSvBLGe4hCy+PdCvNAL8lO8SNkrV5RtLSAMswEgngQ8KuAmpwhDQvc
+8w6Cjdvj9jm5oW+8zwwZUKddztmuWjyaFnq2vwjDRzF70lwduktL/YWydJrYnTV
gZjmcqqyawHj6Z38GA+MWOccDcdunQMzXk+BP+gZJp8KTIUfTN99ESPDFCVR9vlm
U1sLI79k5BK/thEF+Q1zPtYd36Jzi87/bCOcS0XJBUmqyMFONcPkeDLHIQkF2ng6
ruVnJM39gBsOtGqJqDhxlraLGNJE31nN0pZ+1xERI89zcYZxQ5fjeHaS0mzs950L
gtKKVjtJ7bX1JFBFVckCFfUMDFAKwRWMVPH2wxa0kVIQ3tyMdG/NPf5gfawq7kOr
QTVES5ql5Hx7wqPswZ5z9BM3aDfEYxuoj3gom2AJPWi++8Ve6YsEk6vXXRSsppj8
yxZZUaE3D3LdbNY5KFnhInXrndToWVrFtzRbCP64IY5QpJZessexzdTXy5h3g1H/
304GivKK1IF1J/S96HYexHAQBzZVgT33kI6U89ffD6adiBQeeFlNHKtRpIjR4G8y
C2KAg4CWzOoLbg29wIRAN4BsevNyEuGF1wVtuBaiL++87CDWZkTwdaL+VNaLlZ4H
odZNt03df8YqUGUd6jS3aJmDWYDEl/fwcYOhkBqEZ9QJ5SCakOhZm5YIhucHkfi2
rwsz+mMCSjRMn3N+nwFBCVqMg4AD+z8d5r/DT65oKu/QZGUGkbz0CqvYGWA0m4W4
2QyrR2q+6zcQSI1+zPZn5xAdtW5LbHFYVka1UDSl/Lfqq1yVSdH4LbqpXaEarU9i
8bmaLQCnR6euxuc3aaaF7wWCzBXrqi+DuDTf/0+V4NYGEPor1szZkbMYpG80PvPK
6mPcEFzOcwGj1NOmZiHRGh6F7M+omKzQdUnBhQHmLiyrCgM6njDpIERWvsYU1HoE
8Liy1DVnLxSXKtit5bPVc3G7fJYjjYUOGbn6RBs5ldlqYPcol/EK6gTxTzRCOi8e
Du49VfvYYK1MK0w4EpRAHfQQtkqeUdFTtg0PrVNkJiChOphiSgiu14i5EOHWs98j
nkQIJq6wumuF2RgqiqbL4laWS6dbvka/FHAqipxLArNGv19aTtKuuujvVxOzSUDJ
chdQSS6AxRjGlQk6oMHCnaD7Ckl+dnTOFtbFijoS3NEXCXFKRDB5mTmp6bpZ6RCU
sURf6k0CF4YiyYtNnu6QcnWDmbdfcgqNFoY6ouLmDOIE+eCHlreYXp/dHtI/cxWK
jC38gqsuhmpSKISTAKfqmJWwAqVIa+xJW+n4mfkUS3syQtrskLBie1DeGNylKBKa
dsKJ5RA/tEKjVdynF6QiiGkJl6aXFNrXScOUW/CJwCK6e3aXBzLPnde/611bKz76
JAfWcaiPfSPQlfq6oxu8hN/QY9oOsSTDOQbPZKrvudkUPHJLnuv/gz14A5EigTw+
0mvHA+N5biRRtgzM9vB2hANYPUmB5JBzwbHXqIMy9jgLJnhJzv0P34i130XnrwGZ
eLYGKTBcYVM8qQ+oLq8frWbeFh7Y3u2PNeV7yaczfMTof2xVRnW+K5HpS86qxQFZ
PHMUEeJ5Ejz1df5P8t0XAJRAc0Mk9lIYqj9FNNKzGLKVck1XmRWxmJhRE6R9QTpC
thTdUDqlHu0HVdNIaH50VsNwmLNO3yztEr68Uon8hMVfcxuXbKlIVlI3j/E+r+AN
suugoLC22i6HrWqOSB7KEd/Xj07dR2LzuFPr4MSCmsKcqDvmuDUoOobhYUFkDyZj
Xl7IykpH5fCaNVCZfQxPUYJFW+eAQWxrTnb03wxZnYxZVk1/VZi2jBkRW+b6OC40
U5CGNzYFEbiZjkFW+sV9fEzMrbHlWJZp99dJS7NYTQ6oPaiQToFF5/s+SI7MaIvL
htyPfVbaT64E+i+Yd9zC6y3wzzBgB2UECoxmbhmSTin2O+d8enyA+vkJzy0Wi1g4
8AdlcUJKu3Yl5Q2M3RbKy5rEjeIpW9PyHalx12AFC9UOjEkR7LM5KCITH6SevJm2
yF3ZJreqfaN81x5tOzE3Q1hJLdoyejJF1uXQmt9mP64lNOpfpX+5CkYSZsRY0idM
3oDyxcn82EnRi7xr/TLcfr4p1R4xM2bjNv2ZcFrl393aFwRzfQLWivJ80p8HCqzE
nfYkpZTc/rvGTQzibJwxmcUqFTWQleGvuy/mC2maTg2XIFVPhi0OI50P7KK6PRxW
49vEwcdNPCvbDfl1HeX713stFDTTRP7JY+F6oGvqKFPix4jqnlUAOxR88gLjBPHv
a99wUaMXteiyu9jov2hvpxGWjc/vU/aIvK5DbhyIq78uWBzGojx1NfeastVvCmXs
8abvcuzD+4HOHlingMQ9ODCBcJ4gJkzYz1ZTneIhhYcXygqN8bEdYmjs6XUfZi9U
hOUrzjcyjTYnIt9peewXPBvOGG42bSfi4CBgwHPpEqzio0jFH3mxNjEXhOBsYgfE
cjMRETJxH++KNr3lgFMMIsKkU+Zs9Eylt9X9d7n4LSVmq8XHupj9tF18ukZEzxbm
5LA5WLJRTzy8W3AOwJfrtEfkay+5urPtAGA52sjJeJ3AZZXQLzQirs3j4g7037+w
jibNHCuqDZ+p9gkmItS06AFsWuiEnJguctvzkYDR1pAyQ6X0F+EdYoQhwuhAMalD
+PvKDCpp+OJSm3pFrSU7ugwyht+DGzCfaV4F8D03jJglzCkjLxRIZezlnDYyd2RO
5YaZqsIqa2eJAwNZ5yTJ7hgV2AmdC7anH9fh0fiBC8lZyocDOCmGX7PmFf1YKytq
dKAY+HglX1sMNM9VFkNv51TE1Q0fdSyFq9M5VqHFlgtzq626uRCaSGVdwYxjma33
qONBOvcdVW3F1MXCtpMswoqcPAYIbUQt5dawzZ3KdsfQAW9ObvifIrqE0hGl4SOX
HBxOiRuwUU3i6BrTc5Yj85INAeytSGxxAfsreI38hMTNn6Ojqt7wyhP1XxHJrTFO
NhTwX/z187QIVc4sZeZDOTG5nUV+vRIAGHKTNevPGZurJEQKt45Ca08tc8pRvKAx
CMti1HdNl4Um3PJWPafFBhTmBG6PLMOCpH0RPpBK6KdG4ZVLLjFnGDO5sAGaMMBH
LmfeMf0RJMewyT3p2kGcyz+V4WltXal7x9qzbS69xStIu7nYEc8T8LrTgx4J914c
0p9fn/HkrgYl2KI78tnFiyNEZn/uhzo0FRX3kkVGEajyq9iEBoSfB0A5PFkVXd3o
l+12SlHNM+wcc0Y7aGoJBA7d6TlIzbWurz5vow2nNMOO6njrTGj7ojAh7n7kAKvs
aVEv9bPO1i/y1PETZrWuT36o6pXCLtEojTvoQjxd5TuUtDblU4OdEkDyWJqgN++u
Wyb7IUfM76WHbe2WQt7RxFeW6wVp7w+tUaKqYXHQGTwu3HrzWRWIj2MECncK5C1e
OLQWPBuP+fNI5WSYGazZDO3VJY1FEXjp9/lprIoEiyS7mNGw9Bl1Y/q9WbHY8FxC
XBW/+SL2Un/1psBTSMHHOK/5b4IpS/VtpwQmUA3y6sSuaaFI1vd/LOJMbyDTFaUm
/dJDGPVSu5tFmR89OS+iUi6zAoyiC4s4tgE7WgycVJFFpzJhFGk8RsxhOQwQxUdc
Kmr1ZbLU/jlbOAuB1boCZqxTM4JPOPF63whPykgDYZloI1FD+8IwoNSPG8gzU+AX
xgTRLdvFvJP0FXLcBeaGjPjxYHgxjU9WcWtEZFXXITjE0O5pdk65BYDt0YENvjFW
Ly2JxO8qD6uLOX8U9t8j8my9cTi3UeWllxZ+qYvg+QabHHSBv8EVW0VVZ/tA9sqC
yowt28iXhaWfczW3euAzJ+5GijoPn+UH5CAM0Hkc2vs48+/gZWtr6bL+oOElb/ze
91SliMWUqkqJ8EWliKYGFJSy4iiGbtPTD42NCxon17u2KywIe1K6C/Ze0noQv1vQ
5ooDO9pF+8i3fYewtwDkpXAlGk94Ii2pHe8+z42XW1r3fnPWnAgKqh9wHaiKiqc1
g6j/fQyaXrSFlBxpl96cgNR3KHiAvWApGhguIRdBoGL2oK2ZgwX8xCte5vR0l2ja
qJNQHVS/xfsvaNAuWRQosB2PLFi4h+iyv3rP7iMFyL/RLp0IiuPZRVUEMqSsxXMT
6XYcGy9W3jaCIhgp8ZX+RErxKFdg1hS2B+e/yPlU7HYTsLYuOUpQeL8pAMxAg64h
6tLRqWesVDIcgxR4FYJkx/bhvN3Gh/JT6SfEaR043u5O51TP3y4Lme+5JZpaU0AY
UIptAh9XqsCh+xAEQ0AP9RaFYPzvVKHgZPa9MgqyVQAVBuBXONWkmufT+ykDS7es
gazqeezUTl15+2VbaoeIvQPl7ndyJy7+gewbDDOOiZ7yhYo+0So01ITblmzxgGqm
KW++HFJ+z3H12MPewRSYDwOC5qMAOH5QoCmAxyoK7yCxlLNkFh7dX712NAi/qTBc
Viv46d7+l92Pqj0K0qmoI6zlflYX30yBqOUHLhEjoEbevG6+rYiJcHdKHcDhgTEd
88yqG7I85xjywnyu+6XutITvVhgdmJhYhd2JN50sw9pe7UCaOIR0lhFqufNfze4a
7sIfgWbJC5WwP5LkcJLZ0gz+Nr0+3xf+DJRhQOiFoeAf9yTyekUfZtNlRRNcdicg
DZ2RMTWhjG76T+gKCQdihrx48byYmFeWFJJn40XpVwJ6LJV9h43xwlXS04/hBpiW
Ao6RRWgt/xD8VzYyZ4A0Sr6Mxvdbyp4LNe2QircVPbJOrPcaDZUyfvas03syLvZg
z99rJZVbCSBFvcD3o8ayB6Hso6vtz9T3Xh/HVmMWWXjL3bVKm+hlN9ePDewDxIgI
werAQRIgBsF87hIqHd16/gvD0vaYgD9gDIyeuR1tPdSGAKXmdfeaZfbUjKHisMz6
kxcMqmcPvztY1kK+PM6vemS+aqRkl7IddBA9e6UVY5l7BG7pP/Xiq6YFW+O6etpa
a1VAaxZuGU3XcFvrRQKYsZfl1UawTDp8wMB3F2qyH3agJcHFEwekBQh+6ml6Ubcl
y2A0C19Vsb2Y3UvDHOm7zzcdH4JFs/3ArsOmJGq8WMfohNEsaz5mONeHc9OdeFve
CdOPelmnGvTfHzjleFXEdBkn4K7wTRRzRJ5dAg/foFhicG/OJ/1pURUK5fNhLEFy
nwhOiQc7pRnDL7J3lf4ZyLDaCsGLTKic7ZOSSVDzJV5JAePwFQu6d5T6iBYSY2aR
V7krKjIqywUoJUSXBLK08MC7I5GH09LmTQtHwbdL35ERxZNtRGAeXiMoDCL+7ydl
KVhflhUlroAGtEaW9WAzH6khVZ6I5CAvtrdg8MeWDFyh2HU6LInkfPjb92ezYvVd
ONqU1I1cHsOO8twbd6nTDqpyw0koeyVmjpmiMXwO7220sBBE3ETkeSBZJx3PO7sz
VmsJwGA17jpCL/PPOxGu8987TzkelbGNxjyRh3GoLVIraMes7nZM6rZTnr6/WSJy
AA1IbTwXHIAVawzp42FgrhDKm46tr7RV6yBi9FtMyloUJA1fI2m1usO8lWk9DqZg
aM68ctIgqhzEgtQRFCqo9C2KEyrcpHudycPtDBBlP42h4aWgywwgBwEw3H9iFKif
rIvxYKh9A3GM9HeSdc/scjWJqM9x5ETwjKEkyHewAwcF9m4WXpiVxSG1qpbsGh+d
gXwBHYaWkTdvzW3G14ZvDAWvSuQOjZBe+SpY83RxGCchJIScMhA4EurnsAvmm2BJ
nL2CKNHgGbuD/UV4TfG44vbv1lqCQy/ieYJdudEgGUIyTL+x625s+Kzqfox1ky4b
mM8zbqWjcdU2JL0f8JWIghC16JfbK8jruBL8GDpOrNXANe4dmELs6mZE6e6LYtJY
rLb99r7MsmtQ9dxNBuS5YQR37MZgK2HA0in6w9CwTfz3WA05hSn74AbT4t4xV2YD
fG0NtMqVvFM/THWX4n/5MLUzGd0nUt+axERZULMUgttOMTB3IbuJQVZbb9agG15z
qG/sfm89veYC8SBVd+k5Uah6XbZByhYuxCRDOSftTjvUIVsXT3Qy7ZHGPnGpLLn2
aSl3EdFtX6whHGlX0kgJRdCBghXgH3mZLf+OvSFQfn68b2odRqSRCAdoaSHXbkJ5
dbDQG5wEoOsuJ3UEJVPWIK6BLW7bq2S2eRJ29TKG4Tou6CyW1Nud4OupMvWJWYSP
oMJ0B+Nlp3Aq9dgbKUo/I0IgINdlD6dRFpZzqIGsRC2DVLBkgc7DOsBIugc7VQXh
ykydMZFG8s30ZRnjO53R7q6mK8Ek1Emk6z4//C3fhvk6aK/9nK7IHh3icXwVLXYI
QgNLs6XUQY/G620+xZjbP1NzKSXZLQDKjtowTdfa3TzHqKI7vFz/GDmpm9RXz+dZ
1dERbPGxs/Gjsdzyz9tnO8zyervgUZ0c/8lRpO5ZdUQTR4ARNcVD34mrbpy20BPK
/jpMN/SbeoE0KMD5p0dZ0FKF2nmh6Y2UYARwvX6nin1sAJbARtXop8vZzu9w2+FH
n2q8cNvYXTyyf5n1kve/EFsiPlQwrwpa/D3xCReEfWDHzd+ZlHj8H38cz9UxVa0e
vitGkhhSwsaXL3ytGtt6fQxUe0Fucab8T5ydrc8XRgjAyd6moRpgPVvh89FgtM07
R1epF3CVtTAkk4NKT2wfc77q5Eyh8xVVJ29O5KmU6ALeX0Zuv+PLQ18TRg6aKX5S
AyXAuDcrO+nMdNeqMcAqbBWiHxWo8ebg5c7MgEYPqX1tW0twRMf2ZlRnQwTBD0d3
/aIrNDaA/rEcXhGTiIPBYxxB23wAfGK3/cWd7HZl1fs2leB2WNFOve8V3689/U2j
iOeiuhpmOgkM4YkUDAEeLYWr4283ewgB/U/tvs/O/TDwlu1w3KrGDvKCjEtGTRXQ
K9MOkzsc27tWEmIDAICFLc1tDozQs/xwUG1BoQOJMqG5zjK/p0A5mpmWpXpZos2/
vvHM/2AO77CzOchuGOwCodHH52DOkCpeNchTIhrFmllsDuFYFBP0eTOe1fJV8BMs
O8KVsZftO0MGOHjNRx9/zKT7G4wt3TNs3tb1ibD5yQWUneRYhbU8f6qrmKFQfwV/
o3Yd5Q3CLO952jZm5z+EUc1MrsPpGbpGIPuNGdL13nNij1TijxSoNbqSpgyKZxcZ
6256gDd+UDl7/l8ijsCypCBRmTejG97CRB8Nka88BOv2LxDuCluuRRhIkd2FtEuT
ZRkCflsG2L8ImDKay+giWs04HR2iy8ExJ3bmHC2pIfc1pd4w5U1Xayqcyb45uQ/E
JHawVqTb+MPKSMAd4dSyR15XL9I9qbeKVR0sZZVKJ3ipJN6QnMRULLWABMuSA8wV
JeOnUBBnwuZErTz6XIjniRZWv7c3vZWZ4PrNlexssnDJnMHeWi1oRTOcN0XAbuyl
BZduyjzwcvvWk3X7TG7SpA4FUUMwEmtJGBLaLQJM/Gmj02bMSoQ6+OEw4XFWX7Qz
fhsDBt3Oogit1FT06P2+i9nppbI2TK7NaZnEBFAkZ4lR6gwO9kgW3PrKZhfYyIMk
UME9DX3vX3/TsaqMFGLAgvGmXAiPgzabFs81qgcvWJl8dR4pdQXrFibI3IOxvn3o
/aACQQMQRJskN7+ABaZ+tWqZr2yMianGQdo7Wvobu7k2pZTfxffp6bsv9StXFjSP
A1416aXrbAZrqgse0SkEcfVM/H6Tc8arncUaKcShUJZ8BgZU0PWfxt7lnOjo00+w
fyKddHJRI/PN/QuAVgSxUXUeSjvfCg4AlDrZCxJNWfIDuZwAD9Ath2seD0PhLw6P
di3D0mXiPpMihED8zkVNd2MLdHoZHRTRmY1n2iW4HqXIOqenMx+6o3pYRwDHulaS
mq4j9VW44KNVudtd2FPM0SG+1LvKqSxldm5NbLTJPMLPeIurFR2JECNSsfXgeiZu
Rz/3Q+MnI6s3r3xBSiN/235UO0911tl8w7CFGwTgs9g/T4X2tq3/hgXUG5/XWXPf
KcxgqmxLLOolcPmZu504vns7uZUdN2KBQLMJsKrYIE+ZDWKOXpKIgp4Bz8CJaheP
8xq6I/eKF99e5MjwUp4ZP0yCkWnmSgazj4+bdUVB92CldzdOTuNanVhIrDUMMpJH
pCj7+yWpOSVTd/jBaHxz6KLiug+b8RVSaw/UqtkFr/bkbRKcDw76weGf8Gdl+VKB
PMPoBWzRIm030t3GNzkkdphIX9WSLgirAxPgV5tGPmjG2Kjv5e7UiSFoWBxLaJxv
uKKsUCBLJKlReh+wKlv8LfdZKsyELtxv5JThmBIfUAEUh1Vfh4gA/jklIuS00ydk
7zJUGD7C0cP7Fo4Pi6angB2kk8pcxH2zIjM+N8l7AR8nW04JrzlJnqdFBflDFjiU
JN9UrCGuh7jEKjTd2PyYrWwf4c3MKtyscc3bmKQqGoKu0jYBb22vQt/8rJMYWryX
Devgn1tMC5yGW0GH2d/Dv5gvJRrX4LUJIA5NMzeTmU5wwKaFM7Brb9ovgaeO5WiT
KkE06nYTaxULhHJm1BHaWclbXHGNNYMDxofNWmfjDyh8wC3pN7+TZK1Ulmb05JO5
uhVt2Xbp7/toVnegcjp8IRX5Hw3pSvscgKo3x5Vql8ZWSi/LWA0GH9JknqnpID/n
UtOYGaJeBKLBloEYt6Wa+QvNas1N81UFJJnZC2EMSC5LhptCzNWe0QRIPpClfuRo
mHPS3bfiLdd8M0cgaK3GQ92sB8HZVr9GpXNa6UpOQd3DbpV2tY55xtKQjkShro3c
2th8e4aIpuvTWOoQ662dYnfmtHojXqAFE9fNbv6dGOMxVRqt3OvPnvHmmRH/3jUh
vJdij0JnECIAFUrpxGC7Y5SYYQn+PJSj+uBXz8nsTC1KqzrvOJ8ZP3vijD5WqYOX
N+rn1AiqFmkZieA9au7CT3A8gBEiSlkggE1j7kK8o+4e9VzLq8g7V9uq4b1zScp5
JsjSVGa+ZnTTZFZXjXxnZzTtyhVUQ8YBWqYHl0jN4RvKymps+6H/+efVBsECNyfd
IaUSb0MJFwwiSWRXa5RxYOBVM1mHUsuIYBzTjXPlVn/FuNE5Vr3W7si8ggKbPzxY
vUR0QjXU0ZjAF8n2eEqAhnwU6lPuv/a/DxVegmRvHGys3A+/GXNAI8d2KcCfaNe7
lhwpXqlkCBfmql4nIxu/xWE8LuZ3AkUC4lOR0h6fH2NPfI+bZHgSFB562/2EcsZy
BHQANakrjWl1MQbQQCuWNG1wkKBj5hobGgiYmSGNReYkjwNIZNCI0XASHMM+OIWi
MVoaeAOh+q0e/YPZ+9PsOM4Kk+TcZPsqtbMvzFr2fd3CWlG2u6V/n1mR1VjQ/ixA
r5EC5Irjn0WOfTISRxMUcWwen7Nu99itGohmi1KiY2/7TC2ZbcfUSMRUg3YM5Usp
e9taPX7D/LRmWXQJa52oa0bkEb1i15YPtgsMj2nJvh6FtuFsEAqA2JDOCvTqSwZP
vpG0Vq+EIUYmvcTpWbMFU1AvnwdOqZ06T59w5eyixhIuNdQX4Rb3oiy5kfHy1bU1
ZEm3//akllNFh3Bs7AL0OTO7TLpiodMTaIJ6ErDJKoId79AzUFC5mN6oLYiV0wc4
ObJxFewiKTyL4PqpXRW0raKtA+lHLYkzTfSbIsEwuz80SGJ9UdBh0TIYKIOVOa3t
Dm09vjJKAcRqBUzsWjgTsRyiHTobT1xVLjSiKBkM7E4WvrVdS7/h9bkqTvldmxmG
slbmOznhbiEIgmveBtacpX8g9rPygTxHKdHP2kAlOxNnLJ3xyJMRMaFMA4mzhwQ8
s7imyjKwdWdkAnXqDJ9Xq3VhXiCLPg6ozFVvpPg1JkV3hy11J/iOAkQwDUpUEndu
CSf3oryv0Ji/do+ZJOjyIZdeqS/UDuOs7iaEDdRJT947N9QxsdQyqxEuRM+sWF/M
cy1k9tDca/6K04yab3+ZGx1b11hVmOpqVgyIDlyac9Ef2B0uuj+izcd5u1dxGH/U
ZEV6nSGUCF0oXRkabS+OfGVMwEaMJeQHiodB7sgGmrL47M4vtmW2VY3DSWCT0PSG
FobRMszNr3QAr7M1eLNJOOMIvs6SlOLYXID8HwV697wyipKdeE+MZjebNfo+k0Z9
cnn6P7tMbBvV8wkTEleus3eGeIGylc7XS4937otAEQCHQj7pKIAfvdZkSMeQoNbg
1Tf4FdHxpIX+P81EWt4jYJgPQV0TQUQFFazpeTBG8GZcrKoeDrqLQ8cM38nzAeNm
S9bOjs0MGA1TYsGaYYJLmGEQb88YC0JxITSEHjs/1kfGdEHQ0J2x+JgBkUlA1NT2
pB6uCRcI7KVOt2MxSE7vgq/ISWK+Zzsy6XgwsH4kEtfc+NuRkBTbA/LX0XPh60XE
HJcJeJQWT53Cv6MHM92YFGv0t/vLvj8hrolVJNXwZ+K+0rYFj3tOdbbahtr2Mg17
UAXOwfxo8LHigLfQOW34op4PouGzQ8LGOVstrPv60SnHRBLcRUoFlENKCOvMoHtd
OCasn2bH6gD1WhHMUkUfbM051fAxN3rJD3rttc66k7sGzi4OFsbLZARdhwfGDOvv
Si1gkOjeFHh85dEUA6858Q6Ak/pLgIEwDX332mbNUy1oB7gLyofhKf29rczzNap1
n05gf0iutnlOgU+iE/fadXiowhORy1knUALX71pWaXKdguR40vM8RN6WURApDC+9
K1qOxDaRIRTM09XeQ6FVQr3m2GUKkzqL0QGwTmj4eQisoFEbf3z/rmGk4dAXFpGI
/dhOZOKkK8vICl+XSZfU1T5D0St50TJ6Vd4p6oXfrZ2JZzPGmcHIwRlj1F/i5Qfg
CJF2C0KjiTT9dmOsojMuajlqoKhqDgsMc70k8cdDx5QgHqJI6Dv6G5t51sMVlh8p
P380N9HGiwZuz/yxY5zwvtFt9hNuqBl8repnc8QEHPVmPu/z52xCrwvMKNnDwtQY
J8ukp/ZXiUUn46pJADipyszbYgZTpoFkKFn0W6FGGET4sUiGhuHet8nOgaKhO2cL
ijjXqz5UU9zzNDoG4qeedLp12400F+FttLNYvpu78FOSXuglHm91wcO4MoPn7PrH
ecJcxu53jTIkyiAtnb4c09V4XGajD8i7e2Kd8AAtYO191T9nVbGRxqQg/HqSnihm
dewqhnv6m5yIKQ1LMiWlyxHH/XhCel2ipdIbLcTvhOgq4deMXEl1+hd8qQGvFCcn
Ns8ieFGgGyLzwY9Ln/G1oTDRoJbNEXKm86a1hAb4CG2a21slWcghwGGwvgmzX/Vy
DXgsh6u5sBJrSvLqL89pbmTflU5gCGHwtIf1Jq1d0ExvJCTJQaki6V9nww12n+C3
ce6XRSIYCpeFhUiQ5jaWkUryPJoissbY/VFme2oKfl7ZG3+kH7Y4gjYbmAOYZcK+
FCKrRkrc71iCrWkUtD1G9vMmW0dRy9Lk0oPgrZc27xKMSzy8Wxe9uxAUcIOZqBf3
iBNAi00z1/9J2Q/ZRXdgeW3L6bJCfl1iUVlfoXAJYz8oGvApWReuliC/GaDiIi1G
RJO1ba6v6W9NQNIj9iWtdI4lLQYB3/vyHNyd1jKKkAGIjgS7e/EIu/yxqWfG3bda
sS/2ZCp/e+49kBxi3TjFWm6VWZEM5IWzQkCMpv2hZTeafwfYl9SlgYeWTa/m+DPp
/RTGdIHB4jpgNrEz5FGlfLfH3R16W3n3R6yIenOf654twAjztgElo0UkNLspq1ex
7Q4ZCy1y9bN5dEqXLu0ox30zF66xWYQhM/tvaDD8vMRWojqkaSRPsrGQYYt5rRvb
4oLQM4I45fDjgGEE00W69P0BFZmsLJkJIw3mxGW05NSzcYSI6B2MERsOFQTFVlYL
XVd330Gn7FRLGcfwdKtHgSKlOpcF5ShWY9cfErviGSWu6bUvLStwQhfTb/vO1Pm5
VnroN+aliJJLqH888hhB0e5Gp0sw6mJHBHk3+/+5gdILpLFZmu4A8XyM0dQNx08L
IDUJgu4OOzDtscrNKlsjhW7ux/XsxotBO7ZjG0JmRg+DkmRklPTPjvwzMH1g+RWm
TfHtpkBot4H5I3QADQWUFyA4IwwrOXOVD+jsDDKgRpi94h34MtEpUEwvsthz5WhS
u+RSR0EKQiCbNI3jiBpZ9BdveumGKuUvsDUx0Kz2NrHVYizGuTjRH5M6RFyFGhzX
4XhxFcjwMxiA42jkTDiR4cdNqajUKzZZLroAztcdLF4cf7sRst7YLmWeUImTGRgN
EmMdGrwEwM0kcUmDhSWI+sT75Avu49RJlhhERD6qNonDgR1tAYI3a7y9jQ5fecAF
nN8j8zAhc6rCitEukng/wD97zanTr1ez/xGtJjd4qC0ls2X6uLYSGhnYumtc3sRL
cowo8pcDHEMlPHGhcVyYNP2EXAeBmCVx8paraHS4ORfuyWESMxZ6lWXjXu/3w+Ka
xWRIY6TOAMxS2TZqnimzJRVhgBF/V8WTQSzDcmRQFvMUHUZ68PbGSBynH8TBmkwp
W7SDHfQiSkNdL8oMn19O2SySUFEATxq3Ru6z841b5Dv5pCQlkN+fMQtgzrP5mAPc
dEM1PZZzNxCP45dzItqnWXRdwsXqX1Y35KFfJVfm8FWUoF+/nJhc+wa9EhSsEZG0
FXiZ9m0CSWI+lTCDn6PFc5PjCJL4Mg7N3xKVXO3m9smP4vIeV1aAV++tluzQ5kjB
qv24IWRi0lSbcMVPQo1BU1Pg2pZ8oV8wA/aRS6X6H2mHV1vQXDjSQJ76jJYGVC7i
r7rNThu763LXaVPXysjKtHYXHQe3WjMAGfOtfOHnizTHZE2Cixh15xb1KyigDlNw
FNRX4bAY1Lx6KQMFbMhzni58wN4vkfuaxmEXhHvXFB+qk/Z2feimzm7o1MjPIYoc
IfoE84qjYzc1DSgi7UERHY8MUWNVhKEsOuIBGvcTrYh55lHKmaB7ZhcSzGIMjh1m
zjqwGkxmv3EwnTsWbyQvobKzDL6ytC/93Oi3OUNrGM0ujY7/0KXgtR0FjnIC3ZjB
0S/7Ykh8UB5RHmvSRI7B+h7gNRVIeIyhOCwzXekwacNFsskQ+zUSj8PCzmMX36dV
Eke9qM9A1cfFfk1hdd3JueiLUspLbiylPEYTmsGeWhigTnX7pQb5GUS+ZzDaMEsa
1cZAl6TbNjrqhyz/l/bAbgFFLO88YblycVgajCNWqHWUHJwWb8hPmYxVlGubuDNg
zk00mL92pRy1BEA7oKtTnkgg5LhZS1WlK6Go4cpZPjxENK97KsUTT+8CNTKobnZO
KoSxDMsMXv2SLBa3UAzKAfNf97NpQETAFwNUve3peayap6nDcaENb7LyOOLrRRsO
ieP0cFZE07CbjrtmEzrct7ZE3vYoaKeaaBwuRz3HdAxVhhgVJFKKBI/QEa4vDQQ1
0plJdJUpq8Es4RJ85eQXpqoa0/Rg/waxzA2S05Uuge6aU35fk4XULmmKebIhdOlE
YXiUDdV3KPGu6fdpkTyhbF1okhflOprJsPLPTRBCv8Dg4iVDi1tR5P7UO6SmfbRN
49HhAu+72575o03e7EGIZTtIFCr1rwyXPdjI5DRrwZDMwKzjty5uEVfyNJjRSkJK
y27ihKFvhKCypfPFJ/hrkJTEDzgJFIIQoSDV42KqxlRZXU/n9UAYdfmX0xURbv7X
ILq9sMcAnFQmNSQWo6V7LchnIyEwYYgQw3UbIqDi0U3S9ADX6ikBUPFnP2SSZBOJ
UpT1o+d55sve31Iq70BWYDRzotVCpjSmQirLcvOHHmU8q49C5AdSHgZ1nAv6P6rg
LVaTrre6MdZursG4+tMrPgNmUu+uRy5d+uEi8f9txUxoWrCfQDls42D9LS4wNbNS
FD242Zqgnuv8qEtGu9FKB/B2EVrTayaMPUfRgNh+YZ6X0FkeWLO7RttTEi6HWnCO
lwiByV9baiY9iPkq5YvN6s9c0lkk9hKZ/RXgd0vl9TTyC6BTNWxY/1CbvQFXGqz8
Ki0jZEEmONQ7bV4E9G4RiZjBQfPqN19NwpjzrId3OxnasAEia52qrGd9Hndrd8of
SwFKIQLMCWOGGWbZcC8FftK3+wCR9ac6p8Ug2Wvei1lfZU527LFKznclabg3XAsT
iOl7ppd4pnmM43y12zjS78cQjwfGEINQBuoDRr92xRfnGapH5Yt+sOp+sD90cyAW
+WG4Sq8IpCbyyeyukdKHD4Y2XXUwttjaX00cp0I09ZyXD4NUVvtLxmBMB/Qx/wPT
S1+VuBR62skSBsmndki5NqB8k5d5WLs0dgKrbswGIvVoMNxgu/s6qgw8H7FCgZ2j
6QjnVv2GNNhUgWVcRaenaTVN14k/GvT97LuJJ+ja4hcG2mZUs17qK0JBxllCi908
Bq+gzdG1Hn+7ZMcR3kGFe+7v/YEq59QlmYsmHWwxYtUdDCZTRFO77eT4bkPmcnCv
Vpq1BbRBrq5gHuzi3RWA3eYVG+rtWC5xZOuy53RZ2/Pp51m1aFh1MBmTPaMBbPeN
rvgh6nJ79mjbHHbO5wpvj34v8yzekbWSxOQlrQhGVFprM6flNh/Ib4yp1N/6wUle
R0xJB79l6x3wfQm9YJ8iTABNBBoGr9u4cRmEN+fZKwKeftsbL0EkrKBBDrXmF3pn
SUV1qjyPXd3X+/DADjf2b+Xtbyr26Uvr6zfCnwGCMEYBT5lzti9EeE2OhB6nBtc7
3amoguftO8AYezqcu0C0Qax8QpR8WeZRonWp/F2h6NhFugy9JrXcWDlWhuKRGJWP
6pXtHlKuwLk0r6sc0Y27vRpVhF145Iy8NmP8oXTI+aaAOPY4f2EeOuGY4MiTNcPA
xzAE8FCpgWr2TGqW47x5Db8Q0NYYsDq0kzaA2jMus6Riqxk3fGN5/RpFx50Pn/xG
d7I8Ex9JPf0UUV7sIgYj70BDo/VvU3Jex+WBGqmxd97OAbP2pEqaW9sb8pi7Kp2X
ZAV1QW7rzvsoVnFY/GxgyXGBpLRD7QJwc8t0kaZT/mrE9gLsdKwuOLS2pIHriUDf
5QrTVchBWPbWyAdwPcf4S5yN2y5roUT1u2xVIrQsMV7L+Io+CCvcuCjlDXPDoMQg
qFah0zGDvB+eoUKc5bXAUH0KXLumX37XZ2BjCAm6SUVgPCDjWXJ8jbxieoF5jZht
O9OHoED0Ty30Kejj60RN/UC6rroySvgT+fj2bWTA9ELqHkS0Zr29ef3a8jKTbJfK
JzdXbyPvk1rBWZzvceTjBW7iYLIrd5noMyBVbpDqQRn8sdjc+hDVqYwr3CuIGe10
9x9eOODDScFDfWfWpfIh1eBbO7GwmXuhtNmzDCIe3AO0nEG5xgXbfE/NzciLas22
halq/1iXgHmgxE7Jrz45X3UTpZSGIal73UcF52YUmc+yUUrCQaMaTokAaY+JGUNi
JEV0nRAvuASChv+n8WU5Yo/Vfe8kbXM+Ff62NeouwuPDKdP5lBnfJmbwKHml/bGF
R228Kv59Ixl5cTzfOrvw0Qffexp6yajhMq8I6kGFxmyPJh18LyFepIsvP1vmf89k
exPIvtfHjRxF4mUNlZlDQ3s2RQIXDrSG5fUC0w3Bad4TMhLwZgp7GoPiC+ezZNgS
1LIoZ7xgc/9x879BpeVyABWGnxLjFQPyDkRV3q7Ka+Tgt+gJ2maFKs5T6nArIBAo
K8jCjPYEH8OpP3v1RIiDkCxiWTUywKe1KEOTFOY3SX2CNbmaDdS4bVz4X/Cy2DPz
9N5qR9TZlG5IApSkLq1ao6CnzNol2w7WK0St9EABXe3dX6RLc/7ffJqissgkD+Ew
ZURGMuiYH7Szaj/R5Y5pZnQmtvl3r9a1KS7ubRKY6TxuwdhBLgZtm5+GV9YOAXJn
wMjqAjYYXsTMRUtqzsjhL3qXioRmPnagHO/a0FaT0UT/zKt81NZ709P8F5KYw40z
GkQTNkYedth+dfND7uUh3yVebqYiBsi+dTgqz1V4hzLEA4ZpoeUCbuqxtaJ+mfYD
vTt8LzV6cUET74ciINdV30H+gb5IJC+o+GEIutxtDeRHSq72TbtKCdXx0Gvhy+SN
il1X5flb7G456l4NwpFCbb4DIG2+eroQ8Ky37M3DK/joP8z9fFgTkpqXPfYpIq34
kN8/u5Bc4JDiO4P21ub9tZYL/UDsxIptVa0RV3p4S1Z7GXqb4WjDe5vl43vIVnzz
zgB6FX0P0R8Ip2dFr9gn3TC/FUV1pSKgV1IemQoFeq0NH+2C+qjJ16mjtXCrRHIb
U0QAJkRq0hUt5peYg+hvRuUQcZmGSrSU9jQBA/ptG4BOoQ2zEelUZ71/5RqT3UG8
SXFASZ8HFz8d/o91+PQ2YV6q1k4wJsdomnU89tjHRpbSUJceFchbzRhTe1bsnaJ9
ifD1MDIc8JeIyOcpthTWLPKVE91kNExD4w5/UpELgaNDNP6G1qYd3QV7MlTrBivx
2DceVezESEIOxCxi9EWKHmJWCUFgzIUFdrJCFimjk+35uRPkyXal/ne0CARVH37E
RyyhvMg+0/ZqXdA42y1D0lEQaakTONisgIqgoTCdsskvB4N5D/brVrYAPEdg0CIK
4XOoxvKdP1ayX6C7HiWwDCHhys5/qJxIozg54HJhmkE8ugdYQyPrIYbgyoLqYSqm
kYxmQKhP/DSEWq3DwjoM/6MLQgrmy4i+rR4Y6gSsRtSV1huJR38uU+k18bdT1LEv
Tdic6arI3/eNfu15KueSeayWNiv0zQHRvVOGMBIswn/8svweiKhTN5aBAk0PmCSv
gp++ER6PzX1Wr343DM6vbkE4vb3+uJf1EwRjFDtWTPsuwWak7kJdFkMzgCaBvWGn
99H77XNzTyaW7xzAXThpCllJRSlYFJiBSwzOenCj5AsHpk1Xdw/GUyGxn3Uu8c+R
G9r7QnAo3MGDzHXsW7svrBlzpaEm0akgedQQjd+aaUIIAuId6q2mNHu5Rod3Z87J
KoCGwkM7uhmFLSXcteAlHNLumm5VBHcVnkXMFhr/NnnOeSGqrWThdnbMRAR1Ldx/
eB+0ZshAHFL7569tXBouMD8Uh583cnrat/nZUEarq3TZh8A80G2baTyCQZcVfiN6
QKK6QC5zBxEZoIb8xt7PB+f1ytQiwfcZlvcXzLFTtUmutnemOr3gGdNglGi6gGkh
7tQs519JwYXbPop8dJuJC6a14kvZcmzr14OhGbXeYrdgwnm5By3Q3N+Uc3ViunFZ
t4VUw/QQlr9lutnoRKwTG4C45jGZ5vqDea22j1jXPYOHgt5U6VbRGbvawaT/wBDM
GQw/UJ7I00/PPW8mVJ6BCYcXj2cVYCDIhh7pgXRIdVFwCCw5ERR46CV+NmwrMAPF
6jlzC1povv1j4ZVtZl3HFZuPGhuo+VkB7Kun/Mj9bE1L25myQfI01qnYKCOiyIvg
xMTfrNG9nRxcA4umAI2XCf2mqu7uDS8EAsSrsLqdM+ukRoc8rpuE3jiCiPqGQ6nd
LXlLqQrlSzPcDjQlWyA8cQUYTicE+vB6CGwzczgtWNpLnCvqKRoLnzVMCm1NrQ27
khiRXfeZN+Izren6u3RYJ04s4Ocswu0/jpLXh0t+GE4oJFBfju5ntI5VJVi0kh6o
0qqUYL+ztvrSfsdGSnw8QjX8d0Jy0YqqWpEhSasKWx1vWwYjKy0fZVj7ZVDncnb6
kgvO91eWqVzCFEkBqLgo+im4Io6VEfgRTmQ1MQ9A6ebxTgfMTWpWakAgMxW6bb11
MLn6PAXWGemL/PXKCYkwUXJaxQUko5RiEmdjIEgLf0NX1aWEvLyNp55YBPkySczT
xGtFfRWje0jZLlz0zjNLqHo7/wKi7fW4xLmrefhcme+c/jJuEzbHYeTJYZNYT94v
RfQIgos8qgw84MGutYU7FQp1BdRAAqfqmIGjgLe5qIFY1CrDownXn9yV225SSlnH
2lH+p8tkR1OoFNKnhbSoq/8tuCGRQnNptMF8wRFOKfFPwWF0eyXTIJn06w+SeREp
iIhaSxIXOBy+GwYT6v79Ju4KKMNA83pq+1nXfidGKHpU3Jviz+RVotkHlAaVXXDE
9VBpvQ3IoKAs+zYgPcOZ4LKBiRbNT6aV+8HqbfGSyAY8KXdotbRMS74O4HiOKI5a
hNcAtpdhCOcZ9TFfqulFDLF9AIFAMNgdVUKck971b6CFAgUMKub3qNsgI3HhqL+w
LJx3gRsg9H3sht8CtEHuPOi+JoiHK+eiMr5Lzxj68TAgwVmH6yxtZ7TZ5QeJkY8b
hmlb2NWqTQTlFfXMNYCOKLjXMFrDAFRLB7zUKCx9rBxxX4ekwSaZMyoe7mdv0ywZ
OybsYkenYOf/E0DpcZDaEH+8elo/cG5Y5Mj4L+79z4JRFT8J6Bc8rLsIxWkbRQXZ
o1uGcfY6HZ6BZmPIn9W1ROyEgLF8SmjKt4VIElDiGAjDAFcd+F9woouqsPPcyAqL
UK6nnaHArCN5AeKy2qL8+RqBZXnSmS2xr/aN1woaTVR6kzjUSQf9/RifgZFHeteE
nGeimF1sRvsy8q0wkj8tqo/Pq2BU5tKHrFy1jvavu6z3672f0TNJ4m9ZVp8xSuKn
UPOAIhdcSevVZ/CfN/ooIssX/l9JE7Ap08txpjFUXvue0kS8VbEtiRSetbTU+smD
VQiDAkFeo2zo81cspNEyFXra2wpXmBFJDNlR8PJA7IDBQGKYN02EDBAYWIBvhOBa
YYIxN0G1jzKdA/irx/ihN8RoQ0wOSOeCDpvIg0smhUEUfCHcyqQlz6gk2M+Iud27
D0Wrnz8JpnGF956jrYkTDekPrdY/D5HdUxuAEdySxYSBPk0W26O+ftrCBIOaraFM
xX+nKxbD3GrCjYnmyRz22adAn/ZoN0RChj9E99PYalSqtGnquihQEx7WpN66+W7i
fqcyLd0PT3bTlPejDf1k9Urk+LpYZ5fsFRmNbIpcdi7S8HO8NF9BlPyY0O0VUWZP
re5spMYxbLpRY6vtRdbiJ7scyDLCF8Q6gRnYKakvIleVjeV7sxYUIggVPp1Lzitj
BCf60AKWKUr4CWf863rXRk4F13DjtDYVrXXT7kguBC3Ho1LvzS+EV0aTjbwIOzYZ
ErcpWyfW7NfrhDEYlMZbHf5VV3oNiyZQui6+xa8MoJSiwp13q0eBcEyP32p6Nr6w
RI9S2glIr1hXFK0SCApaiShkw74aXt4Pw7XoO2SzVYrWtxyZ81cs8zXQTPn6wPQH
kBo4ZUXVC5KVhjI2MyObzZVXyiXgJGw2EvMsoNVSmER56MRNqOsJU7dUc4zLYL1o
Q9TKLp69iCSnAHiYvcrH8YiaINT9ouIUo9mHnKbaJr2XAa/NVg0bo9+o7EyXnxD/
Cr8EYW+zCdHji42CAESnITdHLBfy056P3jKjZFBleheeIGb0hHiyeaFdDghudyn1
YOBzeRKEUENaPIy39ey5wMxjlH84tASsAhCekjA+vVT5Mv7q64LPe+AD0jGfwi2F
EedEP0y0ESPDy6YBnuq2L3BGxyKCedbr2DMO/5ygQXHT+NAJ57d6BqziRUBzN+YT
3aWbf5S7BczM6n5C2Jrj/nNeDvUgXEvOttzqlQnQMCzEt60NXck2FCPioU2OFoO0
eaM1XZZImp5M1ygDs7zMuiGSpVsRhP0DKZjGpuIteemEdRkoV4ijAO6DizS4L45i
o++4D4WY0o4LCWvcjjVK9doH6dMxpUH+TtYdVL9+4Vc6nQC/hX+cEZUSOzLJICUy
mzmvUIPuGwtxVQwYTRbUeKt1VJksiKJgsGvBSR62lnb5fgOecM9kKR+B3+Z06x9y
niW61roMmARSY8bIVnkkPkFSmrkDBdNzQ7ynKQXrXDIsfTv6F6DLM8A5F/S/riU9
4HWwTA//KZ7PlmDW3vzZiyiVZAlJa9PpZogVuS3ZMBnoZ4a21NDpLF82EmBxqWA/
ovJjVM5KOZRRYQJFsKdmmbNScdemBzFI+sonJTvUiZuicY2Uq4lkx7GxBVgH5e+I
DCLj9OtO+FQBRWdl1uBFxONkekauQTAZckD8D5alWFnb5FI2hKbqUPdbNUPOKERT
xLi7noGSduz6DFnDAH7Meb4aDIUzKuf95Sp3lGpLRSkoWWb1waUQHox/OLBFHxtS
F30KFJFEf0Gx2467lRuPEtT7ORkOdPqYle5fNCQ7+rW6rwQhPBiz5L5+5o+N0BdS
d3eK6oEDiqupT207YVes7dV0hKcXz+HamZMutnIiV7Oh5s2RqCUjctFfqAQQ58md
FqOFkCquVSkBgubnCM7sYO2hC3YRNdKb3Na66HawjZrcC4ZwCDr9uT6Qz4/X4R1T
PwEQKMVqF47U2rnQMiX4BnbZu4GPJd1Z/RpmPLUZK9o/OHVJx3VTQlh7wwpqJY10
0lB5K6Wd7mdq1cZI/3FYpQw3Vn+p7RVHD5XqVIltNS/Idbs8n48Ct5jl+4YMb4++
lEW6uqh7RG9YxgyLdjXZ3d+VDnso7BGfaAljQxrIwiTFCYAA+qj+W2KkAorEPP6e
aT/GDsh5dZnDnvWB8RFuqCV+aGM4nusPu0T1CKgEifetw4wqBqMJATe4ew0qnLcc
bUrn0VaE+Hdj/3nyFIHzMNYeceuyuHizflzDOi6fZvKvp5+Dg2fxGLiGVRHXd+u8
JpBZkyNwpVwLoQ29LkRMwoTu5ezMCu8k6+VuEkn2ZPt5tCsrWOofSGTsN3mbkKdd
uRrc6sZQQwWMDdjFv8ipYHVEdvUw9JACQ6mqW2n9SpFst7aBKHiS/BOw/wB/vzy+
XQ6QPczRfQokjA0hGZjs6R8WlQ2GWzkKopy1CHMiZax9+S3NxurOWLOOIzcicaGj
dXwyTqzuvZx1fZwY1K1B7bK2/2zEj5n4/svSm0CBW+rmYX7a6iTwt/y/0Y2WABG2
LFFjQYUOVzbs+4Qc9qRJpSIIiLoP1gAI8FRrKHlcxsApBnlP4PW5SBMJiYi+hQ2B
Od0jl7kmPPPYhwDaqAkuv5horJcGe8rOt3njrBF9qVES9D6Pa2j7Bi/wsLbZ5NYQ
c/tSRFFQBrMtr5hHti4WOSq77wcpzaVciOjUo0/vF3zZvNl/wTFYITsv5bgkYlc0
NA7Ndc4ZCb77+aElMdAl+HW+bej5j5Z0GFargd6jZHMDTRCe5mzfRplnDFQQefuZ
CnUsVrYUhUp3cCVisWMf4F/worgk4YJ1Kr12Hm18jWPDHKZxHDTI8cOTTM1pNSIo
wxleprQf2TDNn9hcAq7CQHEYlBvshif8aICc1t97Q8TY+5cWXZwyy3vrx7oxXoaL
2fWk1iMBMDGn7ORW4G4izm+ubC6n9K8w64Jv7BiWUqUtidz+5P/ORgUnRqp1kDbW
VsinJVatv7d+zaQkq2Qtloph1+Lnbrs/I/+1DtBtobLX1SSVo13J5MSihOr0Bn4o
1UzPDUAKhWhDHwMD9yHOoGl69ozAk/6Sv/3j37Nt0031PYUMOH1livnE++RYIirX
iL6L7p+EkwE9MN2GOhmHLmfaxMmVrQaDVwahqC9lgPddk+0ePCi6uhMCIeHgWMHj
7Q/IZvZGb7cWLuHsRA6gDrJDZi3pBkXcc0rIVF7w5QLDRxdLnnQ2LBqxWw8XcWwO
lfwcAsArBN18nwy3u9tRXsJE8n+vPQj4wPz9fpVZlbQjHWE6zOM1xJvqFPElS0Li
a7L2SruG3KML6lLph1mh39qMoM9xwOhqwzJfv8L/6w1x8hEA20ZXhzBk/Jqe305y
DP+Q8ZMOET6WY2Fi2wxxR0L9uRoJB4uKWd5rcaeh0zcH+JWqV314pBmMmRTUxYdX
PJkKT9AkzI0A5Mnfqw6IMLkR84Ak8/6fIE9J4aRiiqnMMC1MRfDNup5wbWkSHYyp
Y3HzcFkOwZ8c+XtV9+dcgUkKNXkgtALKVv6G5yYW5cDjHhFwGI7fpJ7gYhWRhmri
W8LAz1UeJAOPB4uAYU+peQMZ5Pt3L1VNnjW35Xd3qZeYNqif05ygLpAV9s9tkhHJ
3L4hGF4YzmVNwvBC1Zr1n8QLHqnP4Cfa94WAmX+GB6V67L+7JctaFUIg4z9abeXJ
R2nSLiRO2xGpQfC3z9/dsdI6Xjp+4usZkWRIRoh0F5EVo/wHK4+REK0nmtaaY5ja
FjSjoVM7CJHx00DjYlglNQxkDJo0iFG+7NEk31lwQ1dJKJch6Lyeg5PQ3/QeKS3E
w4fW7LD60KEuylpap3ls9JzbQOfyzkPqSYR4wv0bzRnmKoN2jM3cev2yw52C0YXM
+zcEVxMd3kKUQs17x1m1OnZCS9WBij+juZX4IjKjomFTDSQuETkwHXMwmAgPqiFg
5eD+KlU/Cqmn2j8i7ATleIWr+UlSS38AB0XwW9U7VaiDQrvpFclRfSYddkSRhQ41
qoiwYBpUVfEPgEYfHWqC4t6js2iueKLTtPgDfj3H1WPVOG4x1gq6g4CC80G6Cqhj
n2/GLPDsBXFkjrzbgU2C0Y9u3Zv3nyfsluDt4EzIzYM73tLXKgzY2I9yH//cmabs
yFlOGTCatrncIoAy4lF+3BW0bhEwPlXBUwSzNMdSAxZbh3LUxERznAN+eDl9S92Q
klLBsKdP8g645OGTRKwO+95MpgMvLis6UpJoIOuMvAbQjsy4xR0/HR0hSD16FrFM
FuxPTtgegy0VU5bi5qHhU3M1C6dgaRhqwr6YQgUTIiRUP+NBw8Jk65jyBB9A6zRv
bIUMA83XRezHI4oJaPbJN0YtpiftZf9Z9ftbkPr5BVjqG70Mqvu9/3KS3NdOFuWE
+NaJQz1ri1yku6sSs8AJrwOQZvUqg+bs23BvOeszsU36tyqWvHVXhlSPOAx0bCfR
Nwh1P9hmDJ6q52H8St291bBpANeuKI2NM1X/0iTZwjpEKKtdqEm6/XXRL7Sqevcr
Yary6Ekbo8vcba2M5Ma1dC9MaXQwE8W/vkCBu/N3n/CfsrrBloXJzJ6naTQc67D7
dxuftKCDWJb1korm7GgANP/6QPjvtUycOSKgqae6lcQ2SvJ5wW4XaHl5/JZ+5X53
4jcFzMeua/+oSW8X3HCFTN3NfQae6fF91ACksxs39MUTDHF7ZwaWdeJw/OjsjB9N
to62aleXGBxfQml/3ocsvzoMDAQUMNx1yTFbGxf9WWXBAOq2FvCAY/1gfFLgAJ/B
G3hUrRQrj/yE6J/tl1XkJlEJ6Q/Pn/a94KH+F2wLJWVF2F/HHgR8mMbkPmOraokX
OvMXJ/1GMrSdm5rMNPVPqkW0XWaN99LLdRUwMNwY4ZCx9FLm7TpD3mPUoDwZZ2EQ
L/jLdrQ2FBho9eO9X/Pt5HxmtsFZOhN93DY4DzKV5PRTNtmvrqQuTzelOMfy82Il
/iC6LE37DbHOHiUAHRBKhpygwpaSHHi1aG9XEWNr6uDAZVaCxAfSGhPr7WYyN8EP
5+Rp3J3XT81vgVxQCbA056AW3QHC6oMq23QnGGvJKaCcTkBZIWQCP/uUOVUnx/P5
shCkwzmWU3kJ9W23ZMAv1BWM4lNXiEeMnNyOtz37KoeLbGrDslDGEq7MCI7I2go4
ESt1Opz8ge3oscK0Oyp+gnVZMJ850/ZJJbm875XRov3hDRj/dRleVoNCarMTRjZ3
Qf8fdAQPeUy6S1idkJiUacIC9E2rCcr1/M/jf9b+5w7A5XESzjZDKRU4+tkdDwko
fbsthiehKKx5sNPaWijE+/yovXF/CTmDQ1Hp0VKaxx89VX663M5BAmAS9VWUoreY
HcWupz2uXvIPt3JwQbaMn78ck2cSwD/vcBXXlXrD3IJneROAOTMVsnR8VRHu397g
B8Q6JAY0AMzn55wgJHpMxjlflh0VWvTc8Mr5c/fYkO081I37lmnXQjk4nhEdIvuD
GjlDsEcpaytCPjSl3VypUMewwKloBzch0iROwvU9se4hQFNMG60FDXKrhWCPhqFr
eLxxh2TNpwEwE2ozhQTUPd2A/h5dDrF3CNzddVtjduPobf8UyGUhxF99/d0IBe0J
XyF7kd3U7kD9cQskxSVcZazkcwtnPhVACHX3AxADWr5TWabrTwWPGn1bhrqmjPvV
PLnnIcOSEb92i0UXeUho6YTlKvqzrY9PydPx40o2kQeOA/JcLFoZkzhEvezNr44F
kDmjTJVpPlFPEpYj5z3AcgcS+YUduTygeXd7jVqM+FqMafrN4TL8rYOU9ti1hiwb
s+2AyZGkCMR1C5zdJsYRMmV/aLdMvh4jN2WyY5mdzqXpRdeSgoiQ7fqkYUK6mMrY
pv+hnhH7++d1kBy09rtb0JKBn7ey0fWzzVbzq3AufcvrpoCqTTw/CmaZJYt0RvdU
0aj+ucdqH9xSrPTKCAu8hxSzDTzhIACw6nh85WlC/34rdNzrS0+JTeleFGUOmhzE
WuZf1yvcmJYepaGH+hvSDpTyCgV2WhJzAbJ9UshdAulnPkb7+0svQ6M3qj+cOElX
v8RfXTAlhELGykQUOoWEqpcNsmHmiZzxWW/a6WH2O7GO/R2O/dzfzBRnWTdMhOEt
kQtC8xQ5wpLfLuT3QdQORSMkpD5zbXkEfIhsX/C57al4iZsktXigXRbpBCgCnujL
zdOXT9MH/iHsz5TkC8pmR84OHDlLDyxj70Vt+YqXH/JwyUR1UKAoC+9MXVm1ivmF
adLRK3ZYGGnHsazMKB0BD1ft7JGd4twzIdpqR6Ps9Za5DyjBSb+PSqhpQx8AXCxx
uEcihFJgIN2c72eT7jf3GZHrKzlb9vZNk4AMslMpNQnrUxpEARqZlgj4Tm6MjaKW
OewSr/xJ1EM9sirACSEkiJ+AyB1Y6zeQQzWS9EaNwxQ5Tr/Ky76lvzVP3aYD/ayv
JPHu/ZZ92hAy1wIlAbzL9E3lAXusTjCfURH89bPB+QYUxIq5/5KjJfOW6AKn9jFm
B1G6CvGofDI6oT1RPN3D7nWsOGq2tqOKeziRr+E0KQ5tdEQSvLvJvrw+5QQ/Uc/L
fMVfl+Il+IgFtIjmo2IUx4NsIEmk0HOZylCbJF3efNH/EdZBuPA50j7mPpPT0Sb2
YGs9PH0W6HpWt6KEDkYcWprcU5kqkvUmc1pKr/cUQ5WmFLUg0e739clbSY7twxme
KdDyMLDX/EAQeGHf1Xu9uXDohRYsQSXmuyhQzS8MoInAFdrBksl2sfduULMD3QdO
I3VQXi/zaiTTOI+BdhF/RhxSpOfSjnnBvuuch6iTbxKq5Qc+dxJqm1N0ZVwcDcCt
tfKUo33GkuVM7uubjC16T+0TKnSnmVt4fpBptGejdG6Lud7fFR5zWEQR3PLPTSCo
aSgAcyn6gV0n2r8yallRqxWqjb8GeZ7bgIKXearsERgUNEm3m7Iifa/YqKj0NpvQ
iTAIj5f6PPTFOhyEnhwYh/qcI29LjOT9IkmOPfUi2hw7bddqjS6r9A8Ck0Kfhzn+
aiJkC/Pe0wF28eYpIolZwo6RmaeaCF6PCNsx4SV8nk3707yDyc4N/KLpwjuUVM/M
yV+1eNml2JI/NOw6trGAPxuntKAKVQKsJeI/XCd31wSt7NCmxlY89bDJOoBtX3v6
A16nREBa+oYrCZy0udYw23EVZLOWJI/8vdYlZzd/jhfl2KGjeEjEhSGR6kY8J6ER
JFFWnUHr+kpJ923twODYaW7vIJBQ81DiA+LqKlMXdH3O4Fb84zosR76MDNwCRtLB
6ssNBCaPspowUvGvW7KDtb5v4T+ebuHPEOmLMwD1kpAd0AmHrDLhpjpTaDR0UEpy
NwaqtJVbNvNvJ+T3sMXEj0Qa48o9/qJhwhjvKiIWQ8+3fxKP0T3fpKyeRNIAM0N8
zIMOtXDYy5dazpvjtxB3DkSIvWKW+dTMmjCzqQZCJ9cQj6VxQFkajfqGfVUOXeaG
JJTGApu0pyZcFSbhFADcbWl3SRN+bqkXRuFiCMABuyiTanPYTvIb1MqjY+A+TW0Z
OlkjSUUrJVo3CMewf7CIACrVtngpRq1jqQG09Sv2m0F0MdUKNTydTg+xPYJMK45d
BR5Y7chOePty5VfQupCOCU3rubqgmGGb9m3DE2C97X4n4r8KRjxI5rZ4uND0qL/W
1Pk91GIB3fSU5ST6sbRBgxkRg8mFtgHX6rpydWk07JxdWA0xCf7UD32W2eevc3Z3
Z5ihpxwXdyz5FIXLq0YvA8QZlzVdPYTHtquz06fthb0XOd/KDF1vl40FXM7ezedk
d8tgoYQMFs8qDIQhmNAgfEpQ9GFZ3rVOYEuCT+UF0HlPy+sYO4Fa0nKFOLjKt/jn
Sj2wvZY32KuhFZ/ONRdE87DAPIa6QeNumdBiwiKr4KYuHN7QOSHyeu8SiufAq0x0
nuUoakpa7vtx76YU0i9mT1FrLjTGyodZL0DbFHA6mzvTHO6tJWyobPBi70lALBFE
8JVIXtljTPT2o+mSNuf10gT+grtOqX92Puqg0bAP3lphwKqgizgq4jlV9sioB8xG
ZRv6QUD/kSPjS6fEu9vL9t5GXgAQPFexzdMWf6SqqmyN+DKrgz97LZ1FtcGdzwWs
xvCDFx2YbyWuBAMgkhNareTcY7isiIAg+9wJ0mbpJcSSC2NPMpfKbJoN88wmdumr
6smLx083KErUm2w7dDyR699pCGTs0wDqIPLZPR90MBzgXG3l8E4Fg6iti+yPSSGK
qVF9rUAs94PEJHaidxyeV6DkoDwmRco2K5FODVDkBzIYb9ZcGJIeIlSsxZubrjPW
pEB1MU79Jk+5d6EK1PUYg4pYNMabBFdO9jhGU1HljT6EYkIrDsUD7Z/t89ET9SEb
fOR5dmutQrG7jsF68Hq98fvUWGuD4IS6RrmzIYD+VQQYODJAZ0/1wsBN9kns1yIM
Z3OtAV6xqZdXi7ESOC4YVoX1IteQ1jg3zqmc8q1ejHpAk60tME7DzaaXMJpHnmuu
+BtqvdVIDJ3pdqR0yYUtJneA7T1vGrOEK7+Le6kLvzzINjKXSaVR+T52+ozs8fv8
0oHvtm41PCBNu+j8lGfVPp/6+ZJRjtsh0Rbal/0BR4rOvlcndwGwpN1a2XOCd8SH
ukXg/mszCwmZUX+u/MfBinvOfpMp7bnG970Rhg87jHrtISuuh3Ls8muVRFYuqKpO
mR4JmwWV4WyUnmkvPoO6ZaR1VmtqktnLTSXkHZc2yb9s6tbovMWFrIl0Jt+yhnbB
2I1XFjrbbXEB0RScIiiOek/93UfSBCYsL2LOjGhUK6rprSXq+10YnGCWO3X7c9xB
nmfpFawObIQ061AlZXaKBan/wxZmQyZef/Nk2tcPs5jTiQTVfw9Via9Snl8NfRQh
DmRIIsqeob3yczf0NE/iQdRm92ggQ45XgWDtCXu22goSqtgoi6wXF/sS5IEPo7gr
+vz20CZUJj4hPWhZu2Z/Z+jsXFE8niIQMdJApRxuBs8AlOu5dubxxLrAmYdxvoPq
rc/bi4SIf1B8l/oJAQGp0j/JWPOGNFthrP9Dbz/DbDWWnDwI51uFWkI0P5X456Rp
DStvlXbj/oEAQBANG6EAic3gcXjLYMFrj4hImuOxTfdSP5G7us2JRXSJhpeqXKhu
RVmXUvCJxkVbSgMW7Dbhr0wyb1dFVZnyuivdPSpg1YJxPtIXTsZFNznOMY0I/WJE
Svx6xCrFsNHEuXFQjMaf7zwUDTKpiq0fJNA03fb5CFz4RdvAKzR4DsAfZEfTEj0v
LHyQIE6XJz5/c4+AM/MfQcAFCtlBd92999f2wrmonsBCHZ8BubADayYuokt/wRCR
+H/JWxSdpGsmPoUPYVEm+ahpKSCjzgtLNPkBJS39VjYVoJYOXFSw9kPX0UwwFtfJ
ARrvekNLojlt0d/FIKgGYhk59FAnD9qb5dHKEspUvXk3Ts6k7x8HQGHHxtL5B6bd
dRTqP5UtWfJ9nbwjyJlWtp6GoMNdxmobAMs2rrZypZOaUAOZHNsi2MT/o42PKP6M
yQpWn6wK6nhOvAuZ12CxdyhtEzkRE2GUQgPlGcV1JoTLJ0w5uagwY09QyE7CwnkQ
5bF8bNV1L8gXnMfUJF25zMtSUCLsb7igEzrUe3FuYnhXw97XIDxgCm+mYxswbFlJ
gTaqlTwQj4GNr20Qrj7jPYSuNsAt1w66+2sPw6CjWM14vAori+bDPXI42p3XDeZH
AQ6e/6qx7wx3Pm+oPA08n7vFqzlj0O7bZZyp635xHg7+7w8qnIVixNqT3NL2jKEd
nLkXoryxwKsPSqKVpVjnLjPGJh78cGOpmw9zmkEzRaWsGQBUznhkqscF/cW0+Ykl
IvA1BnIMUpwwz6qRTvobMzms1SyclDe7MyqzKFOzsdWmvCOuJuvkVUxjUgNBuxJU
GZLFxKXrJnx3vASmprQmV4h3oAT/DHEcdRwoIe8g/a1Ly2DoGyjUg5bK9dr/Oi6l
aqpXUCGvgvk/GOPAjjtNcy9DC71IK5CGlOF1x1PeAN7LGQ9iG0QiK/vSLczjeIqt
zG806vZJt4JxjYLIT8EvYBj26kJXEZtn8MGCm+ik02nAm1WTfu716fu8YZ2ZX2QR
Gg1j+QrmweQP7nQYBDWEgg4a+cDQLqStp/nqxvtFq7uLLixSQP366lxieB8TSrKB
enh0RbUg9lQKl4v3IAiTucMltEKXf/zdnDRgT7qwx56RuIVHrzhKssTIIjeDWmLw
y1nWsJfj1skAMIC+aOm1Un5qm53eGv/Zq44XRlirNsdwBpBEjb+2bv1iMlp0yD9u
RPL5uwUPtq3YmzRodgiO/qdjv836bQTZecbK6TJnmyc6k3DspKD76PgRaJNOuiDe
Srv0gpbE8mF545V6y+77W5z7oUvm3oQ8pJQsBH/2uznLbd02JIqXODM+wewOI9mG
yumcMPXx6TA0Gc1Td6qoOf1Remw+CBX17a7yaGjtwT2e2NVYMAT4EuFbPBuljm91
+bFC33qmgJJJHrfPlhTHTgdPwdzZ86EXaSYhQbV5YaYFHwh78oPWv++wBBdjLkXK
K8wvSP2Xz9A07Ia2yk6gqx6EaxhI4XzgPmnk1L/UC7wB9Fav4hDr48VuqSFuYwOX
5lqv/W5CxEiuWtCT5PooTuV5StB4FzK6GE5z5SEIlKnkdp/aZUw8B3QI3NU7H0Xa
VzqKlvS75v8VnHvWbcpRit1tmpW21L5Hb4tHjQP4QmtLCRDwKb/pI7Se4fewC0W/
fcsmRdh8hNlheO7Nhs39L1XnxDbKJyBMKH0t5I013kcFSDJRP63C45Wc+Zl2gwpc
5EWcojaw07I2iMxSK95LvDHiA4kmxQGHNck30xVWZTUdr6Aa4/z5Jll7zYv2tccD
X5a3jOtwO3fIPfCQqM1myamjd+nanJ9XudID6vUZvCRWUWvVZbLB0vYzgC9ZaJRW
nUZpRHsC3EzGQuaXr6aqu6e0jWeKSVkT6GXXTTqwqjCiYBJQ5PDKEuuyAtweLxI1
qR3V4Jb+IsSFqOBhpvIjILs9MdTPWzcb9QDjCjvIMsLmIK/XGvwslhE3WLwmyrkx
bEHAQz5fveqAKqzB772kSt0eMkMpFb0+Fe0Zmh7p4fwAed2zW2G4+FjYo2UHVuzm
zcMb6+Q0BJmQ0GPWjLU+9roSDWYHRe5dtYkTq58ikLgKUaJJl4Nx/v2pexnDg0OL
DoCGz7wckKzdOjzbQIDkmmoW8GAWzH0pMlRckoAwbLwqFAc6whxaVzeQwpqUY14p
g7Q6I16m7dzbp7pf8kZ8CMQPCFmlp69CSqy5Uvy7ioziwGQQJntIRfcEo1ozapou
nMNv2c2Xhq+iSgzaep7N1j8NYXs/bi+ICGFg320kQVJaYT3U+CA+byo5BND+x8LV
Fv7p0HS0lCaaYgO4zC1O5cl24bkoHwey6eZ4FWw7C+TTSPw8ccOQi5leHiHZFZ+5
mELqpPJUoMKSS6o/5ia51fn31uakiF127pFNz/LZ9a4+1S20ArXpsbxsxIEpkMhM
Z9qJp9drakgfXM93gjFp57cJ00WAz2w0nb/4tR3MhSwCoTuZj04GZ1fTg3tu+cpf
OGOcQwTsAst7a45F92C0cCeDfPYF0qnqIAX12Pp5yB1ArQp5GwBJ7gijGYYm+Jjw
s9tI7vDCPnNkrJVIhuIOKT2zovCdqcKAFiH9efqR987JeVwaxHYiWp9O791ZpXKA
7ViD3uOktfLBEYmTFoSc7o199BN0UvtfScdDmLYMIdyyIXE5su7KY7U9IEGDMtbW
R0ZHcCpPEJ8flbwN3l00SpWqy31Z6mNsJUZeUgbSjGbDMKEZcL04i/KUMKH4Aycz
G/5b7dJCGoHG+ToalLP2uOyQOFNsdbsZvxjxgFOMQ9ex2/R/BCz5uBvrpva7BHqV
RquQCF6KM9JXoyHt6cWe6+PSKdrGF0lpR3WRSg+g3GMqsfS4PIrGq5WHGd+pnMWK
22iOzwjz5zegG5/6BWhUG+wSBz1y+9oksIN4uy8Boh14vl2ZIniZCb3Gs3LXyGJS
rsc63NsmjVJIYBLVXAggc1IZBFSM2iJCEF4Zuqzbeyu+UaQk4wSH4bgKrTXhS5+E
ez1ahc55BMhcKq9NwVIOMV/vRNweNk0BQpO050vh1DUgX+nMVIbfRuX261plOwJG
MxtqxKO/uYfYcGVi7lmTQT9If8m4d6tjiinccyicZWOw2XPONkZXI1IhsVNdCse9
jCgTnmsr0Jjlcwsgo/eDcL/GY6l7CrZh823Ca39EGD3Xw1Htp8nBj542vgF7edVt
rJLjYc+D9MtB0j+yUzm1Z3BiHd5O5d77x/tlFl6LSHG31cp4ZXgUTd0Sr9qpJC+s
CcSSa+3OEoRxHjuyOsuI4bbSDCOs7B06lrdpDxx3hV5Yh7MEVKI41MYz6AcpuIx3
Toll8jMO6eAqcqwveYeB6r8T/q4JqTr/a2L0S5XFw97uoFh/Ik5c/kIAEduKXX8N
HR5/GNKXlAzWkh8zkLi0m2zgH46K34Rgj6jcb1ee1GGhKnPLH2jHp6zfGopD/L+f
LrUof5rWmZXNCOQOaCQog99RgS3yZy/Wv6q4Yf87tpz4XE2GgTzSLMFqYXrOMGtk
U2L5OJU07ZfsMU/Z69WLWVFdklGQzS5zQ+vKdTesGzDo9DH1xDXmLzmJ0UAGrRJe
niFfocmW+sEMAj6pWB9+F6tGF2EjH0hGu8DN8wbpbr9OYmDiVRSFaka3joIxohHf
kLmaLhJ+v8Maq851LDWny74awypwuHMvREQJGAdpht7Qhe8AxbZviwbQ5u/Aisra
fPPWg8ILGqrAeq88cfck73AKl/QOWgTWxFLYBkzP0sIJ+UgxorU+FvnIaWD77Owo
MjbAmVgZ3R/d+7tIDLvTN49dx1wMCPPU/J6tzmUqZ6dnFT6bPWOP4+2NjQI2Dh9Z
GAjtZ1nzltazHwmy40sW5bvRU3l8O2BhoCnI8cEL3FdN21tWFujdVyLL+NpYV9c8
mezjg6tKgHTo3ubA4TX7ZxroZvtLBQuU3PtmfMqgiKGoov0sbPdKc7ZlsVT9+K+q
s4R6IyOOYifXvfdBllA9RX2w9u6oTzXQiOI+LemQUvxsKC/XZq0C77jMNFElm+Z3
JEC8lUH65N8bDnioq6HR4N25F8f04mtNGFPYtG2PgUxjOwnre+rTd3tKyhEbTYOf
uMEF0Rbm0pDtz1yzuqKMtDu2VoJ54BhLvNbGDftwpL8ipLEuvtq3t8gSKADfGJtH
ebEJnysqUscNBZ5xL5qwnPs+FfngSuGR43Suew46s0K/4IiZQeUYYNuJ3YLyElXE
6PxbRIq/GMW7DlrusJV6pX+SLua5pkqWxNnyhgk25Py2K3y+Dc2daUTjvMZRup6p
4NXZswUrzvGoyRxmi+NFGVon6EhKAlAFzMiMnLHO46eWGXovyPCJ55IIsj9mACZO
dBoyS72MdeOxNic8F0ohF4WruivkXXx8dIjHLBHybaGnZ09lHuImCx1s75RQVD86
h9g4lAhz54BF7HsBXS5yT+JskCgWuchuc1kXeo1iFj+ICyIDw9gCgwKo+ToR/kZX
JJsj6ZoaDpgrvYAJSEmdu6HusFDZ0BIKVGjAWl9V39TIfJ8twx6zGB0qsbsN7MIm
kMm1w1ac9W6f9OXS2xEq9dwU7G5cgKB5WPTvG2p9VIHgEH7DefiJVHpNLB+B742a
KjQLc4dfs5Uo3xkehn1WAImZfaUkiZzoT6Z3kUMKbrx6dQ93j6lPXUWHoOn7h9/6
V9yP0gvyJ4a5DAJIgQeDEdwRtWAqOi/UC/+No79xewJExPfNhsRDB4pqELDF7Xoa
Dgm+INepAJiYhO1WKHL05Ws7fJKC/tvBYRkKzI1Mq0MucSriQfoMP+q7imwDwxoe
PshNFUJiu4p4qjedno1Rbd5c5ldDK3OUkx4eNA/wR7kFOadqDiRnKJ/WEkAlOspN
NR+stxEKa+SdiQ+AAHCScLbvmQQPI688QxoJUTkOPa9hU8TME4XrpJBFJmpZkmhX
J90+j8kKucl2KZubSC0/e9kUMsa8zwdQm5xYMrXOepN9A+Q2OkIVinKTpCOoc+Na
XbX1yVGOW38v+67gphripfGan9mlPcc21GG9qajgv2Ne+TmzIDI4pVIEVemYBegS
fMbMpHXGgVofMEbKobvVkAGu9Tmjs9+SfWfDqQgwn4srRz3i/lqjsNnH7N3lRoB2
C3KwBiFxXE3Llq3acbXxkex7hpLGLTbV5PujDbWQ1SJ5dktObPTRex1JDclL0zs1
xjmBHkUK1scRpAk730S5qENXWxBKY67TVgdi344pliI+34pTPdHslQ4v/RzJg9DE
HPJMM3UbbyqPRpSyGqXf0HNyFfCz9BPfCH66Eu1LGRv+qELXDRpfWR0Dm54UIwNJ
BcNwkpx/nUh4qPMe2A8pFRT/0fXcMRhf+aLJEttz7xSqULvZ1C+sG1FDWT6dkGH/
vIb3w/fRuJXtb0CJlpUAW0iy52OED13H+9abLp7Ffy7/vdYyqAUZpT394RTscYm8
QJ3Nj2nDoqkwSI/hMkQBXKEAD8HwnFoKObn9uxqCFCDspxqexyvC/LKNzYSKWmMe
gN4rM4/RZe3/q/AMHsQ/u/rXdgN69lB/8GdoMjRxSfL2lM+SJTqqQvx/jZEFmEG6
HgjjqyJZW4h9fQgALrkkGhX3PiriFHkNgDCY/K4DlMIBwEeKmaEE4HQLuA5NzSNU
6nr1YggS6KVlK6pN9WLxd8c05PSE6/DY/ALYo3stj48ITMD54N0Yp7W9lKHXeCaW
E1LiM+CdCKnEl+vxrxjMUCDmqJwwKfCw8MTvOMY8+QUcNEeTGDK+w/Lf6eGSUw3X
KNIeYl5le/rj4PNqquyfTDZ/7E1rPXu+6vDtrjss0n5UUnaEDG35RYTenuG/ihzD
Q7GHeorHUlV0VnsNFpC3M3rORNRxaq2KGUsbb9G0f7zULasIbruycOyB0VQWf44/
NZ0bbaH78sxjNspm23R683JTKprEZWWuSIj3kFEp+k91sDQNweD+zt/EyZyNWaaF
lAgzLnBD0Qwii3g6wroCQsQQycyXSCvsoXEWQcx3snWEmju6HiUC3BJdVD4rLwdb
Ut+NhCdg6a8eYxfzeO5ZT8F64yyzW/lS7bKxtint2+GZUeyIarxCsCe+3PfLtxyq
tsfUsYa9B5M7F0JnZYvL/8Kmr1xbb9qmBH9TQ2wouVWfvnjvae/GOKCby0Dmegtg
YWAm7H/3yrnc+rwBJdWmRw1fofbOeMBAhFAviDX0GHb91YUtIaZnEYEqgM1QeAOj
7/0k0NDcF96lgM5eU9XF9wU6EAoywomBHu20Pbq3VWc6LLWp2hLsDOuzF4565BDB
Z/skSP98VMUo9eeRgdDzk28dl3Sa1qgplgnH7Cz7L9hIyLSz8ks1Zkn50SzbrQZT
UNLOHiohEDnHDfU3CUNy6jfb1+zlTMhHchzWQUSOMXVG/tjRscIpCBSE7rkJs28Q
SwYPAiUWg9igUvTsWfv67v5JvHgePmAAchaRpyGK07b2bZqXTtZ2X8KqUAlTJIBe
YZS9iocT8ve99PK2OKFjLmNXIuqvwsGMfyO2+oZfzEFbo/BveEy7DgcXOReu2y1I
S71gxH0gaA4ZS0EtdJtlME0UvjwPr+V8zfWK1bt3ZpCBOhpzTYvP6JZOr95NUV5k
jJ/DRbd9drsGYd6rlK2pLW20r2ZnoGNC0uawgDQ7DXwbPvkClJaqEZoCNZ6zCOUM
Ab0iESUXLj1oShGFvRWmLEwpZ1wsF2xpZydswZywO+PGYSyY4aJXHcOnGt7OKDSu
gEiEVzBSJl5mkA8a4eVSfcBK8VAfRJezwkgaX4q8LKqZP9TFcAph6bt7rL9ioSPZ
Ij3mPCcnlQiS+eHKQ5lNcqao4NWvfB3CGmWpWU4B+JbCY/UG19MsUM2eswFar5XG
yEsh0P9pUtNIBwyck/8NDAuD5+fMci1mXrkk0TsH8AHNLWS18Fs4gV38U4RFGWhU
5DfjJVmbEk47b2MuyvI5xf5RBwAnq9cBF3ICWDaFaCnHNIc77Y0/fvccueC7Sl9t
tNuRc8g+rwAaL67ZiqXYVVhmhrKc27ra4pSB5ibFrgXYZE1So24K4tiW15yxfCFI
GK1JeHoDNpJ+z+N+GB9J2K/FbhGrE4yDeRfHkqWlMQbNhT3ZILI7RHONVwwlRN00
Z7botdb/1+6Xtw75uJGHMwqzDF9GxpL3ptg9x7s8PBJRyi77NuGioR1XaenHh/5c
zkA9huNqF13GnM3/LzvR9eSk8EVGTLMJAYhActQ/tcsdyX6ytIrLrh2JWU4wkyAB
p7UuNErhGtDUKCem8o08Eqbf2X1mieHilNMu1SJ8uzIH4YuSdHE1ITXQMDXtXyzR
8YzEqTrky/Zj4FR7GnfrpF1nZqbjGaLp2WoPXyqrlwjv3G1e1Yrcte88nA9my+up
YxMW92EoRgmJRFoRtZAwZgXv0/+JwwXs8L3BH88FGnb739zmkDZTBPUB6VohKpG6
DOwBNK1FFL68iOsFqE/T5p8oBVdJbsOdUxZ1fiKKO4TzM5aHw4r4qDBD2IC40rDs
3w9ogMCAM4njVp6Fom+7xXKIiItBGRNDsbVt09cOMSafrlpNqSdUPamOBgIhGqa5
c3Yk8UkZp+3qw8x1KB5idO9a2Wb5cyggh3qDzM56OJFORIdlnlDsa5dw3etUT5Jq
N+qVjkvYs+wKONSucfwCBopaoMYfcHZdJt1Ne22KZIH8uB3nqUAhImZCIufpYwtI
D+v01Vlo+5WDRimiFwH7g+m0u8onXfZdbQin/13pUhIL1cR6RKYP8vv+Hm3ELtel
lvX4sDeYM4Hqa5icTmTMCdGT8WAOQvN/kx22PtYMEF9mHmz5kUCWSVoZlWaYPxvg
TW1ooQeeaqnB9og4FNGQzCCFyk3mje4bgdei7Y+rp9w0oJVaXq5yYD5QjDOhvJ85
oO4W2ufvPEBPa3x/RUXRWy/Cv0qzK7C8zmSgkZ0qsE99rW2JvR4jjy1SDtdP+/6M
f/xQgzSUY90Uz2z2CmTwk/xbmGPh6RMmE+947cQD8P11hqKDOsSfZPbMUUcM4PEq
Ds0La7WDdAKfmog+WajDLCL15RKk0IcPUVaRavhBLASLD1OMI29MXd62t6Cp5LtZ
b/nx68GGDvhiDiRr5G6oh51VKGzYswHA1UPBHtIZnYao+I1cYjzgEEdCkDFpDwAJ
Z7IX/nEBki4c/olWMpCpeqH5lMAyo9ha3rr62nbxPuboeYH/BJQJWAqlVuWIoecI
7dIXNg5AzFJEt+QGDk9lQy6b9BfV+5oJqtrsbDqe4ZDKf0fU2zwcWOqtrQRBR1UM
QCfEd6BzlTPsuCRF3Kgyz7qDUT1d0g+3lVxuKCxyvylUZ6FonHM3f+bRzQwnVkTt
GyVc87XkOp7qJFdfVlM5spGD5A851rNFZsxcgcPWuyX16zWvyQ2/mmCLjyRIUN+N
BKGYSF22c9nJ58pnyaEnxJh5Z02shwH7QVgNpvUpNhbTGQB3256oP2MRfarbfFIb
Wz5v+EGJ5sZjMlz/uoxxRYyCg4In65+nLBr7QKgY8gJWX7YQWbQvkHLP7AVmArqT
YFzA+wDkMkc8wAxvvp8VRH5A8iOK675oSOQqWZKDhRXFXBzrAxoylKN5YNHxx7XX
3yC93VJ56br/4Of6Ey2A359+rWle9PoC1A6kjLVdQyXkoNd8VyOIQrHHfOh83K09
PkQlAcigm81cXM6HTUV9NV2w88vqvnJlcw5IGe0BlX6fWzr9aiL+qOf0nojX6N6j
Ei+RKkI32Q+Q6EJpbng0bFL+2hl3x2Auk0JfXKJdCzISvjaKmO84un9NJUUjd5ev
/JKqjSYCDij4LSNM2LymKXrlOPdzw8TkOPPM2flcTVEMzk0FKk4mMjJayJMfhzfU
CTREyGuUQRjkRZy4EqKzXVREmxdq1NHEJqw6CTVRG5XXmfNED3bAfshnHw+WuXpD
l1ira2jkBV9HCoNC29AQltRSplYwnIOhev8by0mz0QuCFXd2Z4La669SdahfPczE
2z3SErSoJS7ru7Q0+Gr+GF1aPYmiEnRVRN2qcPbmU1sA8CsqawKFNwjQzbVYI9kg
qdxw9g+tzSjhys67vWJo8IhRLJ0/kln/U/nK0g4oCHCC+zOZxWIoq2dGEqh0T4Y0
vYIXzHnHLQQiCpIm7D1SN1/LfgdPOoQeYNc3F4AzQaiQ/wMcuh2aTJtCkrroY5ic
zDMcN7LAIDSU1J1yuSLm0M6mlNnjISFsLSz+gBaJzY6BdTPPgyaAT/Rpu9qfjfCZ
XHdBlLLPcfe/ICf9V8og1ySwNtAdy7X37Ays4Sck/tg7hRfT5tiV6L+k5ZTvxeVT
i7vqeWsbDW/X3Ty3uyDI4Wgr/2j6ueOfSYlrp8ouxrwHycBG3JJ5Mj3p3b+bQ0hY
Ki+tTpe/ssW6jtSkReB51zrLCloV0fFsFEOoUsOXyvvHIZnqOQp5rUz0VmW055jK
wgMTvp/OaFIhaA4ogywSyWUTos71Q8zO5ZBhf0+0gGWIBLjd0fV4b92vcsMqWxwx
L2JiGWimqlwtHTe1YnCyDQfNx8hkgtTGoMNF1kaY+brpO5D6lGHVXljwLjrc9ZF+
u9u8lfHSSj+KSmLnuGf9lHeKXGV6FQniJdp9GkxTU8SG31LPS3gwuBMIbiLos7Of
VbcpNuWNSVFVKbb/8lJ1MZnFifcKVrhgFZ6LStCJfnOMmP7JTHI8rli93czeo3Bl
dT/sbieLgWjMi/ZzxOm5rWMgwepK3RqtWGE9yHU6Mx0hzVd0ocTZGQBqypemAAF2
2tQCgQsBnPk9aVw8hqaqDh9g77nQ6bIAE/6g6mTM43QxPtlYFYjROHHaxL5sg2RU
T76FkpbSkreVRR+qrCXOi4K6FOWKmoI2hBu0XYATGJJ/exMj6BMbyS8fqlK0sdCh
l1pLFuCSk7WKHzDgdlYaBrdH3pMSZ4Vi91wDocur4EFtjVOZGLv5+Z83fVBae8s0
QVXSazZGiiHc/1NogtsrlQ9PU39Uf0yd9Wg3nqv4EFLG/Uf9n0S91vzdmsGjct2t
U3xMf6EtA89c+cenA9QtfNhWBITLH0+0jT5lDDntQZG9qjn9t5p7Gc9QX56lObNZ
a4aezVdq/mp8QCvxINN2uPgUS7BXGmGFp1F0uA3o2XLqZuwOq4LSvirkasme9788
i2ZChtSYkL05KnAjPK+p96TD7E9l4jPfYa27tzDGK+/D2VCL0teuifO2R8LggqwP
yuSp4N07eJOmCjwKxVqfLaawDy94PcAXT5ZmXbCV/aPgMDJ4Jblk3L3JoGsHXqvz
v+SgyH6AX9WT/at4VGrmZ8/rPMPeWThlykSmoNV4hMVGZWQOiYjbgxvxipEFc9Gz
tWJnqwz6qFBLHH/r0Z+YtwXP7ZhJ8LZXWG3JNw8KPPVXCK//+EEibwudVF+G9PAf
v1URU7HaRbJ8Pt99EnFyAnaBvbl9lCIICMYkAl+Gh54i6ZmVJu7WZdlHp2P+sXCw
fUEy7ME3jupq9C6ZMkTUbYzdetpybbfBeRSG3qSCEbezqNMzPQMXzHfjd4JTaRmA
jgKnEpU/SPzRKIufVqG1MWvZAU4tIqgQOV9jDgl9M6ydRrc03arlLK0Jp25BfGCH
ubX4vdKjS+/ZDG4mHSG8pZRSmrbiQn1BQ88Ilumu8SQkTcS83utUsyo6rp4d+oR5
j+k3ROlfxNzlzvsyvl8z9KHM6NFcU3lvmpdolVcqNj72T0jYWUX/7LBd+Vm6EiQL
Saa7TTg0ooZ44ptEe1G6zc6L7NzgxAgrYsbS23EmIvZezgN2mYRkXhG9cUvrcDbG
AMXrHQWiFaNc/eGcAsEWEOS7NdhU4pvJdSoIgZnnUuNcr993aUk6N2oNpKMzbWlB
FI/MAz5Af5TI7JTlQxibk3rECIJ6Jj21wvrW1M/cCB9IByGM4Zpq7+vAOptF4886
4IwRSHyQ0+bbItAHJXIzPr1L/zVYk/ojDcijwGutfQ0NcwM2GcfssM8U1sORxKdc
GwJxH75v4l0QecyWUqfQ8PTy+ayh7NRIRPIMUoiXnwXl0mF3OFV82pm9NX1vjzgs
0ZwOqVJ81DWpeQFqz1V+y8ILeFV1Y6/mYNLEEWJj1zvXMTnmNDNzQ5T7jURs58pJ
435YsfUdRoBq4nbh/Sv/mrRwx0A5sKm0w6r+R/usxoac5OMsDj7zs9Xz9egWWhf1
a2/GlUlBrKdVbpVkBwEm8t6aIZAH0lIywMKCRuxjaILVAptXixAlR4J2zDbg6V0z
UtUsF7lq9ISyKmGmJkdFpV/bs6ob3xU0nKDzRV15Uk9ZfbJ4xSsOeyQWz7CVyKlq
l+yAXAOsSFrhZXsy/QK39cxhk2E6SXXzLNm12tvX0icW3WYN9pWrsFCEjYcLk/xF
sKrtyBfT59seojbk33hHJgL3/VRlm54XuPKt5kfB9vu4KohCLT7BjsZnzdtnD6cA
PvmIeULc30Yp8CUAyBpgDDAtZGrpWsQb57hohMwDEvFHutVnO+E4l0nHhTZnnATW
xqr8hyGgLb4nnHGMeaEPBCvHwNeqKlvns6UKNCpSsq0yWP06ln61JRIL5rVTbKqV
+E0Yw4hTi0xfHZtwDdqcE8dJq64l9Epm9zfbNOEVApTn9RVx10Egq/bqNwwXZNgX
ayBO6hKO8UCL7YctccXXmzqPJ++JuF27szQaols/np3Mgn7U/cpAxvZMyzSlgNB1
6etY1Fu1aR4EIrufFiMcgdOlW61VwJPmCHWlLOmOnnkx1R1R18AdT3U+j2m+8yyC
SdWqovG4+lgV+xFRqyoy1nuyA7vxf/q2vS1Mt+mcCZq+DT69JLdOUNwJhJ4KuqMW
kvROtrvYzF+GYVvhLzsATgVbbV9ZyOD+oyN+FhpnT1t5T/Vf0PgPeuMmBzL0YvTw
IWorwr7mOvb7w22xdJtNva1qm28BMMn4fRKmCTVXRs16eF6RktTRPtQg3ApMJGGf
fmmr1FuWf9DfaZEtIA0jLY7zOcZK33gUtSNuxaMcDc9wk3ffmIbB+G+kFt6SQxqm
AIALWF70s1Ke/SnPXMhFzCZvmEtqaVR/MN3rqvgs9Bikwjb+W8ueXeAZSDyExvP7
cOQr3bAiIX5YE3a3bQ2+VtDVZIDcMm/SvrJUrJqOGBgLaOO37Xza62yuKfYQfn9L
mWpvTT1XYGIc6mUolO+rphk0Y1NE+9pFuwtVieU6TkRsdCulkiTghpvVkRarTFTF
/ifbR0+SRkfcT9iMqlSyZ5ykudb+scWZsLOz1akt5PYtGQ6Pokxjwl7j0efsKae3
7Rqn0DYZ6fE+t7SUIjKWXwWpbEXfwAPqNk+ix+od3/Ix1ULIwEF0ZealkN556Guo
kbEWUOanBsDDZzDR1YS21xKT1/ULl/rTa6nb6Ohe9WLZGofs1ITt9lHrWOT9iWft
tP/mNjvyJ6Pt/stDbKcmYa/HHnlxsn5ElBQ4+Y5PEWGEqpr6WE/p8ZYuMp56EB9X
ddHwG7BBfdcXGq7PdPccxjgHuxETSP5txboIrN1UV9euShOkYPNhXarZB9oIEwl/
BDB+aYNYnaH9FzauFeNf1sPtiDmhpTblT3ROomgLAx2Zi7zxgYaOmBjegJrwdASB
xM2cnTgU11KQSUz1IRDywaYf2JxK0pqDyndjJ51/woMIqKG42yZlJ04FxGuwsk7T
vZOIa58UC+AcaJCPAWSkijhIBWZkpIbTifksYuMfPMnMNAK7HIFDoQ+SArEbdUpE
aYs7vzygAY1GpmuhLFhxigZxmSldTXbXfKziGNdipoJN2grPEAR56dX9bdFoqYC0
QxIwzmiK2PJ0rHAd4fpNUFLOYDcI7EQ+vCe1PXpxEZJDgFxpB+FNOSjAzRXyt8kD
Y9jH9aq6V4PxRE6NgF/pGhrrn66GngRfU/UrPbkKsNhCQaqtu2fNsCC6GVzyj3Yy
C2gVfkth691nX2LhwTlZAe9hi/VJKNl5tqhjljeq/uS8HjxcxqflVPrPnkEE7qQo
D8A5d7Id5vACM6XN+Jx/MmqNzD8CzRz/hA8yiARqWUD5l8Ix3EWgoXgpjIqtX1e5
yqBTVRO4jQvgOhyjLwAAu/WQ+Yv+qVcsTB6sNggf6+FFwyclPlCtkAn6Dyfa6s1I
J0X5/Avxz2LXM2JZrR21UViEAGUKoCEpVWyEXciODqqoeEfWMsWwQ0dOzx+0WOJc
zf8IG/rWrgT2K8lonEJiFbD55UqFoJv2eZpEo833+qIuEIpAVZltuHRUNvOdosP3
Ziw5Pusbi4/K2rrDZydHlLJ/o7UdszifVMdeTc2vS575i70aDGp4CbR1By0RQLt2
/k3oJM1sQVGr3BFLoBxdLitWIvLsdob7lvcobGRK6cBGkCw60q7xpoJ2ClFF+PkY
x7z7xvzr3lTeZU1k1ibE6hYgKY/9X3jf7nxmuukBsBtdVwfW3LOnONiGRiMPgjZM
hWTLtxjbBBk1yzHZJIapuaIrI2ZvkVpd48UfvMb5kf8hpQDdaEStlEmwabf+Nqyk
YvkFNbjIwwCrY0R+1JMLVFd5b/yn8pafEA0UsAsnWZhAmD12KYpxcnZFvzZskd+D
+4FD4It2bbgqH2K1bzJZ+duVkIrXnmp6i69qa/tzTMW3fOnNzTLZgnlxNnQ5P2Cj
zyXYCVJH4bFSYQFrlNAt+a825hTw9/OMdjUiEkMLPiH7ZrM+VgSajRRE6X3yPeh4
PImMSzBxyCjADnPQv8cFWd1jnSLLOZ/UHOO4V9no9ukoyqm7LhG9nCSufPzZdpYr
TSFhz+B/Ujm45dF+KYrFPof5ntmEvmUw2DFAYeR2GVIb7dT/AJuQKKFrxarcqXAT
t1Cdby+lo30ie9ZFKWBLW+65eBudy8mE3RmR7nbKwo7zJqE23eCQauZI9lOd7hKy
GJeDbwPDiDielv/v6On9DaFmvyU6E9SjiRCGwXRC4xjMWZ4Y03pMyjjYPzvf+hAH
Oo9/e1GJ2wdidh9Broauy8ZzXEhVgW+GsOzjRO/JKInXrnZoBin5BI4b2dtKQTtw
LtHZhtwTX5MmuwkkmqNEkdjeFY9KNMEv4dds36ebWXbYuBvafnQftiRZwbNOsBbB
FbBDcDBVkBGhLKXcZpV2/YnieZ2q/crwt1LGGrY2NOT9E35nvKHtru9aWPRUNv5b
jwLnEEhbgGuAhSm8mo5JFgRfqnJtCyVakSxJnbX8O0Pp02o4VGw/AO8GoyHSAE2/
9ITtVRizquHnf4oie8/XJH+Ev6GkCuy/xILIRTY+qYeoDLUIx1zNwzuj2NIobZ+y
+Ex3gWQC3K4e/eQU9tCZrih9mRI5z7UpWtgWlenGvpn072njNqqTFLPR8mjPoYfV
vcrjFgN3R06o7+/xs3gcTXVEH7TpOaOQiGAa9dvSXYuTjbaLjofnixh+iWNPE4GN
x7s/eKmGaVuwOScBt6JIIVLrDV7efSeBeKAhg1d7rF7EY/vul7vuP8EHLKunQAVb
cTTvFFar/ZlqalEmU0BUUi1mfuEvdgf40sNkU69OAnJ3xt9UvBveTWZZ90ApAXcl
AXWYxO5pbHVyJkwlixX1dgR44Hc32GRg+BoF0NKRP/Xtoeff9Ygi7K/EjRZcghLM
xLL/raViKah901FmkQxVFcEV6YOh/oPNJ/Xwlv40B745+eNsjgm98zqiO1TYUVmg
0GXTeijCEevdOwWP/el+6zTMGF7NmlwnEZSyMkJW9j9eoeZW7cVBuKM0LrTJW0Yl
eNFNLG3duXuBC0rIXMDpXLzPly7FAUI/JByQPU+qbiJO4mptSbVdStDWNxEe3QYm
IRyAzaPDR7kNb6KX0EJCN7iiWMQBD5bDSzdHdZe/PPg69dNu56QN820qHyx/tNP2
siqPCQS9XQdbqIFSrLLvaC1LPOAOF3m1Jdvrql2Vpkc6xzNy/gkMT2IAGbPd5XqO
+YAyjf5SuNF8es0zdv5oYNxXj1ANpH75++QMnEmhjrq8bIR8CpUnZlSjcTr6NJu3
k/IVTrPf+E93TA61kcF4QRQIGt45z5364bfOlKI5cTjpyugQnxmDasr99kk6rlAA
R/w908i4YuFh8+7Feid03YDouuIhtDvju3uIlKI/rPRJbKN7mKUWgwThC6Mm9q+X
JBo6r3z5TG5c+fn2+oYgwv7nXpbATsb3fbwI2/Ccb3FrH63EhxPJ0kx3aPZJok/j
DmdhEGEs/rZKbF6a1PHh3uzKacFPOkhwaSIqDwuZFDNUnt7LIbVIB6rHnMjbXjeG
BgSRNin+Y+c8IpCkC4YITaNdVAZVyXqVdmWUxL3xfjbjIxZ5MIE9o9YY0fenM8AC
YNkde0R+lGso5XpQ8wl77z5yKMAVPy+uH/xd7If4DzMOGlEPOzmpNq4N0U+PRHhD
wC0Eo2zM51Q0N0EPyYagBMzR+Ede40GMcUVkMldy8YkNUoW+qhsnTvcL7kpBD/+R
E+YKCYYvJ/k8PPbe4pDQ1WRUPjNZHUjfEPS+WmQiwsijlj9aO2GujZ1eYGAl9E+h
w7mhf27JmP0VqkyEURnMV7JvIbiCtX7oXfNIyc+2mH6fyAOXeGx4KATEyDcqR/hg
sYFE0r/fS1tPzUv+3UwhlZ13+ixXZ55hw8p7m5ynLSZd8p1qAmXRCUEUnPlfZ1oB
AcTlBBAzVJFkvIJtZTd351TchunJRnFCZjcrph3lFAxiElbFY2jSonATv4gf5chY
eXyuMPgcuYwHbiRszIktzdtTv8vwN91pRIsjZfU40kNWeVJtA/gwyr38eYugYnDo
JhizI+UCN+qJ4t8iesUGuRbVxSjGe4olZTGXeD0jc3lTf1tX8bvGvlTOLJMoVDkh
W0F/ICLKmoDglTw2chnW53JrtZRGOPaEczIgzag6jEkEhhvoc2bCQjS+5gwrlW0A
cKfOrSV9bjTIpcBvMG3Xjrc/g2xSYR8mAfInNDD5UugvqcWltCszvCbGyE3WZFvw
9Moay82NnzFPkReHTNzEfbg1/lmfqP8qaks5eMHJbnAAmSQqIDxbttP3roMDw3YO
3mhKRR3UqZk+1MQOLJNDJIHYVYdWL5d11vIIXqC6O3l+HwwnSiAIPDTSKHGB81oc
Ftgy6oIwzvU1iIUh4w0KQ6D2On07J4baEpptNhBRBmxkpMh3pQcXsRZRM1Jc2cFN
7nkBVJLy/+PyHZzJAEYgnQTj3tR6ztnEdTh8a2+d584TjoanSr08J+QkTfE6lODe
7g45rSXD7O7G9ujRLZW3BuuR3rSZ+bGmdGuHWAWzd2BobuLgF8H+dKL3Cl7Yov32
HDU5YLGHsf+EoM/4hNdceh1FbJtGxyjfj5gnF3Zvj9MKQUN+Ym8rRDmD4JOBc3dO
9zJX/OXhgXmZv+JJacECRGgiFYKpyHqHSAZdboDOHfhqGLTsXEvWE2TB06z9VgQ4
BCXQyLxlhIcU0mDMb8Bl8xIWvEX0KQOGjDAyS9Pygy8XIBWs7bTW8rJhvsOdyLOh
iwJRmmqtyes+8ZHMCD/TVdENXII9v+ZRMbWUAagorCUi3x4PsWGZ+U6VYrTN3Oo8
y85mvaNShyu5agPAO8/RIMwl98BFfLqJiD0dZvGyDwjRoSQWtS6mSjpaF1wDf+6p
s8uKwtwNOlHFTnLtszw0NdRxAZxh0Wdes2MCpNWgcE8F3+kOTDVioM89hzhuuTzg
IMjxc3z51SmJb7y53/j7xwPOnt2ScBrA2q8dlx4QyrezRa6GX1nAKJm5ezhpOvM0
QvCI9yLHtIV8evP6xubTHq9pzbSkjZQ+87IItA2/MJbxqftFQf4bHaYTvRTIIRI6
B6Fwwt3EdWk0GzEarn6fOUMAKxLJAk91bAAbLUQO2s5+Mx+RtSjQcZcK1WbXw1iP
cg7dPP08iLS7IKcfgm6JfUebR08eC70+eKagpMeJV31mKJ5EeK9HRPlIPKuOSHGn
wk5jBA5PnIbkIiGmLFWLSLB130cXSFjMcv6o3JvstxNNcp3MCSNFGht4CZ4/ltyQ
x76lzIZJV5H0OVNV3SoVOsZiPvMof4s1JjqSwenOkVPXp8YwrdFk+MPKU6CUm9Pw
996XuHT69akROE64nmdMi40/qMBXmq6FwgQpi3BR8m9yvQUGjEmCngpxNHcQX1hl
u3XVETXO637GFpjs9gbmYxZK03G2XYoeljKyhsZf+KQVtykfJPgKFDy3qK/SAK0Z
qIrGnZpjGLNvFketP7LDX9vzTaDzEUcXw1Ffj3qS11rEovpHVcAFc1tnlSPaX3H8
k8tWMYhEA7Q+u+uQGVvCKdwBNoC7tNy+tL6nK/ROUdTtJQ1ZGfVCC5NRU/rnyyFo
wOvcczXnblkVwLvTEXlmEt1m4DBzFMbMnk0yvroPbWRjlRBI8L+0X48YG7M6eije
oloLREzaGgXN45FKOodp0OaOlMI/exxIHqNvt6SOYk99HyHcDaNhNeV8MtuIuYnW
8OAh9jBwYY9u6jv7OigYZilIeGCDSYQM8Jtz1iKBxZY5saxHzioUwnoxqBfmjqwP
sySv6sd01M0ji/xIUdmMLwyIuqC6n+aCvKQI3KdQejmrP8/0eX8tC021LVF352M0
8A/VcBOgFLcC0Vlz0iqmDEMS+a0eaUqnnU2Ziq+MzbGggQve1wwvTMdUvukZCvgQ
eVBeFklNV7oeqwckhNTqFS/gCdDwTADQqLo3YuyjXpgnQCgdIvAxO6aRE1MKRc4t
6kNEq92CzCqz8X3yhtVdBCJlummbiMZmGSvEVHHq+cqgRXhFfW0uhtipyHNcur+g
2P8saF3/pOc+edrnhBCzLk97WuMCwS5yK8KXLZUKuleh1MU7P7rhrzburSx55wrU
eBtGiK90kTykFaRYHQtxEkmsCgMp145iS2DZlRso7q8NEewWPNPbDr4SaqQEhAYM
rkzmihMlVtlsTJEvuhWHJNF/CHW00S/9mCTqhWDCeIAld7wzb911FFsTzEoanziG
ZHCIK4YJxK++xImeKLQJtA7gxCmeBZzxME0l94+17DvtPbVvqy0o/SehMHN1uLjw
M+n+FvLFmMlHWebg8bBFtIh7jkDwDhuevjZEByRjWeX14SKN7yh4cJ6DIatGPGCs
c2kga2zl/jVvhV0nSehg6SC4XTCyti0Jar+FsM/EvZgp7Ly7Pb0FrCZZtWYZNF8h
3PERESew2aAIMuqrpcusz/6hoUX2EuWYWtAIoItXry/1YSBi04nGbTgx7U5xzamg
5RS9u1O+Uh/a2Z/+9K43jXbx6YA4Dk5N19VNxbehOlTYF2q2p/Oak4qmg2wn6T6L
LNy6uik5h9fmqrnc+UvLKCdN12sk2Y22k91Dnrk7viMqFWlu4enb1u7e7cYy5O/L
RFysrn3kHXGXyHcDEw0b3JfNer8IBir036uqYN37DyjSWQoeHTiGYE2dqQk4Wcdb
V6Z3T+rD61LNqcfV+pFLxd6RziJx7KyQfA6SA7vpF7hXECYeD2B5wdSIa6WnisZa
sqhJ/f59ziSshyzh41GiIRGyu+Fq9nUlhyt1fkI23pVCL7w71atgoKfcl8AjF66g
bWXAjtm65eUH9ew9SUEG0l/fwEdW7tTpBXs3ToNaE+nZ33s9Dj6zyeCnjYQamAIq
aes5IWZOFF6SFNj1kIPcbCaji77lyz31icoQtpV978GZu1vHksjLSbGlEwJL/rxp
eN9/x+ltofxIWlbACRmM8A3j13Wf8jiy6OIilDcGLPvOBENeX/Q7ok6PV3wBkvIg
eWc1qtfwPrIizojAuA/JWf4UKdQoTVkm1pYGBphzOMKPzq+WqDS6rW+HPgTw5Iss
C09SmQ7V9Zp3ny4rCUSnHPB2a1BzgGXCE4sE15wNIF0Slkz7eq06DcSfASpGvG5B
HjIJ7pTIP591J3uxxj4n+j12PGK6bU/obFhlXl/nM5z6NOHuLlgP1VDwUYYCuUJz
LAtVYG5NDYzmfjNAHKehU8C5o94M96nNldgqRnJoXiI+Ooc5ExLeSFIX+R39IUej
WA9UVmvOwl1c6aeB68bl/+t9gPWw//7avKt+yZk2N6Kj+Rk801atsU+1kl3UhqiE
GZN6qN8okedOlbsdsoBomNVmBqymZLrsV/r0XVAqw6G4Waer4yhbvFqvRS6exTx/
krG1tXhaFSr1KW6ufvxD4LA6WDaWEcBZDEgYvNAa1OAJNMPvjSEkwfvkClIqKSwh
7m0+Og4H+wFzZuAX96M7h7VLEzKze6gkDnBYp3YpOWx2mY6Atg7UIMl0f+dfB/i3
RIRuqATuGDWiTpfyhsYNJpAXc3KcxX04cLi9IjTUnQDbZgGV4h8p7p0homXs1/fN
/r0Jrk7jT3zpTDyFaajJiZVRb/p1qe3wtYUXA92SCV2EdPN3bJllrJSLqK5HKi3v
7Oq7k7bnDu5vNsfKTjoMuIAvy2JQtwOrsZT6SU0rds98jOzLQzjRtHJaidbuZ6o9
ilBIQbfhjGNQC6puHniScs932u1949Uz400y2Rwe7HSSEYlSVZ7Fz2ARvR929pAu
4kMeggGFuj/icHJbKmLSfmdp0BX3hrwt02V4lcrZnDAkm/EZu4zbVzyuCZ5nia2k
5GxY1Ah83M2DGYxAxmDUWLIN/vixJnZOgjZK0YdymODBvfD6pnbQMRJvd9zagh7S
KRPBWFq8eEfxF4X0y5tfAYMkTRLBv+gkxql4liIb0BZHqF9kgrxTd3dVwnSHZYGm
fhn0CgcjIS+3f3ftwO/nsCDBKQxmmAyVX6tF4SCzg1YM0gwE1bNdygpD4SXXnH6H
VE4ISMSj8MhV8R1fQ7Cc63u7legIrpexOmwn/n0eCU2buVLI2vyLk3zcCTGx/hw3
NqzmyDh0dK4EJ7LfqGoRyy/6YQ99IL+nf2U6UPSKRnL+pljLaHbz9VRBNGQpIwHk
dqfTEN8jVqeCDZTRA5PU5w4Mf8dkVzB8bQpP75ZGKfEyAkwVsKNY2rE0bvXw/fXa
bRBkJZMoADHaVM7Y97gN9VM9VJ290wtDrT6wkSEw8MEhR4wM1qzpJQQDqVYh+0jb
2n2inGkkGGFvXROuZv30v6JRD7O3Z4VjGeLWrEHZp8hvIoEIifpcjxYTpAvErxf1
5Pc8bpIkIh+c1CpbrOUEVoa7YEllJkhJoRN1ti6hZ2ytw3tSjlzjAQgCIDuJpqqN
8iz3i096SYyMyd74q0orCUXxsvvaD5j4FqjTcnQiLMo10o2g0zeBUzZ8FD7Y7/6B
S4qzGIYOCKGT9gv2yTq4BViLG7M5501IRcqbe6DB29zCIlAsYnH6kUVGwkOkvoIi
aMcWuoyXB9l72vD0MWmajzSNb9umozol2PcgZG/6XvnS42UVIQ1MabaFgq1Kb7nt
5VyBCANhLUYPsqlsy4+tgfSQifnScUWEMb5hjLmzZXKYhYa/n0fIM8zRRBgA/nBB
jUW/g+JpC8Xq4TCiM5HXpOtk6B5AYyCOmdn3fIjn1dmsUpZ8kDGKj6B1xiuHzhgM
orTV61OZQqDBt3QgFZ3/A40adzlS8uFXvJaYqXD8pQc1glEx3l8hAWu4dpea1vq+
2SXdO8dQGcOsnGrW0gihR6NwbHc+tReKv/HZgflgG8A7q50Y/dtRXwldgcUYDRgN
/4Lhy6iEoDlojPcAztGPenlOzYEDu1i/hZyBp16OoQe59q24kh7eba7lbyqTiqeY
khk7aBJxCh0HRBC6frmPitBPlsAElZ+6fd2Ud6YLm44r/hIR0sEUrxciNzyZBNbU
hap1mtQyXq++8/ktg6466eUxxxIZzLhr91eQuzY2ODW1WsNC9f8y+h4gKCoaurct
W23zy3NGWi/0lm1wf828tzG989IOFp+LSXRZtDVlRtUrB041HwjrwePQ1YJvb7ME
XTsAdH/cV7l2sIx6wQrjT73HXN63gp790hDNHiF1OQbIfZHZajGlLCcYr5+792my
MegAFjWHPrm9oQ8QOdqwy6WRUGFFhXpOr37mRCJhGasAPoZY7O0gnRs7M4IXxObH
Q49UWydVg8/SomqZs+PUPji0fdOTNCsMXVmyblCqSOhUC3uwWybo+AyfNHqk72z4
KOtZZKEvFacYT/YQrJOcenMIDfCXuOWEMdUQRUxQyCZCNQKsVKuqE+WW9TOz3PQw
5f8Yovgraz7T6BenvH9r+3oPLkJCjx2gq7W1lI3Yz+Q2gQMCze3Bu1Sf10R4cvHb
JXnMMYzKTW4RrqfD52VOykR6tEiRhHvKwOp8Wi17vliGHI2K7GKh9+G+TzWrlp/F
bKr8dEsFhTbP2O/c1dwVodVnudxYyqBVkNxVlnSFtrZACJ45sKnkfPkttJ/oycOj
NjQ25Lt+jpkhMzHmIek38orpfiT5Qr64UtgNxgPmXgHULsC4gWO+4fl2x5leSeXO
3Dm8wYejC+FSPBZJd7a+l8LEDYEBXUNT9aazmSkyUcWqyov8+MafFc2aJda6Es3T
a4T5d1EuWHryyyadG9Os0ehUaQWp6MpfSeCXIXes68csfqCIMbcgNceLq92HFLmW
voiwz4dmKqPoHpfTGncQIV9Asnztt7G+uU+6Fi14q5emfKGdP2OiQi9AZ+pGcM76
ZoTaVNYUJ5zZqRizLvUvmSu8HB7D3Wo79S2CEOVhnBNaSRzejr73MayhjJZw1IFC
gZSYXcpUrb0NuJiMZ3IOhMN5Gtad++HJ7m8bunRSPTvQkwj6ZMvvwCpLP3x6oBCx
i/DL9hLVKdhyFvR3Cp3uosSokDm5obmxl5rvrEDoxvJjnD4WzSQUgWQPqJPjt6gw
41UbVFfl4iVv3vo5qIzyKNBdVBvs0v1ajewnzrJyRV5NYm/hX2hrc/Ylj9vnUceU
wTH4uBnz+v0HUNBgrIr0/pr3c30BttJRO6cjiEr6Y5bWzH4v1NCvVh7m/FzeWF1l
EkrCH4uXqhFrGh8Q0ua5O7lexNIHdsr34CPQUWO7jE5ttR+jSqrmd/6D+tY7C95N
hIst1gCw2mD27YB4AJ1548My+42ThRVZgmbzvr0O2rosYYBPfSbwGtrVhFVTcWiE
s/Xomt7sHgzuefEcZdCrvSHGkXqOR1mYtZUg9qwg8+SHQXvw5mPtAh2HvwDBN8pc
b4TjsUAFkMGV414nKsGgA5f3J4Weo9bPBX6C3QwhwwyfHymbmQp0Q7T0lPWSxmUT
CRF6ZEa3qf4Aw3efgYq9KTaFL0MBfeDKXi6CKTLxQYxvGc6dj/UgAaAOQTtP7+g6
8zUV+7DZh2r5+YPFuT/Yd2j1TYmkLmQ54nO5fZep9ZZhafD/q4E1fdEp9m/VZ33P
0SIppHpHyvuVSWJG+1iNFh0WzqL5Pw+iinSMZmRmADPmxfvZswHyxWJ93lE9wu2Z
e1HCl5WINarb0/0/dBxrYYFjiKEJIjj/kZbpyA6CpAAZ6Yg1SfQqmO5+CsGUoAHS
jkN/WkQSUMkBNVTbnMISTXkBn0HrUrhhROxP7wFij7GnF/Vnt0KeU1jh+FspfRk8
q5bH8N3SOWw34u+Q2gF9lVLO2yghqX4CVpINPW0Ax3kUy53x5OohPNBXyHYrOJ5s
08uGWAGwP0Xl1DRy90bo11cZzv1J9xeuwJTw0Ubw5NhawfrXZd7hwM4GSpYd/HVB
3ohuKaThUbqKErZlWvqgpCX1EGFxOHEPfjbSWZadrC9MA/puOWfpGr9s9z4aF7ii
JpZQGGkT7psEe3YhIvK59ACgv039CkBcheQjXYG+LkRbghk0k37lTifTwh7isBiq
slugAKB2hzCOtBTNuEnSdahDZXzDepLwv14fqDH+99IogheOy1be9gnibQakzMzf
cGGZfuam18uK8vIzVTvzARjX+kZwbe663X00yPcwH1pyzq4q5m1WaZuNv0wvl3Mt
jRLIaol4UWqGs45tbcmDdrLlr7a6QUusfEhOza5HSyLZfrS2H/mBxT3trVjKy2TW
4+9aJjNNObIC6YC/MAmGaFHSJVQrcBL6TK+fDNLr/GEoINUmvwc+CGXQcpmq9G15
a4qFUIIXOdlXqs2G883xLkMiLehW3Sn17YZSLljMD1hhM8yCuX7XzZoQiRDC2BND
NIG2IrXqmwc50nV7VNtOCJseIRtebLTrgmxnOJlfuagA7tr+i5mNkEfPJZitsEwR
6Mv4rvcRFUb1XpEZAAefk5Su/DJKq/AcZydSo2YWh1PsdEaODw6qmDbwqIh9NR66
fi6qcQvkNmEQgly/jaooos5ckCBWVW4JGch3HepQ/hNVuLQC7S/Bt4f/blx3duE+
rPV4RFTnKRHowwd/gdH79n/ZNJe83m0CwqOp2KbCB5p0uBfD7rXqSlf8kuhRc7rS
hD+6WXLpnZiyN7ST+hZFYDc/0o+tt7baxd26tLkN5Qa4QS+hX+lrlkMMOUCB2tjn
8HY/AOhTh3zoZCRgJFHNdaKtWn7sSUrwhEBoI6EAmUHYznUTJhMMTz3232q+ohT3
v3G3IoLj5SL9xbFNkiYkfxbJijuFUqJKQmviaH+WSGTUgg83gKbEFZnWAsDSl7B3
LnY5k5k2ioMtqMCZSi/gB0eILpHLVUHQN0f1/tLYLEkwjoNLDODxLC0t02ORP0BI
nvpguHau7Sf5ZUgstcivQAfERGkbH3feGtjIwceeFAGAoCH0i0hTged734bKSd2a
anxmECjpcSLIMHtQKM9mCydheVk9DrZKMCJFna0/6fQccbPPdyxkCsR29NB9quxe
VfGUAixLoex0wU+NbmJ6lFX/kh/ulau0puq3Ivx/el00IHVh0DKq5Y3+w2WjPLgA
cqPMQchIRALWzuKRnmbVbzJSf6+bU5HDG31DXrpH/XR/D64nBXUTRJHupNc5iKvy
C/xy64HcmxFzUV67DE9UQGsYgU7pbskIvb6BjT4ix8AqE/QVWxAfdg2fYne6VeXn
t4yi9ES8QfLElI3Qj/R57V3/fGgbv/D+5WOjL8RigHIismpiyrGvrn+VfCLPl+lo
asNrOoFzrlevOWDtvZvQdhR0vZUCPC8PzobjZEzRBDcZGstTYZse512Fn2dUIuy0
kLv+hYzxfyapYbPM74gWIL8luGb5yvfLU4lA20Q0HjlPV4IwCTAW+7QorsoJx2uM
SexJ1YM7oLNHDkBe/wUX6mqPZdvV49xYaMxc8jvbgus1t6NnzHVrfYbdfQ08OtPR
HxaFMoGzITiHceU93FwJNK871NmBz1Yp6nZogqOLFwMvlkXZkDGRCNgKxuWaHbdr
aBymPOAafERg5y2RN75Zz5PAuGq4geHyBOpdXvS/5Zl6eib6qH45ZCXcAFQpx9mx
qVNrZ1Yjh1RonQyw6jm+SB73P1OuHdOJbtXtghp+qBVH12tmZ86Ez2ZVDa6QGAd9
9QqVdCNocgVOR0ZvOpZiYJ2oOicqyoVthsucRwGqBPxCdPxr9TueWPXqnwX00EjN
1pv6zogyjELzx8YBWIjQNC+4koOYxIKMltyGf+y646I8gS5yGJSLHK6KRwWwp84E
i7fMlyv7lquKMNjE9h/z6jTGARfQq/u6p1ctZVCw92mUPni5dqyEYHCGnLRmBGLb
qhzYZ3peb201jqKW1PyO/U9WKa/Z+0Qkz/oNGW65AtILZi4OfK16Q5E22ToVpiRH
MXb0FYG2B64pxPcqlT1ZZvS2gHgKML0fM347s8sNG2kj7/GQUSG4Hl8L96HxwkBQ
pOrVq9mJr27M68SeyPR/gGJv667ZRdQcI/ZPYqESPU+Dc8Z98Jm4IQXf48DVmZw7
BWQ3L3ljgMvOaUy3iqTn/2AzHFobI2RYKeAr+yTPcXA0+5V+EZV3zEKXFlFybNWT
zg+GSq0y1AKdc4R4eKPgSlRL/iPB48Jj9kZS7cG9v0nqoMo15cuxaQvNRwfpxsbe
OzkUvE61KfcgY81HI+PFDXtORiJ49RkseLhSBwDj3i4m8KBFzGaI4ijKt0iufoyM
9NldNepXpKDrBz97pmJUtm9qypanVV9dWUyyEppbW+Z/uorzycAi0KM799nb23En
Ns3q9g/XWVGPjc+5TDSldFNtw66jUrsSK0CmaVwcoVlWzEYfC6fmDyzJv88fRhWh
+6VnTd6jGpei8+P3IA91JEJ09eAwN0hjHbp9O3xy3xYgvNmKr1IWgmcZ4V4drd/L
WEnAX5WInHoxF+djrqLKOjC3ipYccanUi0mQu9puYZWZY9G6/ejA/iNx6sbxixmA
dOUpQn3IEFYsEddUpBzjqPB5BEbGvtfG1aMwvCFJkIhA+IAGfQfmZn53RzoNKtp/
4qG+r416cvhiwjmX+zlU+ekfJvxIRjyJDWh7q4WVIg3aYtMA2Rqzfut/WFxnfvHH
RaLOZKMdUxTrDu9YpcIEvSxOqOvfuv3VNF0qPLJ9kNo8MNc2wFR6DWtJkxyXTBr4
2iLtDFLRJDVS2aNBs5oclkV0yRFhXh6CzEI10dpjuZD2gbYVCfza+tgA8J6JoEcH
LKal0OEF4laiCb2b/NKRWcUdl4VrQaJHamagOtY6H4pgycA+mpSyEPUzV1c96jL4
sdBjeT7iLtb/RZGQBYHO3nu9SkmdYQcQSDMvaqnM5HTgtErr/VFzY8JV4psihF7k
RpVOy3QVJaLtgC0IgGor/Gqmv7MS7jEyzSYN16to7PaUlHroTR5AnH8TQ28CO5VY
a96CBIAZaRt0KT8opyHXEU5fwXZeDyml4pxD5jWKxQAsHMUYEhvmcutrTugGxFNm
RVy7ktNTfcziMPDVZ/PujedHvQ8zyY6FqfcJeNMq/95/5W5hiwzPyeb/i9pP5UTx
I1YB0Yw54XYHkqqtb59WWr28XZFMX47IM9x7JnH7B5P5JdR+8HdikUMLlLNGrQX4
R/dLScz9kLiOwDKMUuy/EAso4tmiwhIKftXjy42ELy69vqXVmH1xGB8x8zvLoCkx
jpemuuy/q/IqUa5OgofvMtG0D/F9o5y9c25o48GlCdmLZXqkZGpcMmvU7kcP/d0c
WTSmHMtp7A8GMt3bIRyogGJhbBKHXOcRfbIawMws3zQfitc4wdImw2iFYFx3CiWm
fJ2bruuMumcYKc1JL0StKTnofpP5yKBz9dj03rHZha5ssWyEUE3fJ5GEHXrYdDuu
kKg5N1OXnzEqj4hRty8jfczr7fpzs6q9Of2c7BBrJHSq2x+FhS+jD66VOEiCUdfp
H7IP7rMtZ6YXWd0SeeXSqRd8MtmuRO6SiCvsLPFIjN2/6YzYyCalZmkm5pK5Qbeb
Cn2a/LEn8Jmgs2IjbUwTLr2iTQ4erJcSl/IsucnWlBAueR8JF536x9Zje/32Xlre
EE8vysi1io9L8onGbatgwRBrk4qANBIVDKFJvpbl1z47mMCWXbp5ivAI8G10i1ni
5FV9sdU6TE5MCwLmPY7RMv3td3l7YtfIRkYaxiWLbXQVbgdmLiS/mlyhjy7LNKjq
ML6NtNqrOiFCZ7MRPkERMQfh+R4ONg52XMZtYpj79zHaSJ10IapctsEQFCelmPKg
ead80XWtz3RugPx8MdawUEsPMNpZuP9X+S0FGyXnsmhHomm7jEITshkCxK4Pt4TS
S1E3nvr+JTq8/d6DSt61xUhLbEJ7PGnFduKMQksi0KY1DFAfS/BnI3EmNHAu5f4o
uiEFFokYhGptPiZtZ0NJLFQ3oCWq9e3e47bECfhC4OA4TZ3wzhxlCzP+s/PhCQ+5
dyaeJvBmUD0t0Q8JNHVQqq1wCJJ1T99PpF9/WLQhCwyyIzJfKYzWQEqc8DMcxwaW
mnPZUJ50/GhxMUMAyh35LcB7ZFtwQc8qt/ci47GsphP+84DN18ePKtp9arxXZ1PU
vMUdJpLW1YdOdU9NuLbf/G8jEqxgfypaC5JC4OHl3FpTkdXD7MrIt9vYS0Td/ndH
oXUJfSyxhRQQao0Hpp9+25aD5or0ClomgmYqKiDUCdbe5jP/BEBbFonXp9cOPjBx
kis11d9Gb9E0ybA2Af210xkA/hCcBdyn4p/DzWy944nzCsjlJrN/UAoNfhvkF/qi
K+S5JFTsYej68Z+5kvCn8cVo+73qeGxTaqZbuC/EZbDNKb0rdh26Q+TxXswm5VwX
U48Um1mrtT5DVzlPGi+h4G8gvDkcIK3qAqvLbt31IMIsFtjBhM0Cl/tnlKHnOceI
Ky3IlEeDg5SxA2Y4jBYcUh3Wm67avrzhAv43cXlyoblNi7YJuvWDxqYMzQzD9bw1
CDzpuLwhnAZ47bTjh8e9KtL5v/4H07vvzpk/7Veh00ahai675J4nKogycYOf/Qe0
V4gtWp+RINvniijQJUajVcp3FIs7tkZlpfF/V39jg9BZyrDCBZhc1EUtu8HDEf5Y
OEJJpHbcM/mv7VwbgPo+/v/LTcw2SGxCMbBgNk56MdJ4rnhxH4Pc0CAeVzV1ITYH
XHfSmKPiirTfl6payJTK/UTjf69ZPzW0hHqL1lNnXisMs0lkQmEs4v7Ey39DI3T2
R5PciOPzip/XIZKLN/CVrNp/BeHcnKRBy6rz6sptm3PUGIxfN34ORzz9LbhZ0VQr
R0pkZFICP3VEbpAUH5/x6lQ7lsp0lLxXcoKKTXEGmWUXTuL2BDbaluI2dDpHGkiM
s4LJqBGDJbCHG4ykEtMdoePOriTX8vZHWT4OUvdZy5FgATdFuW0NoCNnODbb12BE
`pragma protect end_protected
