// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kuQ26IqhNxPHwCwejUc0lENqHMKO1zeBjT5v/qXCDI1rDPvvXQHld5v2yYWviOfA
qdlJ+K4jGwzlTSnYcPfkbf32qIFE3jdEsJchr59CAAROMqW24KDexNAGCGqXEiQa
gJOR9UGerfq0XfIbwqONjMiRcNe5/caauRWvo7oYkas=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9008)
lQAxTSnsVyxSnWDUWRVYsoKYgMqUuQcGzND/Dklkmc+YnuXGW8PJTpkprSHRTFfc
6NQ5ru5j9We/TimQ5WFh5pJMyM8WB6UZYPRzzWmCOi6D9Vdjhyy/Ir3a1wMMY7Ap
yvMdX1ZtlcyCU3cwgYSC/lW7zkEquwanNwFQFFtCRJJW2P8wNEnghkfc/Pf/PmER
vIPkaFJsmprIezJEYZX6JUTTQBMQmUlnBie8tBxdAMAHP0sbAG/MD/mu4Wh7RWCD
rRHLhKDlitRKNvpJ70CuW2Pid2wOFfmTnknzqVzlTXTeou32waZWa96qrGMfOgA2
dtDSWcv/fk5cpR9goaxm6dRVJQHwWOv8Ey8wavMLsDXM72mxTBG6VcarrDV4sxLz
KQfXusjkEUzr3bmy/YcHxenUQ/+ydsIMmQBJlPs2OwEnL3Pligay2TuKPhxkzmFY
HfU56Bo9fgP8vxtslSzADj7YeEvWXVPZ4lC8xd9YcviKB/IzLFsNSurLTfQofq6Z
Qxj25XOKaAqxo6zY1r+tp/sP/GJ6sBZwoVV5fV6r08EWJxBincD5t+19ZHfmBPGe
hRx6t7mV3GmEyeYDlpNkBsywGZ4qfM+noOg82JT9vLS6EE1CUxebs3UIyF1kgKRD
RAQEoxJB33sCQd30L7nWQ5kX0lvOhcyQvAo/Cqp2i6lc6UtLfXadPJR36rWZ7yNP
u2OPJikZS2t/nEwNKPcuil6wv4wNUri2iS+2Px+3fPQHFzd7dxWSPQpcFzrD/2W9
izM1ddhvCKl1EWyhsZbADh+G/VhfZJC8zYrmno3h+CgazL70hB8rmoFhbSnnFGmd
gkZ7ejB5Iai9/xDvTDKDj4m1vlIMeFAE21By+po8B4KMBY1f3yleKFnQ+FDBJGsZ
ifA0GbULfbxxbEg68kKwKyvKpC/iiixnyuQs1Fx7zpPypoVgWxC2f8OkO6BtDGXb
o59kkqvV910F9t5L6KzrHWe2TLsffwmr5syLfqH5jKrwyr9OjFXVQUYogBTh4fdl
qv8Hpt//iZKFfFTTnk8YDO8oZm79J9Z9D9P/Jy7sAikUjEs+7Lw4Q1PbozwAdSMo
ibaWqtO+VUglWNHCaprtZedDV1J2c6V137/XyWPGOlAJPhCY7I6pgQY0aafQGyi3
kYzudjX3VbRx/1aUZUFiKgazSa5GdxNfDkPltOrQFxyE+WAWYmRfMDyK4B60vq9a
PHdKhPI74p10GggicWScCW8QTYYK/96hHRWL6XTKjLYhR4DqptHksGzmCewBmwxQ
37VS3wyL9PqGfruzfBwIZjYFj98Ktexa5ZHx544Pn9Ajxmcq0rJSH5EAgaDVqS3L
N5W2ZFwq+vcMlso1psAOSSc86Q9YV9Pwifmh3Zm8WoFSq4nBf34NVl/l1e+nK2Ne
MrMOetPa6hJqzUhdeOuElZgAOJlH27effxYnwkPXPp0SSDEjzMroTJTGnYFEPNm2
2VrYbnqhJS7G1Ehm/bCuRTzD6UzeW3gj5U8SvFQav7o7B4imu31Rkur63WPvasCe
xHudd2y633wJtujWZ2SasKwIgWpbBrCPLAdcmjWtYyuannaeSPzsa8M7vl5Y+SPI
yA+rL9QVzXCby+aGx+Jr9buOMk28oSdP2tjtBrAQFsz2+jsVIab2qGBM8c4TuETr
z3sT8VFXiZZYL3zwS0zJW0trxwpOffXsW7XQOEvfDT2uhubqYsd9LdHzuLmM2SUZ
gs1YwfGLwTfjqvp1zr7suN9ayjmvyR0GXaZ6am1gd2Hj3xGHxT5f/QC3SpK0mTpL
nVBzhl7Yupn4aZbLiyMohA18QTerwygQMuwMlPw9y6F38Zhzv9DlycxgdiruuiyC
CDLvfpvTMX4nKUNRv8XSe8TQH6oORdysFqJh8HaqQW2FkYXbFXceF+eDIWtUma6x
G1pKOqJJu4asE9i27sG7i/i+soUXIpQhoWGm+/04xXgU867oiDg1JrHmhQbWAdK+
KHb5S4a/b/mIriWaQW5Yty5E3T4VYcBOqIJtC5wRHWXSYUt5rHtLFPGSqdg0qCQM
txmNk4K3il1QunhifdC/+qxE9UbMg4CGz4YuroubvgsHy57iJnS+W42OIwSVgQnc
k4fohsr6PWwWzCPu5I8Kw39QIcPEOSPhXDgsJaoPax6U7/ncVN3ny1DH5mUG/rkQ
IyiO2E5jTC6QtJsiDU2AzIM22KsDuRBebaLu5pQPzqp4M4sGBZtEFR7Ki8+R9Xti
FUROz44BrM6J6IF8RcyqKsequLSswIKnj8mhogP/qE0ZsUD0LgQtYFWl45kN60T5
7ddRjPPWWZOaQu+79ZXPjU6Z7KzPgyROL4jQTf4eFYL2umtdsqX8Pbf7P/rK0Za2
M66YJwv79uNp5r0c/cTN6wAbl5S3ALOn2iLZqphxLcKK/Rb/vS8FiCLvukbIXmSy
ds9ZWty+GLSVRm03Cjj0/9uAXHgBqPkza2nB+4/g65q/73V8mt2IF1KODWcXicmq
C8iOBi+qj8V+eWi94XvYR12l60rurzPDn+al/k3FIgAgEKVYm2coSFEUEfSwvr1l
JQoA5d5hN7qggenUUZ4KmPn26qaCgSYBLJVdoqoAS0iEOrwf3vAFUfGTayZIa5Qn
tzwJF27LXUyJFLLD6TVFM8vlzigskKWxcZZH5Pe014Vl2srU5GzK0AydvG73YVlP
0pOe13ZMyuCj9NIuypoheemd+HbxqKR6sJHB5+mpGJGf7fjTCfF78WKfEP9qhSvp
+8lRDzBsnZ5RSmG4AdWpyaC6gWoAT1kA5Wxx9BeTBblgvuVlKhGBq+fsSjoAf96Z
dJvLtKsMuN2o2yH9ZsIc6adEwfRSJ1SH/+cO/JHTxK6Otyjoax0UqL/De0brwAB8
kKrK1MkY1j8xK/+8JswX5Iaep4yR4H1iyzsyVgmgQu94pcq+cew+koeDpitMO0/0
c7gUkklOJR5AxkGQbKijLXXq1P87Aqtl7klEVTGuRo4QxSe9a7KIUZCJG/xuSXH5
8bqdzf2lZOyEHO0rWJ0rXmfNcHi2eJR2qA666NmlsmNFS6dUxUonNoGQ7VYur1dY
lz72mX0Yu13H2LX4FiJsJIZgxuniRTlr88viTbpyHxPLJpZZm39vHP4EC1GW1x93
uGM18rZSDdZ6IMIykjBTtUqgEDYhEW0n8zxXyjLIqewsCNUjUGJuMrUvjgaQlR0N
AVcUkWJ21dZg1/IuHLOjRk1Q2xEtzR818BlHGlw+6+HOYU7TvhVRg98QKQVVFu5Z
D4OQvR36LeT/keG5ILCxtHzCvL8XDKjreflt5hnS9RPKeQJB0wQz0stqRd/QyvOr
zc1Q7CblU0/o+D0Joq44MIZ1U8OeR8oLgBKHoXTODisCOJbFKHPgD7kFOq5+X5Jz
aEc9NRjESBKjhAspPleDxz8BiQ401SPrVwAG7mtxaihISHcY3+5GqyvazHMLXwpj
5es/XQ8MIBVCJlFxU++20+fKeBv3+jwf9KcS34UjFzP4/+DhrPnoiyn38J5HOoxN
PSiu8yfTJ3tDGE/0KWr3sy2e4fv6FDx4JOLEYySxWqETxd65hucrDLzdaTdJhFCm
fDpM6X4vRGLr0XHMy8m+hYHLu7piYEvUXullxfimQOWNvAvFwBHpt0F7gl3iKRbg
Glp8qwJAjSLOkiSVSFFhQaSk1iGulKNG56uGPWCrNT00+2ndn3D/XpSLYgStmyF2
0Jj4JqD1S8QcM8x8wZVvHTQs3ch+8tuKbbuNtvHbouQAUF3UASwcteO4VMBv+BeE
VAL8tu/O/gi2mVRgJLrfhDUISfbtLvHMeHeF/3H1FG322KelGF6bMGWycts//OIb
OzYoHkDOJBpuJQRE9xKLHrT70VVgfPvX7468LUek08HbM+GF7czyAwYCqnFqKLt5
bxwsSg1K2phAzmz8GXiMJbMti0w5BdGEcHEE/JlXqUFN/vU96yn/gJ3flTkvHd9M
bf66eABHu1zn+OiOINlyGBdikKnfpheqxosOKq1t7y12oEKh89D1c/HAguYdkito
a+xgTWdt5GZDQvJhXa98AvGZ7f944hHC3DNKpLlmBUVCfbh7ulv/dGpnCuhVJBgv
7YCokLyO9cKvAnliR6YUzmLisuzUZuSr/FvGzjcQHJ1X35+O2P7lDpck8s3JkrdN
8s3TRjf/IYAjKiTOxeXXYuGXdqu/TJbYz/9Q/K7Lg6s+AEWJcqLMv0uwk35CpmRd
RWHOOdbE1/1/UKf1xJDheCzY/ICPrgJHCBGq2eC+rSHawXzhgdgnFjRjExZ09+ir
sJ7PmNSV1krdqpNH3DkyAdjK/L9b8PcC024mVyJgnvv9pSvC08LNN4GkC8welf06
I+lWjWGA382/MazYgIKJ/e2jdklRx2TZI4hc2rZMftQdUaGoLVmzvqMpTT5ZoAL7
gKwu/NDJshjpMqoOJ6JpDEgS3OPgbutZhJvYFJF8pru9CeacmwlRsjHjUkLaWSDQ
5sDUBI3voS4g0Zc7V+YLIdJb4JWkXwFUosFY/bochMPnW4iYAaIt/F0lS/22W6kf
FFA9UJAcJXfkU/TQwMzmg0CTesNgd4CiAbq0LTmO4oJzTVhm7eL/S/nbwHyIOppi
rGSOkh8OPYBw/Wwzv4VXOBGT2MsxQ+apl/Do0AYy4SPDP7iPyu8Jy3TBglijpZgD
f79wsQ+G1nuKvzDjv8NtbYgkXWBGM/hWuUFEVGqwTBer82CXWJ7zqQ1gMDP7Zuox
pMYf7c53N25co3w+/0d0I+O0M59gBjptFK3FvClUP6BIsihmj5B5xc3hejNMZ2fC
MxsX9VdyDLALv76rXUF0e1IlSUTSSirf+hx9j7bN4AJQd6AIDMH5fQyRoooZmeLm
kAKzZjvp75Bb1eVvPHEyiFjLVZHb5erELHtaFIqIegLXPz6bGvjZuCK+jt4uNhV/
Q47TfDQUfvdVTWt+wSt3+KGiD/rHBx5gzg4Q/a5b/01REL2ZWrBa0VkjApwVn0FY
Y89YV/4SqseWIub/7K/jLAwUGibGSE+Y8Me+a0cUxUo9DSx5FT6u/X6IUOWEjnVP
vd6EpCak+z0K1RZLji3Uqn4/YSMHu22Qh6XRqgK2X613/LHTTBDEPHGQ0UYIgUWD
n0vAtguCz3WCK3Fe67335H4y0pxv06d/5eXGtk0f4T2rF8ZnHFlsMp2ZbwZ8fTBk
lr6vb+GhfPPHs70aqpiXTDNi4plVEvpMWg60z5n/1jgI9uyamh6VqEzghF/TqsBi
dmGPjAa26XzYWXVdJmmDN9zcxxCy5SILhw5i43c79rB9Pa/KdRo6NXTKIjbmlvHI
bPwPFdg+3DXe9EiISbLlsy6b12wMc/Un+bdOB4zp7muzdv+BptqZrKWiXQxMYKDx
4EaiPWUVEYUSLNT/DiQSnXEaBAhD2H/6kAHZlvd7TDSgm4dt7dmfgtWnfHIPVeXJ
qCTKYWElqff5Qe/nxq2Ht6r4pexLtyvlK6ZPp3jKHXHrXc3+ZXAWjVq8Qeh1WaSl
e7sYCLYyV/R4i9a+4OsW432udasHHTqCoh11DY4GdMey8/xCOR2h0EBKChgXxn4f
bZPj2Wca0bL/SLRn+GSSrG0/J7knykPCOUyrM7FEabQWrsFBsa+ZlUsQxtyqULVw
U8gtnI2gNSqLHcVzttms2tz+NxheEmgjVpTvEiJm+5L2wvoYx7mP9eXoymJ1Eq+S
5pCx4fhhKE3Iq+CON6Hg+cW3dO3MrlbPSw3UVG6qyQG6QI7UUlT0+Kxw84ez4c/Z
HmTie/AavsrwInX6LiWb6NBmpKb+PcRy09bDFFjgxtQOB6fgF7y5Uofw/CKrEykG
SQJL4RjjinCL+NSF4SJKkFUlSIBEvMR9jI41gri++D8yVPZWgC5R8foMD0WHiX3p
T1ISrLLqx6s6I8qibuJRFaRaWEHyHZwqqbQy7VX0qx6eL8FbtywMs9Q8Z5gixzCJ
K5qK5xDFYvorkcfuJKhg20URAOgTjFJpqMNRBg4g3ozm5HgvT41jrbI4VLLePlcN
4Or6HEJDkIXWelfkqaaNXh/Dw9W3ShHxHR/+3f7RrBL1NF2/9uV9IqGPmvsMHsKu
vPO73uUxvM/PuJauxgSGPI+/qiT8BkjKa+qwtDhG9zv1L0LJVFKBno7Y6Zfy9IXc
Kfg7BUCB19bEBbk4K7aW58m3xcB5lqC6QSQDfey1HdyaaM+GZ/AzAsRFkKsmYrkz
W4noIOoMs+e8e4pMEUxzx1KIvN4f4zHidANDlaBvIsnfsseHbBr0+cEYce/gj9+9
YaP1HUUPw/i1pU5BQlSIHMPABAzs5cdUZebeeLyWYnWFnsi5dcI2pMNi8mt3m8Zb
IZk2M6QHbf4GJxIPJQpAQpoHLmhIUvgnzq/Ohm5SxFfVuJg58fW/dzCWVigljsIP
9sFpYG+j+48Rlz+vi6SLw5L8x5z/5yPmnLLFpEbZyhUcBNQKRv79nEZEt/Cew+Id
Jh2pCkGT9X3YWW9Q2Fewqq5DD81nCv8XmEyKgQC0/h4b3x62BBL4NFcXgdbWhIL7
o4smbvj2FsD+an7SBLHL3AwjyGkHWBmpXgh6wdQ4M38QckOfnAcQ95SV9R1n5kq2
CldSw0a0mV3klGYE1Y5T1uM+QXEAgYd0TZIj6upUWw6y4UROViLLbCHV5Z71DeGu
Jd9QxZI1V3hwfGvHaiWF6h2Tuwwsra2yoo4Ig0tVPE+LY/nRvA/nDur0l8J4gFnV
P8y025kknxjBRcqoN9cz5AyBr4/iVLr0N3CW2UOAxbRT3T7GlASrTXzzaqxJEW6u
fiE9fP5mJh4HqpoKvAqfGI7jrs9cAZUPzXNzrlDu9j/WtxJShr9yyHnNp/RftqKN
Fp839TPUqawLuufrD0ixKPXBu7vzSW6F2G//jSKLYaoZ51duGfKQu/+GqQhkAxlA
XOh+lcZApyhLkIPTSd5OBtUlX/iMK4TuePuTFOg74WW5VBGTIMWCABLpF2lKPtpw
wMb2Y5/Wlj9ckOGrdIVI4LRndgaB82rldYTjIFIXZBDuJB2UXfGT2w8oebjtwK3h
L8KDLambrL1IpvgdH3F20Jk2iDIsDFz9voGFi3q3vtCvY1UzMHkYoVHTfndci47e
h734e1TnK5VMjI6SBcZufdhJ81tTZNvx/ej36rUHnXyuhkyHmGtKjEF8FUDicosJ
Ce7M1Ao6o3edJKnP4kAk+X5t7cNCZ4xiVBNpBhLyGEEklVrxP5R7olj0yP2oqVeB
yns3ZA9Ycu5qbnPYjMbc7pl1lBWaWrkBIIhdoTrVJMrBhJLjbvX3vOxFpKVPT/lE
5FKeBydM2BBMMF26n8929+VR4cWdJwKnYOXi+Fq7cahvMVNrrO3BwHg57W+hThss
4LyZtbWL1XjeMeGkrG8iOIib/aDOFobxPHo987MefRXq1mFM55Xla8ih10Dnp7HJ
WW+sPgyfPwpEq/6DiU1zZ/n62AwoKkbYXh7eVKcjzY2niwEMHYb6+kVKZ6z0ba+0
GBFMTvXWhpvbjsRvyEWh4IS4YFXxaZeiAlFI/uggbsJjRXpyDnzkz6aSowxCTnZt
HVwp0sKnYt36X+avb3LcHr0bd6GhxciNdALTHMSGyk7TA2lkrUS8LTS6nU/yXcCe
C0AC03t9+X67pSZDQXS5uTFyYhfBh7rqGvtXqwNCzs5nn5z/KyxRG3ra2MEbqWm+
0WddAxTOhyTZowQvwgyXPvr8290xhGl7lNfqA6mIXdndNr8w2sB+NJSPzVtQ14K4
dm/f4sDHalm3IezjxFXVShWY+KSxjEhbpMHPSCRwYT6s0O9IDEo6h1D37Lpy5eAK
12gEEe+AsiYT4ENgMXIxjsJpglG93s7yoXBm5UD5sKOPPqOjU9OlNjg/GkktZag1
JKYJOsXPFjebqYr2IL8z8+wTr/MmTZzQq+5SqusvOfVff4YrSWWpR1TNK8EZSgRO
rkQ6SiBZKR5qMdAaUBYozp3kgd3Ip1aVLp7mV2cz2ovzEMB8TfOfvYDO/cRjBH5g
r5W9grrpRAm0+IcA3K90oj5IMZPlzqXaRNHihzSkXdjpG2DOVyIuXMk9NAYn2g8R
C+pnFuitHr+JhBx3QfIBSsJpyjTS/QwqJ3fGyeDqtl7BcsMpanbW5ECAkPpVIZ5a
b+tgc7JQ0IfSEUYaUQlc0vchXYZ5N6yL/JKF27SP1vAZqvsP5Th7s/3q0C9TrVkU
apIf2P5OD7aKteamT700mfM4E5VuROyWqosI0JH6aqL3qpEfHzJeHz+8cCd7ccjm
0F45wrHub+qV1IwyMYkxqJqyMAHbATzR8HBGytAHaCw4NxRH6WRucrKRuT4Byy90
2iQIIKxjpFMrFu+wnGPF/d52sMGj3WhvVnrVQwASNyUg8lZuIgnIR7fxZkQ/70V8
U1oAEl+HGBoaFJq9qHChRJa1CVzKrtgkjjSlbCCm69Dv1LtYat60kcJjACcyliAJ
S1/ku7IlcGBi71k+dWm2ovYBJGxNL3WMVIDKA2o8Byg4VVEa6JkTQWXNcMbYCc+C
bkM51+uJUtuW/tB+q0JyNsl68yvuLqrEEtnVfVhuxGa3P9GeeK5E1vSQlg5ZAcMI
sK5NHgycNNvlmG6HdT0ybI8u4GFC1Ie1GOWT8wwIt3eXoJKTpkajSTOv1WnfTG6m
RBqsX1yh+GdlX+banteMhmL/ZuFtgvKOO3aFKF9nn3Gj5Hpe7z8QoTof/YTWxGzy
VNyg8EkSHUELGtaGF9NoxpeFPncrsVSNtpPmttESNJmXOuEiHROQyqmPE1WmQ6kV
ZQSbbZGyn3LAYPwVv9MeGxnTRPjBpuBdB+IK7CQzcVEpydiPuCLAib2Ri/2+Hj4y
lzjqtUFXT4GDBoyvs4Y+FuWbKOclUomC8OYcMoRu+gPUVyJA8hevBt5Ma1Njx8E9
qDvijgceyKLppBdCgTtHzRKbdiJfvckiXamG3y3S5VW5IMSEsj9q7qfSPqCuSejG
u/dGS+l2RMCWPzDPmIV9eeyEqobnrZdyE9Gv2cFB4ni/Sq8YjvHvdnDRyMKbUMJn
WLK0P2aGj01/2nm0mOoQBlc6PYPts2FP4+45GGlAnV+/qYxU0/4wY8tMqDTMt1AZ
mJq4AgkZuzxCgHeSiuNGId+8c3KVM0KMy4buHMH4CV/cilB+6ckWxVxK6Rn5OU6D
RuiNlSLYkl1BDGx/Kd2N0I3CK0bTZ2kVMTf/bmuRQFPtftCW+wQwPoiBtzByLopF
aZag54O0HN1Lc7WgRuSr4AxFZEEdITy/jjPcWXU6kmr9f0CSxf1B2wb5Kh8afNQJ
eZucLBFTdnncUB15oyaJO/qcpaeXVzjgLcuqilnA/x3KJxG5apEAiWSnBDO4NRqr
dUZUq3UqdkycXs6P3dI1+MTxqPf3GO5dV0HbX+etpxjgu4r8fJTOpdVifmqVeaXh
z+SsAp6F7lPEP9cFNQzwMnVoB7q7qH0vEt1+li+toUhAzs9MbbFFRjAl+KViTali
VzmPAsVBuyQJSEg5c8e2w8kLt3YwAwIFmIqfbWLkeSM91hsVHBLWgQa3gC3NVEh3
TW4YrdOJcPqtFb9c3yB3t9Obet8ejA033WmFvzdsVXleADxL+m302nwe2xC0PiSF
b9qFw194R+/06POfIS73Ct8xs+k1Ad6ayz9OEvykyY7MJONed5F0+u0laIdx98a+
QKFMD9tdCGLEtkNgm4GSzDb+6+XtCveiZGmcOVGaDOCRkYzGvz2I83BIOHMtVwKE
R+PciremhKWgZvPkMFznYsV7Ynptk1y/2NwxQg7RU3+z3JHRxgvtgJA+8G8tGXNB
q4FMJjlW/C95fcTHtbUlQFqcJAM4wlx5keJjc3zUDSLG41djGPokyv3npt4ex5DN
8r3UgTw2iFatYcU4gius7W55U0r+bUhyABQF9fyrVtX2IvBrA8tXtKdjVJ6XTeBn
F3jBddBlDaKCxOU2IXBeBiCWqNFSy3ff6/W3OXutv34u4YIRK6nZj/RV8URjJvdA
1Cc36akhM0A0XEp3e/ku161b6TVe/Lvo4vKJbvljkl8GuxqoN2WFRddwoowsCK41
O0fzf5cuRvKIYqFHVuztp+PsTgrHN0KX5ABGnvTgL2NjjpGvmhPrUA4DnmbjzUlX
5rO9d8mIZrpMzNyQAKiLqZoNP9TSCQ4mpImaQZlRxpm1x4XTo272GcaIhA4gNwBT
nKpvw4rDJGCj9EtWvhFvy8QdqNjscYTh3U7RSjxyuWnUtXzXuucICeeAH8arAC8y
0/4msJNvGN1aeL5v/tvuq98/rYEcr2VXhPwfo6zd9RPYBhNv1e4yfulzd4Bg31lF
j+6R/RThs2uN5GX/zqs+n1UVhDtj5BrYMe2odmCYAbufOHy7aRKLoBBc9cVvjj69
H+6bqLVNMH+oq0RsLbTrg9UVrUJXyK+HHL+fZvh26jyVbDM71Cffr1iYgDdcLWMg
BxwUr9Q4vBcM2s9gEExJ4fJs5UcJjbbovA6wNdg5m1QmQhhhTZmeMr1xHF4x2LGU
RScisuz1Wm+qU6rgqCp2vcwAvNupRWS3E6snbqUPOwlvTkLMPVpmslfL6wNhdOmH
LQ2AAv44WgZCZxd75HSrItviQASiTM1UpdKUxG94buE2K3gr9rRdeBtII55q0Jkl
gmvkoEI0KEDKxEWO0T2r9o8pqvIeH0x4wUaaB8qM4OW2FCQJmfBV4n0qm3OUjs3H
5cdNHhorRjItR7xG9sFXvYsTKoZBHzt6OQ675rJJKkaHSIdzWfariO+NBDiEHbjI
Nv7M/iZDzu0AkMfIXEDEOb5eQwPNcJDY33+GBcmW5F6+nS0AaK1gjRXoGqELSCCR
qaFNSYBV8PRXWR3Wm3P6+zjR3pymIHcIm+FIFEksi8Acwm8iGT++AfTVCtTvSleQ
HoIlqwyyeDeD+9dWm0nYxfGLM1Yd0Dg6LDTL9K3buBtrLL1RFaOy/1tar1pdHL5Z
wSAZng7Y5rQTRVa/lGux6JtdqKDkwE6ceiK4F1Vv7b+vAKvy7DjlTXsK0yeCrEGZ
DJ0B6erdaM/EJtbvsJBeb4JC+PkFvYG6pYtK3qEk7mvWW2uXAbwNdkUDOmZmyYyV
1/8tbfzzRV54NzbPrNW6NwqY2dP5TsmcgcT2nTV8LiVDCE5d1lLUjYQuy+HiG2u+
CliCYS/oGjorB8fr1aTi/kWkmmDUCGTulx3pst2q7OiPZRlLuJQ5JvA26My1u5dy
YO9VKo0UdTx5uZ/LhOYbOjXfA6oSwUqCImfVeoMaMs6DHLeHhIsl9D7jjqjoYSFH
cQuTx907xXDCMAEctj82lTCje5dxaq1hQOCpT9QzxBkGunncpJSahXwHOZoQcq89
6HPlNekn1h2U6XC6RUtHJ9/QQcGSaLCb+1vUoltuvwbV2AFZeCqJKqdH7JyKTJT/
1GmGSFm8D/dI6EKUuKOdX8mmg8JVJ/hj/+GcxF0+YbXP5NxE0x7VNuPFVzeYA7WP
CjR2p72qxUpuALAfOaOTwJHgYRVUinNY7WWGwO8iefa0rLGB+398UQ6NohgN0dV0
PavfD19+pHMyjbez79jfxhvKc8YbGRkcPH+QdLD2YHe7NHDvlmbX+Vsn/kqxDcDi
PmFnRLDcOCPDYeG5i2JZuxaShn4/vpQNI0vcfjj7dQ1YiZn63RQ8RgWuPV7fKAMC
WcAVJFMlI4pkVA7nckbUOOX5b+AAutswnIqnesw7NiZHB6AOVs4YLnsKJW9Zb/YQ
Zhnu51jycB1IBqbmMYA0Nj1/yEsHghJFjphZWjUEx04Mbz90Vnx+RpWoYHFmeoke
4TB51E3BYxaMf0cEWiF/zmgzBJfhK+Hws/8C41Tr175nKLTxRxCQZ6IAD+j0FJ4T
wF9eavkc4oU9GffGzOb4N6ieFLdLVM1bfvvUEyJY+zkrSuQ+xOWegsY8Dl8MYQYf
FbfKIdQt9zpWMY95J6DsvN7AxBTQCNtSCvVtIU1wtZc/01tlAbG/IUAbEEeeVBdJ
KW5cKZR8afCbTtJfycOsrJrl99Gk1LvQ34yw8tTFl3w=
`pragma protect end_protected
