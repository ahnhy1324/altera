// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
d83O5gNNLyO7OU2ibDXpCTL5VaZkHq3oeckNKUFK0yESA+Xtlr6JIBwMEKwKgQ2J
Bmv+DmLaxTpAt6HXEhI6zVBd+A4jGZwD4dxKu7diKpJGX1Wa+2KeIYcXjY8s9HD6
domXfIv9l/Gb8KYWgoJcVFJNaQ5BxDtaLcwi1ABxMmM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11712)
GEYxnBn6NGwaEfiMs6zZhpFkJqJKlkLUemj9bvg73BmwfaLW3Nj9lbZ17CK9aXyP
JR+OYZAVshcUq8z9XxaaF6UEoQbTQxTaLTlupLYCUspzGn2TLE5hktChJIG0t7fF
enaiV35m5isxNL6gGxinjXzWABcWd55nM8k6TXJaUoFiFjVQG1Rotk02BTz6sF+W
8/HHH83Y3KbQ8HHxquBQoHq7RHmu9PdyU3odwSt+cVLIWwAB75nt9oO1xTwAkAif
+s3VhdMIw+ial9Ui0fr8PPgycKEidCBnmpOJXXhODr4l4dHyJM9vOaKrItX1h8sC
UyUb2K8sVq318JO5sIvT51rPqSE1vC8WIuh7XcgnRbD3zw8Ef3mVDmt8vTkrazSq
SifPMK8MreQOTjF9pYiiafXhsK6NoG4wOGNR2FGPde0SIvK9ZNoFsHm7rPf+134u
3mB1y7WJ8MmhvBZTkDuNQxAN/x2pkqOvVMF2nm8VXfYtRK+D41DPhzExxyGK1BGn
CPyfsfgkgWmeedLOfAIBrrZ26AQj5f3NOw8UdMHqGnHLHSrY5AjqqfVPqXjDOHEq
bqfyrS3Y836njhfp0+28eYVBsiUnAD+o1/FtBbm1MmAG0VCAawdBLWEubMxWmU9Q
KrciwSe//Np0dzJwZpM+mzsmDD71Zy1hH3bZGkHcr9pjhEoFbhKwCzuScK2m+zrz
aIT+bIkPvGcA5vvtw1zPWX/en+XLW0n+DF1VtsLCiwGc6ygcx7Y56qVEsbsrf/ob
yypfna5AUuRslNpfz61B3tuU3MCvvdQG+BFibBx/8uEiE86NOEDOJ4pUZKU3bd1u
FyHWo9+jijlEYSnlXZfd5H5j9b6dpXLQQHKEjcs99ygELeWiVIIAIwA6WAqV9qy8
Yb3UGekGZYtK+swsRLvrsDPJ9BYhdgdo7gMJKJVZaR9DdAt8cFUGcU8keKOoq5Lo
1Y4OLOTG6DjvRSN/1idFsEU5Zove6bOvusv7XtEy5DfIpLw3siD8JIrHvaeTIByJ
oV8/SVFim83k9/lZSKKetC5V7LepdGrhPlqrxdpBmPRjMlkqRoEg7KkmxFqUwNpq
mNf+ZBQKgAHqbxpAYVwz0pZF+YUuXvlQS5aU6j5Ly4YLdMdFHkrf3np1Jm40hvxB
zHEnAbS/pgv+mclC99NeAdWUpu/6oRnoAgdKxnQVzjac90oHd+hDSGnWnZrKbr7S
RHJw5GaA41neNbwaSiS5289jJMHqQ0prRBMftMGSB4VGIw4fnXhQxoqntLCDmibc
tItZx4R/qBfEsaf33uiNz1yuhG5ojRb35MWs7m4OdeoPh1z/b9b+I12bm/8pVALc
95GusbHxJ/aCVW9R4sougrN8fi9MVlUTJ9NN6Bt4aT4FLd18Ldq+Xjbo/D+CoQG3
5guETHfG0q5ZlQlm3UJu1GuPq7ikC438F4ktOvzv6pSLt5uXhiH3aOm6HP2T3CFL
tL/E+6YOoDJ6gFdumgmnItPQNGlxBAeATccoGm5NRei2yVlKeMqrKSeA/rDNa+YN
KuYmIIkWZ5YR7v9QPpm7M4IQQxy34Xez5k1s9dyqDL6sKIvNPGe3POmrYRT+waMQ
sBnFN9dSz0DKFjVJoMBHlMsWrZso+ALUpmwrHxd4D5e2XD7+ejmvNVD8he6HZGPi
TdPf6yfwhheyzWyc/WsJguqd7co82IIS1q6+8nVz34bCmP0T3L2Koqltl/1ihKwc
VmkSaJ5D6OdAy9GCm08AsuelzStbSZGNBn/gUuUcBLaxZ5WUWTwQZbf1g4lQduoo
cHVUx5OfdtsamLc9cpXsWo5CVseEXWoAMGJ6uX7b6QmkoLd8ekTYy1by054oPCND
rt6Papmw0XmiSSkaSFIAJgUMz1t/93oee7CvoMM4mdR5V8fLPCK83NknKe3HCi4A
vQIJDGi91MiD8uIs4i0vmqeSeXARi8yEHkyWzNNwOUO6vWCRPmssVXJ3CMOpduUA
1FfL8P2F1/VVdCpCZsefpv2VXvAI+SX3PAN48E2+voHqfitZvVlYZcK5UXaXwEIe
ylUKAb5CramNWZ3JbuDd97YfDii8qBeQfaKGme3nx6sS1WDx2wII8oPE/I6arwiJ
d/+PYRdRDqMPbB7n2IUGUKN9yEdBdNogO5v2YWtbTLrQuSSJFkyFS7aTfMxVzxXB
lK0x2zniLctO5rf13lzweLenhQvUdhE2IFzP+f0fKUW45z2ee2zdeGmBKZCnAgdQ
kLh9o22svv1jMmIJduXYSs9ehkt31CM4xYc78JTsZ+MxcWFBk6lEiPCeBQGW5ogv
YjMbt6Rjr5lgDWEaxAHcFrXronkhMkTpsQn9Fvzr8oA7/UiXcaPeUBYwagIcyDnR
k08iwwyHd1a6xVVdG+N/E3SKak47F22h0OrEXJANj41AldBbhkC/jQvXnSuue/y/
UIJKQC1o3geujQnjRGvE+oPKFHoxxrUfGCgDRv9L0Kl6JWXDQ/DiKneCFad+7IjK
FxvJyAOC8mQsY+4dhlGCfddTc+L7GrJdtNO3g3YMl9l6GtfcT6m6SPZUPmMc10M/
hD3sVjRhp+rRkpMTrJmdf4w772d0TwiP7sjCRr3gF/1UfkAFz69//msKYjcqp7YW
Zia0qUFMYwhQ0FuxOdwECdRGalbuxElGE1UjF273c+jU+qo007hv/5MbhEJcT1DL
g0aZLN5y4rPYWuu1Jp2ky7kSfxf54BRqs+CsTfnKG7JmpCdyzF/q91yTnIBOfKbA
4IeZJMxN4cld5vbrJDKqPzf0eTTzeWRxuz55NXEYXL6z72VaCxx8VI3DyxQ4MQwm
qi81oTD9f6xmmo+lAw2eZqDqQLPY87c6mPHaAtE+Hwt5D2RtsAc2Qxx8APwj8G5c
JbpOP6g+rG6eZo6gHFipiap55l7Orm3YgrYomyIWa3foBBCsvN0Etf3JuPpb3YMa
pvR48YzFpyd2EccQe3tnf7bSJa5gMn1mQwoiIkF5Y2xwISNlreABLdZCUajiU6l9
H9TdsXEA6nyyRfH7bkQpRGef8T28DA2KcHZHnhFCO6md80EE/cFgPLc41a267bvE
WoSWPT+nZYFol1LsAdy4pJVcQMDUyRi4+sLThV0D081DNDepI1qejUUQGp5tHtGu
Pss0nNz/k2s1pSt3J0HEnRP5cIRPZJcsBcerwTTvAk4P2BAzjArEv6MqRIiNf6up
g0vbPyJq6zmnEP5S+E+PHFKU+SKxYS7DynJG+HBV5h1HFnAezAqy+QbY+sI3Twxz
8TGU+WFtq9l0b6BHwqpKy4cGdWKdCsh5GaRaHWEzeUabflmAa6HOB0AS3tUVbdZl
72FR5UWQQetpZPo8W9Ycfx6OViiwuuZRb5tPbhpoaOiOgIDmVkcxCuxOQ6MHGgM/
q4Xp0ClIA5CTp/NJ2oLpdiDCnL04ikWH+3bXh4OKUWvHywZKdcm7W32CF6X4rnDG
vy7qlz+lyYePXno5jtLSs/r1vlt070Tjs1KoSwC8Mywyi1+1BZjmd0PQF+66gj/M
tz9brxIX/agYtzZhFNJ91dBUjEmhQcyIP62aY5Ftj0mqGxcpGrZwX1Q1YC+3s+kn
ofJzlDZQ4SiytyTrfzMyqP34FX1y+w/PF3ORAl2QqTwRi82D6HS/1plu9En54/tC
kkoPIxejUIa0OauoYINnBPpolxU3q1o2Gz0m2u2bp/10bv853Iv/Ruv/xpxSeS/J
FyuGRrxo7JgP+aT32AvL39cvmkuG3vOl8grNp8ftakt/u8BP4RWZUPGmOt2GjlXY
pcHd17hebPB+69OAhxGLel9aGny+5tBG0d44MEdR/F0l5+M72vraq8YBSWq8mnw+
ZbS/P6TzAzZICWVrot6KNNBi2vFCYZiw6rusvmbgFna7r6DKwYdv+oedt0RnchEz
xj8VksCKyVc0Jl3Xo00MEUkhUQY6CrEP9vkQ2F+WgLuWTNVTI1tKOjRnJ0L6q84M
io+Ywqa6LhoijRCDsbRWsDeQRLa+rqKw0+AnJB1oUIb1y6NpP8S2T5plH1r6ZR+Y
nsLvbECGHH9NCgVa6lU0eoO+wMFy+O3d6YugSMwEjb0lzkwrvYG0LyzWG6sbcVEP
B2bhcsR6WvL62MdtfbmK4BFPFa508tH1+ifJgumUIQY567HmACsuXYDs0wMOc4oV
1HzzT/xn9zsoCVmh9tOnTBURVNkufyt15FX0ocTwrIMpMUJ9YzfkW5jrI2VsKcjT
DFS0ruIj2e6OqXxCg0OLXLLmhm1JcrZtjeCTJBGABipP4V9T9e9yW1KvHC/J/VSn
iAiJwgSZ6XkU/AoPBLwcr/Zw17XtBJSDP+y/LvWs178CCM/egik579nf51XU1Tow
TXac1fDQESCUqnlQ/PaIqhEZYHtygDrT4raJleBgpfDSMU24eN1/z6+VsTe0wid+
05wM8QwQ+BSc9DFsH4wF5Wf5+njjMBF4L4VUvOdYMap9UPsA4NPKIrCZNWdaIUog
zrfUaii+CgdmW1ys0T8e0DDQeYty0J6xNRBn9J2nInH7Bw30KoklNibttk0PxQtL
4vDiuhb2JDz6VMPkX8JAz9lopHdc4Rtz5zghRBl4bTPKSkfyPHRV6TpGCcIujvQE
ztHE8R7IN2Jhm95/BUD+nzoTubG7/au3S6AU6qbhG1BF8IBvS+oNjjBBCTo2MHCK
pvpJMrJdvQYi+gM1d+eRBrXbBvyVxwSoBiIdxSS0uoJopJrCTE4FmbtEUK6MRc6G
USCZrho4eqDJO5j2r4Z3IrGBcB7eWnmM11rsM6TmXUP0YwXGuUAs3JaTRUigeXiy
IlKB68rnbD4xY6yZ4NzHdkqeAIAbqeP6a3KG98OY9YLZXmcZbp+f4GBbYzs81Fpz
uR0KGOplK7oCETRuCivofxHLZtDk8Y2DYsq7Ep1jmK8AW46APDQKESNy43i0LT4E
Vm+yq+yDk/hNXxeUibYOvJBekxCxlDTtGVIXMZ0O73Nfn5h6tEvbjPt2R+FOfrk1
XY4Aq+X71+EkNETbeUdBTLtWRiBvMgpgGbROw1tcQ86Wmpjx7OpbXxpxPXIdL6Xq
xu52bRkLOvXdvR7IstGYH95JmRIA7ZGyl0RjKQcE9YUHKFRiuF+wNonEa3qZB98R
8i9Y93ylwgdpMm67VfLVLdWOAgcDmar6yHvlT6cYGAmJO7EYuIzgx1zx8t6T6uDJ
vhlMlGKe+bZ+taWhX1ZuRtasTaZvwhxk5bZbjFcEuPnztvD7fk219H5cQbeIjXDN
62fltyGFikpvx5733vUjoR5ueCigBwTfQVFZyCr2p360LacKCa1FaKlRZrqhaa6V
2LFnfFnQtDDQS1OSAIxnxBhfR+oGNy7qNSayvNKhN/NTPRyD7zYg9w4uyTxWre4v
VttgE17Nizpz4LmR1QGNYs9LNsfpHXQoj4dcPGtM0Fr7J//Ov8U40MFFD7BrHc0u
xUILqCWaQOcc3ZsCdmOe9rkqlyCjK8NU1UE1suUgHbVz0AaeJjhNy6nZ7G9UcWRo
cxOyEtkOSnDYJFg5A41UHYB1SIL5946zZNSb91vPe1lJUusODkm13f2ALa5XFOwJ
99/f3/Cf4elp0kI6FJFUPRfvkAkRH2oQgJpJzChO+u0GhTdij4kt4vUWQNe5Y9/I
XiziFJ+KGn7tjgPqV1fyOqUZ5rN14bOmgvm/eT3cWjKyH7uRiF/2zYXRkqRQ96OM
s4TogBQecMJLKfSkV1wFHO7V5PqZc51feN5rbWQ3lFv7U6KBXfqRY8F41P+sUhVJ
Fx4lCYnEqT5Huu6PUNxS72VaqUEdns4+F7mkfe5A1aT9vfoZmpHUboitrVSPyeat
FJ4+H3yX6jcASpT3ZmWqi13dwXCStVU2UiVd9pTgxlLSlaoZ9QlkDhO5rOyu6DTg
GMCK90eL9mNcdphNfc3kVeZGetMbUkjav3hwEa/UG88UtBsz3wq4mJXnbs4f1oon
kAgODkW292wYzLP3YjWbEBU6PlUpSf/Cb5vHQgTvTngEoAnR/h3I4m7ZvOx/1z6j
7DkZtxi8VOMchEkpJoyjWW3vuqzjlAQplnmEYtnyLvlF2HIvo7Z29YX919i/aXzm
jGfeJSDZC00Wh68GEXu6zGIS8xO94CZwLU9BTORiIw8xGhVFNEaoM43SfNyV1B4G
nBSnf49ivT/+o8q2J94/ifjT2KAOmvc3X1ug6/37ZxIF5rd/np0nnml6yo7oCJLo
81K8z7R5ghCu1S4dQ8YETmLog9CAZH5KwMYnRCSF5TucyJWTBo22h9u4RYJTkY5N
mYmqWp9Ig1rCUAfSyROfQENfGVnrqUekahBz7QKeNYvUXVzZe2WboNRh+SoOWy1L
l97/ShUPPfcNzEIciEyCRmOcA9hBBiAV/NkYbobY4Rm8f43JS4Qosp5pQQJApyYn
w/2BaxSYYIgISIKZpAnWy7FctyUOtsnptawaGFdXQHZ26sqRYIEI599jGrzjVuWv
pg2+Bpka3YV/p4mnf2OXPjKr93ngZpt5e9/xIbWMts6fmzvXKaGHughwM7yBnzyG
bpV/N/GlK/NwDEg0gNSsImC5Qc+Wu1/eAMkrs+la9ITt9K7wDAF9odbFVPg9nfqO
BPa73RXgjIz1k1LAIDsk25jeomiRk+GpHncpEewf9ZmsAJigXUNsZDvTcPzGb9w3
2OdweASz9cvVuGxTchspptQoo+7NqpB5PSv16ScWCwOJBky/n7q7BsaykVHthto8
Z2noo5CAgOyg/YPQFwtUOXNGnOfBHrmSaKkllGKU2z1QPl6b0VYP+QtYOALUrZsJ
Or+goWYLMP0jeRqkkzR0FrfxEfndMBOmk+dlsJNBy3Y7ILH8fZaWFA4hXeSsKnAp
WHJDlUhLHWu4Nmz49TVQWB3eDACj7j5fKF6JXLDFRFUMOvhpNJzKiI78SQPtZ5Ul
JYJQ0FjjHJ0t6NGrAWOoppQynnZGDBfjtDZyBjIvbJeIyab7KF3BCm7XzxLr/SAM
noHzy2vjQirJzqW2DWENaBaI+AFZkazvk32G+mngHhsfgv3u93LOCZRWpKkMFfkl
kwswl0jkKtoHD/+1DdbcqzLittJrT2nwLhnLSVyLObZCJGOj/Y1cKHt9ZLE/3jjG
OYRA16BMRlq5RTpQ1nfvjPTC05dRiv4pPFpy13k2K+oqLweibK6+WnrV7QY9NsJg
G3K5XQuV2Gy1D9NRwylK9cSZK4lc0CX3Ft6dTxw2kqvyvzTJOaM0LsiOtNxnorWF
2Lu1bCigl/RaZ6gZLz7HZp7vNnufIbvzHld+naBi7gOK4oe33E3nhgwfPLpgK4VI
u+TdW+42A6/QXkLweHc8wZdBuAzR+L0pj6vLtEWkE+V61FxLvRQdvdUsW83Y7ZV2
qaabKFDt3mmgqpSapyHjJJVBO9HynE3OhHaq9o+U3RFu6DWGH8uw4aS+Ov3WxbQT
9A3oPy03GEpyK3RaG1IahvVGzPGFxAqZvAYqyeulTDvnfY7UIB2Xckt5WtgLEdgH
C0nuXkf81hFzJM6EI6UO7qx5Btm6zg3d8RB8RP4jwVDK+QBBZUlTB3XoF4MpQpUh
tXd+CINFyy8tnb0nEFXPjVINpLb6oH4+rpZk8WBB6KNHBdmp++OHzQKFqmKQ5Fca
ix4UmpZ0bUhAGX8n9G8i9b3QpxYmPTNLrf3LyMyy34Ly0rRg4AqMZEzHM8aH/+IJ
csuWy7d3ywygmFjtA/hnnGf3U30Nl4TyBbuC8fhe5lRDJ07Kq+p7QrnTnYA4bKrp
+r6yu7qbE3bAN1aejmp48RXr0zIYFvVvrr0Ifwn/bdGzmDF6zy6RFV5Xl0QXtnj6
zo0Jtxlbm3/kZtfrT5dnfUbZogRXs6mRov13cOwkz7yJnXLvVKE1kQiU4ZbTlt7Q
4+aYu5HiPj3HISLcI5n1YkU6HX1vbzmFVVBZ7M9OzENSRSi1cIF1ErM0pCzBopIx
PctkCVYrRPfCOI1xcvCRNH9Q1nTAFBoJTQr1BCPbv45vqGuoDUndcKlMlkVYvtf6
QVQ7j8fC9HMy4WxaSAGPzJ34EafsQO2mAdjcTlmiOkiOp6bUcTpt0C+EO7c8zj40
JiUegcuNmlinfQxQQKNV2iTvDkboNeS98yCPw8GgwpGAnG2fLaemxqi2o/WZ1lcM
qgaEb8fqO7ftFPm3sR7was250Q5y+dyuk1N//0XVpg3q/OdCjd3dPqE4DOS84P7r
owXg9VS1UfCFxP5WOeqTEWeWK3JywHbT0LuOyWouo9pcMkotK7zU6Q0ZLr0G1Ktg
Bws6Q+xQhqhLhSGHaDWEgkKLtIjslz/08tAZ7fgXX5ivtP6okKSS8NNru/kAflx2
gN+eLUyJCz0xhMfAicQIAny9w5D/CyZD+Z8PiCxlO9s7eVnCKAfCkOBreAt5a/rs
v+j8J8+o0GemuouOkNMQvtP1/Fs2TCdL6FDGE9lhqmnwRhGvq2Wtvihr0lDwF8SQ
gCiS0losYBXyLDuOKicORTCEqkYJTU/9BF9HwIqGmmmaHFE0JP/RH777ZQb6W0bt
Bv85WXbDWQoGENQinv9tYRQYIB8eR84A6VkRTrRryvHfthopElZkiGcM4Wfshkud
JKqw6WN1ZcY4euTNmya/BAhSIhLwfmliQd1EPA967Lde5ngjzJw82sdWUEncOsjn
WYStB0tUf04qmhCLh9XnaKOkn8fzrU3gaRG5SX9tH/0p3KLedOrE8GVjoGwf2vTd
5D6/AtEkHz6eP5S1y3t7yHVC1CzQ+EWriCrlUGH8omlVj8JpELMlla83WsGycfPx
cx12Rb3SdDzoG6FzrhvMIq5vqTETLmOt0Ye58m8NRZ+ZjcqkbcElRb6VkCtbLeB2
S9A0EbgYGNtQcQ4EAp4EL/5QSyJL48t6edhdgNzf5AynpLKpz9D94/uZGvpjc7Fj
1pyiWFRfPpw7HFL153BPMRG07tGYYGil4hYjMEX2b1plaQVwLboH5gZcuGR4ND92
M4za1wgB/9fAuZwz66riOZIsbXEe86s4Yog+oW+HMF1I0ie/sn3YGUkL8Y5bHJ8w
Mo7cGTb9Ohzj37AVBv+hKMaDJte5IB3bQUXxndKJrLa7N0+X+w14dIsxfFQkKm8c
WYfkvzL+ia25Jl+iDmTJHbC12fMMDtBTh1swk0pRsmKRCvGX3bYqdf+CCooCBMf7
KsDLD5Y1QEtMgm33LKKE87R5ArhUQbYtr0v6ntW/TYd7frHNlh7neBXMBlEKEV4L
UnlWn0fKDE+VF9G8hb+Nd5Dv3mdwNYVboUaSPoM++y4L1Obgq1FvCLFwk1uwUiHG
eOLAR0lu7JwKg18kFDmnD5y6iirlgIW1vUCt7kHSVG4YLrCfYUyLgoR8RV1RYCTn
J8pt4eruOAeoC5Fl+1y87hUn/f2jkemMVlz1DBgOf7ieDtSe0xPb1WAp6biuJal+
l0xZbG+ZdBUmgPm0NgBg4tKFZxW1D6t+BpiPBlEeA1J0gAoF/JUd0+vwo2Kzc1AG
DLL3cVHyGU4cXspHRy67nkPIy3ZqU8ZqXVPWALeUW+5+b8HoKr822ZNid/+w17s9
2LoSXzCYBJcXOVCr3lgXuT5KqZMQj3hYoumf7f+ZwOQ3GcxrSYbTn84JfAS+plNN
d5aykRCsYjirwwvkO9GBSgJ/j92wqxiHQQRc8wWzmUq2b5uEEXbWZg9SE+p7K63O
4s/VNbyu1Z7uEDxY6XHVB9kd0GdvrDKkAM4AjntbVlc76xVn0uwzIFh6u25ItDYv
fsKvDeug7IvUb66rS0UogTM9o16uoJAFA4SzwK2sKFE+0gARx/SLiFT3D18EiNfU
kCEwais+D8MtjsvJHh/3DB/U0PhfVUkmMvJMAW6KpBtCbYtr8iUnJcdC8iOyi4cE
WamgpHsW7fduhpO56m+NLAFy+QI0f0PU/8/KcGnLY/a5gfTIcP7tPIoSzeNhQzJf
evyKXta/b0/ZZj93hZFpHV6FglwOpWH0uLD8x72dak5C0lhGRheG8/XAWmvKs4CL
jImfWgnv1zKY9/fe+WadeIujBJargzRLvVwPvkHCSvEDW/O8O59eFkvZ0ln+oCCf
eOkekJhQpFSCBD7PR+FuA70f5T+ldFTqVlF48uU6w0k2n57BHGh7JXjstpjIRXWC
xNvUJS+Ey2fe6briGZ/LG5I9txaoS6TY1iy1HS9q9IFFuz7Fm/ltUXVaAOec0aKW
fQQbR2SgSl+brCMWaqlmKoZUc1tqTd+tHYI36HiJIaeeExVO0UKBvS4ghaK4sLKy
jQQQvbifs+x7qz2n/pMyTGcmF7aL0aqBi6DUuIsAIaIp7qNzWQUFfq8h3gzBsti1
Zhf8Ze1J0fHRpOb7bblMYiE+cjw0UGGW1VTtfc8V2AzESHR3P/7F5+2k8iGE0Xjz
Q1z/Y+5+39BL3cqCGWOKfcavAEU/zZM+rRpElutboDDEvygmiCF/LUz+oCUL32cY
7UIPmLebfsvxynOC0FwdIwa9woi0G3mFR4QCXNfaOKqrtlhyJ3Wd3zvQyMv+lTzE
rJKkJ7lhLOc3E5lp+4C2YNAvYalvQMyUQlI8SVxmAnS5afp6XaiDlM47Ow9sGVIJ
ka0E4KZJDh5HVRh2BrOg7SFrt3GRpcGv4LGppzphKMt+h2rg8Z0LNisz+ZAcq3W+
Fxqxga4noVXKr39nkpg2HWa1kkUktdUMbmZHDyztY4L+vmThJY+/WTfELVZ8FYUi
1GwzH7SegVKfGLcZtmcQKivIOR6uWlhEOCfxrHnuyejniz0jslb0pCjw0ebvk2Ln
FRHn6+Cw9zvypYm/tQXlNAyEvfqaEsW0prZpjjM8kW/ItGSVGyuYLPUSafAxZ6LT
UQu04qtUHuM052nnZc/HCZIFIMuRD/pBvz34hnldxl8JCJ6rjNW9WgeI0U5dR6qB
tHkc7CNufKRF4ucqCCLRVTDcHTFnYNWZzfilRlSHqFKoDwF4bPNIimppltH/gXCX
DQj6jaUmx746YBeFVzCeT7LVt/q8jDABx9qL1SaOnVSX77bE0cJqcH0iY6URfOh/
5L6vqv3uCAMO2GTxVFdr6GP4dxzyCOifzlM1+RdlqeYa9o2UjIYsZSLLEkjXa/47
Kdbix6fw5uP9q41YjEULEsX00DV/qyuuJBkaFrUvxlnr6Yj3i/00xRktmKsnUoXU
2RIwY7x88ntcDqyg7nDLF2K4Vz0yM9htw8HjKUu/Kf/TG/OjYTNpJLYLMRoNNKR7
BL+XhpN8PqXkyC+NFS9A+JtI/f2332L/p+Ql7LuyvFkcsHR7izE2AXoJhY2jRcaI
jBK66XEM0Qr55VFeFQrtH5dkaL8yaNcxh2q0pSXsXUkMb2kfGfH3WPIX1mghQdTP
cr9jrZhx7HkXGIVYKJug1+afbmHyXIDqNtXi4ntJhjrGyAW1dw2Ar/9teqMwI7p4
8cJ30EC31uojfUMcpLCM4Z7DvYBzSrKBPc3ZH88hpYxiDcsvJoGIe9kJIQ4NN/6P
PXuKEOlOPcy7Mcb3/ODyZoWYWpa2TzbfEgstCTVNr5LB+/WArhzLuHPkxx/ny861
aHYG+WYjetQBnhMll2NAE2b9xOJ3uVGS89WaL3SnvEMSjFMskrZHZB/7/rzwCOK9
Le2i9wF00D541Da5MeyIPhzX8UGIPgKFbuPoH71Bc4S1/1si9kc4f7l0AReRk9r7
PT82gZCb+QyQr1NfcqV6Y2U1ecGrU/Fa4o7sUag98y5p8MoRPE3fOEb0J7fiM6Bk
kIzF8IfaD5QfxgO1InIx+8AjvyTFikGyDuoV/XZoWQMjiu8kNlqZ2e33HtxJhRSK
JDB6uOXNJc2aWQjJ1tIyfd9iYyVm/IIVbGHHtkVTHT7195obb8+978BWMT+nSXwf
HzSN9M3vPnBaYT591Ch9rPqpwYbWejhtgUCV/aHocFFUTSNYTK/tJPVtzruTF37j
5uvwshwcbQzNBv8sf3zwyeX6yfD3CR1XNVoAgKgkMJpVERHn21nrn3Uf0gUObBQM
EZu2kMiuRUyVTORu+NB5GgIA/XKbrnleJf+G9XVxb8OW+5FHZHt77E4tUMSh+IdH
6O5dGJCmdHtMiWH/vsTLa/zRuABAGfFydRJ9wGdDNUpKUM26XYxUl0t0v1H5zAQ5
TDheQqQy5K33Tr0ZHajPrbQkqau6pfEDnEqOjcgllb2oY8iuXL073JlGkfABKXyO
0Dr0drGSvRkvo5NVJ1LL7ZksP42V8SF/RgcK56JIAqrOGV7hxh5x5Inz6nljBY3+
ar6Nfrqhp2Ff5LR4E7icbzb/+3Z0oD1FdDGJ22zC34ta/jGgItlVid1neRQeSF5F
1UTLYdcIValzZ+wAKNiKsUvsCXtH9v3qv1H43RLRNfidFeBrKu7Yu8YCwKzPYR1D
ZEX7eLoFuxbB5rZ4BBU84+rFZTsDKUhX2RPoyxzloRaJabGeOHCu5LrVwB5iKG7b
7t7fHZciVlYEZbr8beTBgrKVc6TRzR9pRXQId4eDfrliCB1xsQBa7vtnPrUROJA+
Kqo5AiWya4cnhRXIkBbXQ/mjp4YWdAx0q8y/lhdtYAWUcdMRXuTp1Gs0Zc95jJwU
7Ij2zOlyY5GLmosBSFDfvHxNU38Eh5I4AZuCE8MTCpnLd7nDIGBjU9IEOLJkCwDp
2bOELSnQ7mJqiv3y+AICVCi4GG8qIUW1GDI+jsMpa+sYhIVjRDKvDkINeXWNJ3Jr
4ufQeEVdhxSueIlJVnQAASf8z2Uoj8qNXBMvNVCDAw17wSfZVv7Vd/XmC9GuKdGg
UewXYZg84baWZup0YLyQBiiVbKn+vavVaoUceiFvjnRgoCsMQsoPuuWxIbk9e/BU
ZoQrwvlThz8hPof9yWl8q0eEM5hIWKCBRTenzD+nRKpQNHkag0EzepQryGP/6/Dk
gKZO4SNQ6yykGaWCqKcjw1fRfplET1KlWUpeEcwsm9XuivPZcr2mRp5q4TFwJIyH
Pr6b1xn15csi2Mi9HXL4NHBYMfgYHIXHaqCQNqGoD8ApSTYUrriN9H4jp/89qpl/
HG15xHovnxIRfc8SdKE5meRkAGcgF8Y9UWQ8f82fPoN6w7/fi4QSBEzLaVczSF6i
RPsS1NeaY0LbDFiK77VbmyCU+Jh96Nm7TJ3lv3lLCTCUAMykIXOpTwizoAW3yKi+
8L9W/NM6NFOrSVSwqzJmGp86W/2dyTd5S0WpumVTvk3JHtPSdlXeT+Q9q3e5JLme
CshQM1xsK/L5D04tSp4Dqc4ZUJyP3mUG1N1ovwRtFMJxg6fGAxMQCkPmM4cDk3bX
9khyD+E70qthx1utVlQX0Z7ejdcVqQr67OkkA8UObaTwKmHIXlTniHIY5hRrurmT
ydm9u5groK0TtvYU+FLcxeGIws7AzD8xt13QyQKDfe7mFpFb4JHGtBQaw9pGC5Gc
+ZmjBz0AzTckwdONoKh45NMYS9q0rQHW3E1DpwvdocbCEv9TLwSVKsMGLC2f3KcU
/tVJMzNeZbnrBK9D6acpTXhBzLr5JFWRU7H2K9PBk7wBdP8p/AWOMnOl7hrKriT9
1d6KQ7dDFGJSrKSCDCuFQIjvzbS1O+ufizQMbjtrRN7s9h6B78zy3J9Bw66yOyTX
z4vj3dp5eIaOgmn4+/K/qo9Vul0HzhZcDI2J0/H0QlwXjN9RHVH7FEo+r8rMyd72
zoVcyUz09S6QEXUL4ULMzCXesdZHJxUpvjvHvvNIN7YC2oIRnawTgPXCV2aDTKQM
nd9EaQl3hgPGV+11p1wqVA+DYrjULtBYAdmTt6uTer3QCfWCpf/meTa1spURFov2
ANwb/Ev6m8cCy0mWf4sQUK8xsAqtOE7nyTmS0MF9PFmuOPM+393jkJbOFHRaoDzz
ncvCxKLAlio8cOAnfDZv2q+kwY17fhnmSf+AWAzP547nZg3dPtkH3TmM9lLYv+wl
PZ4liIo6flEGIOlnLHDQERjT/qVeiTcbluLNwG/fAvECQJm6TaaXzNnG5zMzKgPL
yUqydyTCz2gxh/HgiHsHno3jKL7qY/wuxpfn3EzPRmy776TOtuT292dAsJYDLDSf
oty1JVOUKHDbXkD4sSk9H03yRN3HftK1FaUzOpRGMpZxODvCXLC2JssZAv/QOx6c
S3mpBjlNmxNOrWQ36GAUaIMFoHUesWinCHBL0yD2J3jS2X+cjoYv7ttt3Geg5Y94
IvJf8vdydCKfRwkHIamjhvwunsZDtuYZZ8O9hhepfNCCqKgdiPMI/GjXFw+k8JrJ
dcUZWmK3B6vt2R33SR52gBUvo23/mSte0tqc2qyuWBIvQH/OGUMKKxvJgI2zWwPe
DK169j0bK8Y0gvu36v0Z2ph1d0CSKF06MmLbK/pmezFTq3fJwcpuxnTJABumX7Yl
xO3CQVwI9T4CHy6bEsirb5TZsLtAnqWRnbP5PMP1KvBqmOSVfGcVUHteXT/1ifSy
vz+qvVc/D8kmhVyjkK8xK8dRxOp9D1DjIsC7TsIqOFg7c2xik6uKZ1bDJiwh8Tsb
LbuSYDFel7h5cjKhnAwiN+DvFB/RwO3alG0GRtn+GosTUCHnPpMxbphopOe8yyo1
QM6Ckc4zTeQqY1V6ZhsIdhRrT0CE/B9MrK5fReVEQJclQy9Vqkb5udDlM2E3aVbC
c3tWWmZlSEA92hwjZl4qnsZcmvENzi9Bv6bwIQwH4dELceAqBjvWlG4jl7Zq0+xS
8UMh5OuoqpcRB4msESa5knElU7ApnNk6x1Xa+A4WJvT3QkVbBD90hNPnXMSTeNLn
Zz84694CO5CcOnc6cBXzNgFnJy2krl7WPZZGgYdhlcFBmEZ7P615xoIacKcqQRC5
pEodWebROzitLHnKnYlq/nLeeudBc1iNVNU3ryPX1CVDwWYZyEkT0zsBGuejHliI
Eimm4/VIzyos8yAMGL1QyODzimToiusp30Atjg4eFmqdyUASQiqNdBd/ho+9nP0/
v+lIYsBXhM5DvDtO4Vkrfhpgjo0D6Ds9ZVQOkWTmNTRfN+VpwGCa/IR92ZYi3wUr
WFgBdx7hpQFnx0gkt6umAHFZ4WgjgXmIs389pGKKCdfPTM+PF2xE7cungDNOdQUq
IyW+hK9LymEa2Ms7xaMckyKwckW8Vf9PUQWsbYvFn0ShAXgBA3nq043v05ESsBKX
+im6S02IQUAjJcrl++J1w+EaUMnP43URlgbAxOCs9EoCiYSOtSBA8n+2ByoIVRiK
Z5K9gEVtUycY/FE6/HOXm9f31uDRgFNW+6eIVi1lAGttuKRJ4DPHypUamJQ1tUWr
BDysSkpdCAwh7tsfH6FYy/C3RZVqH4AyGF3qfCMp7/kXEEz6YrgEla6vozwBpjTr
IB2n8Vun9Nq2wFYyIfWpcrZ4PUW9UbLsfH/Baa+sU5ldTwfMIr1xvxFxwids2/jK
cjWXZ8Eu/EQbi9d7UnsMZMjL7rJiukf1fQG/2EJZhL1MWzTYdEa++HeZSVqYGoiM
ovfLRab26DuC3lOUCOVjm+ENLoUsa++wgVhFCMoMvVN8TuzmFHb/Uw6RUHcSdX9P
29qoIXx3LfyaLEmAdIxwfH0qUnUbVFQNAL5UjO/atZ6EXyMy2dCkpNZSanZXtd6R
tGiU7ZZ7843nK0hifkTLUEU6cypJc3JnZ3/cp8Xe713PL2GsAto5l+ks4DfWU+kJ
`pragma protect end_protected
