// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:26:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sGGqY9yn9HsaghTS+v27SuLJpXuxioVHvr8jEcFcHkKShw3Xso2fkXUJPEGEj2D7
DGGNdUbDaNG6WSW+9s7OWRuzspKj+qbHMnCW192oyJydRk+5zzoz9vGJMKyWWtuE
YyhZJZq6IqxG3L9p+Kix1Zj2tB0z/tXzUrDy6qDFa+M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 63088)
tQLGKz3JQdGrC9+K3AwmNyBMFz7hGQTPXxjOFdfQEMc3s3bc2ncLSg7QVSc2v3XP
qn1tE3JGBIzMC4Z8ax6TyjQV13+nWtgNmT5L6l/Vms51Wq0VDhV50jL2iIJyMn4k
QELhz9paFhnAqn7rbW0+kwlsU9VfBznKuXALj7CmtiTi3hLsVJPPpAaG6LrRAEQY
r2BUpMMWnrgnxDmgoodhHgN5PwzWpNypG8KNiLmBJIX1irHicap9WeL82h9IbQJz
H1wXDWS0X4D4gF3ZafBdEmmnS1EU3LynuyHD6/+U5mO3nLwQcKyZsVtkXJjf87p4
qUx14brNd1YfnJk/if2h7C4DcpFOXysjOCtGYknqamhvfevuN421WwwiRgABZKUC
Wpl09oudI8MSCi1nvDWzz4HFXeJYR+T98bQVnuM4JrWFhTdg2MJxLmakT08Z50t5
J2aIMxGxSxj7Dpr19MC9WN1ae78yHpP+FCqjiG+4kzadqiXc0ura6CvB7dPE2FjX
IbgCOmIM+XS+k3i1HyS8EKH+5YBgJs0L1Hr5UC9Sioeb55mdmU3+xyqVqmwj5mOp
xMS2Qi7eA4qDxiFRuJYRcv2a8UXBLHF1M1ph+9gI+6XP9T8Jjn/daohtascJcyYW
lKr1ZzivSM3bgN1h4Jm0HuH/pVxfmMlWeCUplZpvmkzsOa/8v0zlYyYs1DplvYPb
GBGUg1ocQWlVQgN/zanWaUe0cCLoGMcmYwJj68pHi4zbfkhYocIEwXcgvrVhlZyI
7o1CVqQ2Qr0+tn9CwC3iBIKC1KDkOLpYuBlaW0Bq3kQfnAscb62vnwzT66SbLP4/
zd9z77NYHDLhekmpV89eiC7GW3hXGHXp3dUCVattLS8K4IGKW/dHESvZVI8zhbiR
+eBQ5poKla/jcCHLkM6bbKUneGAZw9d3j+FAmr5Nm7zlFZf28SnRxXAk4UL+L7R0
XrqJkTfZuj434lOdVJqnTtUZBZCaF88i/Ql86Q0qpIoXJlk7iTB+XCZ3dQ/VgYHo
etsBZ7N08RwcIWDU73mOxcoGkZ+i8NHRiNGPtJiqYZME7xYS+mklawfJNSWRKLOh
CUIdS1gh6xqnsbIsJRGT+F+ovCM8EGpo/KwTjyGoaS/6sRPXwK1b/uM/PK/Vchlp
cgUVzVOJZHM+BaLMoBUpb8hdv9WxPRXPpGQobzbh280QpNcikiwvkR/xM2ZSUbUQ
Uc+OzTjCE7zRlO+FWugUpH9XCx/WGD9fHHs4sAxRcvgdAppw8uqBYPaNGzDWR+w6
3OZjhnrq81hi9bNFnNuNW3QpT17gcQuqULBGLaxqprFSwwCtOt5bsu9tHjBRGX9/
3tocyDdJiHznLRFisaD3ji96JadMRNLSuA0wO6J98JJpyrMzhxDGzuxNJ3a0c/oi
6JbWDPUAV9dwE0Lf3yvcrYyvBCjTurPjtzIz5ZlgvZQgiSPRK2ZUdUlB2Oq3YUmA
LdCbSn3NRt0Txg5fLzG5vdFBBT24yBYBjHVshf3VR9R0lgh7qd6CgyQp0Q8JwG34
UMLNIwJCUCrUzIo4PPKzpQy+pF77whOVuwusttvYEIbQYtzNlXmAvzf/A76cAdF2
d4gQ4WsJd0g2SSsZhF53MLEpcAcL25cta3Rd0nEsgVG6KXiS6wA1CnjVeN0+ml+N
DLQSfA2+Wmd6MMmOCrkq38Z2O7pDcUrsvOoCkQuqDqmWQj2tTwerS5ncgWB45AxP
XbpXxwCk+cH8lQYtiftn1zfhCKipuTKM7WWohngJILffJml9+EBXoqOqk+SEPXq1
/Lu0X5BkixnAVL97cbLDlaWixntIdJ9x11qgMah1qtwHWsD3YX1/RS1Cn94o/Iqp
LM0dJsI8Vp3vy1ooU335n/FG4GEvfjjzXheBv04TjcZpr/pOS8yyJvXomj2ukSsQ
G04K6Zm/uQaRDeF+OB2WXCL6yGOrFI6Sck/AGCJFuzUD4gjoBYzFzimNMNyNeIbX
RHi9Wic70gx5gJmg/LL3VRKWJbUQXTDwM3jYoBSqqQfWgLQi2JTjBNH5uKU0exQG
TTtIhHtDrkSPS1v3a36f3K47WriwOf79uw9H4qlrpt0hwQMm8r8UlFAJejhe4gwz
ge3obPSCV9Xl8KsZG+E8n/p8c65gg/kYmwurs1hQJblhHS+gzbA41/09+FCOuOme
ohpS3qJw1ueDSwly+LaTidhU3host0Wvl/OnIpKTmZgjm6feGm7diq0p3vNTwoXU
C1Nags3SuoGkPRDzjvuwiU6ILAFPZ/AKgMwS0MiSdWuxF5uuHEaLj8IQPAfZCb0x
z0DOvDj8oPmk02rohPw+AUfntmyr45PEPJtZPB5S02UGtGMy7uk81NtOSfh4niPY
/KMkRLy/hZUVuSA4OZond/dpF2+ICyy5xDI9LpjnYNGBR3nkOoxgFtjX7Ga0eEEQ
Z1jnTJ1n9G9yF84iB5AKCbJOdWb1xsaBbwGp2tAtCAAlVqQD2EWgBSgS69wKesUo
zlTGhCEcyZukTtmOIcZjTILoBSpnAX3FwAK0QklyBI2QTrX5y7xQpbDYGTs0jnHN
4uA0obSiWfM56+vk0UpMj1rW3cPJBZn29E/3JjpF/QvIqhdmT15HbCBYeMWlh7OZ
KlqQ9FPFxfZvFmAA8fZkvEmuYsvE8PalGp6KXHDd7cAYlHfYauowlspoqaztTmRh
NNswlvh273z3OnRzKAnYjvaznf2NjcAULo1bDb+YscCgQ88hIoJhPKoUg/zYpN8c
K9ApmsODXi9kOEn7qeaFbftZLWOpI/HqrRZdTuMxk5P4jz2qwrkP8+w8Z2rc4gIL
WkxLLR3wn4aYKfQpM2Sx8UERazL9XqfIJ+YChOywwGXuPEYE15qgbycyigXlo4L1
9HP3j0KlDrZ5fLZ9P00SBg1XTZIu9tBsx61Kj96e5XrbrROwtOB6tnup22CLPXbD
ERHLZnSrwvCfEvqXFX16ULTw3jdAm1xDd6IfuqBZJ+IHXd/PwhfV3ejJSamayb42
8vtU+sfe1RTATxjZb9zmQJR66+OCWJwL4SIsRnnWKgissVPskJuEzM5imGeKxQG4
8aWfHVjXRbQLB/1TSKYKvIYOjyRGU0NfVtn/AJDrYE1BGGpckz8qyG4uqgan400N
z3pcEXFuiX8NtYdaWsXnyRyu20WJhDRwMHWqM3SpuGDfJSmu0N0/PpTnqlzNRMXF
RMwm3LPDF+WlQbKsgTCQR7CXCWssduscgdgjdUKqugCMkdzepXYj9nIeuA5Ys2Nb
0oCc50NpeXxSQwtBGse7FuvKZa1levrfXghMBhMcK6xCeq0M8Tw5fdL8TbQbj+mh
dEc3rs1179b2KPQbZTR1Ip3mYkf4s4vuwPkIbZHzhz8jlrshsdzH/mZRKC0x7esC
K6oVx8DY2y4ebxVLwQ+oOuUp53VG3M9W/zm01Xlm0gSf6tFVbjCbl5bqPH4+ZBWv
Aod7klWqDpi1PUslUMnBnvMF+BPbsrtnTtFsiSppB8ccySkLDvvb9v1K7Kvj5Sp4
jD8He4+t1NWtRiWvLUWc2QVyAWf3MtpUcZQRbhJrpiqrtOBoyDdMtQ3EFsRN0qGb
1A9parBWfhBPNo3YGfO2QKokmB5svMTd8w9FKKz1Q0g+Ue7jDhXntVkHDOB3/h1b
9YzXKj9Zkb8ROZo7EcY8ZHE44C4TY7JfGVZo8lORPn0yyut2jlnNshS8zujgCHwT
hIHrryXJNOJUIitHZQO7DYWiVi+mIIZnlc+vnpzOT96JVfE6BgL9/M8aAFFRR1CT
KG+W4IM4l3qwSABbD0wiJwfEV6lgvpYaY5MisqAWoELbuNvtoIgG27E0mzuO/2qQ
9Da0ATFIL5Du4MznERWJyFF1GCix03DGEiQjFfoggnlHJfOEQHxwJhi/11pfbQHp
3xIVKLn4ykudhZX8Rnlv7RFWq+LydrmodFojoVpeo1rMHoLm5wuBEiZ+Yt4/XbOt
42czuvUZIrBJTJoVaHqtyQNh/Cc5EqUfwuUlYzfzArC02LEzRK2UVuPHJTgd4vq7
6c4yr/QNWi1KM6YaP8LJ+BNh+EtwePG4oz0O20/wZsRQ5C5DNKsrtIb6b6WhTYcp
YASfjOkIYNBqsUepVxVPoLmf/c5YJW4y7/CNxUwVqwmNCkHObboh7rFzDI+DgP9H
vvikEakZM+256zgoT5PN/hZW+cordRND/b4BkAj8wZGdtuHeDZpsK2krF/sAYfUn
ASuah77JH1rXdC8s5J7kxEIb9Mjvdel4Y2iT2oHSVdd/Jo9hDcsmwLciA0hMkWPS
+n9q6vfDexcG4mvfuhQk5bdWkDAgViivHl6g74Epp7gxQz94LK4mYYdR8W9TACMS
+p4tGgMQrKGWB+WllVbzI1edMwHm27BjFFR7r+R2+IwWHp5nD5PlImTqLV6oz4ZG
f0FsRd/1x3MwrR5YXsQnqsrYAqgFxApd7n7qLrViHR/KKGirw+wfstuthk0hUshq
AN/Ius3gXNRmMlwsqTXsymgGc9Sw9Op/0Voy/WlNo7sWisi4pBqbIrDAF+shDolk
Xi/eeIHmIKkRPJoIFV6CWi2VF1EemJVGtD/QwjAHLRtLoqcqrorsd+QgN64a0e14
Moc9cqYkZxRuUsT7U3Tgbb6s2Wclb4zvHYAyn5pLx/BLTxlgOpZ37ren4Z9nFrdi
Qz0KOrCc1EPijX2cHIPETc3ayK67qvPSI9rh/GtffTHpF4dczOvczAueYhNt2mRE
3ynPSBXHlbeL2I+PleNatHVhmoCsm81jbA5WIhbik+iFYsMfcLfYUgiptVbBCvXN
FsBwBqhlNtnyjiscGLSYfylhozlZv1uOLkrk39i018YR2qT2+fnAsMSo5TSfAkAb
Da8HdPdgDB7p2+5rGEguv4IjIj3M2+AiUDR37DjcfHSTidDSWdp1ViSPEKzoqPXX
LjndQIsH+Rf3B5wcdd593hIrRW67vmGmR8A6VDeyHAZV74NvKUbw5TqpyArN6Khi
xh9djBXK+ndHu/JbWaVgwnUlsbtFpeEId2fPi1AhAbsnX6dsDUs99RV4sv+665jL
UNt2EnRsgFBDmqdF+0T2JUBQwgRuLlF4vou1g20+ax/5T6dPekiSda8IDBMwavOU
bmodvOJXYqcm6u9HBSUWQq6B7ajRCWEPcncDjBnDI4X+HMb5Avz7nh2S1cIFWiI9
BU03j8MaeCkf8BtmvlEznJ6BvE8cS3KQSYSFuTBPM08GQVdbaD9/nLnqeO2umgXe
4Nz4Yiy3ec7+3QNOGHdT03LrnDMyp7zg7CT8Z/U/PhsDW4Umb2Z6yDLQn9KpISzs
qtal1+UP0OxV6IBhXYPYI4crQrXYv4BOxo9Lscr+o+sN3t/OC5G1VWxvzasNgnq3
BgykoKs4DYijjTAoTWEiwsDt6SxsGk0bCq1FTRFDpvvLYjD7SpAEcbrPWmyZBKLA
cP+D7YI+tqibT4fCDE4LOsbxs03QVxdeK76pmn2bBdTf8enU/NxxWVYH8lWRPqfZ
TEdNxJHYy52BdLIITApVbpwdx77uVkMvcm4BhW9GvW10HMkuGyK0IbkIqWBYNazm
xbVNMRcqdZJWhCRm1d4S2ZC4voPAODbaektC6bcH8Twe66t2vFWRdF1wyUZbAuDw
+TvCfIN2G0e/1QnM9H5InZW9GqrQLKnGHlNUK6Cfmg5Ifa2KDpFJ95yfmWByAbdK
yOSxRF+kItfKfC5Bflgi7z/zp0Sq53EUS2lcyRzLqhaXNrzyrwLCsrlS54QwesRQ
NtMmjYINDsdLR8OlTbdRAPx5HAfaRPs9pgqnmYBZolOTRiopjTpTBquLdwbLe/4a
0N4dqmYNBYQZ5U01iakLQsNFO7FegK664a+H1Ft+H0oyiT9Kc8Bg+OZ4hdOF5uD2
K28GqSuEK9mQIDhqOR/Dq20AhU1cn5NGwzU1B5PtZbU79AahDUAyQ2Zwvhfl2Izu
D3IZk6OCaFvN8UMWXyhM5H7xTR4B71c5OM5C6g9FF9AwVShXAY/8Yq3O3xGNgL8v
3VlMHZYyRLEKYzHF7/DRjU41YnJfclRPnEUUVpWOr+6YjKlX/BaT331mnlLhAlHC
a7QG2NQLgWTI/Zw/duYu56+HJ9vu1MUblsQVxcvNVu9SkHOqD4+Z21BISd/3p20v
JEQ3XeGS7QVknDB5Gw/wH5lyWqd3/1vcLKfsZM8Siccn7rXFcI/0hUqhiHVbUoqX
3AgyHNRA8rJIJE/E1/TkMzdDZhi76vznl+ahM+KV3ncFMWd7AH2BYHN+x8Y4t47J
uMJrhDinMcC8WIkrx1byqbnElp8yhAhVrE12qzV8QmPMav3iY3jzqfh7keh7rJBo
qZtvPGt9xlPOb59Y0pTQR9cpJZWy08pqMoWAetgmTQhPaMr0NSq0L/0+ltPq+ln/
fJbSsprBhgJu+9KTF3+oDzk0TsG7+273s1CL1nuhrX5tfzdD4yWHaeFf0sTydHDq
GosH0rTGcp1Db3NcqLNepIAldAgujj7sg7r81PY76Yj9+83Bhy7B2UzpmXi5iz3c
/umm4AvEBqoGtlWTPciTN9a9dKdbuUJscUoWHsfzB6UY/qU/GPgV2l4qUV/Jua++
D+KP57ZMTFaRnGMnHJ+ugBMm5BwRQu1EvyU86EHM1nQva6Q6Kic9OsYES3aR+e/y
0YW/S82QLCMFyCKGOraVqh+bMLMjqHJADRY6hP4LH3bhktx0PCVuE9ofLZ4eIuAX
h8HLohs3DsPsIWQ9dqkCFhJcRM33iWFNupCTHUlnLpQhbKPVjVwaeXtaKuz+nPXW
MMkrb9dhJYYSVjbWcNU8Q6SDtcT7VpDYvxA5XzdtufrF1jbMSX9Un+av9AF4Oe2V
lgjj5Pv1j+C8lVrWw/Q0HODF0pAcQ+ZrXd/gBM+leObqUOyDfIrhROycUHOX4BxL
qUhUXATRoO9Nd1ssCYIQk+YwZh4dGnIviYFJyKR2hFGyGOAF3IwS2aTLrnVlHURA
GIxqI90/sApB9+4wWgRK8axeVqvgwz9o5r4GGzZJEUfzmc4Vg52y1rjgPjtn9uNL
PoWuPKl+25iqtfKGf43XKSyo49fT8YZvk3QRSlan3CW/lp4+UJfPbLNXPG46a6Cp
Cm4cpI7ejiqVCKwSd7xt7eCFt2ZZ+clSCclYx2lKHgNCfpjxJr8s+jax7HTbj4iq
Hxx+30fcsUxaU2bzbSFUkNfYiJvz45yBf0UcYsrcoMEgxGnNexJ/7CzQbpEOeHjG
NQlGCQsb1VBlE7pwfAqvB7WDxruKVF1ltODCgP4OZ7C+pnFVA1XrzXFo27MM0CaI
s8haMBHbuV4jm/fEkaKoj+jL5truq+J5AI4xOCzUn2J6dsynLdHgiOMU26hVHCLG
CST04zjddCbbYXH3DKkP4X/qnOCgAJyzCT6cA/tXdgFRHjrlvaIlKecWIxCA/3Ob
B4nc6wqOI1zBJMx5KYr1IXyuKrpV7EjIctOIPJLrsnP9zCzHDXxqTNotK/bItp3N
pS7PrxOR5bOl1F28yCj+Lz4syNYANLcsJAmjBdaOsN27FkWo01MFcyXRznWXU1Jt
nwMxrm/mg9dCL/AlQy/5U0azMeoEou0SOoOuEzBo/gzuwZOmdxYylvaHleTQR6Gj
rfsc2qwYDmczApofno0LarVglMmEUYFxirg4MOb5zi5QYgzPrunRF0gncftgp3EH
hQZmjeeBeUciw0WhnaJPiYL98p7J3nGoR+OysgJuwRjVq4dh+uNuGC1t9CMPhriL
SvQx7kijLiPs9qdSdvRemVd+T+b1GOYsmcasiCXYkLtIADiVgBwSnng/0UDEL+iD
1D7vc+VPabhYLk6IVoS+kWvHBRNSeaOmlxxE7JQ4yzzlhWgTTSZjsjsXuo5hpBDy
4bMWmRK8t2G0R3Ghg+CgTRNiU6ipA0SVtKImbgzYfxsftiX0nU1C4tX0pg1Zyl0y
LOQHwk3QTGszjiwBd2NEx1ZjwGn7sn/HKakwdUxhVsMEsyzmDmmmQIqrR7L60koc
47DuCgsrWsY/D41f5D/IqdnSO+fRB+6HIb+QhxzTWAFZGRoN3dCQ+ALR7Bilg/NW
8SWDxypjR/hENS5LDrpuLDPZ4hWx5e/ldMzfcc+NYKE8WTJYnMcg5VxScVqx4QOu
JLJDRi6jXGPeScUukOoN2KLHayiEjabOFYxFH+64EYI1/4H5g9d+6a+BAxYAW+ZO
sWtl2uLEPhNG1mNjylhPFtKZMHVamaob47ShAgST3kHwBQh0isUpZFni+Oo535/K
2Nzs5f9PGyWaICXfR6jgWKWBoNxIUukukNmTwKaZ2yISE0kCORLzQoz0/cFCZZoS
eh67y1CCX30we2TKy2xU3m48+RoBP6G5Qg+2vlkYMD4K401UQ1gHmQYQJzXlJiOU
MVgMZmP+X0fHJj/jcJJ9TvBrbH4vplaK3LeJXIyzS63O8Oo+P/QrpfjphxL2GN8x
9Qs9PVoZly6ezJDmMAJAivtL8NZmfHKx2WTP860f+p9GpjUGUVEEAoyiFqo42fkl
RpS+ZT5RIXJDANp8OTiZmHUp+z/2tkTu0awSG927ztRifs5aIxpsiaM1HEZN/ZI0
MdYf9jPdTzmjma7tWCX2VOoUQQ3N+nwO6vDUH1GSjVTgHyMokJEWwIf1YfqIfx0j
mmuiridZgobiO6TFMnXyp2gtBMgiQaZK4qY4zg704h3NLM/7o9rItSNzOVu/4Gsd
wRt3OG9l0xzVIomyRceqF79PRYBZv72MqWHVP7laEwAMNmDcQOLbaH2cLZ/k/0mI
0jqFqAvOoRENRsk2PLPUZcisAlunj/maJZ2OCJdQRJwOfdGhbAnD9Vi1/2rLnScY
ieJHksvVNDv7//XpsLdcrcZscVOXkTVf7bV/Hj1PHDQKS5AJ3cUN6++mSTlF8B7t
b6KiVzdfjpSMhbjS6quHB0N6af+eBNSXBnsA5udHTcsVDeO7JCbEGxh/vr2Cgpy1
N/KVEUbJy+6Gs+ZZzX84S+Sj6DLoxR2UNZY9dchxhccc9eTVQ/5dzEncKAHSX8Kg
WlwJaXLBiDxjNWaSJOpVjSnXtgN8xiFAQKL23jivME23qws7WKXSxeFjSaDqw+Un
SS5INANW7Qq8Mfvf4Q3EX+I2XkWNBX2OFE8VczFdRL05UNZKAmmyuT9iBZQN0Evt
ZTEZC5bQxqEErzWHuqhUCKHiYSPmROocteN/Wujz6hX+am3NndFV0IrA7F9+RABQ
YnUKke9OgQkr/8ecMuj7639bce41gu0xYZh1n5Sl+vWgPqXuECAAO5UASxjtd6ck
LXa8a053RL1rdRbLrWUjk9U2EwCivNOA7q26qSryo8jm49pzCbae4NOmxMnMruoL
41ifZ2gcVU3ylVT0TwicRXbBkw4DKQBgDXoZhTPvtHPBDVPOB4F/YpMThNJ8eH6B
2ucHkQfasep6J8Mbv1/X+0PAiss1IoFO6OrfgkSkhk/WhGmMO64rfR12ezm+YO76
Ru8azIs3Hhe4SXvt7/BMDzpmhkqD6q1PzgEQcATUpXz1w1GpIY+JFTeHGRy2vM+A
k8+Lhj5mMVmoawur1YJ+jEW5Z5ZB2HicSmsdH9ab+fBcNp7IHbWjDX6zdt/anf47
QS/imGCqGGJk0Q9aqc/b5kILiQWUqmttXmNqJA9QMg4Q4z2nJuVwkooNz0QTay4g
P+SXwJJke1pXiT0tw3dF42NolbYvX8le3SD+yUYAOeUEmiwikW+++E8rNQLfQGpJ
bc4pm0RvhcG0b4W5ND2c3URbrAd0U6rA9bcY4AdcqA8qpVkSdu0hLwe79y7+1xt1
gdH3BMTmGN+0txU6Ho6/g44ZUrb7zvJcOjIi6ssDjBV1raqosSAzY0Vz3ZP00koZ
e8RnzivDvX7DzGxiHAaF0JgJj+tJsXUV2id1xOcpQFcRnwTlMMBmasip1BSITyYH
zowdbPxzPLA+ifQ5DLGnxLel754R3CyJWYKjvU9zjBhjmBtXgies9Zkf39HToU73
/+kvbxZ1IeCOT3z0UmlvHChGl7x5m6eujAb7TdrrXTL5mvLXPBR1H71LZPNmfMDO
C8hrtBDY4gsiEEkzDGPUnkcoavwW0YKRhFXpQcyfSp8bsSTRPvixdCskMrBoIItY
wNrxsolTk8l3bc4MXD5aTOkqEQK73tIElw4gpa3YXjNp2QOhQHR8C2viiXj1D8Id
+fNexKNE/xmbo1V60lT8yUcvR+3B2GzzvQRzlDrnPjo9wEFfOq9mixGxgEF4Sxgq
duEQb15j7I9kGgA/1GMCp1uAdyuJAby/N5inlcAQ6gdFOmYH+g61tBWlVOlOacwT
UTZGRJT2KNqCI/JuhpBF8lQIDaIG4ZKt6Gyu3P2v8FESBvH+VhDx9cGWIkL6nLqV
8SUijDfgTmGzQ97MHruvuqDHjvM4a4kNrW9tT0oj27jhaNnshAY+u2HGxWS7flJ0
PYLDHDmtAuJa5JPIrMdaZ8pD+itaQA4lrNGcoHHLuWCRWuSUSJ3E/rzyzBxCtVCg
VfkK9QFjDnP70MJh2SxM9H2L5aKthCHuZ6XTNwrF1kurKbxNgkwWqT8LUqe1wtW5
I/lbjFSu2mFQ2ocMISDtfEEZWOCmiMiPGJD3XOUpthTpy4zlnSLnREF/B/wBDxfy
t7dmbIC9zCdDk8lBCyLCYZ+rP+DEsY+Mn1XSanY5KCCdJnUANe2twFVF9s6Vu2Cu
cR/uko16r7FSGb6yHLYEqLq24DbQbD3ZNsuA03TMSJiWJxGUpVdESOLC1CFprVGF
LGQ7qJqUHoI4EbnI0QNNKr1GYB75ibGhf/7824i69rsJHNBejLi+T+WcfEz5hlAI
7nup4lM5gWw2SL6BwGD8w73UMEzgt7XLqY7B/uCtPRLX14nCYhqup4Ri5UvFSmxi
GjOA33O+WkFK70UB95JhLiTj1L7K4e8y7Or7MwpQ0ggSQIvDOEdAu88gV+iO8J06
wlHRlnPbU3Sk2JlZTiGBlXiVTrGcQfCgxYsX2rT2bRGYIQSIyy+dtUpxLw1Hh9yD
/2cFyJhT7esLm1FuPKxm9zNhK6puj0CTDgeSrWoJbkruBVGZ3xv6sqHsJBAXv/CY
jrURlcZGPJjJ3clr3GmAHY/mPtyvBSTuA7jGsy5f3/DVdSHHEDsHnVldGa/50LY8
paitTaSgPvcIXKNZsMIQsc42sj5XzFXS6GyVHQPtw2W70NG/bAGdr2M/TNovXGyC
p9FxpnDlKAJRmvYxFaD8ic023WcSDTuSNK58NFL43fVwvUUN7gaohBE9Os+QhgZ3
B6u0jbvzecA6rNYOxVdWWy4yZYJ00a9d4x6R8e1pU5bF1aahuL1/lOhq94pWLcDh
JcoAobmrX92/RB6+7UzZVH5DhvSfFV0uGjuXve84tyyppZiX+Il4zHOYpJ3NDujW
lPsz6WXdCi0hMkwfnV5Vk4SoW+gJR88V1bNJRxAHVLLfDJBFLtSpqzhhlLz2q4sh
2mGcnC36dVdvuEAP678dfbs9bcKlrCEPbo9mc237oWyeSlS0KIs7aHMZLN3SBkcN
eH7/qnKEhY8aMaqjUQhfOIf0/e+lnIwUAVlgBV9HsGlNnl2GbYI+u2AAL7vbgGM9
W5O/GyX2qMjZ7Av2xwiWe13IF70yZId+/SGUETZoChsQ5R0uDJ2j1IIjHtero6Ru
YnaRc6YTqc8QiKIdJeDHCMM4M2Xmg5CC9bJcLOAWbJGDTIUiHuLTIcYsYVKpjRvl
Mec4rOU8Eb/53JbX8JcDGU4YE1WTNpWP2v8TEGtgZEkvZHVmnPVs2EJwLm4zxN49
cmWUYHzA5kxMjD7F7iwIlxE7Mpl24aF6A+L0CGFh7CTGouDdZSqeQfnj1//0OLrS
23SahLLYBYvqUF4J9yhvsupTaRKXpvkUgwttWJ4pYoWHIJBLs5KLaT906kcLQOJ2
r4UAil3CLdJoL9/C1qJJMS8iNxw+vivLqiRFxXJZQGysQlPAnAbaZ3wV5A9HzkcE
9INybFgMd2XrDacCav17vyu3OSdBCzmoqS22R1vYLe4Mpvxnj/I34CqCF6QeDkwd
1bHGU+DjgDOgQFGBJQ+14ydSHFNVaTK7KMk1XzK+qjvoCNj19HSwOqMzJj+INRTi
1bk4luSzmp9CNR3gUHjHPY2sar6X0gqlDnmNmpNveyvcR+qdzEBTC6J19wzpwQFU
HcUf6Mx/OG1u2iuWTCdUrEJHTc37ZFNwmy6X3CHcKZcl5YjgCNMnxMvv59NIkT2g
tL5i5+fxLUJey3/anWK1xz1/LBWTqPnVLq9Kt8N0eZQd6I/qaVAsjFRm8nOGk4Pn
FZwLpSEmejBT3tU9gGuFDZkapEDuOGUlD3naQEYRmKLURa1zK2eHK/My3LoZcaBb
USpPF9z66LkH+OrROAmGFvLKHgKm2v2Y/iy7ul5qwh4KLjXtCtopyXRRHodYuh3b
Ij8oqZqbU4gVV4O2IlZtepOZN0a5D1XcARimUJzdQtReLkPTXWja+k+zpCRMrgBv
lPiOP2DfDycpWVY2X4EUrzVGVzAeGg8ybejyRIIIHq6z+xWSSfdEF5/nFXGI3vo5
iRFuBuWGPu0MW8n6m181uwRBxIrRYpVpA0a9vtC4rItNb7UpMeAEXnhy96xd0aw/
dsYkp+IfmcBV+zpkgbil+NmFM/w2cCpw8rQs1fh6lOE+4ioS/vjQVJ4+xUm9Bn6Y
FGTHU8aVdAn5oRVd+RMgzYCp3aAv1yY/nM/azH9ZZ4i7O3ClpReIOk2S/KA0poq6
+zJ5BwQaHDSi172TP5LfmfhpnljdMuywOCgSEwhqxi++BnbO5N5hracDyd5KDIM1
JqD03gz2L/iiupiFyrfy9LuqoxmEqXlikJoxwgD/zl4n/D2pxO1ae9hbLJ0bUGSF
Bn5ijCIUMVFFC23QHn/jctdmwVVYeb0T2YRvK7bmxwj5Ux666Jml1ybnVzvZvyUe
WsCfSbw/sMZ5Rtvu/eX4X6zfCCIzqLtMWy+3XQxMRhRD3C7ZhWly/foKQe5aOXKH
2Qjo2/lNA1CrblpS1UOtYhyKvEZIzt3MQM/x2fUK/OF4F9O85iYCO/IpP0SRmRfC
ifiwS9LFfLQb8ly8gWIOrdaIb37ZpeCPqDYRLrIA2mS3rH1apRZFW5DEYUCydWle
LOz5dP4IhoR7sJhyTYLaJNUiwTj61l0PXDGAOvuVsrYn3lqbUTMsfcaNUnHB5qMU
i4gbKe31GKb77iemTstGfl+81ibQvuCWZxH7kML8FPS4oXX0vmjbyR5ruTmIC2XW
s/91Dj/Rg9stcMHQm5pK8mQrh8byM/xJOGs18paZsByjq3xE8FKtZHxYWPnrwPD2
s7fYKTJg9o/UiBVWuT3qpqrpUQH0SJL+/n9FA1Tj2MW0nE9uByleuSQ0EQ9P+UOr
iZpUsZumrNjl+qA5mR+ZLzXkbzu0OhRJ6MHoDcuqiTUkKQsVUWVBEdNm3b5Y+4fC
Gz2VvhrwJNulvY+6sfCig108r0bLkcKRBpNwjz8BUaSZx1Bt2tBedCMY7TbvogwM
tk/33sAUrR9YvUVIuvx0eot6NWTqH38aOvSoelpM6CbVXeO5fQLVyh/b0s8OVXcM
kDfsc+XQEVSXaV5J1bqJrNkkacVgntLCxUBYpLnfpLOdJ9b1+5g81Il7ruju+1oG
Vo34BwdZI+zu36KGrz+E9vc+FMYvlceRFKa6SduDLiPza6vJdxcCE8pXV5HnlGcq
Zm2ZjIt21Hvdj0qJb3dBrmcNIFKDgQb2jOXKH84pDIhGeARDykmALXyLIoWZiq73
juJNIBKJEvbQDkJLmzB8wK79zRegUiJublWNO7QGkXtNpsqceS/5ky/uA6y/VZ1D
1QORaMI+s2vhtHMs5wsnd6X4Npxt9qaBYUzSI5E70LFKyPX3qIZyMzFXu9vU/AQe
t3NVbzBpfxs5gC6f+G54b4BindF1GUGDQkeVqrL77/8js4fX65dLLtXMJuA+afHW
JCsy5Wbcar8x74ry7G1hEy3fRKCdMVen1TL6m3kmQjtuAKpDVlzYhFeaJglBdWv7
/ONWV7qaEejmF6KIPiaApzlgypUIrB8KXs5mUr0+px0bPB8TT0Enj3OVtOMU76l3
jNZnV8jqh0+i7r7FbLPNZEz7B8FriA9klhwoQa5OSyGvna+yzYir4xxq03/+u9dS
XaqJyFPHuzvwjCW/9nyRA95ntg0Q+46HqRBDSekYWAYp0s0N9sUo/58aazo4fzNg
hduyBzNVzsyc5T4I0HxBiOF8ieTc/8QflA/NsRHj8/HkcZVYhODKXyJmJRqSg1/7
OD3Gr07kuB6y4OiPHPRcyrbVJxO5eMnQWDrxCl1+hzzXh749XugvR6JvxJhMgAcI
lzyyPVTDKW6VYO8ECGxCJioV8tQPFwxxvx4j9bVmmhLYHbXbmBLeMCtLSH+f2RgX
lwTjKUxB/bnjtXGA6XTkGxtvktSXoUxwxu3jKV5idP378k7NUai7rHt3NJIRvtu8
YLdaUWB6kOqLIBULszzEcg436OP3OW7E28ZNlBoJafhV5s9qAzuKd97BsveFD4PY
shzVdQl7b2Pl4Xjl/Dj+tJTr6LEQQkuLyp6aPZBvgVIRhH57+Sw0PQ6jKY7WcDRP
PzWifPrRI78UY+c0CMrMAHRXRlBp7ZtbGW3nL1bpf+5FqQopNHrrPxBmmJ7fZw9B
KSE5vm9yvraPwAeyAICnKRLhaESUZtn4Ao2Oalo9wEGZFD+aribXfXBdkn9l9L6A
+5YpOXzCPhQrv47ALPwP7KkWIMyzN4D0/0PgLVQkTtwZIQq5rWjFMG0a72yXVQs/
9iCFPr5Tu48voE7qOcAYCayteFUvq/c9ivfrgQ4SYezKuyNncc914iDsi/gysRMV
nOYe+3CKLp0XqTVetrhAkmuU5Vq5TQP0JPrfCqZcfTxdgK65RsXyNkpr+uzLTBlM
RLGLInVWW5kytHQsRkGjKnxii9k/6DbS95NF3rrlvdyt3XxFDpfMGnAvbPltW1sE
xGG9dlWMW6D8L6j63JxX2niyTg7pBNtsSPLn/mPVQDHts7A03WONkZEBnM8m3g94
WuZw3TAjMzKz5h5LRl53FeN+82Vb5pkmPBuYPbvR5vyj/fmpBH8Kqp+XTn4gJLYa
yOUZ981OSa/K94WxRrhJCFK3wQU+eOKhqR3tUoRSEBf5u/8NUmZYE6XfcKyttm1V
Sl9DKk28NSN/qCRtLjxWaOT2lfGHKOGLcAlzHqF/hbHbcCteOeSjz++/XqNPyfzW
rH8bKQnm+87zfw4be9ljtAMfHV6+EbVHTJo6/Ci61mFtmMF8nGq/MUeyhph4lMan
AIHC39p/TWy99EoU2z/X3En8uKmgtOBoX5otynSCfwlL4s3GKFsY8K/znxGSem4i
7k0Ny04qrTJ1glg74D4RWYMAP/50RS9HeXWC6jwPcJfluQv4OuW+wKWfupSUtOy5
Xg30xco90ZjhreVOCCVEaw/boN8WuPjvpyrxKufpziT0VrMKnv0tYv6aZz5zKV91
OrgPLbe9YUyiZe4h8AFNRzzO+u0HMc4ezmoJVlreHAmoFaoCp33y/xSocVxCGryV
TQIFyehmgb6iqDXGAsW+s6rEpj6CDQaSm7w5aGxpO7mV964TpRrDTTYakCKdx8Vj
oEofFbG5uzER4Tm0Au4guNr+jABCUgFt2aDIy6glNUxtK/Ro4woXs+qG71lQBCuJ
Ks/X70nC4nDi1uVpqUseHb+MImbHNmbniGY0+fo9dmcRQQ5aUpZKJ53fL5Co/NwU
agmmShs29igQh7bm8mJzNBXH7E8Losv/+dSpUM0jaUk5vijP9AROKdi7+01e2cCz
3QjDUzP65hC3P7w25Xf00jCLsk4OzKTL2CjPvqtkfrpVI0fQG+zqvqG4f6T2moCP
idKcP8sEjFjyviZARwx9orlCG925qddh0ddjTNvZ/PAzeWdMG/c4xJAugBRRiOHg
rM3q8IsDsljpXILpXrgseSqgoK/eeVsEjUk6IVSUX5VJtSeNhjJ7qA2vHEOnWmKm
WI2AX+6VGBdKMv8iR9lrcjYoxbyNY748fOMK2YjCeAibG5CKqEULQX1NM302/Qcl
L6wrPXpNK2vjAxMcXIHH2Z12CokUKD1B58wpPeA0CQt/HS4S81j+bl5QYV8YUOub
zUiFkXw73CA9XnFYUUK5IKYqrRZcHTmpuSfbevu/uAXk/dI+RTV3Fx/m+XY40ZGF
jorzcfwlIbEqBzO4PZHkTXozMN5jGy/xWcbcWn/FoH9EJ2iLn9NTKv9eKN2BqLBP
gUFcZY4y79SxqeOuAzUbsk9ACZwRjsXsSRQ8lnlPMGvWtOGOjpAwHYYuh11I5GBT
H/7bo7RNYEliXjsUypy2uUr9NqyubBABLm5PyBBHLZLHcNMRVul9ruu+hiayrAG/
miVzrlGVnuRp10e8a9pyvkVAH0LW85S3vtAtepEbND5gYfAb/AI1M1tNNZdQNDrz
p+BCs/+KDRO1GXYeVpcdUoiISYXSpeq+VWyvrq8pVvmU6Vph/aeVdPcm8M/eZ3be
goOqPQmRbrT+30kwiHrbDJsZLBCpWqSpr6IrPGvpnaZ1usbqp3v01Snwm+uskuOG
lNSFREDFF38dNaElQnk2WgdZG0kZ533GF/B4d4CNibePm92YVmfRI08A+AkRJal6
j5oWGx4nin4Qft9ri8LrKup467If8VjSW3BMDWd6SxT6eeHYcUseLrrPuiohDaJl
4In4ndX+V9VVh0WcmHwN3Onkc/+N56FfZCX1NbpFxo7EfGN3IquT4/ZTaeUBgUvy
CEbzTi47q/bmPoUftNJeB0LYHBsmOSsU2j74NEqnQvnpRR7yPY+IdxDqIpjG4/Tz
asQmsLgSMdz/wR+4abI4P/pvgQmFRReqQ2Eg/ca10s3VZOooMWjlhCJYkTBMIt+t
O164xhVODxPysHVjKnefgujkL46anHARyxQ5h8RbXszZUVsKV62vgAsxM3nUga2V
tVI2ehchHAoo/9PH8PQm24Bmu66iqG8m+drJYhwVd4ACw8Iw41kgsN+qma9UeuA6
8awa1mCIVfcdIGlhd2bWWpaNZ9bVeHgPv+ApZxGRUFLRJNdtazAjtv7mlmiATqeH
eYpcvwxwsp3a9KntnGNeLOg6MSMrqwSqFs//JyV6r80HemWGplp28Aw8EyDMZ0Lu
81kjsdulb4hG3c5vL+DcSkzmZZkspkQqMEvRREUGzup9u2o4eEzB4yqroGFZLJmP
tEuJTjAXHWTzaM9VMorhz0GuoNLPftpaijJJ4upW+bfCH//Setk5PPLJLBOKBy2e
fM/Lbj6d2LJMmq6aExqbhXUHG86eFwSR+DVIjt90hdWb+pnr9/Q30O0+loNjyBj0
Utk9wjsuJlplCEGFdmsNk1Ef4Cerye506++P/w57TyQJ4IyHfme0XVNsULn6yZb3
7qrQ6R0yHFDchEDiFlolCuMTgPF+Bo1zdF0hhq+bVOARP0DORuRQ6Cu2dCOemWtY
VNG2oSUD6SI8/7qgg60HId2au5Bg73cN6GX3ve7gvScAHf1oFer6+1MZVJ9Q26+N
9ZU3Nm0cGKOPgpjzu5SRoAZHy/zsAc59SbJS0Lga+qzHpaAmXjg/g+fHvWjfqTfe
aJxx77JDbwOdp/YGcSiTWPs6gYACrl0eui50LKlKejKC/lGW5Wee1YFzavlZ1ZnL
HqVHK4ynnyAX2lq0SQpMRDnv++y9m4WIOVP9gzOZ0VQ6XD/05pasKzwcqFlwrINm
gvZ4mria0R57FLN1IBBUM5DYwi1rhLyD/YYRbNwF0pGMTxzp//sBqhcpMfIODmz0
O9lyrSNsPKjcsIDGag6ALTYlVafELnei2+THwusF7nVFBgzcSohwlguQGYCZjR6X
7v+nYxdSRgMGNArnyseJflZhRE9MR72RUc8Z8MVbK2S/w4RYM+sBtBpCld6WtAo4
morN7XVlrvbNo7fMticnuuRjdgTFdDcY4YFV5o+SgI+C9NvGVQjpF0X0wr4VW7mc
Ak9I2mS2vLhuZpVrmcrg5SdiCrRzUYTxh05PbcZ+DKkTMiOigtwfxRJpcdRlMrZW
aRFe+nzcN+/1NMFXyok+dANepspE75GlkRCWLrd6A9XJwh/iTluJgfIhOz8gBd4X
kYhU646kwJ/+tDpfHrFJZLS6ZV2xSoQUkPIqwNXltrmgqunr3RWsYc2TT4qEHgy1
xtiCNXBTJu03fxrjAiN601LYp5kea8f2yCmvo4pxDY51EPowRWSTph4ySO9Nwdps
PmxeBa2T532qjUuAvn3Cg0aV705VM82sNPOMqzRAD1OSe/Yb8N0+Ktr2uneu3Is1
3BS9kjB+XOKCdzowq/QAkbv8niFaWD5b+L33ThW2mWtc5Cmutmz4teBV3GYErsBz
w6QA5+VgXP5+bNYGvLe0SGxDxfr1ALW5pgQRJr5nyxv/7LsjowVdyZw4rRQwXZp/
KE+jdrssyoLvToZZisX99cQp3njT0Jhb7YJxBYy9CaTQJY5KwVt+e5qfBO5ngl+6
FSruWGxdp2vFOTM+N36K3fruEVkj03XQNoV4lg9Kjk8djBE7qJxFJCoKMQfCLYrr
4pMgwAObkK8yytePGGLhJFE2iaUphUTu5700pKBVkPq/THWLT9SwFcRfiIEoipMZ
VSXVOz1DXAtowuTfRUp7PzxbuvN2Mj8De5/oFAe7sfleCBVOLcLbvbdjmgRnQrZo
1YkN+Tfo1cPeeC7T6mSSmZhqHpIh1MRP2JWml28JQS6j99ub1HqO62XOvUG+UrHd
83hjDE5D2BhrencZt6gxcD8ZJoJ3/f99y6U0Q3h4LZz2sWyajchfic3E8meh8att
K9N7far8OHGUWK3lovb/WtAw7eX0dd8CKy5LSwbBpcbeTBugFWs72W3/XOlZeqmE
jAN+Cp9n2GQGxhxiKVYWPDTRVho+1GpxhRLBSxWIFkL40zTs+fQ9Eb8I98uszv29
44oqGJfA8grPNLOPEHx798EwCkIBcU7KWg7tSeB9XXVM6rTg0cEW4SJklXyo/hlu
Y1WvgoJtn4O6OYN45eZBXv31mNhm90X9HlrWhkOQh26ldTol9c7y83l0pO+XyJLo
blnCXamQMtxUzRFQ2swhorrLdk1R8I5E/SAJkOG1iSLwMYzVkj/QGOgreueme30f
bi/b2Y4Tvxdw/5kmnz04UFND+hztyPh8RO09W4L7GPc6ENmTX/+yr9dv+JcDzYud
EHhbQpJ8fjvBSaydCcGJLPo0+4cStetSR5Ccj+6YXG0HEBpMOqUO1bzbp8ZVPygY
HnTCnMrArsck8z6wTPJhB2TvR4ea7EaHQ2gdmSZcqW9DJQIWj/fyET+oGgKJ/CX6
OJvPEKzx52fzzOFCXIdJcWHCTWib9HpuN5ghV09eBOCDpNUAmU4ESNPd9ZVhW4hP
xwtCKoGlyM1fWyGwy0IYKaKBBGgptE1hm3Xxb8LDd2xsPCbgg+MnfJg/lIbwOvfB
tfFH5upwp75vPv5qCHxhc1TEBGTIQswG5ktIP/zGZdh3DMBoCGrheMXyUDZ63Y2l
a2wwWVlu2grruRAYwcLW0FmIDhlRQ/cPPgGfLx5pnRo/G+Naiel1JhWOa6vNKyHC
KQd44mxzjPiGmo2Ext8DfXfD6ujPEpWsxWbKWxAsRDuJXzE7X3UoACc5pS0P3bpk
B9rcDbD8GEr+TEOMQZQSDNc9L7+eZ7Df9684AkIXJbkqXezIUZV6Al+SQvWbsvIN
BzZ/YQLLHFpQEskB+w5cqfhH6WslQAXE6AyoMOySROV/ihbLRkcTdOjfB6sQjvYN
4tSAJISKAQgtyqF/VzV2CO/cKtIOEyq7fjtnbEIUQpWTYJNMqQptLhkzljtvy5LM
QPEeLZLRO75u7CWqBmYRC8cldcpi+0I9lCcwk6CXlYXa5TjogYGtUvQNiQMdQiX3
7wSwIer1vDVPAEAeNiGj2c9Kr/S8UR7O/4mdXV0LyjdYISC88UAXHE7Q9Z23cTh2
m6eL8T0MNbJ3k41PGKlzBI1jbAZBymOPXV5vrlfD05Z3vKfcFR/5CHrCoMr9rzm6
w0KFbt2e9hgbmjN4gmjtqSctG9Opv0womwywiVU5vlGUPsnx+8cxE/xbrsUlr84o
60LhRhJkEqyyI0XmY+fT4hBAIsDu21qGiy84xYRZ3w/u5uc7/oUusmiiHoqmiy1e
s/HAYzDHDCfYYTJ8N9DyXKhySXyo9Mjl+xx01360tmz5uytZocy6U9ODPeonQCSP
bz0s07qy2Ic1x/QRkrw2FveP4ZEe4GkBRf1iSikI3oTywtV4Af77xerGU4kjKPfB
bfBub1iBAo3Ill60pnWzBEXiZaH3SD2gwL4vPsgO1IgUoL26QyKjSkyINc74Zq71
K/t4hfITQwBKzA43T1nT0g7ARoGqxsJ1xF7iql0qvDwoJM84fEAby8VJXYAsD2HD
vTAXA4TZeXvmVCHxELLB+2XEq08cKeN8Ix/awVEhsSWGjp2XvkRGsfwUEKPAatsW
kYqw/DNudW7EGyMWjh7D4sKfeUxWNWI/lNhmlQtDTkWUesYK1dsCO3laScptOL9W
zvP0Resa3tgAQI48XMIaqxi/ofxv+5NMmU3zZbPHAzJJsK4nBCIk5MKcn/DNtUAt
lOcUshpfBtVufptSnWG2WNrVlX8gwUlz8kxdWHvv8Sob34Gl7cMoBCjVOa9sj659
Clk/UTbNM85tQ74AVxQiEOxZzrYZfONKNPC1V+w7rrf5xzxvHqVcNB+8N8keihCn
wVc65AM1T0hnOJ2bCSUYrXjK2x37C8bpoTM/ECZYB1JDJ4Ne+T7TFdrMokspzkBH
n4KwGyFQirer+hxVt9nxdy3nSxnzHZMKscEAESPIN7a3qG45Zlh75/2d/UmU6Mua
8w76WxKE5+D6P9ewUckq0fKVnPKju3YHM/+UDQhhXQ2c7y7o8bJW4p8wsWwVFqvh
kBYAzrR5PBNEjSClppLIjq+vbY760Dv/tBuPcRHbFDOn0ktlJQR0GsehhTiVi9Q5
+PNRFWNFEOg2v5Jd8jWAqzLUsPu0ITC8fRQFJyVsdKUrPYMfLoAMpGoUewv9IvH4
C44UqNe4QAkDCkkGIJfvrADqb58zX84Rndj2JlPUhbCCNNUtX+NBMYr5efpCFHyv
fSanFes5JmQBJn9++3xj+hjDclmnn3cbHqY074LErmbp91cXP86nUgE4qDmprQaq
pdl9I/tGnHN8H+/WVzWtYcimpWte4j/KQ7mA3I0SH0AKHzGKi6KsBGmX0y0aNZq6
zbhPYPj7lQ+Z9FRwL49HDp7XiHH0HEr7EkLLIE83to9LV8OBBvw/VqS2hjkF9/H9
TyzZkz93G/Bvdvl0mWsdNQ8B2tg/pK2ZZ4PByS149JplUtUdQG4+7VbYppn4iBDD
FSj0zhl4EIYEO8pktChu5IvUjxlJWSoH/dl1RjmLo8KVLHv0FFXGTG1O+MCGOaey
FoWq/Sl6/kIC/dISKLcGOvj6Mmfpw+TW5Yt91KaUEtpKVMCaobn+++cUuIzb87wv
u0CaQ7xlIiNRio1MxqYG3R8Hd/O+VuyhxS6Bdcj8MSF4eXK3PiULbXG43e6/TmfW
CRBbOwcI9Kq8E3ZJd7EaEyKSs4UMTiPRFI39QmG/+JMMsdXCQ2CKlgLRA/1U3rDk
9qM/OMppQNDzsXvAa4Bu2Gi7YEtmbJJIOjbcOttykK//6b8AbO2k3qN+Aqf+uhOX
aH1TP3186V/MQOh21qJdxJA5nQ7i/uQV1CJsrihZsQyc3U385aioG1GWfDKPacww
C5cebaR8DPHj5J+xvv5O2wCSlCiV8nI+LSMlrlkNB6/2AqWp4pLD2yK5IJ7F27U7
L7aJkmk1wc1ba4XUijSHkaCXPVO52HXzt+sOYBCBUyqcGrvq6yc7/8fEeD57xSR8
06j2aaaZJNSLsxFbupbig55nq1znnm+9mYxWufkRpRV5VutJ1XmQPlsoVLkkKDpZ
bG86CKmftUadCWV4LQa7zTbMX5LQYQ2MFMdat1LUFvjOgCjQcnPsQ0emCQAsVYo3
uz9oICTmqoqGTQFNnTS15FPkD0Uafa+nf1YBqTCyOdLWPkkrUNyxKo5InEz3avBo
ZWnoA1XGILt34FDW12nmSh+oJ2yPsXcFCGjWQWdhH3owBWBoUAFlw6Xy1cSBwJke
LrdEMTeHgxGRxITEVtnrVHZHSmneRDda/kPtxuF38JyFfv4Q71rEBp6dStUmijki
hXpRi4S8ALh12gMeSLV+C0cLJhrt/JJTLWPS8VW11owZwT8N73IilwLRLywA2+ku
1P3OxCRAH/TThPoA0nx9F2hwtKiSIUcc3ezKvUDJOSeuE0krgXXB+9AnwiaaK0SG
0mxfoV0vc9xIAYWX9NxIlBlbuFRoerMlLF+yne3zapBR4l41jc/CC/Fcwfhk2CkC
poTvjYdLEF8Ys8xwk0sE7UmkoEQGj4M/ToCjoEJ97hMENLsWVAVc4SzH6MHaSLGx
TOJQHMRhPwdpusYeS6ww2mabX5YMgNIlyEGvhJB2IYoGSQfW38mOZ2qZaJpaoSrG
E18gvUPOxjDz7ztbhiz2k75Crrvr5r1QU51rv2MsPDXNxN7wU2QDFiO1c9KHh70T
CHtWlqghiZCBCH0Tj+8EgcxTIiFFssyZsS0AQf9MHJBlXX03GjbguIfBsXCOcJN4
G5V8VZxkyefh7Mle815DFCKNWMsdhB44lDxRRFkqUo4YQnYem41bWuv3kyvdeYOS
vzZ42SXBXkpTq/t2nStJtNUpJ9q4fD+/Fqwyy6dpFQqsB0ofFSazJF3glkU6oZUS
Udb61/J9bKA2AY0etOyyDU0jbO1to2sFT06x3cwSC/gVoKTAT+Lajzi7UqoXvshe
Ne6+mLZo+NL+mf8mFdHnEYjFE39VES71BerYQ6m+n8+iYBCYWI2m01qPyuLJuxSl
nSCVsOQgseh7VTijsy8PbK+WxZVKA/5bx/a4NPbt+E7pHgpChXZ5lW4h4RsLVNBl
DwFeO61EDJamD77ri/V46aKbwOCpc9h+fx7/my/OC2+sbxAYH52B/1YS+4dDipFP
L/6+Cgk07H5jXIf/vF+7W+Dxc3A9QNJI2067AbEBOd8D96NIoSCuHnroYmJ2tbdw
TCiXmdBDJj7wO/R5kRUEcoJRMUlvfrq1C7QQZzarUf3fsCSLMyH7ziT7JHQE+GvF
FmPcne7UVaa6mUIKfIRruFk2itJnFFuQDp9ndIjDI3cPGPE2VkESYgcEj6Rg38jz
qfJGGMtO/PvSn4WzP6yFQbj9zvovbBvLd3cAchgIKHb2y0O037Gcf0eA16ibHdMR
zvsH26A9UUcUfRNTUe5k3LK2hAGl1TNQPtF+ZneYCUp1jxeNKkez3yCLhruSgPIY
GZ8eo08b3t3u5YzW1vIL78bHCMLv/qCB4bn76yPlHhaRGKr24JNTuLjQT2mW9UEi
MZ+hWLPkFCmrKSTH0IrZXLl/evEMQF5PnT0TFBc0YCeDbsvEjA6fnZHFe6Z00+EZ
D6ySh9gMMlkN9hOOUUusIhmBfD1Cfw8zqQ40xZoqGPQd+gF/Tod4p6kRF9iLZEvm
PvKhKeH3TL+XkgiqzwxC09OAzYxCnTm1KrpW9mipP2mH3lhnOj4vShuYh26XrhN7
dJLIxxHWULGOEWqrxLl+qkJj0kDpChf1nMro1ywTfBPGNtovfzL9O0kVpIRavVp0
uGlQfTwVZMMglfjttCMWRg5NpYgXOnhiJjTK2tEJ3NkwUWMpyiGgFRB0yNbYxfQD
rK0FH5m829fdDu8Pi/w0gydGt6Z06pGJXuCkhEymSdTLWZPV/NuOauvcbOuTjB+e
OZPW1fP1tpko1nhrrIJDy6Q5DXmSNCZDL2dM7FeHfqa7FpmReHDZ3BLH4bD6NHOJ
Qj4BIMC8jhqtpdpfx8em+SzvS4kHtVKCaHfjE7Y2hDZso9DK2rGdI9tT8lJVUSIQ
Jr0wq45bgYR39V18tvzTYacWktERCYPd1p1T4Ggyvy68kM6WKbt0nTEsm0HmmU5S
99znelPh2FcNzrM1i2hA0d78/uREJgneMLX/UnVVoy9KlpnbaqK8cbLKfe2OCzpA
V4k1qeDM8DBmNnUKR/As6vgBJl32ufxb78+pfCGTi3INV2bJaFTQL+wNeV+XWphc
/fS1Y51LhQeItU9lDep7zRKa+h6IkQg3QyOpqGCNHeBYjblnxqA5HWCeIoXoXnAL
FueDHgmrRuvEv7Js1DqyVAy0YhYv/AC3as0gUMuoUzy5GS0q1sYcIJJ15EX33da6
2HoDbkTnMV/lPqsm2ksBrWIwtMkGf9K6Tnp7yr7neQ1NWZ3pFcboDXanYHFoOBnl
0tM0WjEOY2xEI6rbyu0jBnyg+541SFttxPX7DDdl8kgFiyWQXbxYAPb6XnU77w85
7i7l6Pian/kW9m8sK7gXrzj4TuxOf00EQ6opahihOLJxn+pcl+ek1LVlNuIqLiDK
1nvkJPIvH0xx4uqV2ROTsgSAeuVqqMUE/cVK6JxgrXLJxnsg8ZixVeEceoOpoWWM
6xv8tU/Z/tqKPCD2hRO90ZdozvthjvMrC73VzHYCPdopYPBigobqk6K8d5gKuybV
o39PuYn6+Klfk9ys6HOtFA8eOU//ie4QInuwgOdqdNtIaFHQCKQu8y02RL4VCAXk
fnrtPKtJcy/lOLp98tiU7wdKJguwI2/RgX+eaSDRozPNKJSXy31Oaj8IJO34rONz
ZL2vYFLohkWv9uDORmfochuAVrhB5oyTusPW1OdLrqIeoYEi8TWvMiSRDtXEMNO7
jyTbDTYyVQuOBZb32ZACA7WgETI0rkBTodnEfcqkDabgkWjEHaDzhE8q4Yj/oHre
31XUVnNCIXHjEUMScIOzwmCMhhKYEs0bQmUxuHtfNPbkr1wZF6LWDpXIj2Fiip42
z6Si1JQZqG/ylHflaE755GxQci4r8SZAjooUCz3mwfvo7Dgy8CduHXpK7MlSnjwe
r6MpstRV4rsdKmg5M49SMqChk1UsCTEfZvqFN7OiKfnMBSk3II+NanIn7nEEe0Qe
B/fBjShOYU6TQzVWUEEfNk/BK22WSAgeuSYbJzkzSqGn2Cs0JA1JmyUDjYgEJleE
YqT4iZ5IryTuE4fDBbMZ5keyvz2/F9H3YLp9Iu9yji9jzxkx1DB1oBdGmrhdsqES
2zLEYxehFNNLHdn8FkE/fexLOZBRAM1Cq4cgQGIfpi3wj3s52OdB8SyV6E6394j5
lacy08XNJzq11Np/P/ftc+EH1nkp4L1aYP8YmF6ZMHlaugB3pD/O3p28BJB6tCKy
5F8lUbbSedBZ4ySV+ZzQF4aikWAsqR4FFPxRIsPMcABRykUgi5VxdK91cFScD1Qw
ciiK0gxBO1iDQLIuLWgJpG5NNZKSdxq8vBX9xlmt1bVQXTwY1Opin1FoCBYKoxnk
kPuXKfYAvTwaDwit5lB+rZ19w6TayZPWhOcrnD7KX6zWi8TJ4JZT1YUCFxz7RBlt
4kJB944ehlwwTnUEPjEY/fqJw4leT3sI13j3IQdJcOxaFPuhHOVDuK6CoW6ZBXkX
7nNpj85+rY36ARNSGjWHv0sLuvfmvfbhknwDCa4zZORKlSYA4C0AHxn8EBV+MNFc
wtn6WuwqiRphFTkdMFrs5NoAvQK5Nx6+4LSx3/EeC89wAHALCfqLlwElua71ZQ7O
wdPsXyxh7D09hE9JJfCOZPQ0rOhFovMfrGqXS4odqmaXOkT4QzHp2Dei+Lx/NkEn
AjdcM5F81KTjn7SJDoEv940ZLIXZVhJ1gZ8Bsy4ThY6c67/EosM4B1MIWRq1CI84
ZQrjcA0jbtZVPhsLkFeL0mB5IUFHQJi6mml3I7f4vsQEp2IlxZxiuT1RpDyMFvqJ
RkVhFSn3E6BAAeI7zFAk0fwio2uE6CvJKZCKjnl58vR/pjaOWBLs7wVjT0ZT21TL
t80SBEhvZ149RQqQVDzft7mGVX2nte58ePGAWB//9peLJmmAldFznLsc06qzn/og
gEHXcKtIYErWRci6LVty/l4UuyWzrLnP0AWJAQX4ZJE/GgaccRmaqF6M20NryWo6
muKZX+dGzodXJ6ypJ/DxEemnUG+luSjfScUkuUIVKGkHh8+ltOFxNCCyZ+k33PYT
w+DmbSMRDSueBLTc8mRj9TKMUvwU8DegSszfCH1H1VDbG/4pbnME1h7o0I+xBMCG
AhP5ZHW4dAP2K0rFYiIiike4WG2v5uGHya9s+CjnyFnApSEMnLvbJHBtOw+w1v0h
TxkhW0wJ51vAgbDBX9iIcAGgxR7ta9zZzx3VbyrdA3wKEQ7PQED477lDTBr9ro9w
0fT/x0mpt6t6k/KY3UtWR+ioDR9WfPdnD9Tvf2bd+P0lNPgWRGsj+7uXxQvGz4Wn
D/r3PUkLd4C7Hegi9tXWoKgFGIZ9d9t2xUvJbeReVNEKCQg2fQ1WDSZYwwDgj/oK
jnm4f0AZwFs+aVzxNfFJnMtqBR71crveJVF6coamXgC8VTHUPB6bFgu3yv/3TLjX
/9/cE7PaUxYNHEQeDHGEq+BOD4CYS+BcfkNr4vLRTi5FQiNbIoQkvGm7+VNGax9+
E+aCGODZ614C5BJVQb24t5YIHExZRRh7ABBQUSpOSfsD8IsB2U2mX5tYzgZ6IcEm
JYqyT/XxWaIimHBIzcqPiZrC7RbbUFHeA1EpRJLOyZK8JXSWthuTatOcCrDhJFQX
1zzgHvPwl59SDK74P2LFpWIeVSfXDeenj/fvnUjNwWjpJetBCDNW30QX7tZz5CwH
nY+qUbZEAuT8PkVOiU7WFo3b7ZsufjuEB5HHIQapa/DY/wwSK9HOU0EOHEsZkv6f
3D0SgbcIWX0XBkiIuO6qXEaKktbn4lZsVZ17LvT5ri4cnlc18ksmZK1+3FPiFVgt
x5hQhr99Ipr5D9wlN1bfHJJF0fD2Lh3trU7oI7g9MFvy3+CfHfJU1X765t4lsZMn
1JWSEhCMxlV1p+JK0CcayfjAzUCNp0tne6TMZvx0GLPhbkHxo59Re3KV/BlR/wEx
BmiFNillLQGWwh8tR2rFsb0rn0NHLqqDeeogiVC5M0zqLS2cDCC9N0KTtGzwbBK2
5rCz6nsjQODvfdD/0+TdiV9DSXxsmpoXoWJIjcihxCrsjVcwHNvXdTIUh3DBUlFx
NKWzeZRvMke1FPL5nKyWbtjt27XVAAcpChwFVQbnMZ2TN10xkmop9EDvkyLnn3Na
qJIja97v52DD5UiMbULKMy9xoKbpNPObOmTHRXTymOHRUE5fMXVawrQRT66OzkV1
HDJ1uD+bCEvqlHa84pU57tL1NAcKqzlYC7a1Uj85DzrdDAwyIIdB8FOX8olsCNQL
q1m75Pn51kVIpVq/FARTLlA8aF5N5ggt9340URs4hiZrbDRzrQPBuaScl/kjp26B
U9fxsp//VlQ4/Q3Kt7JfwKgDyvHQdXJArgiGEmgnWadv7wfwlrXegc0rEazdV3xd
oCqslMM1FB69On1OL9XsS20pJx5t/26zye4LJax0qIxXFwf/I8hsB1QqoFzTwCTT
98W6uM8foiKXS/doC7csEodHkeq/I7wMcxTfqeRsQN2fAd9VdT9uvPJyRSu8BUB1
nZ8vfFX7tNq/4MlSAOxSSCii1WQEqjOeahWRsAKKU0b/2/GVprO1vWX9Jv6Mn4dH
ar//8n/U0bEJoL9uyiyeBqENmP8CrHHHEa1yeJphuQH8Bf7LA2LtCeoAzwXDz4+Z
daAwJmmsknULE4X04q/Zk6QnzoKIXWbyLw4YyvHqCdSgvy3AJ2QwH+COmJ294Vpy
Igq23nHtQTQM0ac8beoxKR+v21vflt0pmeXlrtQAobbB4sqHsEmT04xl2idObX2y
afaotsf/1oI5m3R3REECBKwA9RG398JbxRmIUTyouj38rgwh8Hj+IIwBrqpNP8z1
mYNrQ/UAyVzpbraHo1liI8/NB2k47F7ZGD8X/YPQTg7jDDF5N0MqmrutnA3U1x7V
BsT5Nro5bSRhGq53gEOw5gughfULMqpygJ4ZG9TOIft+IwHEdBiU/JKaZ94IhlKi
3I6MAH6CO2YIwn6MBLitoJjNCGJLFPaTmAa2lyz75XnAtoOv+N7/4m5t7ssvF9iG
FYQjayRa05wIn9Teb4hv+0GgLXKSQGtFy6ASe7Kkwayj2KLcFhRhu0JUM3jSfJir
g0xRuzkFmTSgsbafwTsn4M3G7Hcb8CT5gG8+7MiggYfR1TdFFWHufnOcYQqr5QTm
5ET4/7xN3g6owDByKroPepW/By0jNgSaHCit3IwqjjKtqCaF+HFOifFHmOD4yVEb
WRMzkPJUDrOALXKp3cSnEDeBSOpz1YxdkFkWGbTM7SOol4EbXMT1OG4fPm5wlX9A
XvL2ba0SL7t1xvzc3ThM5h+LY1uqY0PHx07aQAf7Vy9ys7VRt+FsBh8B3cnTaatE
dsoq96QoXJfinEvR/ZLG5YIpajJLlpWX2Ot9CpLFQXfd+kJ79S9a0d/A1YHMR21y
hsYgQ+th1e5/94Ozq8ouXZxnuQx91xQMiAGAuRqaYIPx5SdXk/ZE+U647yCDiUdT
nI943Pn5URgIv4DrgKb6bmHX6x5cVnmkiq4bdgN1EhPsvfdgQFri0MBPb6zNNBdl
xjB8gD6dXDGcsF8hpoYlGO4zo6nDE+P/c9V28LbbFcfYSfilHPz6ycSBEfOKkEhs
1GQlck77YuqRh5TUE/K0fGcXCuLK9pdxBWyNrTalDhOWp0YWo0fHmL0AxjSsAnxy
jyWtjIMkNWX4Ci2Lk6epu6x22d+pSg8qlWPIIAl7qLHe55RtKQPnG2JACy3KrpkH
rAupqDXGp4+wL7H+7ilNwdg0P6HDrVTEFc4E67CXZjaM/O7GyWCIO03xDXUTOIm4
cXuY8E3Q6HmLGJz43RUDZfrXS5XBjMMyaDSAaTmTJL0o3YwuNXoykpm/FktVOeKp
hWJhE3L73rUsx1eEPetpqrBTXvD2vhxOkBEInqT/vdQxPWpz7aFXFBOiT2SmvT9s
IuFq0NGcjKZimqLwY6PTreMvNqu/HOHLTall8EcNHHUrMJW2ZsQ6XtB3oufJ5zIw
09vK1LoNSF7NZrHUCUU7E8YiJmKxNjvkvn3gi05pmnaaMyrjthA6IyXEYd0hjRDw
O50GGw3mEZ17ObMdL+P5m12wJX1LgCnzupd4KSWPMX4CEwan4oHERhsSZV41xD4w
353e5rN7/ngP3ZdqHWvlTgumrhnyoBwXokoGdovII3QZfhJL8g3J1/s2az+OiKFz
1+sgFPDKnfV9LzlvXIwp8Y4VKpCUXW/kEgKHdkcFrv7kDjI1NGpYINIQluAWE+tC
/deJpr/2IcDdURZXwIVMOx/H/hrbWWDfasN4f0Uh8V9FB3ChQ7mIvK3UbqvQIVwj
0okIcejlnAiFbpISE4M9LvpjDbk0SPLf9dICTX7wb0OmCYA/TR1J/1IaG6W3MLUo
LqV38HkKxKzEyBHcqPfiFLvtJT+D9GqyDOl5KZA5alzI0CNR8ramDyK+hsb4Ye4G
9hGzpL+HBYDFWdU1S8ArtHCJuxdskOGHbLG7CDmexeWemnD3uKvfZIfDEua1C2B/
NfXG49wL2OBc4ZYyzrp1011j66FO6cOROOkNp4oNO2bhjwuDSwIn/JkDzP4wquO1
a+iCJ710i0yOuB7lSZpcfw5sDO6QSvztYMlut5edGbhWRQHNv7XOzzSPmRMCh9bX
LOjuRfgX1/Kiy2B49l7sYUOtoZTGtGkXTpeUFZUL+VopGvH7YHkkytQ0AgpOYqSs
5DP+IDFEPt1ZVomt4mkQti2drnOEpdEZceKEY0++zV1+7comqI5FpzZ6LT4AdvOr
mBbtRAaP9IwKHRttVA5z3TfF75wacmPd8SktZL1tDxgjmhteMWGt1mu7393FwFAZ
3SlEYR5/L49Bw+NarEgpgegGfddxe9mnCHo7OddmUoZG4GWLMElzw3PEqKXJWFJA
OZB0CZTp+JNHTZxPwP9/zxe2bD8meFSXzi+/Vx9yry+ZDhBijeHwcYl5Y3niuKKw
mgr1Txg/r0wi9gG4Tj8y0FnmXWSYwOq+bn1MZB4fg3Cpc1su8zMiZMxRMv/ucVpy
CParSvRfjVMMbWZfoiImgTP6vYoBXxxyzaFGN38klgto6/ruFUY3W78sy1nlYHxv
9lNNBh8dMipvboii9GGHeKp1UuW8AIVpM9HG9zvfGH0/xiUBlo+pTYWtlVkhhW5I
0/aBZSRLFL7TxTJSHwlv5/IMk8FChMHFHz3LUjLtznz4dBLYyx/BRE0STUxV+6tX
iVkfO81k5JiddY7c4EbL6CLxX8/9x/Q0skI8aB1fwZ4AKuzUa6txFfrcMUIBKnx8
z3p1RNGrBkAtviLvegKKNXXDV978m6mN4zhf83VH+6t+oLsTrQGYg6JsE7iD8Eya
DHOj0ypxehHfRfm8AMEOfonbf1b7m8zGeWWXAV3jUy/aGY87RYgPeXlcRHkQI6zO
nUvZ2oBqd/HujWf22pQGihHaSiQBVsEHGthHqkYovN548jGOM6k/5ODR8onZiMQc
tIULF3lGspV5Vxjj1upZFfTnBK4uCzNiIdsSSbR30dmdOhvKK7vM+Vh2BLrIneT8
26QNh88ap09Ostcqiy3o+rNFYXII9iBm8uKzjf2hWXjYCZ1tXlytkpoaBObpxQzC
IZ6xey+usE9XpQGkpbpSlD02JbV5armUebpomIpvLaV3jB55S+UwmGIPsuz4NZJv
Z+68T6fCGH6e20kWOY1Wpgxpkq46pnUkwKgg0guUfOcjMDE+LJomB4WIlZ4LHjBP
/Fn49rn17INLxOIXiHqchEC6oe+1O/O59ZnNOZB0bNpGchnkfLsEN6UDh219I1d+
bFskmt/Xkud9TXLXE76Kaek6yr1oyOePqt3SWV/4+O6WaeGpuyJylb/bdIgR6q4W
dLBWQKGteDi0kFVXqMMg7Wp5Z3qC0YjqdqkjZTAHPbjNJlgH8mXbg7nPiot89xFC
azo2HqRZPNTqOW2BqyrbHATYGs0Xnf+l8rac3B7+nOKBCvD4sKKV2HqhcLjAy55g
iSv37qwSSg52sjcZ+PL6i76Ff+ZedFe4Wg+pYfHLtucMGGX66ZcYVivUhXqXJ8ws
ZsSzjVJB1QkCOuXmgkwzx0oRUPO8OyrmAJiKiVzmgjlbyI+HmFeKSbhQbQPUozYY
xARa69gz+207K22Wn3Rie1czut7PIY9Q77hiAlfHjnXKwu45r5lnGSZV6mEu5KOK
mfSZCqwvxMOogFmdaNqWefE6KkxqRAbt3pZif2NbzUEmyNC1wQ097dISqHVGnell
gVp8IZD3hN1312RPRWqCBUm+lJL6cYuk3z2aErCpYUB94PqvBhmeR1JVPgGMzOGs
1BxvHQC8/ygF+SvEH649Q40SfGFcvyvFQRTUfJqQhmpB1yEPJ+4qpBlkv910ga+R
cGAsGwBBXbylFx3axuwaYVp1KAFRyn4NoHamlGt6zHyZ3KLhrcBuSfh7/a+6s0hi
9BOAPipRk5khEXMMZCUZkFjtIJlekeQjfqiATp5Ra70+LBiBrSydEvsrszLBwADZ
Qo9U2stdDWhxNXTlQuS+bIE2fEuhpmVYA7OrQK5n2wap/y2Ibohehg1edw1BBsKg
7i9uRacT2WWqCd0J2YaYsooDnh27AaE9yzpMLdqFP8aT08fK2ZmHMEBwklDIQwzo
ng3nm4MDsJ/aPek5qy+ZjDIVQp+XnlScC1WpQIix/MTmck7KhSUCNB1mBsPeIoF7
1AzBiiDFglGVDJQI22sizEvqDU+kMTppo3LVRfQbWsd2Xcx/kpU3N6c+L7Yr8Y76
WtfIOK32eszTknjptjuScShxAECvm3lQsy+vOOFFxCg7E0q86YPeBevsan/3O4gK
WpykI3xAkXAldi5qtfnMY4Gqn0b020LHp3WHwXQh8gRl6asJXhVKv4OGy99cm2kq
fTZml05RceA12cjMsLf8E9BtlYHExcJ5NeC6TpAR+wFQ7UJvGKNqUxPeg75smvha
oeSOypO8Nqmx+m5d6PecuQ4SzIxC1INHSTorWwDzMAO29613JLZtTKs5jSjdJPrH
SMX+eQCW6Ckk61QCDJiAdYhOShdSMQD079gmi7LSwuK5nCSEFRdue7KeYHYTDy9B
A9lmc+K2BedCs0wiUs0v1zywFvySiRMFjeEA2HSqzbO1sNDIiiyhpBcG/k7iUIJd
kJP2qhJjylOrW3OMNQ2k+KXyqV9T3utNxnWEouRwsecerbrSY7O33iqXKpIM6Hs6
2xzSK/IxGvjOc6hGdJ0DlDN/Pi+V/x4WhTlHQ7yzbB+nss38h/4uvU92nnES9gsT
W8+OI1DeqlosSAVHCrbvbmX4iRwIkQpYjQb5OlWwklPi4kiXha6m5zLtiYNWikd8
JV9Qg62Y6bgki/UflCqh5D2mq264hK+MWo/1n5cByH18001QEi9iHWk7ns7Z/bdc
PhN66bwZqRskk193apphqLjde1wI2+cwd4q9+9jtf+0VsWjBwzrndZ7DCxA8Ny8p
UlHlnOLt7aYaFMTDod1EdmV3qq0n5HC+UuX8nSyvRRqQoSDcwFJLUTWct+M0ZN/i
ga/l1K5I7DWK1LUNOdkcxElGXy8GPISoYlqLVkdftAilRJ+4a7zpuB/BKGJysOwu
joJKhB16fUgqYISQlp8kfGCpeTJ0+IOCDY5ZeD6Kgob7TiEJfgukC9ER1acl4QI7
ZRlSS2m/5wFcDdMCgO45/H7JuIOm/dRvPqDQi3xjXDUIqGDbJWA9xpqM2ht9RF5O
Lc93wVjqNyhLORGVrLdZmjQt6ZdSY4l0H2gzGVFoZ52EWz+aRCcAK8iqJxP52pP9
us0CT2auU/51OWc6EyJB+PRRz28VnYisZYuaYjtI+UHDBF4JWY8Df2gFu5HDfBob
7+fin6RYrfUlBwveXGbjoM2ig0gubma+l6E0vyQDS6LoMKLpR3hWVTfJEvlESEZD
VsdfTHNt0covjPbrEljFpBG1aUxRsfnIbg8Z31x30KFP0fWzfkicsvdHG4Tq5Rsa
whlPIVAaLyDXM8zkzjvSD1ZbaqLdviTgznQEiQPIUFqIC/hzhX0NblM6k26yNMAd
qtbnZfQ3CAxJmyxtPNv+n5gNmKHe4jIwcx+aHWO8heTv+nH2YEzm++yEIxesa//L
wzADPjXgzNe7DFs3QAitrIiPghQhhvEdVzWkVmjbXci1BUsOfZzvkVbhTlg5IdC+
CnU9ce2ysYU9qaUyJvEwVQxBaLa1+kyERTuzdMm7o03mEeoWPXSguE2KECH3Uwak
XKYtdzEaJ1MQO67qat+oYCk+JEOWA6wCbdO4Bkcc0YgrrCNJFr0Wl/MqvLocL2Vf
lde7rKJXaxcSUQ6WEBu2tftarLnwwZwkXOHVUzaVOoXwKEw72y1Rrmv92daWih/k
AaEw4w+UPuCqjF1fgH2w5r07+FwRnyHohD1LnoCfu2tJlMsPjdZvN0XHPn/+srwj
lPkqKqlCT0YyY1r0imrykkkDmZgEuDPHb72aYG0wD0kpQ5yYgUlsv6cs2GKAooWL
WMKbPiUBOF4FFFafpPwXSD6ReiEUYu2ySJt8UnL0Wn4Eftde9dtPvCCEZZRLNyqJ
1kFDsZdyh1SJcieEhoUSTEKQRB/lBhcsziECGcQnT9751AgvpwfBp2zlg7IHdEDo
3LpOImer4C8JVIyBY4OKz4E4ZoULWT0Lxmd45AaAHJNq95V4GaGzp2ElqRNFmPtE
vlLlnpC75uJThTRp0d4CqFHo/YdIZmjRpYlmQcYwMYw276Kja3XaOQ1eawBj5G2V
JZ4Y88hANXwyGxCOJQP1qeMVg/q7V27XeyAxY8Qk8eyqBZRh5C7TV6ywBlYBKdpz
c2xRsTc8AVkT5+l7yT6vFAndYQ+id3UPCrK49rVAVRhQewrt6qpgWsj6NU91koSe
/CVdpJZJEXujKcCawXbywrRvyyQxSYl40/pVcniBef8ky2oRHRI71uvtrgYgcQRn
l4MTwH2olWB0tHRIB9az15EM8m11o9kD+Gjzb4PVEoUZWyrc0bi09kbVLlmjd4zh
DMxeVPG30yt5gbDqPzSNpKeLi/zIU626uCTVW7Bl+4xcEHkOLbqRPIR9QpSebsw1
tsfZNQC0OxbVPnJ/mJtmV8G1/OIDAXBC29Kjl4ksZwzBBpEdKuPtiliQtJC0BdaH
Kwn7CTHJx3Gp/xMebt2bVVNxA438Uhkv9o6O28RyL/1UyCc4xnM4gY0jA+R0lXAD
M6zho67q86U/qguq+nd0SBgQczZYqTJ+vVzauIDhn2Y6PN2IJ0uMKk35MACstPMN
LD/9WLiI7qiC1x7TKz5XLI5O8dH1bwbKyBoPlDn/gsq18q3nJ1hqiY/EGukth96N
FP/mtTMkkDp5qi8UIcoJlHZVOAEO0E4HeIkIdYw0KvyXoTyYoXJumJITLEviOUst
9b23uPhpIumma0qLE1BlB6gAB4HnARfna7LXk8XNXbNgrm1LzKCZou1UDSCEFQkm
7Oa8rfKTO2mRVL6kR47p/uZgDobteJNETKu9k+If7BMTvbowc1TOkRuM3YvG5vhp
1N9a7U1SY5dWC6SJqugpr5RD8Vny1J000X+A4RUn+BVq7nT17NQgPnH9Nf9anJdo
/dWiwx+yTqAe9YoUuYsuPJ+0H5UojPODFvsZt8CQpBarzrHKoHPwWWfsIAmTFGZp
+EiIDlOVtyvZB8sLegvN4izoqYRBeYtcapG/QEcCwArcTo4qoxq/MA0iL1xd3s/h
qP6zGzb+4c4FvQWmAYub4IXuodFPVWQhxXhqgJtDBqfZEr2A4mlM3bdUGrKwaKoQ
Uz3PMqfBv/i7XiQxB/nswFRK7m7c2OiHmrilbfdhIcqWObRFu0TDwi2MwvmYTG+3
UtbLqtn+6XixwkB1pO2/EJDAz6ljjiTqQkddyENRKOVeXzfgJ5Hd+RUHqIpgLz1U
uFmfdZRcvE8l2T11BaeKD2mXasSGs/WPQfwVKT14GceV43ulA8ZUfbI8usuCkl43
rFkOtV5xVR1UVv3MIsd5Z0uOeUCOtl78zy+TAWvfJ4S8ZmvqrmDZpTKz5phl/t3l
OOS4B337CVM0wkhWoBeBBI9QsYkgCdPvnXJIvHY1GR77bJTacDIboQDfmi1vV5rq
Ub72tyfCMIV57t3IRqxAbcQL4uR3e0bfewdQY8gE3d0usYhGysFv86TNVmoKsOQA
XSnB8xfuWDSIcG1rjVHirw8Y8Vyr4+QTy2XwOCzhpCzw+DFqZ/ZrqrkItmFHOFAp
zooXSfg6XRVVTHAKMNDXrxyw1tSQMovaZ2deSnyvBp/Hiym78NU/m3Hxe4SMtLcL
xSKlsskJ8aDWtY/n9gWYQuThGHVjJwU0RzXL1rXW4qcu/BEW0GF6UqZM7B3RlCDI
Pc/rSxzCyWxLJbdjchKo3Q56cHU9KKyifmqkipmArWhRfe4rW4dx5A0ssAexK+Vn
yw6tsrFfj2ZUorGD+RI66aQDwjWeojRste3EzdfGQ5GPpg6FPOhQFTNWOczvrs5K
xHHejVzX2mbin9BadeY2sP/GB23C22Uv79cSSSVcbnM443PRkzOnDZQT/quGYSMU
dwHZHHjTVcKT+k8ChKpOQrJ5EXll9fMBIR01VwaU97epBW5E/jgFdQMvk2+1j5hk
z1gNBgRexB25azyht1kHP6wraQ8aPRzXEwY/jYdpnOm8MjjqCkJ7aKu8j6AA8PjD
11wJdvm8wWdQOFOj6xUmQ1pLXSJk44YloJsmLZ70JCzL8acZbuJffAAeRSmOs8qK
Ac3G4zkGBkcBKuuyMhxnkKmHOGMVHRB8Unhh8sMsn01ohKHgYJA0Ytk/j7yhU7Is
uytMenESsAB88C9MVdrTn5DPswSysNaEt8aCx4ODs5DH4fNLOpbUOmxVzEbc/VRa
Zf7uwhXsfrrTteD/Mp0/xj9ALCD1CEvrEoSnnvat25LGYBUwBOvujDnLAtefly3a
Br8EzWrOkIon+oY+blXVxBxgLO5yfW0iEOxd7ySbb6JYeKHcH5s2qiINPrOsdc4R
8TpjVUSJG0aWBn1pR5bYZH3J7hpO2k62mg4p1hlU9pQ5mZBCLdmTYCiLe32MuWHa
NrBEh6+RaAu+2ZsQXyVoWFs/fhuT0o1roVCYFK1aIy7yuES9ylxTOMYO/Qnqjr6C
RjygYs7dbWRzFtwzBH4szfqCQjTJhL4ompNzCJyXsKmBjWox8DB1xhUhgjhtfJGN
uCBp5sSYF9Y9a1yOW0+P6oZO21RjDXdd3wCAqlSWhCyqf9DM7S57jEtQI9nqJ96q
NC9i3WHmky49iNheLXLFSjFIiLotx8vHFiPc4USeGrdmoyBD8fKQ7/Flqr+o9uvz
SWQcNufbUIsJ9y1Ug8fIPdOvevcgMGGRnb4y8Xf7PvGNE02zTIpPDaztEDXfVGse
mtzfa4Ge0P59HV0/DCpQndgAWUVLiaW5TJSJNRf5fsQm1fURXxnIP48unPysjoAk
8lwmz6vP5AtD5OLVqS/e/kQtIpmRy3s3VsJSiydUQgYDA7wTh4yZL1+6R5ejdNI0
VALZ4SonJY4Nyo5meyZ/Ciw2XiDvTYJU4dvd5TyzgoS/yOSUVCKrl9TpUYrcn+/5
lW7p2qcid4d38rcnisc/4ScXik4xYYDWRl9or5bZstCtKpi9/jRi0nCvupeTxfCS
l7gkXomiMGVWDlxf0lo53TXeU0wpClk1dKLr7HEwEGC7/exns+c3/ZH3FaDgq5s/
xJTSOgEJsQWv2rLYDEXwhuEu4XrURYvpI9TwYF1o6gklGAbj6wvxm+ac6x2MOzJD
FmDDdRzDTnXgKUgTgb7JQBDQmQBt1yzYEshiUDugrsP0nDWuF3vRjaHy9e8uJI77
DJOxwlrrWIk8sWIj7Fj3U4J7xQnxEJP1TzD6Fa/rmkHEuVSFr6YVAVYcm+FCYBY7
9JUHNTnh3AfAkhBbuzd0Crskxt0PfKSfcUdFzTQYDBItZLqqIJR9+iqY46Vr0yC2
WTayhTNJDNMAADgVdF5NZisRx0HMoqhA0XuEse4Z21lDym7lf8rRcOquCkkIXNdE
DDLB7UxECcvUaZCjhbjasOs6TedPuI84VHJCojQgiMtgIg89h8Icm3e81cZ3r9nY
iR5ceDlqq7nXRMg/jItagj9meCcYieIUjip+TswmtJAd8U0abIGcekYegP4H+vY4
xAlp4cNcFCTTTg+C+6cXKshPbP9B/6GUVJzX1gtt5V6PR/5IM1oYkFrkf18c1LSb
Hxbt+N2kmK0v8S5/QRmymTF3jetWWGlHRFs/jLeDI95fvXUssE+0DPK9+xri5w+y
6h5JLdcJye0WIAjD788LLeBXG7APXFd0MPanbhxOOYpA4HDSlf7qL5LpGyFE1zgy
ekCaGIbxZqvPhSDzImtKBEyEeHBZsI44RlRSKyGujqzWc3e31In23pA4JjjJD7+Y
LdisvmZqi2YOv363GFiOFsLM+t0nCxyW/UzqRtk3OkuUI+u8XccGQKC99RShMlV7
G83saKYZiv8rrB/O+xurKGJZL6oxVN3n45mGUj+htfDcxWdLIdAhcslyJaEnKw8X
0NBIJnYLIGQdKpZguskHCKLqPrqe3GS+MbJeogfs+xRTRcAkAVNFeej2IilJ6gQX
4s/nH/3TsnOxJxiZjyAI2LjvIfXz9iT+cFsoUEKRX3C/csqqPSVnIkjkrjrV2SXQ
KL+DpXSfJRnv/rfF9ijaFr7hVA5BzYLYe05WRbwJn97I0nfroknluf0up1CbG3BO
+sfgy0W6Wwiw44sKSFZ8nAT2DUIiC4/VFJ0myTFKAbtc4I6BGLINzZ1qn8QVGYfJ
5VuYfi8/84pOZud4TpaTRCu0mwqmHrzDL/v9XW4Y5qtDkbtgyhHRkxtcuj4V1Qop
GZkdg4lZGAOK9+Zc8JxlmRVrGxnEMHSh+qDuvcrosyoWDGTS+UQtU8J7BpEfcwng
8drdSAt/0VKriHnKHSXKBdAiWhpD9PQu8svpvNeZ7NB6MTKRM5Q5v7pkGI8zOdk7
MJEpy111Vp+X0QpsFT1aR7EZowQ71GPWamS+Ldy1dKmLiw7Fuw/LZTPrAQBslj9L
VRbV7hn7nQpRDIi6UAHSGc1zliaqpFDBtMFUAMjdf3BnnOa3r11+U1vmiZg/jRQB
wdnUPgk/qSJ/3822hZ/uJhcjn/nVf5Ghbv+icEG5a5etwaLTIAKK8XLeaH6K1IkW
FoEIiGMSqfgGLMgdvoorOeFcSOudczCjH1zboNWfJPkJS0MTIA9JoDaHlnsME8u5
bHLuR6QfXwpn7CKws+1FD/h3WUvs2FNCg1/6wNn2cytsZvPRu6m5g43ZEltNTghF
WDshBH+M+kqM5wE1FZ5G6t4oiAMiamDEHTFvC7ccwIsAlvAe69SPrNuk1fjKjxBX
1PoKX3unDpIfTRzX9S65dJ+pJB2b4Mm4NFPXhJiYzffKv44l5QgwdpGAuLeUmWQj
EZBIcVe3siYdpULkWnh6zunJQp0yKHXm8ARwKx0oszoc5A+dB3V4RTfPXsvaffkz
XEFncvR/YkhNtNXyV/OBCb62fPhI6Pkh5kwZKzVmfyS8IYjHP/S5gVGWfjIBIzn2
AJ0irgLEQZ7+t5Ij0Jyej/lfWD0XSt42feZHjxOHee8Hw482274ej8yVvvJR9DKc
p+F8kv2XahM9SPCjcrI4uTWd4XHCCjDGZ/4phR6OSjpw31hSMKgP4OaAF/qA121l
Fmt+kF6JzDkEz5Ipz/o+JWc5lrAT3kVV53ccvWf5zh0OGLrxoh+XMoi9ZRlZsQka
5TlgcxnUB3ZSyxExJsDVjEIaOx92NruV8Poqxjdr9nwkcfO3bqi/DJ29nAmH2U3/
NH3WIooDEqbH4m7I+7IUJwPSSRdcdryUaEVsYf0lfV/8sn0E66ZcShmYfmXPkoU5
Va4jmoI5lxYmT2x1A/s9GB0RLnpdMT/J0b4PJRVViGinGgbUn4iBcSmDnAT/ScPA
SJS3GyNKb9uv/LA/wKnmv1Pcfz7NQ7t1uI/kesT7+wTWoKeZmzeFBrc5xpNCB94N
akyqJZzaenf8tnAxsGsY3+nYQ9CTlo5IyYGsrMUAvZtgUfXhTVfhm4Zzc2iM5FAC
Ykx6t6GH7cso9zZ6ALq9iTAqxQk/p40WCwtJkcmwz4ilozPPkNAKyrb8N1ZJw1n0
Zb3S9O/IGEZhCY/NYrOloJwYF4BIZmAz897+SrPCOtAAElVHTpUXSpo7ltavzAhH
uARdtiRvoLI3gzn0h1MpzxpRaWVM8q9gPNfm0VYw9nXIADvJzzuOsRzK18Xtqq8s
81PO0glUGdZkilnHGZRvwWZ6oiGt/pRA5lvoj90fY6RBiYdplAjTzJA1xNOMl644
jYVH1bGkTyTvFMZPXmTxAu1yQtIghgbsAgXpv7i/rac9lIQlBIOCFVbvK+keXRmU
5TpWj6bvdSbKoWTuNoxLRJqWgAgzerb48ykuIn91U1aUVK1vLgUGWY0+Q0QJZhba
63HSxKYlbJ0NP3U3app1g6l9htuv84RIqj0LUF6aVaK7wCRfJkWvx89TGfFcFmvY
S/O6O5Abb4UJ1kuYN3zOw/AX3cpg6Jr2VUbfnUS4cAV5adDjZaqEjGz/SshT22ze
WqzadFs/tzDXP9SgrWWVLtUcuhCXFbF+0FaglB8wlBC4GCrKRThehFD2p5fkn4pU
FCOIxeh4Z6Jr7r14NZDtaaUuIUsQnpJeLXxDKS/fVAhUet3NOcugn/X1679Zv5yn
N6IRf8dlHjgvdfMQ0enoZ9KRAbeHiNUqkdnOs32Q2vqOmuT5MXHUiBC1YLcQjLAV
Q9mQB1oY7Ky2L72MbtvDi0yUtEzllmuv43/OjRDIIvH4igQ3wKSBcC71nr+p2Fg5
AGcKHrBO+5Q6UTZ5sm7CvKTI5tkMLJYI1yIH4TXO+j43oA/UQ3142sYyJ8gmCK05
dBP7muybLEccZjG9zyeBFmu6q1Ux7kSjVY4tp+eCv71hbQYYG9K6k/d0Unv4SlMW
8cfRxWvDs1duF6sBZL1LDmnK9DhXi+yqSqGve87w9bp2WTi4HD9MJHFX5ThK7J8g
1VO0ozR3kLeg75EJ3L+8dDEZ74qA88tCL3yM3FY30mEi+rUS1nQW1UN1qrUKQIHe
4E4C13YDJusyN+3Qgf7sjJu8+BCpYQbIdJAf1laLqySZWFXLP9SixHBKQAan/aii
AXdaHtxmP1NLdan//+40LDTcfOMDzu/l6vHN9ZGlMYf0KP3Kg8sg2lXOD0qanUg8
EcEi9hODTf0erlEj+TcBInHW/f/cis74YlMESb4MjuJ5hF4EE0gyLeEE6maPw0DK
UvEnd4ohaaiPsUzADGUg0exaPzJGZKAhNH+E+U5Q17XOzTt74ZSwl4EwDXUiOVMZ
ShD5zlqXhRJJe6iAOrZO9ODqmZwYsoKBAfq4S6w9zyiZP+iEOpu081FhwcNiJ0Y9
Vy3Bhc4Fq2VZfvxCA1WV9ieo0AoIosHe0zNn4igmtH4jaUnUcGw+iO7VLCsau7WB
twpu9Ye9q5NAmLonlm9YA/mVR8/iNwvvOtDc9Ez/o//cfHJD/olzwKAZtE0YluCy
ozBGf9HeqHM4LZQQPnOLwbXQ0Jw5b7AiMIENeQuYhEj7PBMm6YanqtYZwR5UMZVC
wyTjk8hW7QGnLZXMKLmMMa4ncK7Bi96CgxzBA56PXUEEl+FqGN4tQKawDcDBAwTC
tV3zM4nAjfmXv/l+Y5tLvto91I8/FmECBgNJKE+k66IfgEXuFvYejNnlR5G+lT2F
vQE7TRFBnwU0GzSKI1uc+CgWguDXbiGpTZLnsGiU+K7LDcmS9VLX2P24zLuFT8z+
n8zLCPlAS3p6GfBgJppciwG8NrLiT0sZRdjt8by68SjJi67f49Ir+vwDgDQtamr3
vy6PIEHFSdapCmXwo7DHPZgCPHIQkszXxqWcrbtaI+cSVhCENp7WY/o4rKlG2NIy
5fZEMC9x5A7shwEraK7vt36OdJo+K8Jvh6Uog4QyyAcHDJYbn0ZIVHwFnk6zWm3b
0+s6Ktmhe2FIei80l6B96aEDyVHfcUH/WUOH10UfIea79JdF0VfQ0yCiX1ImTlvu
Q6O2QQJ4q95xyUO8cl33paY+EJe7PPNgVb3tkNHpw8wxOl9Jya41Sm9rkPC+oNtk
GQ3MyE2JyLCA+FHmjoa6YysGunznOJFEgY5P3i/0Vi3njSF/9kVBaksn2AfFNZBa
8BEH2TmoH9riDmBHUTf2LVRte8AHs+5AoQZNJIP00xdXftFKG2P4uk1tyJBNcHWX
gc6PdB6wnOM7SOx/E5LlsVxFw+9rLpl/cwdqwGxNo/B4SZXHSoKQKV0sB5jut6+W
ISdcJKMePh7n8ll+Icmkye9BPJq/v3QfAB/9A8zw/lSt0MoBk7/QiiHWksj5GRLK
6Mx3S/WYy2zWGpf6RPKY3kbkKcgFUTzyex5VWNv/sT00sXo8CiUG7Pyn6VkWLwSs
AdRauQ2hrqj+rlKoJOM09wFzaEI2Ajf/HWVy/ITMy6Mj17oArNujSlGCns6GnlZi
Lsq2nVZHlwvh1qkMdksnDf1m0/EHmtGCAWzPo10BAKmPNZVTiNOrF5UbAQDMDVZp
4LDXxx723eHYoyxEwtp8eTMV+H1Vtz4jMHWlyC4Atd0M7iEbr2OvJ6NeAIV781X/
6dBQ1Pe1zfzCcu9BQo4cIYxU4oqjHXZJ52hxImq9t+6SqPP1y1DBUeAxb4MygAJb
PKUytGCHpUv9Vo568/a922Ok0fabbKetak1tQA/OdjjA8yI0TFmo6noW7rpQZDPf
xIQp/ZE9Rw1huE4JuS3lAtUJvIXfwGZX+lnLwp0srw52h4A8XA5VPoPyaimZop2G
X2pqcnmMrEmnV2xFCiJVaYjhfRQvN/0aqJ+t5tq7xLNho0SrpSK7ZxT5uFcRWSGs
ICm1fmebKLLlxnsCLfov8fyOiULbhS2xdJEDIM2Hv24bK4HiJmotc4oNGhod1Nnr
u7iKcKqvgmNrxY9LV3Clq6aCVSce9AP+L1f8tUVY/REkpxUeLAALZf366AceUikT
5LwJFn4iyeRboW8zHzyZvFmFy3dcpJM4DV7Fq1FN+7ucB1Uv7dp2CQAclM1PFK3K
uFL1c3j/8UUQX4VHTWNO8wnKi74+lxb3Qqjvydf76S1KxQ6nyM6yWP3XPXkykGmg
x2l1wMohRb7z9yZvvlYCPgruXo/ADvTlvBD5tOwzL40kbi5Eq0hfRHtGNP6JxGp9
PPxxYDkkr4GrL79/tucBIFzHMhtWB6u7DB9F9K9Flx55F+CyR0YFR2C6fulakeLM
YHe4+WzYxRzgf+rZhm4X+ROQhjEiF89vkT7YH1cpVhufDeFbZrmyyUWm44SkhONL
Mjjrn073jE1/aeUemWZRKVpMWQg+GMLgXNcV750dU8seS7jwsnysmdtPaykXr9Ja
cqliNQVgY/7H8zQIqLC0MLsvkfD5JmiBHhSdvgWGI1Sua4kFTcRdAe1U3+MS+cuY
QJfCdVAJHILimfIYpb6AkJNJheIGGs2nkeRopiyYyQhCaZPXCTUh8Q+Z4xAx+2n0
mz5zZ/kad8IxxAHC2On/43NhKJwexuYEE/X9oemhuGyDFrwhzil6Z5vEqT+Jc3Ca
A+dNBkasPJDxVXR0WRpbznQ/Owxiqpm5G9yQaz3WU+tTWY47FpnD9TeRONE2aGAG
dfTW3qbOxgwgBFFwF1qcQkh/EPTLUl7GJmFV4Ebzf4Hqc27o56qBqH3BzZ28dOTi
G3w7VgqP8x6JW0K4VlKVxcEdD9iNyPVkqFto1di8FAE2l6TlAPk4FioCRFklZJZy
QDU4sYoImoaHQUMFEyim0IH6KZ5FoVE5WbQ5RSmy3u+9yqDkL/IdegdJ92tKNW57
fmZSjM1OeMuaG9JXbpnvYIWc4pOkACsm61EvGxQUXqVbfLdIMJFqCt/fkW9tYmO+
OeHfLuo/krn6qJJqh3HEC32y66KLw6YLs/Dyabm7MMCAuk78kMWkPYJ/VA1C8fJC
EJa6Abx8j1COye6gYMEKfSHVSJ6/j4as8BI9cM5Cab6qDXtxbp42kKKIkgZK/YvA
ZG7Uy/1ichrGNAFB2rczdKLAYugJiedphMUlFUUqJwkSruLP6rFg9lNw7rjrOKUy
cmqJqbJJ42UEVuC7mNvlmS69L/UDS8UcBuphbfsKX17zeE+uHIvIR8w44Br1CDyY
OWTGnionzYPI66yBA5Z6Mmant1f/4BB83ObJs/laqHXSFEM1vVFeARS3cWKuI3KX
KpxU/xXy3OogwjqtNQC88DTFuw6mw5+vNVoKOVHhTYUivpK6i+YCXPYBrFERWYMo
nLXtcdIiAbmI+w2YKZTyZZrL/eMazKPC3X/jSd7eY+89+KbT0MhJhnSM7gUuJS2M
RBfiyHTE3dC2bDtorFhSpw4rrEyCi/405NCyHH6lwHEKKEksFdIgriJgs1LFRNgG
1gw6x7fdk+vVG2RU5odaeNUD68UYDhmD196ZYYz4TrXZZNaN79mMqpvS85tW0fWj
7wl3TkAPk6QEkTHegIrJxSe5p1rMfoEDJvCw+qmDvaeRRxA45p6QHxc7yLYt0Ywh
Thsawk6OmmuU74yUkXCvB8c94j8VxOcPLnNAMgzN6lPtNXDfVsjDhaCGoyGeubcc
5+/G7rn+0KChiwj64gsPtiuFpuzZQEpZ1+4huMGKmNUwfs+2Zyewbn9tnLfSQrjx
CL9Itp7EHLQ6ncO1R2VIjpLKiM5MEDMmMU+Hvr9fMsaq6ywJEMkMRvx/on/nxcAI
bjYX9NuYdXQqnkk/kKuU5ryhto28mtqH5MA93LRQ0gT4ggPhk2PP1Ybdy/tF0fL8
8hCNH78QcSbv5cDYoJuHWGb7b4NeXQKHpwYezEDBshdp1UwdoG9qAiO5Ttb09lU5
7idGBFTDE/9EoD7i8FcQC8rEj8X1W/KVY0/enExRJrRQ4aQYCucOVMQ13IiNyYwm
X961+9IHNd6gsSAn7JgUmq3aNLdRv33fX6jLUIfofKaQBzWRvd8xjbA0I1U9fvmr
dayezAFDUkSz+RrwiGVr2tighBhBjlv1DVD/Ms+lGD68gEyWKYhXg2KXFfVn7t7H
GynPpCk0ZkgSUiwkIZEAd8WBaygKYmvz7Vaep7Bt3J2Nha/XaG9dOhrNs4djmhwx
flo82A8JYPuT3oPy3hAHsLK8IrqGhD1DgjBoWlzLhuZnwDZcwa561kyvj3A5C3dS
zc9Bm1E84XyqBR7Ua5RGM6frIoV3AuYHu5JLwexlVNECYRQl+bRAPxWjrlIzPChs
7P1BwQPuXfjW2xATxmUJR0Ly1ZKQY5HXSbYAkBhwDPyWrqyM1aK5aNd/heFvAX3f
ILQxYVLGs1SL3ACOK6y07pEU3FnMkvlq/wm+5pWwgJuEZtQSafzy2E/jKLemSvP/
+Dr8u2W3wA9AQ1LwtxFTSo75bUvFFqzUtmKFv8IWA6pUer2TZ0AZaWBCuMrTpr25
9LPRULt9i4dk8z/OVbYqZ9RtKEC9HIPWskyf+CntEh18k0POrz1engJk99Uo6GEk
2SJbfE7MeVAX0YEifdGkJPxJ+nKFvI3a7XStP0d5BItUMUYk39uk/8DKGP+vcjIj
YrXWz2S7b1S8JqzLtOetxK84AEdRRSd/Dxvcd3WYWTPzXnNUfUAuX9Ce90pTyt6J
gfYIgTi0+wBBZNeSzJjAuNABbOuP3UaQhZbhMOpIwI1GVQed/sXsbqnTe023nAs+
I8A5mMaoO3htvP/bdpHfvgu1ItQPHOLVOTRuapsvzt7Mw0xWbHr49MTnfvewHkVD
6eCzIKcJ2cRwv2yuTXHNAU92ecXNpyPpXv2aD1KXSRs8AYxtwnGGSInMRahi6hE8
Dw2EwScQs5YR+03zszzhfkpciWsP8/U6IPbeurI0sAgQzWAjb1SIJ4JFi1ycVFn8
BqH5u2fd04bXTNHybTpVZyiFmev6lgbfuLW7S1NG7OqeLlFnBSf5LkhfYf/tBH6a
wZRvhiuWFGavyrW/LhoFoPyGOiMNjroia3Ev347Y+zGW5PRDj9LM36oFP+wguFrc
DDxbRUtm/woV+urT50TJ4ZDxHPspFZYAORzswta3ATFur4UIYO3h/hByDOlh94aw
aOv/52zFeGofKyPKVPCFzFIGU2M+OyVhAZDWe8Y5ebr5CbWbH26dhCQm39aHt6q9
fi6fbAz9Eh0SISlHu9VeTkP3y/F+W2L9pP46POGC6vcWYyuEFb1/9YHvEXy+902k
FicqfqY+O8UJ0GNZxcFglsRp7rlGBMObhTq3PiH+oLCJf9QsRVsjwRg1quYNqeZD
rQIxgMdTo9/C0oI9+N/2aig9oDNYOsLXIJM290QZZU2RrBGyyf1VKGiOzaiK5KOd
Ei8QrVqjkUNvjSWsQFbVb1aPCzSt79SY/PUEDfkg6C+zU1SZ5DPSEowZj7q2EDXo
cFI6cZRn3dCZr493ie1W8e//5YDgmspBg2K8itK8G5r1DCWQUB4raLndRCt+BNXF
zWDYdWg0B2zpEjB0AhoXV+4iwPmwI9Ea6Le5ClGsbJIlVcULDE91/Wy9Qdx54O+b
5wX6zCCrfaJWc7z1pbng78j56u+INFLQPRRyau+eeTkO7pBijKyWX3+gN1oCxwS1
4ZiBEz2hbcQ+tHqk0wn3bQTs4goz3Kv+i9jIzHyMWkYCPKm/SA4MJf4JUsXIiThw
rDoKenOx7YxMrMCBpjtLeac3UIalW0DqY/3FKPvQ4c0ZPcBcKVqUDceTTL3DhIko
Cp58BXiAedJv7p9dnOR2Mgrc4jqMZUnsuTcSW177qCHhCUl0b5eb5t6W7BJKhtWR
MgI4cCgcigEnpI4LDFeLgwWHMi3mlsbxHfWrYWF7FLxnRp/L1rPYgE1JPzXfllG9
KHAVVr7d7/t4SZG5MtkSVTP0EUj62v01f4GYQkskidiCi16wUZx4TUJU4ZQcb3/5
1ftt6TePh/+iiGvWbs5VOAIHjk0dujbyU8friMNUmK+8HRzKPBX0z8cXfEYU0Zau
+hZl6nJ/0naexx2PaPXZPIFOCC0syu4dvRq/adZKOX18aH/RKspQ6nemV3jWSsB5
1VpMjqluwRYEPpjwnx881rcbH3Ro0QNZyYbSlQoEx4qkcpDBJ6h82aTzFBEFHIAU
diENLB18x57JiFrt8P1LUoDlI7+QqIO2kbEoSCzG9mmaL8hNfVlSx2oNtMTNTl6J
HeJpL0rVPX4fptH9iz65P2KOp535bf4jJW1+d69fsvPPJlJX+EJasQWeWKSeC09v
ArU9d2bjxT+sS6xKxEhXRwtIgEyfzaWwksZqk6XuDtUYxXuRnhfknsn9uFSFvRtx
xCjZ4hOEFeliFfrMU0aiKKI8xtslj4RC735QlGS6C8PJyyixc8cE1fTNwPxVsThQ
lltLfSQxoVjOanhiEkI83ifKHBeVKpq847B21jXBHgLgi4f7a8cSsJdWY8lK96yU
k0RAYhVVDdKODquVLroWxxtlbdNtrN+Qw3XrtjfMZd7dvscuFGf7qXpEvYSPbYTv
V3V/QFyKgVtNcDSTvvbNadu4sDPotZp/yTPhLFL+WdzfvhdyjnA7ABxsjoPUFFn+
5O+ZS1gdKGDD0KYz66JBeXsjFKTOE7tHqB7ebc/GHBFBus49JxJfTCdNk7WMNikI
UXtNPppThEx6XmXiKR7XGertb13rl0XabOB6drDERZpQ4TutsTmNvO417c0Ylp2y
MN47OpLm8tD8gAL8AYpDpbCkRT+U2oQj5ax93nwgNDklz4Zw5Uaijd7BEXEdjmXZ
2+4GoUPho2EAIpX2Rb0BSiaNp7v6KiBc74DS581wbnFxkxWPLQ5D9lZLgPhVC9XS
04Gda+GAG+l0KCsXvs9HqCJmo546EO0S+oiB3dfxBGCuCsxnNUlbMRDWZp9vanUO
YMRR2xsQ6NPrGmonP2f83EwL9JODPj9XHxWbmCN4+yamtZ0DiQ2p9YUTzMjsSdgC
3k6Av+O5OYA3FKVZ1UAk89oIpvhhe2AV5yhK9DNDHdyZX/a/ErWG9aK2dOdPABBW
yvcZHWurRc9mOkxHQ9X1WbiJf/bxAeaaYX4iKKtXH4xemudPFNntXplGCJ6bccqT
RSfdQ+gyXowfdBI1VElHrA4Z40F69Wj+pgFiKW5M+uBegK82gKjbk6eEtownN0js
8mQEz/P6fccKKyl86wXOJQ3+YZFGVuSFAmyk7n9V7fDLgnXIC3r9fVDb1cAlVUSM
WV+pGfIubQYdMWgw3OftKhi7VRDu9/hoAYktt2W5wmVR1pUMMq8XxoTxeDQ7tC6k
lQ0lip7XynpH9at1qX5r5uaGqT3ipPxF0hC5BCShX3aPHa8SwB1uMUUffwj+fnae
Ksxu/sYB/KsiS5DjqF8yejAJ/0N5nh/rfxjI8HH3EKE4UYq8/kyHLhlVNCSqFrDq
QigVgyl9KXBTxFtoYKxZvGPCaRiXjXbFAFpWZ+xvB3TGmP2QBg3Ei14aOpZEFa6S
vn0q1s8Yn5SRpGvceIIYX8EcuaFvHyU+qfeqc/va/gqheEm5Q08xqPusqlv0T3zV
g54B6Ag+TkSzYaaCTW3J5gEeRkxFxOY241aclidGEoq3D2hpQU2Y51lSpZL9vdAQ
T/ARvFTU2J2lFjodQKD+/0z9ZPgiPCgKL/GLTIDLopeZ8EherrO13n4S5/8V4uXM
Y/EVmE9bMZx0312C6K4AUgkiOaYYS7myJJsGi8wTuVaYDY8r5FU0gW/WKE+u3547
8dBYnuf52SOZn7JftlSSQ8VDyFhD4B0rhnRhoQ/31ia6dlCLmEVZWMUpBHdqgo+B
GuPh7DJZhWOc0CmnFNbiBYwE9PqrNWj/hqxEroOdYFMdXyF1Z77zoXxZE85MODyO
DAGIkYHawzt1/U3zKf9BGxisQIMVY+0E6YmtLqdELXQmFYxVNkdUEx1Ak/+2vC51
Kiuq4F7iPtj85I3rJhE6IYlcWQ61e92vJfvQnlFldL+c4SxweQueoJdo5SgL+4CB
kAS+H1TOlVRkK7RRe6XwR9deCjyHE9R30tBcrfoN0EsD/nVcijn1gUJs4GBmnHWl
ABSQ9CBYCQ4/17ZRPG2JcOpCnU2l8fK5UwS4bY6WLPfmX2IbtGSfUy7bk81qnkWY
0CCfxwxCOVXGduv4qqpRr3zc2533o0HVAhEdrI6AjihQidf+jfhSCnto/hh/1b0w
3TzMFOyVGBu4NOGRA73QMJUMMDfev0fA7Tz1FBALaPwHTyPl5czwYMz2gghZ+IMX
dbFwOVYc4/PAd+0ZG4y1Kdby5cXlg5ZnoIac36vX5IzRAs1P0VygtNS86BPkQeXp
BwowkTDRIlRPBzkG2TWktkfRNoHwF+l2yySVWKyagEZSrbITUoAhkOaUe99Yp66t
mJzLe2bMts61XQOzdU8ta5UU2goOg650//Cg7bqS/MnusblbDMQjjh0sP19SjvMf
Nszc+SDFG4AycQYpEWCiAZYFoNYmacsoTj4/3aTKY7eaegGi6cSfW2UrRS/KQ8nC
Qn05moe1uUL74iAObEKiqjIHoRJ1M1zJSIBse1gwFffHrLpqw7IvhU/qBY95Tr2N
WDFG8++49jq8OwWh41z3WUL4H1wpeS741RNmaUxze27dnv/zZ9riIwWRHuuZIZob
JpyZ4AOjzOdHAwKepVymFaAwltY/sYYpB492WNWGyAuIizy8VSTKtVjrrq1njxT9
hkuIvaPh/Ocliehfd5750B1VTMihKAtJbsCiRnbtKLjXPI06STIZrw+NkXfiEy05
rXR3ue2QUVZC2G47V/oKF48R0mL/9WMsbIrrj8SnZjpeVrzZBQoyV1hHHEFpMANX
ws0mXvs8HsdF5gfMDF2x9+mP94TWcNa8Nb/LLP3ynFm77R0PcL+GK9wmeWJrnuyW
tCsbjXxivDwJlXndvuoQ25e6qCbyELdLPv86d0ef3YOLvOwYmwsDPC2tvkx7tAvN
axTKJ1YcwuytCxP2LOisHNtbfmOnesoXNYXoIEhw6Oockv/Z5BV51rBMwITTW18Y
FMw+8cYz/eDAN6ti3Ebe+lHNUJoo8x2GNLNnhmOKsal/Ysl5Abfg8Qbv3H8BfwJ6
pZ1/Ww/sxYYThAwCPS2NS6beUkuCF6nWgJQQ7yZfhRRN2M/cXiK8M5iXerewBgLt
R5ZCHq7dhXm+tqjeq4/Yw1T/aH/zrSSXVKIM84vywk5kzrS5bhxyyFsC8LefsXx5
HVD+CXuHdeYBOz6Aqineb80BlCBWa3RCtcLvtC5U7SJmNevLh5Gm7hUgeB+ZoZiZ
5OyZgzxpdJ+mckq8GPxmTNE+IOY/gQSWON50A6yI5Sd/vHTIrGAZoE93azR8JvBY
JnJQFm2gNevkC/stf0oHPY5Zp2EXaHFbNyO+CTHXcGnqXVyi4YRpQ9Lp94l9v62W
0QYaCk7BBLWt5VkeGVYvHqvriTaB46C0lpSB4XNqWKKRw7l6qrQyGjtE7v0LyXPp
vsYakwwsTHz9lsc5tTUE6GJBjWEX/mblRTcXvYU5rYIbnJKwXyfM1EA96SACV3hH
cBVH/SFJ3K0GltJFbEiIxZGDbtUxipiS6+1QUNhut4GcKSIJ7KvwTRghtKGl8UTU
HSX0W8G8z0ssSTywurFMinMRZJeh9qf62Cxjo50f3/pNezFnd4s8p8PTYoEUUp+z
+hQDR5EjbdnyHsAJ0GtXDh4MF9c7PK8qxxj+2dJA68C9XGjoeyOPBI/FDo0B+hdf
do07qPl3Q/+l2xI+cepHI0bOfEPDIRcQ5gZm+8x4iybj/133jgz0mRz8lCtW8ZQr
q904vy4IXItI7L3wSD9qvD6IN6rZNKcJTdIQH02dBASjNOSFROVkdNBJJQUKWQtt
AXUuuZ/o1u7QXd/D9uGzkBkFhkSuRFc6uvmP2n2WaiOb5A2a9IHN+M8nFf6YLeBi
BOhgv+agHJsGIPA9/1VVCZVOI5hiAaC3Ar4SmYKcIC8Iegwm7fmNZ2BXrgEBDqRe
5WrjlPXqNw9CvXDzr/0yK+7yFDVLAtT4Bdrfp10vcwiXelLV/sQS9p1jlhIl97D7
2iNY7ulh10ZMUS28MvXSnD4FSj0c5UsojEXnzDczoc78WGppoy/aeO6x4jIkHq0m
b32XHzcAuDAB3hf9WFp24MXxnaVbEtKzmAME/cqJn6RPXsJky4DpelXmYYLmguHk
WBItZo62r2o7La9ycxMWh/ITDVdZv0sLKX3zCMpz3675oqGBemUHR3rVfNb6/NjA
Qwa+zhNbMf0MPY0oLiCX1FoSQYPWQeLuIIhv2iKoNu22jTWuOfTAp9pGdp9s4aKU
ppWp7i7n+dNDrZzYuR7h5YixpaCrHpqVxp2NNx8oMB9gBnzTs7t6W7A+Uvl6ftff
GNMfieXT/K6MvhINiG70m2C7baLUUJmjxXBN8Cavh8agusSsQEOpdieVQE/udN8p
6A3iFf3Gs0Dz7/CD3MKcls659RCUOeTlrtzHZKipk0mmjydQ67ZKqY10cdX94ume
7Vurh6EMtNXDratbfM5vjiNwRwpMiYxi0R1yQxYxSLF/WUibO3GoPhsMfz30POZU
VMMARmn2EJsq5ahnDRFA3uJsmRHjlP4EbbNRsb1uN3GRPoA5gkAnPCpr1gGKFmtE
UzWi8CB6hDXV4JIftYlu8x33VKD0WmAAY5OgT1W8J4aCdeIxUbQVdiQjoyml1zL+
YwreCEejjHu5a9Inn5ZuK6l4YmXrydr75F1DmtNy6IYNlgdZhJaTtgdfro5rcN6b
5VP+vg8w/MWjWhTWc+bp2u7oh7IDrV2X7l0YiAyZCki8KDOEhVSg8u/fL/02of/O
r9ALB0Mw/kxfeNSBezNW+K/DvikMAUh2nCVXo2EQhg3urmjpuDpnBgOx8K7cy7MV
BpOzalJRAGWEMhtj47Rm/P8+Ey1pkc+ZiePvd7CQr3DNve2KdHai9Zz8TkSfvbkB
xbLf9SnoT38QoIeoOmWuzvcowyRmeUvVNpjHwQ9MSQyWXgC2UBcuhOaPpaVJMOiz
vkI3hTp3uhf4VYQvd7Lh5+Xuhw2L8OQV0xthhVDfSoYarir60uhXncqIciDrSCXI
i4vb7XN8RCbLx7APGIaddxfyrJHP1UtnhZ2thLWiBtTq2UwOUr6RNOVSIU21ALaX
vrWFOozFOAb7I32g6SLertQnZl6Uqk8nkZ3DFTF5PPQ1ZvjDE7uwG4cRbvJVL00U
1qkEVT6GC/s3VcYCbPC8YwfuK0dS90vatky6DjWsz5SebY9TzHxOnZ8bf9RGWdnS
uzqpvBaWBjrcLS2WSVxsJj6ypTLsbZy752Xevhsy3kBRsPrkfKu3QFZO2JnPjRp0
ikycl6t2zqonsV8MeWZuMW/QogxwfcJdGBCR738X6iRoCLc/C//7xamxHiHKVYLk
6eyvsfTp/jpw4jbcL5t/p7GCJK4Lyy9B6PmlGgsCWY1UTJs4iCqD8B3Op1ISxw+n
vC+ip6Y7XXr1x440P3Vu/z/zI9kiTLTEp/1yBmz9rRX4meUpf0748hGJ1N4FfUW4
GBqjNBP8o2zEiCckXz6MYZWPwAcF1H0VwvIwyMwDs/vmd2I8vviIBECZlG9krPtO
V9EE7XzwBRm//fJhm/HOG89L3et+uwsk6N2kN+Fz7lCEy4UizDiDCrGV/Pz1mCiV
hD8BlYlnh2Kimfnop1y4UPA3kEoeaAaRifELiMrEHawPQ6AUIYNE1dY8YPZc2SKf
9PGvjrD2ynegCSfUCHRHodZH8R8Uq7S/c7KWVxhg8N9tQ+zZXDvkRbz7tdWztVt/
Xhr2Ed+Hp9/cnTU6SP7F6pJm95oyaX3pnxqfobhaGabS0OS6y9zlOVBWXcR0+UzV
izUpmSSf6ibVoJ3CpZJApQsxJaz4T/2xRbZNVTpXCq2K5j4ReDjcbiVcDLm8n4bR
xZjofonT4tSR3H4Hga44V3A2hc4PQFn4RytU22uwUkBb9qyqU5w21PIsL1qixSkk
EknD5uJjyOhEDiH4jcZgweDntusKYzVpb3hYPeJXaqLS98x/diqX+xynAbo7j+dn
F7HZ6PDQ7IwrmskYyVTn429C31xA20yayTNHZvJxazVUvCb2An1eCgPb2NoaXJ27
vUcUsgxmoWq/8RMZ5Tpq9o4rImYCIHiWpFRZ9wslyk0i5qn93+e9tkxXWmK2sEtz
SjnXwW00mqAhmjU9F+BMAFyyrbBBA8uyUP8hIGZ2rSEq5E/hA5bFLl2tMDynl0SZ
zMobNuPBD1+E+cOnIzP04VZz1qGmckJbQD5lSXfl0JiYq60XcHJYQ/8kYR3498lI
BKeZHQWmdrK4yjz3YATG7E8mgT/db1wFLeeaEevXos+8twk/pMiyJ/bv3w80berr
vsQGoJGb4twf99xFcfg+3MxJwNCR70xrCK9zP24DKEh8w8NEf+wml6Jb8mYmgL2N
8mxEum+Tz1YbrVkWJHf66Tzk9xLDxRro8Xq/FEzGnWe2f6DkRGNm1WXkQjeGY3BH
lFu9a9ybXIJ3GLEsx6WsO4cBuMh64nQihuhVz4eK2mWDCtFOv44aaZcBQReYnAJ9
3ldzqAps5Ziy3tMTTJmsGK/evMIIjX08hxYoEFZLKc/MgepZKFjoScfsM0YboSj/
JuNYlRB8BSNIGBSo6021YLv5xzXZWGsMwfcvPcIBDyiuTePHEHU7J46X7Ngvo6/M
PGLLlN8vNuNxAsOg190yMi2hhE56hvkaJWydORZGWti8rYwDBnmvTcwSH5T9e5ef
pRJ52ZIXEjli9lXTQismHXtF2EPeRPVLPFOwQFfS2XWm82qQyME3x6OzHhcS9I+p
GRcQY2AmuvRQZ6ijkgU4FY3Unvv/lErP2UIHy1fJEaxpi2A0oy8+04Jyq6JL8UGx
XaiBEMW3iG98amMSV/oxooHrEnQQl5PIY4IQaoeUH7TSMbcZZQc2qytnwURNhPfs
HiC5gymbONPjbMBcphqX03G93XefhiRbualbWd0EHdfsenLnZCEflbrjaNXZp2rA
XTvah8lvrUxg0qHsOeQblinHJyAmYDBhB5Fj1ETyJUEryflOaiR6jSdrJSXQtwIx
7nBlpm1IUCei2FST3bbSjX+rK8eNtQ/jCXAxVWGmLgTxpdqrrAAS6jFKabzyXWm/
wKCmgjIfwpRFdPAsKxGPJmnAKSUYpRaJj84by4rTjdgVULrM1sGg9kAc/LemRtop
HrLGOQ2HyAfC8Nsl1o5mp0fxU+o9S7z5CrZZUB0BfrwJ1NulHcB05idP4zXrSZJj
bWG7CpBqZUSbwmHTNYRN+CMTdcwQ2ga2q+0hC5uP7+13x18QbxaItxhp8cc0agq/
8PlNo6YpL2PGWujGsnDERZo7b4Zeev0f+DMvq5Sz4R9fpoieSdg3B1dYs0fpqeyE
Dc/f0ym8qKxJc0b4/WfH/055lBlNsUz+MZhWIPUpOysYmXHUGk9PzR+ZaJuSyb7R
+O0Wntw5xZwDkMMXxTr5rhxLCQl11pEDBifF55KCErn4NfSKicXUxC+u+X7/34ux
yuNbWI1wM9UB89vHSPHvo4t+aWnmvivVQKg0yUrexW4/j+J/qLf11CuJHVTmwUTI
wIj0GV7MK0Gk53Opr8JYu9A0KiXGfjcUtSxMGAXfVZrp6lp8M5EWxmJi1ydl97F3
g87WNV5bn1nrlAg14RvJwnt1r20gl++Vz2N2imTo97knmsRfVshSYfAooNVJQ5cL
jhiUQM2hRbJAerNQxXsZYGZjf54FjAbIJAu79BT0vrE1vkctlkV2cZBzkzCCTUbV
84muPGoTht4LyQ8F1i5CJeL5JTmO6csLHb8W/9IkzfLbLvIhddBTR7Ztq9CtVmVM
2ewBceF41yLBJg8Wu4pGdec9I3H5R2tiLrg4l+2WlmotlwKpCGa0l4hVG9OQq2GP
dqQHaMtXOAwGYhP/cp5Ks4Kvw2twzUZsKkKg6zFoJ5Qhxo9zqa6syGvt7qAfk/RK
biJaBJqCKZ1G8HjjJ33Q2RI7HgScby4d6rIPn3JVraMa/e4rruIYHc+hbc/pBCm4
Y6zfpbUCWyXiK0jfq88boDPv2msTcGs0P6XkQzjRpwA0lMtbam83obSb+FyUOZg7
grjwgfKUMYgCp7JzullWDv9TQBv5ZOW6Mzwq96wkKgme2ruWW+InG6I2hhUVBQ4V
59xleMCbHmT+KlJIlrl15rP+R1W26IrfSmOdgX2uxvvZ6xMICb4xx6Qu/EgJI4Ku
5NP8CvOmzq5wc3cskyWyAieBXiAM3ZusbSG2XEEsQ52u3KgPIDqg30uyl6xenVgh
lF/t0UARAU77hlHBwcOH9GKB2yuampNBglcLj72gdCMRCp2aKRUT/SaCBecLbzi5
XeLPgyLn7XXiat/WQ6cLKqWv2X83NG5HSsX3c3HiN9oTruusgvorehdRXRHSQVR+
rU3GuSrTGsSGcUAY3e/YQE14GOm3rKgWPJSjN55YSHmxpK71af/63p2QqFFTKwYq
yHjSnEknxRqCjcso6DEY5GsVNpE/dB/QQdxam6wE/uRNXAI8URRz6ogDHO2rZESb
eyNO879GHvD4L2PgijBOy8HWnAO1EqpJ/s4e2rm+reErVwqBzaVaGJKPHIWwAPUT
kO+pvTFYe+0FDUp6Hh8gsTTUmE8J+LkvY0txdSDMgvQ+MFi58InpnR/ULakoBR3e
hau3bLlZEzWfcz+0Y/HkMmCPTAjOA5wNZoZ/bmzS3NvFa3sxJHr+dSLUysPWUU4Y
6GcJKc7PCy8mVGZ3Y6Irn+zHWsf24I/L9fZk+OvUi7begzifmOe26ZtiPkv/JFKL
T7Tv8Io5z/zaCYXoJc8a1woByaj53WTRNe2b8DazCYHJqVu/sQqegxgIZL1QC+KU
NSsHCsHZfFnPP7wgkxKrBY0ow3SG0NRaQ7lyUtWS2wECzMx4f2Ul/GVm8VfYJqD3
QjWHjy7QFXkMpS3sjHpHlSOKfwWWaN74IvQ7KuhmPxyWBMbNj7PYL40A6Y9aDiqN
nnyj2c5o+qa/+zA2kKBAuILz0oHsIz4oPVZ3CkGHK+89i5srNjTO9wT9C5ytj2Of
f8P80bxB7uzq/udHR286XenV/soLp1XibMd6TZ8U6Yf/rJRCbbq5TqIaF9IH5EN9
qm6Rgbr1NbaIjCpZ5rJ3rbV5gWQcPX2MF52kFzGFH8XA710jDUnI+/99i5UclaaQ
UAZ5xNHdmDDnbDkouZT3R2hIAvI5D+B+DHTYq56hqpSobIuxsh/GcBsCfwYD84A2
d7YMv+25mp2uGqm5ME0aeCvhjZkyMIuwbGwVqYfhMzxXX4jCjTyQHUwWxxBU3O1w
X+gg9LQ0ZlEcTVPtgknZK8BEUXm/EyA6t32h1P1oODusWLy7HOwnWeGmJPJ2s55R
wYe9JJ1h5M1DDKnOve/PWVsahezX/kXoDn3tSkt9iAAyxAzkuqn1gsRguiwcasu2
lsztxFySrDHxS/TRTK5lXIPwblN7JiaKBUWM4uZPNlVtoIS1F2OIXBqJ+Jceh6c3
3KDlbb4KhT8EwgM1C9ExpvlYUulWHiMaz1hIaE4vOH5BL/3XxrDPSgdR6pDebZXf
hNGmBaO4Jrq4MT5rWH09AUrlJE8zjJN8a7QLz0izgLK3S2ORxZ3AQoStCtdEPvsK
9rsVSk/lb16Z4Ut0cyyO7/ilA3pHC/5GRyMdeEOeYjFkS77zJdR9ROumKaO05DBX
D5xs3nVhjqP/7lTOvRjUNYAwJaJnC0B8Rg51lM+GPNszyUk4D0O3gnSC35bpEPNJ
r2gO9yH7Co1ydisDKqo4OWG9I8l3R1vHh2K2WGW8PpL5graCNbXUqsp+Dxc+VE8e
r7ppTZws9PLonxrTlrPfSROfqPpanox1ZBN+aqRfvUF+ystRWhiSb7aCiF375zyh
P2dXB1FtkM2PnOpmcz94A2yeFVp1ZgiyGA2qiWVhJkXKbB98RL+qUd/IEl36Nt7h
Mbd/4FbYJjqnxGZ6QINGO58PkFrHgQerjiM0vFP9wWRNpu36isv+BzyJEynPeJvj
+j0qk62WHv9/PZlMySDI6wWT0/Mh9VCKNQ9fR9+DwwLVbw5v3nu7m5FvfL8+K7wE
m0EmymNSg9b0vUO94ATarzXp98dpmkLpmW1/mlkJGEt5KkgvoDzLoZwdj30WRO22
9sDm/k+wALw1lmD4GRFzZz3J7eG8CDhHV8eX3O5MBjAbFWVRpwzjzzUQRqbrLcOz
5v0/9pQhWcN6RVXaFm02K3kDivwU+u15ZycCroL9gMfN88hwJnGkwOtey0H3kw+3
p6hYaU3c6WXh9NZsrgWAC2qZVt9fzx88aRbpN+IhYTMTYRM6aOIljDXvvaRrTdOt
9njyMwaQcbhVUda0ztKNPZIc1rwea0O/C9t/Enr9YuLKhGnJpKJVm0SXovQQsNmz
BFRPN9bhvIGrNTUZRNmbelbjcl9yysHbKF4Gxr1ol7MycJI6vC1Gz2+aFFUgkfbt
pwjnhkarmQysz2puzkTJ4W1CuVcJaiuQI18HpSFAcNkzuudqX8ugF4JLWkOLSoYg
/2asTEIsAAP7lLaiole63Yck7y/Td6cI9BitlvY/cwp81Ab3CZ15pUB5Gtb2boQG
8jzMYuE4G1fnoBUqE3fYCBV7boE/Hr2EAt4HsRIC9TtHAL+25czRq02KBV2Y7kVX
E7F1pzBYgHeNYY756xaEqzaiJxyquT3Iuk/vSeGGRCJLA813VWRKybs+o7yQmDwP
/chUh51amfwKkcxIOVcA+Q/wAwGb1LZMlQ+s7Gcufk5RPkw8v8wLjDODYGSXjdKt
UveQrAYAv8WNP5VEKX2r7+BVWFudKQaI8MPZixgjVXcDUIYSJGa3X7TvcMqgi6Yp
XPoVYS3X61grGmUAXySFsDHZB5Ig+L8SqECUrl2L2L7Qn/BWhc/vCa2TiRGRwxk9
IxT7eua6IjdOU1xooAd8RhoKNcbu7kMQuEaQwDBxvv39pHpHq/d812d5WAIta84H
ptRFXZCrMYIkIDPj9yy++3lUGAmGR+NsoF3kZwypGuMFVFdoZBl8QwcruP0AS6oR
iLSxlMbQ9opFA+MqeJ1eh7xesz5fFklTAaECIZ7wHBiTvYS2WZnCy6aFqgrorAWI
DO8yxow5ETqxafPAlpea4kzXL4NWLzTAy4fAL6wRFbikBFOpLyX0hBwqg38dk8kP
Zivqez9t3X3o9Yz80OtXCTfO5peT9vEWadDknPu+boDtrtv2HbEOg4TmtAgOtuxM
HvCpbXIca8NVyD0iXc3lv1uenRSX7CNHe00ff/JMJPhac1f+5VInqfXbxnA2V8TL
11YOeQ6osgjvR7YRPsFQw4xjPh4ni2EfgNk5m9koQiJui6AxNzTJSCg669aK9E/X
+TjKz2ZCr7KoSiUhyHk0pKUQ3bm9eoJDphmG1a+8RRwQ4EfVzD+OdTJX5PH8+ZG7
fwc67/E49ih7EpuwQJ3jclq9aOauMT0l6+yhDmPxk5DFi1tB/kptTOOulpa83z2q
Bss4kkHcyPf8xAhOuQOCmnkgZV70VyUG5MaZegnuAbbfDMty2mRyjmLqRPY5O1S3
ZaTOXGEZEvrA4JMR81GtjYFTtrkGee8ckKYbtsVcZQqLcMWFcPiy2SsrOqKwUwdl
T2v2Zxk9RNBFWmfr7mwXicgsEa+7djhLF5nD1NZ3eAxGPAX6lL69MssOJ24O0Weh
ahvVkXD19uwq5rcPvbgW6yVUOPaeWUoFYchm7IfQAXaBRf97iZdPqOudYWgkRYKQ
XHTPDL+Qap6PNUjJfQ5NrNpl2Tl0LRgnHDdrfBYkWaFzikQWDZ8/2JsGxkccxIZK
OSP1lJv1iEm7bhXMre807buPuLUfwFPGdbbZw5T1Yx3umL3EofWoH3BA6ScY4WQt
NMcmHbDoxUDi3NFpcfoLEBRDEi8WkMmnIgoOyqWItnEMpuV2Np71EViP0uh9yell
8rOInT4w9buhhxDBCLnd+uYaPkQ60qv+R4TnADJfNIVmbtScfM/fb7gWQQ5HN8te
io9M7qsx4oSEBU7LNWxoMzu7QCmGoqjgNpftqo0sztcvfZ538u/1w1v0W9MEfItl
fZAF4S6R3ii77hZgx8DAFH4fWalbuxq9thDlLAHnAX9qXZZnIXnFuypSVbhwSq7f
qTbMuhnYnf3Dhao9wPNa/QvLR78FH18GvsbYsixNUKoBh0m20KMC/FYAJggewUcr
726rx5PONPEtzdEPGraFE6rJVVk8HNw2y6DlQiB8asJfH/af8zPAHp+JiyZVQw+T
n++8Rs/iHu4vieoEUznrOpRut1U9SB6A48yEQp6ukg6MWqWGC6zff8LZGcaMo+4v
8/UidxJ1IbGC6L8shtZ+jUvSTeYRsqP/VZ7idIFjhumrvJi6g26GFYVlJ6dm71op
m3RyANA9SRz5ihHsD/qOREuKWJ1+DaYJmaNJyV4V8QA4hl5kY/fQrnY5YDjP56pu
hm7bFRWDWe2aGmwT1Z9a8f2ZwHRUBnb0Hq4GAXU+XMw1M2C8VXnnzz/Zyx0BAJQD
ZOReSGXkrtUp5O4vqv00DuVqBbZlwBHNlCnrqiJK9Kf/r9HZrh67qjsqeIXR6Zva
kh7l3Sxy6LyA+Gmzf7KUXvK8VfJ57o3KX1WUdBOynBCloJNzriJTM383U4xuIj0+
p+yHCsZuvm3fdWEceLkHitqF8USKSGKUma+6yIxypE4xpObqrm+LxXjpxNccLL8P
N81E+BfUMznChW602mG68rkOKRZe4ro8Cd9scl6JnclgBhVSnwjX0+AwsojBhb4C
XgLeRHRO0NkGx9/cTfu+Znnd3r1Ew89vOEePGCeuIxdB5BcPdXGlTB4Ri01vhbBU
v4H7UsXhVCFfQHbQTjUf+d1o5VwVDHX1o00gCMoDiHI+csHNdqK6SQdAW2bxpnKz
kN1kj1pZoY3TVqWOjvGy7wLT4w3FI1/nyUy2+vQb4kJHUVmqhornP3SplIznVjGJ
GpZHcc4+c1U1oYVRAP3BoeVyrOdE2nYBtU6BZUXcffhhntbi/WsTbfqPmYPZPrXU
j2FMV08dSZsEW2xBZGef/g9XUvruuMTzngGphKU+X0NyBz95btEATsRINbXPbgif
5xBBKToVNb1BBgb+Eh4/XYPb1ggqCbbjQ2KkvWmgWrgUM+0SUKLi74t20ZKfdqHO
H7fvyFvc5UMapHrgRFO2eAIgo9esLadmY2MmsXNRgbdaXboM97Z80neor/u2sy7n
M4W5Wxju48OaomRS9CQ3jkPZfxxuO0VYGiSobM1i+e3hXmahwAXpog7+2VnTziij
83rOqoOu6svOf3vpEtzbxG9JVDMp0J4nl2LK3mtAb13EJN2Pi3KE8hM/0Ct0pTWR
DeQPVnqYyeZ0nVHp1EXYNVBmn8CrLwe9pYPURkNq742pW8/HmJDNmdSgypx8jXHK
6aNkKLsYrAURxS7mY8Juv0C9qBLaW/PZomGhVSUMv/2Bo20cMl9K4mUrS6Fbkvfr
i/sL0YSRK4b4P3izj5vbfqqatTRfh+wdeOK+MCLppmZxn77bTJjVgZpaCyrF7LeK
P2SrBXFbBEeNc0rWEzojczWEiRdXChtlM2ZD82Gir56MnxuELkd4iTUQhnGOj/MH
0c0+0ByfxVq8hf/0P1+6VvjiGWS1GFQAHZ7bm/+KYoR0NdT/jKmm598oUB1ZWHS0
2cD8GwXpIqHpIwRrBaqZjCWbdsnnRVYO/o406agJkB293/q/6Yr1HWI3kJqm4b9S
poa/7dnFTs14u3WGam2e6o9/zO6noYTnsb2dwDsQm1TtV/kKrJ3ZMtd4kCZK259d
rk/Oi1pI0njxtTRDUTyxEoKRlvgOer0yImaoixGkqlmoaggvKCcWEoI6k4y8izD2
4hc3k0AgOaC1sp5F30HZFapIf6OaqWLFL4g1KP5oZ3dFkE+tsQ93z9weaT97NHmv
l2VPtbhF8kF52MiOVNOEyTTL9UbNgbb82LOIHrU543pHkHJgjvPELY9ROucIVSow
XtrK7aMPasrXMw+VC1Xle0v7u7WY+bBCsNoM2mgp9gk+g1Vg+aksBsOPxj+5Pd+g
FUWNaO1cwmrBezR99SK89YjSe4L12PZbDD2SpgXR3OXEW5E23Iegx1F5vWDndqZy
Aj8KamMUxmkOCLU5Wivreqy89pjc8KfVUevzUhqe4G3iD9pLl9qYPgdrn+Vk2cW/
AczERLsc5h9vXqzVVg9ucroQwO179Ti3IDnLbaXxhkWFk+xctPioWcuBbZ1WOuvc
CaPVPSFjioEauAEFXf/7/qTDpeRrMqN6Ykce2tS4PL5f5QRLvZ7U6ZtdyXi5Egy0
pEmXbPKZDJnmMJZXxzlOBO/CgoOagbasYlQwz39SsfKScQ7sYVp8G+AuURfFbzVm
UFb3P00nTupLw7UzqdhJiXtFoGm7PR/n5HIUChdVJPwAREQygEddMIRfJ17Y15PK
CPfVabTQMvo4uXEXl2kx6qPAw7uIzmKCqwT6yMGQ9837h/P0I9stJ0wq3HvNPv2e
CNBQVDKSizkYPehQHS4hPcdo19jblj1YDIj6Lu2XituBDAwQUSh5t07KfQWZNLSk
yubawcENxOuzfONWSb600uo6sRpZOOqVWMxGDFNN01Emy4JWQa2NTlBb8RzDIYyB
irgSPceNhcBc/O0TzyEt6N6V1mZZJBRdqPGHaTn424plNDGuGnn4/Npu/vRj6VdS
rERxPvHTMmzVf+qUAhE/lMLYcp3rVXEl4LqryQ5Bt5Ya6H2U0oY0cVIp74NkXYY9
S7yCoj1fhsiMynWx5SLVIh9NyRnpz6q7eStt9Au/NCSMvIVZG5kKyAMBMjI8Xijj
3LMnn9RVgch2YeFqwIP6Vo+fTIyahxBycL0QImv+NyR0LBwL0gdoDvopC5HMbHRr
6DYL4b2sZ4J4h5rxDgyhjZdg5f+s++/jHaj/YWrkRUDZd+dIU7/hz+i1C07Zbqtx
HokIkZiuH3bI3/rdjbBeIVmzW/i02rWvb+CYVV2bPrQ4bNNK+Elcu92qpfUcZG6z
cU7EBZdrZa/dbMEg4SzejvGmHPn61ZoZtgak8vkpHwxmj3twUbUjLFMBE5VZVePY
AM3rXXfIsTdyMG5K4ylDb2+qxe8VvZFqEMIrR8ncpc6fRLDao2a28uvXRMvnTXLl
c4IukV7jTQT30MdhvbQeTcvHtX82/tYAHyDf4AeyyqQGSxBU47Xa5hhV4dg/l7OQ
Lm2ZxJmOweiqfgql7E37lcsI9BSlI+5Egz6+lV4jPywfs/vz2vVztRT1TAQCpSfu
f3ue+xNwghsGPCplDfzAhx2TQOevv1QR+/tX7x2v3UtYwZX2IV27Va5w+miQ/1Od
e7JC2Xp0dhKVQ3qslzghK3HBHdnpZYwm8UQMAa0WkrroSu4pgeZGbOJhKBqSjEVg
y0QL6vpAyb48j64FxBT0kP5sxmuQeqUD/tULdGe6amGkz4e6u/34Usc8LVjyIaBG
J1kVHPKMISeOZOwZ2WFr1gKg0XWCBEB9EuxPY1RB9oh76w4/O2u+5F7Q/Yey6yBE
4ugRMKLeLFHxVok4f861HxV/F2M0B1ofiqozm7YXLpqutiBOq9N5YK7HwRscccYx
Cd0xwJoZq8AG0Vi6Lq1iKALHioWdziloV+q/LbWDZdmjWy4Hquajb8fDZw+w1ktA
igqFZD7OEw1UX/LC1Xj9EcrnXJ4YtzP6BY/24XmxAWY446W7ZOd/0da/6Co7K4kx
xbXBHE7A54nnL6YFiILyvxtu3mCgP1l6V4f4t/s/3DxZXz/7kL6PcZm/Jtj9Zf/E
r8fEkVGmN6EYrOzm9RIJwCR7IYW70Ngr+OxCF2UhCKWShuYyUjDr48VYMtyPk2ch
FbL10xYyj6pVUifl0aN5GNS1WRdkwrB2hsGKqF/JHiDmrHJlSG19JHSPIkrnFKs2
oj/+SoCaN9NuZI6JB5QIyrErDoRFeeSOZXv/PKBwG3hI552QtoTZyHFbyue3R/Rv
f28izANHKunBneWk+JOjiJF7bxBJEzpg0A7Qlb2UAgimvUplIOekiQs/6lomuCAn
fOmVewE60AfSqg+bRn2O6PiBF7XJr++nbab5twcBGEBLSZocmXlEtNcfBDc05sdA
Z+yHQQBtGIZBAI/NWr6j/H0uwhXHy2MIybDUE2wCtlUIH7sRxXTNeux2ytgzobFA
jqU52LxEvlIn2edS0XakSUcVCpEHfZaI16L2ok2yStqe4Xh8Bsp9sq8mcTO0ZkLC
ANSfc4YawajaLyiY1Td0SJrZ+W91P98kareI3R/AsZvJDkoMmQB3bchHiuAMkCWb
otQkRuEf5Ed7N9cVoex2xbipAgiPGlX5qwWqSF9pbdhwKw8xBl++5BuizvRh4NO8
4ih6p+PEjP9xqGx3wBEhNvVsW5jzXf0Mts3PcYjs0BgMQEe0uzhzbg8C5jaUzTsr
6bki0xsgM/LLMFvd4zgTx8nb9vCP6gXZxbl91JW0FxoAqkgGl804XhyXxUfiBbAS
9+SHyTb5zTANbi0A+Kmt1kAgXJOm0nRqyzIdP8kBq1f+tkHrx+BXLKUneybC/2yA
2Bffv6IMqc2CHgebjZA41s+K+JHebcwLL9+beqTyKn2UJInux1h45S1TOYHKCZLR
n+VJSgSPQOlaPnl5LIzLh9ulzwkOLejPz45A6J9YIYgk33OLFIBHDtPno8wAlYDn
Vv0LSmsYBNnU+s/nHjpaPpG57Zklw2E3GYwEaQXigp9M/zHbsUpv2XZGqyxXnPfA
nF4jwOdpjTZ2X8IDFD1rIVPSsqQ1BMj9P/h4Mqljl8Fmds12NwdzvjuMTifg/ksR
K8EdSW3Yq19V/+pjGeSCntfVjkIQ/yHcZBPwVR86q8C/uX+BK133RygrY0+5LZEA
LHQ5vA/TUMpuUlx5lc3gGYXesEZjBtDvHMAe701vy0fn/TdTZQp4J138MAvBlXMn
qgwfveVur1eUVkTTjKXesgdjYO0U2Wj3/LVARm3WBbS0L63l+F693EgxbKa0E9sf
zT3IsW4SO+PqIamiyjs6ZFKGxak9pq0XdZ4Yiio24IL0er/NksgiOpuL1jiGiIxf
Pp89FEPqk6GG/+ushgrEcbVc0g/aBArD2tTCZHL/cHLgdbZ8vgCoXEEaRTwoGCW/
uddHZAI4PdMFRIYbK59B9ZkuUYqhAkX+rDOgXvgSUzXkSNu85QaagIIa4mzKcrRz
UAbW7EOMMPa1s9KqSSJ+2Szay4LSdf5URMtn5BYxUxqi+XfCBu7kclVts3RyJQaR
O4pqQGcE7lZrvmec7ScNzSCoJDdLZrjf/brxrrfpoZjKs8GrMUXVA76nxomsuiR2
dC4lO59p7vjbH2Kflrq7riwccrAnU1JZ+qL++6yWR+hCVzqMGUlNsR8bawFmwRaD
IjSkz2d4KyomQa0F9ZY8U1DtqYmJzm9S+v8ohfEzXaWWU7uWmwc3t8mKABHapGyq
Fvm1lhmrpdEyDNsYJDwxR7AsZZRwvPoH0r8EDkacVaJL7LBYG2a7ChP40if+IBPF
IF+ScZktKikiN5ExulOZGDKGDRF3e27cLGRFOYGxZ7oHEHjI6zJ9g2FD4cn1h5E/
u4pIe8qA6gEnhaM9PPJyr6n+BDiFODP213Dis2V+q5PNZU9FTWsAxBaeD37LvnrO
MSmPHYVyTPgAoQbPLzCYbHc9wWWaGUTWIuhnO8V3O4RwzdEEmSuS/6TWegIN/kPb
KllvUOMPjtHfoCAWq3H1q07DOoF4lajvquL+CIXOXIsK6LluwBQpIGAcaU+ud77t
58H5SUx9aLq40xiJbIBc7v0/OfxfsP0+KJVM0Het4pFlxu4hJo5W+nM9KxCdm1+9
G08secJ9copemvOAUp6UeJz5YW0AGMHH+uG8+HKoV9s9pjcOPMlsV9igwn3nN2iq
kyLZ8uRIDJy8GnTfshEfFgsKRJIT4yrxqw0B9UiK8dr6rRejg71sL59+vzT6IIt4
Um+o1WuAiiycpjNFVENiG2nL6fIOk5OJFLhf2DOuvstVzuILJ1y5US5/FI9aMG41
3oX9DRwo1DIrtq1UZNwBOqRAU7m3PI2qyjrqGhWrR1M0tzFTorshotsU1OvsZD4o
8nom0cWmOrzYk17AihIPsGRhFQeNQZXdY4nWAiNNgAtqQvkB/9du0pANSGRJaK/B
xU+3CLQ5jogv6Hu5v4N9TV47FjvO8HOUO96Kz5QSCZkMhvrLKnxLwbv/SbSC3cHJ
2t+ETvdRbQRe01hKPdE70tqiO6IeCCSe0wzfh2OaYIjrwWx6e9o9BB9HUX5sr276
eB1QfkNpia/sfJ7+BxuKMeW8KIg+mNmwZZyj7zzP2pIrKDoZc4xEUx8pvigZ6XiH
N+F1aFlor6/TiNZb5VQGKmSuMn7h6saKZjkiWy3C9BdkhPzyhc1i0dn3CVEasvbe
HOXV4n934R+wExWxMuG8zhVRDOhmGYF+BXZL+LIo15wRfQ9fbnStxsJ7aX2Nxb6R
fJgzT8yxnJ0hTGj/ar5EsUEocZBUtTwUKNtQ9rtt9+om0PfyISXtlA3vuh+Af24u
3f4XPRJJJnwcQeMbd3vZyOY6Z94EgNBW6efP74loH8QQNlpsQlo6dIX9Ics5UKRQ
capHjBFqnurOhwXLnyZ8s2lug5eBFcEM/LZjcMRJ02ZxdUbX8aAolFW55zrfEfut
Rylz9nmKY1/F4vvsxNeM/vaxR4nieurEbPPLb7Rxs+BFSlwaDW+A3l78RMKRTZMo
1mMl/zYkszcBc52JcRW4QR4AINKXJzfq5qMxnzwcRG8Z6QdDyGuDRD7TXsigOXM7
Wuj/3iQraDlwUyQxh4v0MtE5YjzsaBkYWptHyK+0/Y3q4sNItz8vAPCV/wThCtNo
SINN7rCFUl3mYTZ7w0a7O3oyCy/tWH8aJa3POVrPfRAWFyFJf4pS+TLgIyWbaJwR
dbmSc6+t2/gL45eZX4zVJ5GZnzOSE6UYmSMDvojzHEiWJnxOnlCFsjTnZvZdgvlC
f7zV2rQEbxxLuzEgVWyrTeD33usGI2sllevEBplo9cvM0OlYT2la3RCZHk1MnSlh
+DGNqkghJR0FrP4PAUG+CFUnwsYbxZYOR9tryiFFOdaeLdQgsExDZ3XtPyAIJFvd
p+7AWXqk83OnhDJ9S0WxCIOSMEWs5kmeVcek/mh3c1RgNRpMfd7GXXWZy/1j+AWG
vI7fR6/W20heV46w20DjJRZhm1xdzHYCwX4e+9XFwQ3TRM8guZSG4W0db9nL9up3
i/pgLz8s5uSyETPA6Dw/qkiSCFkb4GCUqFrbbhg3yMfr/G+muF0pIQ0SnB7c64hh
HGKHtyyZg0jBDiz4qArJMTI2GQFPPCwAXr6ZzyMzoW7c4XCfBYPKH+z2ZChj1jjE
NFKdCFhKASjVyvmz+RPm7kQvXjcwv/WncxnX6m0qbr1tRDwPDuNFGFGhSMDbkuyr
CpW1T5LJlVknx7E3GDM2fioiVQNcAYc6Rja9nXXtf/s38iRg/ca/9t7EogF8KJhW
ueo5vn3ZllVS12TZ5mxVGNomLx/exerIRtRj73z23zjoY1Ql4Fjw8QMfIiI7lgGW
G6uEbX59qrkEYdbmhuVOtKgMutXwRCVGpjpsLe5HtZGoz41PuLQ2EYVfuGNuvwJZ
iRgISxhUb+A7F9uOXAfCnnhJ58m8UIHp1ffVHuGpuOS745YFs+2MYMPPtqDMy/Qy
HMcdVJPdAmdwYBjiSvnCO3YPoPKzSjHNWVCJucLH+V9AbyxyK6HxSPUQyh5UZlS2
1UamhzBAiKkeIcrWGkqJnFN8A/JxA9VBN+P/kBtfVfdvdHFQ1fiodIXRYy92UI2C
rrWgkPJ5PX6iD/leHku6tJzpdqB5MZsw9RXaKsYSs5ugrxzi0iASMjLpPEAyhKGC
ChOugrXk2QOZIy1OG62ZUlqSoz0b64mgzb+89NdC7DnefeCiU3xMI9EwCK+ggMya
AEk1bKOyEIvG7yP0Wwy1EzolEXXJ1kuRbsTiCKNWaI727GjqZ7+NZMtb5KSpTras
3ejvJJLZmRjhwgElN7CPTX3lsls62zxJc6IEe5GmYyAw2Uaerka92tZXOY6YZlkh
7b4DN925NVkuJejYilVJmhrDaHbkBtNtAfn/XzA+8xkEsbIlMvb9Xs8qghr41P9B
LBnumq2w495Bkd9RcjHR4HshAEGIltbMgsn004nGUTWrGOkIt731FQX0gs5Jckh3
d3kZiVXMC2E+I6kSKpgMe03Zsl+nSsiorCMHomFh2YSyWFzvwZOv1AYO4A9/xy8C
t6cvawflbw5X2bYdfjHhtM8pL3rkQwKSU7QrVtzAp29q5r6/lVnVioHjhpUdMu4K
HEQ0Mh8LIDR6a/F7kx4jThBxwbOULAWwoqnxWDUzNdhPKpGFe6Z6gusHC4FAUh1q
5oMA2BQtb6/d0Bjg3MMv0rWIcfMmr++ubcNYblfVJ/cjxlff5TvfByZrn6gngTto
ULWj/hdYMXrvY5MP7HLYJRMw1IaEqiQ9pr11bm1y2qKxe1NMsTCl/7XpCktjg+mv
zHouqg2jUDba4UrB20JOAvGV+LzTK550/x1jqkjYrqvwKR5jB8fxuTtSsrUnKP0n
EtUEhcTO2tAeEGoPvxtElkR1fcWXeCkfeWLFS7bs0CatDI1ucyrKj0Ype/7RPWRu
mq+yXmkRBi6P5/OyCPu3FHGcUY2O367D47kHJpy00M4BOu41GnjW9kGLmZs3gRNL
T5jqZT3cf75b4mCKVbIVRAV0bXbG0Cuc+V/rsm3vX6oUKIkjmxtx5E8ZQjnr0jDE
lX33ouMf0SuM77ejMAAniEPO5g6ikjOBOI5dyLgrTO5Kz0db+3yu3TqSJkhgzSBI
X5+gXpOzBiurOJ0g2rDwmT62hVq5RT+QHeteqSP6PCUO9s/VxOGEQpBwlJnacz6/
FzIg8Dwi9TAq6wmg1QelGju/gHPiTrNRguGYgnhE6mHMOGihgRs+k8/5K/4LsF2R
6Tq3vu/xThCo1YGUrKQpwvjn9MBHS58LYMsQdNpQiTH+uoINA179uiN3jWDc/ma1
j1/JItmz668A3pspXFgxeBNXzSAoZ0vT4l43Pk25gKtH73Q7N0cSa5nE6sEVKbxe
wZ+/r8BQNbIU3QiCiNGJimv+n6popjwfyyB2KjTOCvozHkw2n9LX3GHnGsdwhyaU
kYaewAeZrPQlcW5+X05qWyj+c6304FM+5lK0HtlpmKirulL2dTtL8ocLTBHDR5sU
a/uFR+uCHe/aIfACkY/M11VRY7r8svv8v36P+I/xs0AOxbKRgOE3E9zZW2wjynK7
7MPCrm+ORwuvTMEO0ch3wn9aGqi4yUfPCaKMTZJCSAz5pt1RAtMcB7kneYJovfkK
hZyg8/dU+ndzjNCeqQlPp/xj8gf1gIC7rDf3QITpnQpbC3xO+K07c6TH/4aMK4JO
2gmZKzWsTQ+EE1QUwk7+bRBbTntusoE6LAYGj3JOh0pTPNgCotlM1rtY6JkwY8At
XN8ex0+ygX0MkwBHNtHeT90aBW7+N2R13EuftaB/65H2tIUTi5NQCvgVRC++1zIv
5fKHn4kNFiTHjbHGoXfMWL0Zrts0HXOAm3Lpc1g+wYnH/XoNG4znV7lpHjdynUfg
XcXSfxQbzXBkXJCH/aq40joL+URLeHHPeezbChRS4wMacZWGEep1WGzCNlV0SCv6
iz/weY4HxyF5LT5bpJHxY65d1H+Sf3S+YlzkP8bBqR87PZ2y6jf9I/nBEMMCxU02
BnI+0wg7We9dKlHWKkUJZODIoFwZp6QhiUemPzO06elABuIAVYgk2l4loSh6lP3l
TrxMpBVcg0je8eBb2cV7CaFEy/pIL8sKHULn1ZLTby/7F9Xr8rZ8qSjHTxwSae57
rFe3tHY1ir7MNtsFAtMpz9xViyAhhAJ8KAexlezNKlc3bGrAVsUr6a/NpeN2U53L
cqXE7QpH6IhE96yz1vfnqk22X6sG3UAiq+Vh90n7tmsi0gnXM2C/MKamhhqrG5FZ
Bb96+VpVy+tYDNgspNfkv5twDcq6SThzL3kIcljJjs60T3UgYMpr1kiAoHppxtaT
GWPwOODq8cQL2cuJLzfEcKpVHPNmAB0pMFGe9wHib9+GyWH9zkQ9hD8rQV945D6B
aDz/AX1gqf2iaaitxy6gNL7yZQhYk48D3z4enXIUF53ceNUjvW9fVw4dngv2bCA5
aoCyH9R56PPn7LSHLGGzR0EvQPoNksMdvwTtOedL5SdxWlJ/5PDrlvBtK/ttnCqb
XDXCmeyiAIOg7tsqqFECrSo/yfh5Z/zQcTngQWnMKAmkJbWchfPw8qBiHgbzycPT
5zh65wE774fB2EuXzTiMDR1mkL8nIdCm6WDXNMESg3mpTTJOxz9L2hMBIIQos12M
XpZedHSN308R2KTaMk52DHnVFnBw+I9pgPqt8JCa2e0xYaFyXZQrDhzDoxwUO6hb
YTciVRH6kUMlapDOUazi+PS4u6rlyABpok48/DyNC3tiJzi0bKZ/ikpE0VBaIqrQ
iUduhAE1vfkZHlYwVwbOb+0YQhW/r/hoidGRJkZI3mVyRqf5e6op7ZprUAqjYJuO
4rvH7FrS/Qt0nU+GuQlfVpDF09I9fJQzmdPru0VBuCSn6pLdge5wgFfErnnKwnWj
9PIi9tBupcUk76YnvtlDrvPuhPYn7AgO+lagqlTvFU0wmQ49qb7jdduETRloZz6l
xRj+S2nV3mDf+76Pfka6v7RX5DidmK9Lpo+SZnA5yKdbnh0OKWm0CmHxO+I+o+nn
9kVagEvQRuj+YnuVeBkcKbwSZotPMLvl+dqmcXFUp0J+0A41Mlkvr7PRRIdxlArn
hXLReMC8uWHNlsOnwcwsiQDcMn2R5AgLk2+qaonGVy++EDyWSveBw7FzGesGDebE
5xWaN3xAbbO0G1KL5AlDP8CC/aPqjZ5+DVB8WgLv0Ww+hcA4iGos8a87cMllSoAp
7zHL+m21I+ktMxmwoqAEGfKPVPaJXEV9rI1lFlEredlGGJUze7c3Jp0WYoxy39l2
lQR+REzQtIMswX9PuB5UPkam7Iu5P+AFeZTPrwkiBxb33RAPShW4LNt2iI6vZEHk
SUch76t9KTUkKWpzeqoSR+5Gc9hHHIytTBxsmD8Ev/EBlKyQzv/WQh/wjOsT5LVA
QuKSTbBxm1dSufEqcGhb5+WboFZSugFS4bcN9DIT1j9n4+5X9tDGT3FxRYNswtOT
Z5xFwpWt1XKeilfz3QXxRQIpFim/+XQMYI0YZdEBCn2oRPYrZZ51PICMKJy3j4R0
Qob3uJ52MX2Vjod5zwzAfv0ZXT7IMNaihE/6dwpKJ9r4Z6re+zNdgDuHgAehWnFt
q5e/YY2e7TaQIPeoxMyU54hd8G7Mm6lJecFOZAo97EDV5nZOybCe2Eb25yElwxxv
BPXP6nGHWw9Nk3NMeFDVinVSG7SuZY5eJ5e63r2mUcZgD9vfsjwxjanPvuPpMFry
Js+FsJ9WXKu8qxm03hrObMkvkODjLJrJ9+M3NiWhDergo6DG+tb1aLfryXYvNh3B
PkqLnwA9K0K3oMelq4F78oyeqpet9jlovAIM9pji253YaLoKFd13M/ZV28QNfk6m
RMpEg8zbRZb4IcNnl+Nirz9UldBWV6s+4F8p2nf1Onir7Za9wJeNpBLAFQCgj1vq
zc8MjPSDCdFzwIrAbbZpReFoQssq9BSxehUgBhZcF+K4dmUYD14M85Tm3DHfscEo
lanPmaDtyEyWSbeJ0biDcYTiaL7mRFZi3XXVtUQqvN5PtNzYYFNJmNhUjLWfxAA+
SjQw2LUN8o7Z0jp+WW/vvuMHTR1wIzMRCC65KWOpRDEg1N0qM9/DpMtsoQJrQT59
mKWu1ILbrX6nxeuG034NAPRtihf0oy/B8iRSkfR5517ke03T8achbiMciZOpgjS1
DIIAfsShQuycX9S/M8qWEwLBpc+rzaXip3HpqvYJregPMqrnvKFq1fQgMpZT0Pu3
jESJdO+rbSoPADxtlNKXGZU/2OhVvwd7xTCYFoRWa41ssbZZ2d6oWcsXhBs/kGBw
pUqcqxmau+iytNGIUMJTvfIXkyimpfVP3Ateb2/CGmVahoG1qnn1A6i/oXnmAMFh
pnW8LQ97ZXZKtHTakLb9fxRGFJ5bhj1h9uUt+9EeXdsjLIzwcEMNvIJKDiVrcuXm
fo7KM3AMLL9HU17+/4ZsW6+5OhR/hU+tQH0vNtft933P/1JT9JKAlDKc1HZqOMdO
Fdo7Wpt+aOYDPG3A3xqwX94eQ/27McS+q6nYnd7zVWzxf1od+huRxCKnEGNgi7m5
ODddSL10fFw1e2YxBsySnVecS4B+WCmCFea7ojgQ9xCLHipTHwTc2AYD7S2DiJsO
LDejIhUsNPukpvRq391VaPShfaSQhMtRFx157E+jCJItRp+cdxe4A97H9vOL08Ih
UKi9UqQeIbsXAwoCuVcuotfcX7N0m+a7QyWPwD5nBV6ypYhLX9gLrhHpJFlXrXt9
ykCYeEdhqgkkhigJSP2GFD8jOcFeRwUyvm1GnMZjtdBvb9QOOiBTb9772gCRBmJt
QnyHFy4ESqE+8ujn9I2KciCn1VfrL8HfFuluq56SWyMaSF5RR4Z3i1aWsOCW8liq
hJt45STJ1OyRmLQtWks7KOk6bywdv0MPwlbqYqAoWbQhwOD9JWPQE11+rGIxrWVS
VnvgPRhFljJpj0ZNvnqq6p95eaRTgWdBvxFHc2+3XobIaX3JvM7yknvESlwJFrQq
9AtV9HxPLRp0C/8MnX8FxHbo07RJS96VmrLbwcmPkkhJ98RkOQAFyTxYcP2C9TCt
oJFKkPDp4x7h4SDhEWQlTLLqmKH0wxw9aXH0fqH1ux/NQFKKq0jd7SmfnMFRZHjp
Yhm2njg3Ax/7yRpP7vL7TcQvMM1ExOrWUTjTPx8PpSwBl5117dgma5m11bF789DH
rUqTc1eLDY2dBPLz+vdflY6nna1ky2ugNiPTDepY36aGzms9Rzf7phLkOXjoo9bl
OmtNHRBc/PYi9k9sbY3zgdoSIi/2fFlvUom1UgnRuIv7x7khdGROrWIL9Hr85gAf
WJAKQ4nIrGUYD2AMsv0wtDifSjaBB0cbC9GOaCFcfjiCDaoMtgQ4Jahq9p3BdcMe
cy2xTAVCjSEWeS6Rp05pwi1zBU7BbctQ2PU/G21u66Hg9AbpJF7+vU+/J3fN0eO4
BU7aNcFWSBaibGcvTcVPFPDMY9J6Ms/rvM8f/miZvE2muinOp97+gyvdF9HH1WAk
YHnZ9iv0hGHpIU47vJmVY0UHvbsFVzu09b0ro4tG4KpCUnVTqUp8x1dLrKx9j5e5
nKP3fKsWlO0De7Uo5wjh8JSZsgZXd4LWG4XtaYak/c3Kn99YtDvobqYjvMJQ/hnZ
KyOa5s6s4OePjUNT9VY35i31P9swYQrsjTS+Yg5faZJOQZo5HmAk/HaZTtj7r6Ou
2p9F2vKD0pU+KQdLBfzGRgrEVWcoJ4dt7HbFnwtm4iM0Al4ffoiqfFyHrrBS2Yaf
3ffMFX/MdudsjNYV8lz6v/48IgnyjVkgXX9n7zrPzyE0g2yqItBTnE/LRCsort9Q
holl9cH/9mlBHUtFiOz/YpW5+0M3KqgJ5UgqEVZxYahYzff3nvfBOPQjIQ2KHJhI
kKkRA7SVoKoZ4euD3jtdSFe3AQwS9cgO0jzpk5XFkaNBcbM5/eGdSu7W1yvk+W6v
4Q9FwBuVXBteph62CaFP98SHyMCZspZkBV1kM6mi4Mke6rPcUi56c3mfaIgU/9UU
x11Y+Odgh6anR6eDxI5jrNEwD/ZktohBoTsgYhdTaI/11wlIn0MPGZo8ou8WP7pz
DLLmAI2tRQzkHk9XuHUgZOVLbrfTPFTBeyNizbAIA1vGIGe/wtob9UcpkRvf4XhI
pF1x1BpdMdBcsfgBhF+Y99vPEEeF5Og28nJBJsqC2K/JjPr/0JfiVjeCM7oiDLFk
zhkRgGJckW5sOCkpd/5LfrVXB7PH0Ijzb+XwIOeaX60V9ZYKJCDtLnpz6CS0CFRD
LElnxFZTijBMn5rSHPXSGROj3kog8CrXNC1WvjldoQl882nPJlNPVbyMBHefd3Hs
Ew6PckSGtKXtVNG6Va7YkotsruvLEaK/VE5c8c99PE5F0s2jYS310ut5HHp62KOF
TshNm3qm/pMt8P3EEcehsuvxFlV0pT6t9oiddj2d6RZrlu2w2m07qoiVI9wgcLuE
HAx6ue/cMyivBdzvmVDf+q3VmKOxd6YUb3931KD4LBQufFirWBM4GP4MS0zIqOlO
mXgATCdcjPYU1cG4//N6jg4lAz5KVnieN3t8j9VSOHK0uhorUmcHcK+QCdnAj7Bn
+B5rcNpAy+ynDOmRG79SFfQywvhqK0xhulymBkN+KmZcx08cp90pRtx345UatgtP
G3CJGzWZXNA4P/qLiRN48z2y6e5owH5jcDo/yFUHR3xe5yxE3EPjXrGA9rKAFwn9
V71MsrzTrhL+r5BAe0KY9MPM/FJozT6jHqsgNQpPdXeyDy4ZibpfRU1uotv38RUd
e9V+u9W0j3NkU38Zd/PGCT3zczuOhSt55Ia3ZAdVRog2iiAkQ49jbMvq23kVTkhu
9oavSDPI4QkCZq5+GojWCruat+xttWrK2FJUaHNqYx8nuQzSgta6u5BBB3/qY/cP
WU1FI5Q31IqM5919fgXaPD6iGDoo8fd4tC9Gmd5HTtlKwXx8NYLImkZp/Z9lPlO2
gZnOmEAKATXqL31YKPWRlZYJpBYmBvmqsgRDwNhWE1jimOCGGWhSNn3fZmQLkgFJ
9g4QoiaYJ96267UjyYgqPCAm7Kg1NnQptlXgdxJFUmRU71imFLufWTxRRTfURGFq
xHaFoXatF+TLtCFNp+enZoJoev6lZdKseQQPRIAR8hSwtuyYEiRjsZ8tMwfGNRfC
/rVgimPUzxibbmZFV+CaBv049qh54OmvfCVNwZHd3D4iMPsM2hNdPMFgnbZjZWIh
WCk2LYgrWp1czJ18hDx6GNdiVxnG8ciCk1pxdkAip3H5L49uoMxUp6Lk5TDgh9cm
C1x8np/xbKLb6z/e3Y5SljK6dI2Yu3dZ0w6AGYx44k+4FW62/iC815dbhnnTWh49
Icve7k1HlGOvqG4fi+gB1LSgD5sPs17dygUVfcC0AzLqo8mlOD6hTuPtNsxtmmq7
shoTQBGh4Xn1jZ7jrczLWPB5PlDqAvEmPhlTGdvi1FVLacRbtSIOEJLl+9bKSxK5
KbyHtMFJE32Ex1B6gsEVA5chnOxSL1eUDe3JGJmIIBllc/ZpyY0ksMDLpVjB++DC
IjaOubHcrpOwmhi2m4bVGPllx3HBBzPU2W2IRDIlj3/j48G5PXj2XPSA8uYLb/mZ
XJhU2x0c8kCJc4ZcYxaipeae7bilfFAA/HqUp7YNANXUym1of6dchVerO+Y6tY7H
9dLroHYLcKLgQeHzWEFoAYJYKSHwDA9zbsSnc6U0FA1OvOHultN7aiv5Yzbxh9or
mCIDY4WDnR+3qGphBuvRvJS7dH9sU9Da6mGZJcRDvY+3DCpQkOZLngI9JE1Pg2St
aPWt6iCX2kdf907YDE3gwUFJwaYNRe0wSg8GFMMpOF18LUT3YkIgr+a/hOfnB2bt
lPn65MqIfozFoPiprGo/7rdbkAWN/WiITqvOrjon+ldIx0R2kvm2ynp5EMoonCQU
SXACiUtBgYxKc1+ESMT5+9J0T/u3y4v1fmdEnBKghZ5UwdTd8YNDqmPvvSrzdpLL
IGg/S0IZiy7egzl37O4yplH+iYO0VRuwtroKjRa7MLJ6+8vXQ3lr8tt0YOFgEwBA
RnblcVpQjlQDwtuvdlxj/UJfgLYY6q4TipMjC32CEZfeN7V+YJJsMwXNBts0dTGI
jheheISs78UooPPiaHCtfeieu8GiwG2QfO55JtDc2YoIVXAakocKDyYadKOjcErs
Omyn1CKYL6CGqhALJx8/jDH0ODSngI+PRNwiur/Dkzi5YklsEydnx8f0w73f6SLk
quEkzTLr33i61jmhbr6Mxy08U5Pe20f/NgNHuG28lMwR6264faMCoZ9GXYWh/Ka5
ohKWBGtNhNKpy1S7iqMZFAG0suHiaIJZyAQkOoFhWOF6Lpx8rvcI5Em5Wehjer1D
ukmGUzZvldzcUuViQG05nUsWz6MWeMr8+M0Pm6SMK26ZkzI3LWTRj5+u6gfMR4D7
NV24UTf3KHcsVAVUhnEOOL31YaogHUoVSIn5uktyO/SVc5L+Sv73ZwQMdCsFWBIN
E9N2VBk6Azn6uGuWjqBkvt+4F6XYrqzGx2Od1LMbSeZMKUr76lekDwLKvG5crDn3
NUlRXA3HBHHt6xQu9l85r1BUZaYn6rjO81rl39wJ77ecD92fnwZeD2dgiVFqV24v
0S1UMRxKK3KBEu0qklNTaACIqEmGMIeSMor4FCGLRsAAclWtmGuOyVW2puYoV4d6
Wp8VJv0t5W1S8ci5iXRb6ZFctnzZREhYuBKQoHyjvDC90S6x0/dfkMRZ80TIfTVV
DEsl6iKYUg59Vp2Z7IBbVoO3YvaXxTolXAZG3IC9zK5kt/op1Uv/v3pz4bQIElqa
CrJQBLl4hUiZ4PNoq+LqNaf3qKqH+Hts6PSFdmU1soAcBt+b5gD+E8gYPO0LAuk1
Gzu3tD20W1HYoN7P+NGSGHjc+aEXGQ+UjtSLsCZs1fM34L96DLQCYBfiDAzT832o
LYTgfpNdR4iFSyAuspG/59nnP5yW0RHurtNci/v+DHHApvrizNDBF85FE9+zrxbg
LFZSlqf7l42QbUrLt3z46zfeYRVM9PSSiVr+++U/7dAPGWqnZIIH76F3yfUEoJsm
Z+QSd5d1teRJvhOXXMpskA37fmARHB13TvO7pM5Yezc9w4EkD+p+MnO7WAC/D+mQ
vOMFvV1SvriGV/hwd/4oGkRM6l78auj8XXbgQ48hGRDaDv3by8dmHlaM4VpzDFQz
233x0Tb1Mc+6PYQdAlRjDtyfnPLz/OSJJIWIU2i/v/5wAUTz1zkmzOh8kLklIKM2
ZmRVIIceWQss8800QbHLyjQxqy1BEO4QHyBRIbNaSCUhLtNcNrQZiybbwpUHHTua
1IIQAnTZhn5659ipTNKCv8w6okGJ13XFIU9sge92BdePMrqQ8NL+UnCYmzuNc1fK
hBjSpyZw8hlZqo8iCiAqeQXTuiBIXQP9CivfOsIdu/+A/vPgX8bszzsC8BvshoSK
+JGNPK+xtsQ3JrHjSPWslE/1+3sU8FlGf8GKU4en7wD3qgDvMbgiP8G4debyzz+a
KIRqkWhZl4BF/YVzULfYq5Wvgm8YoeLT7Z1RxTGAAPVK13rspZdYoWqgD1OiYLiN
/zJjoqagW6An+Nbx7Tv/kkpB7bu6PBYLO1WJ7+3Vmf/fVbBMtW2TEKFzjBfUxzjR
wzzDgXVLOEs0dWiWW47vdJwYDMhnZLsGcXvEtPxpObxX+cfgk9xCODOADLqxZFUt
tkqPvsahmVVwugbv8ve6ZePdWaRZ67dcytxoXMhmpNpphXRiPzeq61zemjoWJHpw
u7/surfpzOB6jw9od5caOGgjD3W9DuQhNwbDGTec7zkMhOX1EFTzgu25WuKCLWQL
luCbOBAVV9ROQtCctBGYJQ5HoZCTPBfx6oBYOcWeTA3dKlskvXINrNKy518YXiPL
apJ9l1PdbTTZ0y2eo3W9JPzABlHJMOVHKtBqefU9GPExzhKoiGG+tWGPMfoLU7Ae
49m0SOdndiPcNTXv51okoiaIbtCW9YEUvgtMvuA92NUfSGVTaB12M5jy4R4xgTZ2
sl8iKIFbBVZ42trhRRf5IccP2ykxC8zNLMkizFLr9Umt8rTV0If0ClVO91bV0cpu
0/T2yU/0xbsTidJsA8gpdpElJx/UZZ0F/tstWmHkpc8wBSkuQFf0qE6BQRjaSrsE
+DnuNQkss7Z21fZguGZWpd6zhx+d1AVIqkkPVQPjSSSQj/fE3ycfkCNjMNDmCDms
nByuAnKkz7Gkkp3VKRj+H1u57Kcz7lPZBjJKSW+yDs23dqNYhVgIytKbOnWM5Ura
YgnKdSVyySHLx/nWmrwTKM4WOOgli0hnJUyTXNkCwqAeptfHh5Y83T5bVEoOolZT
QjcA/hTVBiMQEWvNLN/kTAcL17gAaZbUor9RDjpovnywuBk9l9f2E7eh5u2olul/
cb5qog06eBqGd2iJG/kW5b756NYQttqyX/ROKp4J6t7mmbM8P9Aei0Mw520Qv08X
3vpYE3MeXBvBi2FoEZFxr0bA8t+9EXpMqM36GE/ZGbuX+j089j4dtsHU6tAXhNkp
r0MijSauv8eR9oXqZbTgUfGG7qChnhDVLJZkxsNWuER3HORYZvSJH3MBBp4cbhJQ
rAimQvG6Ql3V3r/Ys4eiSaFmQTiYejr5jvthmNpjsALL/SJUo8LueO87t2XEAZt2
ad0IWEhURdwWPjFW0Re6RVl/5v8K4MJgl1FMqp3//3/YbzY3WVUL2tsTmcLOX9EO
C2+WrFol6Psy18HKufFxwIB4oslqBN8mJWEREniAlnu2LfVowuAyhUgyB1MnRUZ7
NT20z7XnJu/txlB+6t9o1sq6dOFD1qM3XgXtPQdvW4JHoZct5j6+erCx4VnwOLoS
Vh5w1hsgkxzYRl+Ii+Qvyw193US+oDrBFU89KomElIdCYl+xSPazZBVKd5aFo+V5
pqeVxO34AQrtj+rTpWqgMEwfXMY4X2Q83apt6y4UiPM6l1UAXRFe4Vhz7T2a2xjK
hQcjKR3AMM43q28f6XmFezb58e27ieAc7AcF/HbJ6hJquOx+pTiRMqeQ3n49GB3J
IPKjHI8Nov2KbnN464KYZmybuvkhdj3w9sNhdrQuaN8M+CmgDjWtMivwwdNjgc4J
UKpg5hfeh/Lj6Bydmg/askDOSNWMTzAMWHHOQ5AX089wJReq7yfcWjJ72dnBpU34
MCLH7hd3u6gpQlpfeTikCujYtb8YIu26FLGZO2eEZmQ4v6ef4NG1sGpFywyOa8LS
Z22LhmxdiUAQY7FOnhNvvG32M2NqVe4VfFNWzndekX/bLoJoES0SRVFbORffMeS3
A2Ra3U3q0DU8YONCzVgOQG8W0G3Fw89+LtrSPoGwP4Q2yn++FDOvyYKa1/UAK2Wk
UThIhJPF6qsHyiQ0BTeXT6DFsppaM3/irM7RL8e1Jp9gOaqAql1+Cbrrex29uzD1
l/onOQNNVUSa6PbJjAihDgeM+7mwAbLgUmjmMfUEKNDVG5BSJIABry8IGDiKZeTz
DdTmZplgyg4kypErphi3KL9ZJzA09+QfNGkfl8efzRikuJZT/qatRfBs4ZM6zrEo
HdUfmc/9YtMQjtWY9AStuEAmwQ+R+E0/LReyzZpP/7bWo+4O8Hg6ryJ8q9/5bQfT
/G36WqkpCRQjbu1mVwY6/9MA9MhYJmthdYwPPydcCMgEp6NrTnCgKrL3Ob5PMh+B
VmYl4KcYJXHWrAI2x8JlL375WFh7avqzPlLmirrHVwuHZ1zc46Bk4c+bW7jyzHq6
JnNVQ6zU5fPLfcZrrOwZklxRLmsrGYcfxUWOvU4313FTYNV1NppM0j/pGWFZCPPO
vYVqoGRZUxfFU1GOmxomS0vV/HMvh/PhqN0V3+p2Pt9OmyE7DxBbU+96NIg0VeKL
10zoiYE3dXPcbyrVteUCuf4kiP6XCP1ueu9MAniAk93fpFbXvaaDBbNiwJFhbEXV
OCvSzLrt/DsBjy58EWXeuZEVvra96GR1MoGphsHrHu+fPJAXpxHs3+U37oBdEyaR
I5CU5XqO10ckkea/Tknk+vl1Nwpu8xNxuMx7Py7rGEgTON1pVKxpIu94nKnVgJ84
hoPMpTb6OOJHQt6ydF7GXh/5uT2H1r2URruUPOatjmepPI9JxgmC31hSAdIXXDG2
5IXPusDclujgiSAJgWolcvVFTZFkbpGvJ6rbYyJutiM9jQbynhSJT5EeM6dZQ8Ib
n/eQY2EKzZLH7cWgZEmiKpBB9k5Z3l1qKDUnLj2sw0XzypE1JOZel5rOBA+eetR2
6wkHgrChTdzLfPny10QFKS2HJDyI0QPmKZ9tTOoIqQL3M2plIE4jqwz2l+KskAXD
BY2pX/q/3Cx2SpElnVtkrqDrYCudLCVOmgkbv4VppCF8MRQHUwAVMj/zizbkOiKo
fSIQr8CT6UhxQv7hk2b7PKeFvfVGcqIzmz2m1Go05jm9/v1bzDK/YJ5z524oWa6g
dme4tnKwzfJbKwilsYMQZ+Gei6JIBt/rixauGVX/CLD+0DOvNr5fKAk8kOmaoJwa
d59ppNzVgWhoP8LjDmqnZr6XPMdn4MOm4+14XisFejlEoJEES7N65G1LKlW0lKXk
/60LSbyIcz8n88moTHeoDfqV731dfSfzvmG2KgOn/1HG/Cl5CqU8F6SdiHYCNFlD
ZPPFjyCQzzNNStSxaCnZvVaJttp9NaPqHoO8SDbRxcmyTO38gaaBjciOLPAMT52Z
solb+2qbbbdFHj6tV/Unlnh2/BNiLwPQpyZnai9qF2pclkKNcDUg+sSzNix1sUs0
ZYvsxWikO+IpjTUap2X08cw85RO3+rh8WUkIqTI/Of6awdG3WqGPvAaGe8RFWiEq
jt0qgMegmgYwYqBd8w3M2eCaM5QZ5q5zCApDXWpj1UzKKXJIdxdnojebcOwobTUM
bq775OiOWybHtCh0Lf7b58fFQ0D/QVq3aU6fE3jmxZ3XVCUZG3ivgmG1PJW0xIp9
pabJueh+5HyAWdYK2bqCxOF0JfGPI8NbyrW+8qa2x685EvPRfkx28wS5+THhXBGo
9TitqbF1l2usfajPZij7sYqM38LwXuWQ7ArlMlhvtnbyYM7q+zZFyYxnad4BhCNr
45wyKGWKsWQt7Bo5NdKtmj4b12uWgLtiopxUH2gpwUw5po3oTVNPZXnlf6CZXlgT
rRrOQgABq2ZR8QVScpHgkP86JyM0rKl7yF6xWI1ri0AEYFp3D/jvNtoFcqdLAQf+
TJIOJ9j8oaqvWJJvEWoi+5OZC9COMIqMadvIvWQ3PyOkaesGAnYv8n8xWoN/s6im
U4u7roWB+Hv7eCLbGJ1V46rPC6M4mr0ncRZqiwPCXYCdio5D+z7nGxFqTvT3feJG
aYqavh8VyhDDfTJ/NJxu93mcZZTaajdvms5hAGgjOV13L1F8nOUuolAVFs3jbRrZ
wy78OCq7J0tSbU0WNcnvDBISKxRNmhm8PoqGz1ZkiJEmToVQP+EAav0MnSUDLSu4
Q2A3qQByDFi90FK+ykjfX/7Btrmv4zpKvwUZmTgIT/yp/HoY3IAY/kMATMy1Xsx5
jt45TqaTKj4ycRtvH0g4A+xvMV1IDbHSL8m1WGSnW5ck1pUrHI4df0G2fZmAQnF5
jxDRcPIugpaYehgdTsaA22tcjxuMt4VdyyZ6IyKAgQ0f/eNvpabhqWKY6JRUPkJ3
v0HT30OxAwTVhlBVYPJ5SBlHwcFX20hL6TlIZdkVog6Dm0ShVKtY6UULeSZkvmMg
PAdBXT/HuLYnrJkT2WBqFRuPg5FB9un9H7707Lev/y6FRkfZ2m6XVNWwTbDkVt9i
w/ZGeWLQsWzzW56mJuYU3jjHEjc9bn/WSXjUZArJg5v2LpNbje5nYk3qjfYqqvpP
k/9kz5WQIO2FS5uKVTE6Df2o3EwVdvOpolxRGX0L42RwBb8OYN95CndaOmiWZyQ8
KTt18mV20vjJxfg7QaHq0B8Tq9ynk/r8CXErv9ifWUcveAUc71YOyrh9GKqyzPbz
o3aEP1KrxmirXoNpx9EaeZPzzo6jGhVdvW8wRRTdpcj1/WyMdegEF0j6cujdrp82
Wkihj5/PrzpOF7qcHWddx/+JkWGG+EI93FCD5OWnvbiQZxIZchbSEufpcFMfljjn
C9eK2K1e2adIg+/fqhTK1EmA2ixu9gafL4zDWa7d0E+H2q+ODHyLSoFFOnOcg7wB
LNv85JFdvfNu/ERwfdlT+QMlJ0CB9UEJF2ktcklTXK3eSXdoAGjaH/hHe+JrVOuc
0nz/Mm+W9MwIae1gY9Z2bDs5Vl11NlVWUid5odWhvBVq68uoV1bri3Pq6xoe4561
HYWuLvVm4vFGKDh3kEyRqUUAJ+tSGyGQGbX63CrpQL3swfYChmjCBW8Gv0BVONje
9tIE220bewD/6ukED0x6Fy6RUVtDNo/SZ1CMMFHO02zwyH7yGO7JpVF2oKhNefxU
JR21o8mJdqkyHBSgjhYd7GROMP4VWVoFNWpu83NEp1JbdUWcdxWy5QvBwqq2mZAF
egvItwPrhQPMdtvvCkqsUfzXEisaJmU1se+F9I7wLal9E+ITYxjaBrQH8ShNMP9A
v1BfZGcIvnnm2F/SmhQsJxS3qvwWBCiTfvBUJU71gXfSECMxArLxDw4tne/EmHQP
OAjPFrk5VCXcfhKT0fgBBnSiRcKzGrna7PuL0UG5wduJ9fGiYuQVAaRevXFJ6Aom
jel5q04+Jy3ndJBmdVUo/4cNBACSKbXMSE+WiNPqPtyhzuWu9G0IQN+VzUIeHJtU
nlaWvx39UPRu08mbTaCrfBNFN6DoHfvbQrFu8molHVNovtGDCDvvIAlpn5OLU0FX
DWPFeZHlGWm8BYScZaGXLEKBhDgDL9eKJ80wsfFlKj6srw0r7loLtop13pFSc1Db
+lrYH9AdnzAD+YHT2kokgv1dnQ6TnpSXmA6DWFKAcaYEVWyOHWrK9UZjFTf58I95
M3t3wNaazfXFL+658Qfht8ato4mf2FgX8RBF8jDYybM0xi1WoWP3Q7e4DC3izx66
hWXAWwnMcx0+bw1p/YUmJ9IKtlt2XHHCzJtWruSs2FKP1WyPfRfnGwzv39e2HG2r
2ejKO2jZY++vQqByiHcf+WX2N55Sqwg3z/hfuw/B1DdaeIOJMNrdXrvEF3UXKjVc
hGoq2GH+dhuikG5yLmThe0uVPM2JklI30j8E6vLuUY1zGmXrUOq/5UvmcI52Svuu
d16GjARyQDqhJ9ummz6lrVXG4v4frx2eTc3sb7/dOgcN5UuVXdQyUWgyYfPfSAZD
lEjRxzp73q6Q9OXuJh8UeqCWaYxELFoooKadpGCtvGD+8bEwGOPak9a1HSp7oiQM
IC6NtRFB9iFLv2RMdif7mM/kooGd9ScWf2Anl5QLa5xiN5izxTivgjdfr/Cwagyy
IwB1W7tROhz3xEJDUI/t49CxSSwfCmsX1x3MaY/47Ue7q/QJA9p+S0duZ5XhydPv
e6lqJhywbV8fI2YsvdeJ2AwsIl664P/bP6LPjhsEkswxMyqc5OGGGSawC6hxFUUz
37fW2HipNmVhhG9BXwVRvyjhUuzlYwNJE0o7R0dYvcoUTRw2r+qb94jfFGjwpzqX
91DE94AREVEMapmr+DePfgmMRNtEav8ZwX/HpoyBW7v0ETuFKeA3rsZStHUz3/TV
xLs8J7b/GHlcg2a5mT6dPS7QC3dohjCSqnuvveygkzDX45HWjLvBdR0I0uqnO4cW
R2LoTKoChfEj/hkTqDOcUVQfigYvAGfZZx0HZvCEx0pQuk1+xTYHTfrHYc0sCBs+
YCqhC11QPI2+CW1WFzmzKPpm5aqG0uBSXB1TQcbnGXPyTLm7kkoGPnTXFw/xGRe0
Gs+9l3hrbntPQ77UsEoDFbvISWQC5vJLfJilQ8w6PBuqX6lSPom+moXk3JP2SYfR
O3iFhTOT3OCKoBiItlFR9zp+2Hdh/tehWuoszJ92dffX62eV6OlaG/R3uUwavn85
iZXRThFi/jWJRuxbwAZUMk7cH5DvxmYwiPil78qz1d38vZpNmHoV7Rt8ofxVCrwk
+HU2IOBpwOmz5DWhLeoTBFjCsvRAInqiCW/3mdpLxZ8AfNk4wOzEeHE0WSaULyYa
l1CGtdoXzNLtB1jCR5+QzERPLPyymMi/8+HH3GMJ6Scm4j0R64eKUQxhjtCpdfr1
/pGxy8fOqIXS/kxyy1nsqdcMlYXWLCGRwmDZLsX4eK76Tj8HfT4nyvoXdTOzz1bO
zcap3oZQErXJkxN7bhCa/GBPykZNx02Zn/rKgC5m0zjgz0tWU+8uKG0c1JeRfJh4
fLl0oqbbvBPH2GbTlkegt7kISqdgiQd0k3UPf0kpQa9fOuonqogqZFUmsmEkpwY/
3LByrqMz5W4RS8RmzrpvWa0Vsl/1y5yUFTnMbiOYv8QQ/NJH0h5XbM41Rn/ZqrkJ
AgCLtYwNDxPzaamKNBvabkns5uFJTWzJieDsTKl+X0ex8eRvpHQiB7DkVdPGGlNW
kym4Gc4bkpeVd05yEFS6+dN5vSvMrHMcabVCkpITmG4j9gsOXnNvvGuEdiMLXkd4
V/5fqwGfvlZjzDjrbCu4Q0STsBOeMqnErVhpAvxsLkhdxVyOzT5UgpofQvoAGEdM
AgGhBRfSa9whGT54j15LjFKyX7K4JzLjebjJBLzwi/it3tSjAIHty2Z+F74iIVFT
eTMcIsdph3eJEKNjuCCf8xZJ7E0eRr4r3oW3hhJ1RaCsEfrBEiNI93ykuGX03uyC
CON6yWfi1CIYA8QuM8wbj2a2nrwSh/UQwaOoyI/NHZlRf+4ycGVyn9/5/iLt/tFD
waTEbZVOM9/aSEcE6hEFHWd+B4BrV6RM4Qd9B2P+Hv5WiIAxmZhVZcBHsuebn6eP
bZE25lEC1KEPjkMw4nt7KuxiZ8SZB/7LBmXxf0eZmBs3z+mX59lQWp61xtKMxaop
YCcxIvbZUbnctwY8Qcy5ZcwghkXiS3dHs6cZBOzdRTLylDj5qs4ucnQe0fVAqsKA
M2fcLPm//PTxVqZhXm60xZLR69tjXqbz6qMVLLxlo0Y0hZ2Wf0O/WCY7piW6n+Wa
2DzvPNkQUds777esUwttGXHfVXqJBUKlWoptsaNfGPUJu2Oor3CDWUKbACkqGOQm
ib7YFVfwIO5jueb1sdausFBwQf7D8FQ520bhF0Br7J0oXrGbX6+FRN2nBCPwxpDa
lQ+RB0L9mfznB86/0qJOLKsc25M8o0OcayHpYcPqipuib6rjrCSJn17wpkRKzQJY
/b2Eg+UfpHUI4Um7riUY1kWpbk5/b1E7VQGMGJjssJtmpEmcufqIflM+BZI9G4ZG
9j+VeS5elkMimUvrLqAhUTTe2uqjw5dKz6VUMWy/wAGMii8HrxgfWIrm14BoMw9R
wQxyLPFqOI1VOFo0VyWPx7LXcSKtaYqu04kk7074Ntif9LvKGf0e2qsuojn9er68
ctcydhf5eG2F7W7wXeLf5+ey+Lr0I7WjG1YpqakMwcc/DccBL5+20YoG4PTsbyqT
TO2TkGQgPu/46vNiJlD1wlJnp2TfFB1lc+Ov6U7dbpNi6QDOWtv7F/WlaHJwQJ9I
SKn0RlxBQazByK2gANQusJmQ0Q9DZq2n8lCmUWtrMJfUWL8a2oRxeg3P3WxofYom
W31wCTZpEI+6+zwWMumpTZv1FkXsC6muaskU6tNeXVRrsy77mp85Al7i7fIkDx57
WqEdhECX0eq1V9lgjn62mmIDYvENiCBGl2q8qwIlR1Sy1Hp12AQY3kyYHL1BTdIU
zgqQfYT06fHohk7T/RM7svqSm7lYxq3ctvk4vqgZVQJ9wD8Yk9CkjA988zXZV2mK
B1XMVhN5fycUJlnAakhM4XLP4x9pS7QCPBZlKE/W/qze+dVyby4V3RNb6Ac7YboK
4vkFYN25u71K+M8cditqzOVQDlhO/f3SoaDapbGB2haRSbCBxZDDmHJEF4T1JX0p
bHUSfpEHxFQhak+Z1ISsHw/6rlCU+Gvv5NCTgzXE0ZKPjXo1MBboszI4Ze2/Zmp1
JgtgybQY3vT++SFgX0x4oh3HF/058uKkD1F4ilyOdwy+L+XYXc1PSA80LTAA0YAh
r4MT49JD1j1I50LRMXSNEW+dISsSVD054kqvnnb1hSQYs8qPjEkHAWTxuIs4LhRw
qAW2+BA8fygazaKg0b/C57m1SaL+eTfRRElD6lwww8fT+WB1QA8gohaT5o4gCAEI
12a31YIsKQUANCqVtLZP4fs1oyK+nYkEk/+tVVVdQQN9BhrPxUQNnx/EozQDOgvZ
u4UVbRYRUOmWp/MNDAY6ULRfNs6cVrRRukiPgIIRbQ9a5Kbkzbz6azQavpkOvaV5
51WP26w/dJ9A63UCLctB6w==
`pragma protect end_protected
