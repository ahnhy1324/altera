// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
ejl3YBrKRLpK2R0EzUmnD0ZvI/qK8CiDNubHg1oBoGDkL6AwD5thIvMSnjhJGALW9g31Ov1uYNrS
0SHuub2v21qMw2BKEXw4hxM5v/WDKIyxKjUTp7SD29WE4x9ZZTWo+LLIfBCdESCm9eQh6R9RkxWQ
rQUD0eejG1XKlJ8nHdAQqT4Y8Nm9Tuwhxa16ilhpvs6vQiQbWFMTGOjDVYIpJZth51m7UwEi0Ino
owlhMN4FHXPvRoeV8zRYz9TVftVo8qIA3drdOV69LY4MhBJ8h9KOLUhW7g03nClFhG/4BhcYQBFJ
+JLiTton26WLgHO2qAiybHWEpLUTB/g2k8DsUQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
l4w9w6I1QIYih6tqQiOS2bOSkqApa7eb/cRkY0XQxDH1C8bJ25QqiV0h2Hq+YaNy1gaO08a7e++Y
woaHWFX8asMytcBnUCH1ZD9y2rLdM8OTL9RtDwZINQ7aEgovpmx7ew8XDMFkaB4aKCrrjx9IKHbJ
9Q0c6QSUaKNjFAq6s+s4O+SitCIKSHLa7yfPzRiPRpfF72TaPPp+V3Pt9alpq+PHVlhMK5A2Mn0E
3GXupahvv+JdIVLEVzqmPAK1qgSRM0bHUZTi26JzCwp0jIsa8HNsgftQW8WbI3MnrB7BJGD4hksg
EiWXdnCDQzJm9/HEaycPpvL/FXFo8SyuCeNtmMQ3m/VC2kK8P6VSZg9nUNsTB6bGtvLeqfWBqEhb
aeMY5T66U2tAr221Gie0nu565pPyGzo8ad1puim3Rg04/rycSU5RtztJDgXCLLHvR9UUe+dJ1Jdi
3BiO0jY0ujxKzy2lQLTvkPf/U53Pvxc95xDdd2UdYan0AHe/TtFQ77vPRZcEd/iyOoq6jyozd3/a
xIhBeGcmUHffHpU23Pt6ZIlTI+09syMlXNQsi+UEO4UEa97XiYFd5qqXBO9QNj0khLoct4+e+xNb
BCTo956B1+BvXfFqnfXFSsI81NO0PPsFggf1HIGTyooIwspZgYRDDR5nw0vchkxe+jG9pDO8MYHn
fB1fHZRpA1xD0JXaOfNnzjHCvXzI/HBdVykF76Cj/UansiS9gxvUBTsqtjiYK/G7XUHm8SGQ76hn
bijQ/O+43/4L6RZVzVZBGeVZTc1TYvdMRKRKrirnNuc44+hHcx69fONBDrvejdUaXyE+o5gAWoL9
23vqAF5ZMki5p85U4VJAIMZg2J6KjRW7IY700kzqFSgPeZ1aR80frw/c/fd6DxTrXma31pwFk08P
vP1zh4Be41JU2ENg/18EdQwEVloWWnMbxRB7kb3NFtMb2Ew6WjVeExA5GniuXHOkd85I75/qRL5N
/eIuQ8cCkVZQeDn1QaKQQICP9uXR6GtMuD8hP4CdCDMg/dKU23gVmOpesDcUWOJ02fIl8qCX9Y6o
z06lUu0HLSF3KIvVf30cuwoVao8HeRXI2Q9S2u9n2qaaJDgTAKXVz2MVq+IRg3Pqrw/x3FSM1GJW
yue6LFa1k2/wfGXXKbABBDf88qoIbDN7kKfIIUSJwNVmVPYeO8vhOWdmPwlOeWvBdCtPKDVNDEbF
SanBjgGSDFZBAw8Enyn5Ru1nmXnLlDxBx99gZruDBpGjG9+T58EvpU6obsR6826zO4EAya7m8vIN
apFJCRE848Fm0AMQfBByN2e2ZokGA42OR7q/Dw10kHR/S25zVIwJnEDetojgriCrPvGAtgzVYEKM
s426ratPMC0dTFNrM5MHNPt2ZuVR3Sexx/pwzeifWs4xjthZrOLp5mDhcJsXpJwxQ+M6hqQzc5Y3
dzY2zUY5VUkgbo3REKcwgfN5UWmgmt9dmimSW7JHVA5K8ysEZgTBCM6e7fENo7UYmfGBags+g4DI
nIihvAR4dXev+/J4HRRToWA+BJxFmuRnmgquPKJgaO1IZChagcTIzBkb0ebpMusKxskyfCVQ7ooZ
BmHnYEzYVap9h9JPIn/+OMBhJhFJON4LLpcYGhwDTCELBX9EkvtCsd61kTjsxa5/OqOhcwYwjRLC
wW27eIDwdeM+dRfZKYbl3o4MIQ7nm3jT7daufzfAA6YyPTAXIKc9RI+/4a7G1OJbaRvNOZU+2F6H
1O9y83m15qRW7xrtZUFLk8W2QKjOTGn3dVS4X/oy6Wxjq7tYkXjtGuCAY44cYLZi9C4sm4e27s1D
mKS+dhVYoaOs9jIecvmaYEtD/QFNhqUOVLXVXWQ2xjWE523vrSZGOOXnULl2YnOJh4OqDAoM8Q4Q
J7sceakIOdUS1eI0kS0kGYxL3dYWVqnjORI2cg7aBaukUNE56DkAyQyJjlcuVoEF82NKQJAhxhqL
exbVN3T6r3mbRQCCmAgmPzavcRY/Zq5/Yts82aHfhbEOV9S8466v44efyHX7sd7Atlpu4Aw3iu81
p1SSaI7hQuXzA5JSXjGJcs5f89wWXqsMi3ErcOVKsKuld/F/80bRrBKE50lztmH2BW5zLe7RWcjF
8S6jtKt7NXOKOpK5zUf0b50BnJALw1eeDPQbp7gyjazr8lY8SJGzbbE65FuwQ+8dOVajSYwo+cYm
DB6c4sYJ3fPINarXk7PXUe4bzkmmg6h/+Kw37P3iNPx5xDBBoghNjZiVgOb+QIXjlnTLO4Op8xQz
QIhgVSbR3JWMi78mBlKN1ljRet5ooEHzy7+Q9HZ4e0Q8GGl8hp5HWSYJPp//xbwpMq86np1P+gDr
/WFR3LDEAClFGQdjd34IZo6YGNKcbu+kptbleaYmpJS9L8mFkN1T2Hy5pXG2ctXc6QWK+tTDouUa
7YNAmL7StGQcYTnv3rVAY1P7h9YUFm+/jmxE3wDqidPXely0zyEvAH5p71WciYaYAIE5CNe2N6Q/
+YNSxnAuAo/O21nfIaHJftpb/NsteC8ey2evT6mgsXqMnPZS9onMPachMgolbhYzIFXI9DZjwmgo
IigVYpkXQ/SeuCSYirEnFAvMOJOUkn9IkD5BZL8DgtX7E8kRXJCylc2N0Uhc5KTP71zaLoEhFQyR
78qR3PDFIAe4IBzNGVA+atYBUyyiDiSYpb3ssao6Nq9Pv5pChOv7r0sRSUQmnwMfcP7jyxRBqY1Y
MPmCQwi3QnS7lR/qRmG7zmj6ytStBbKEHcBhKaNnKWl8B7YzQhIsGmeK3U28eZdYjbzzPsRw2C1t
t415ctHe/O75ToaJXsV+/1uNlCNSHX22cj1olOHGV5QoOJkcAdDrxeD05z3NSUcORzG9snOXehjA
GWUyrdRJmuF7FJ5YDZQFsPKKPOgDe3sQMj+9e02VHo5kQxUWIZ6InhgqW63YOfXZ7sgmcqYjkgfi
h9KJjnto1aR401t6cqybUODC3u7jdiTnsV5SwefLGeX3/IOHUXK0YcM192ptbfvv9Q+gyagGdcRi
TRutWEbSqxdho9iAdGV6rErAEZp58uCaaZ9zXPWMJk8x7FICGQ7RGzNntv1XKN4UsR/cymquCZRp
Zt8SoeNoyyn1RadqmLs2Oi3bSWm3vr+8AJYMA/R4s+VMuiG3Po3AhQp4+pndVWLk1qzcwAYmedLa
NmUsPy8bDJs/FXI9O8dnG5fE8k1XfsbdM++YQmYLUp6WxqBWpxUUlsDIupSideiohdE+HjmMziNQ
u1EI+4PP9o76pYT4Lf8EENUErgtN9vGnq0PY7h0D3620Z2kz0o5nAgKLrDupC0VxOpYi1wtzzcxd
zpURckE1+bRh5bA8qufAJ1BVRuBgyxgfPpt+epJliszmigIhxdNNjK9k2bOh4fhFunEPOz/Xi9lo
RPcOILwbeK3lL7OKfy90ZqtTIZvw5Kz3M6d/GwRTgL+9Er82r3J0alEaZ+QGFiJ8FyfWsW97H3vn
wpBFG4ekpQjTaFYXmcxc7KBoa5P7BBmgfyOuXbpio8vkTi17wk7yhRgfX44GZkEqhlwUEwIz68qB
1ET8AI+EuF3paOy498BicPrPDYWTFKe+KH0ZgdcDnwCV3bzcDyuDtwU52GqE0J7088kYDQXFvN8m
LuXLBqj54ifRnpN8ApAtTO6rfr/SxQcCibXu3Azord58I9u4XohJa5/9yHUxWAMv2Z/olYWYdLGk
CZTml/vO7P7rrEXgsi+cBBTN6fPsmx9Pzs8mPZkcwXEq8NU3Ux5WiYgxV8jrpZruYoX9cRVzWeaz
at2wXRxK3jxWLkKWwJmhpVV2rNziWVDKJm2Wk3AAW4kSXugvR+xFnPxZich2uBeJtHI+Bdxhcnk8
pCkopBHH+dRaQD6igCdvgyunkosA64Y88OgReUNV+mr4X4FDiXpWfeQ+0iNBYqbCLBJhrcJB9HVD
FUQHxnm+ASIw9Xyrqhup75AwzgiuefgFR5MUgBQWxvTWbKOPwN/yKTY3CGWP0LzKGyknk6rf6w+y
YE2Nzok+JciBWO3FMaEqHB5wkK2gdu6xOYMsd6p8ZQ3jK6wozVLA7byxeXaWAz+cs/EycfMJQwml
qQoLdyobKVMB+EFLJVw5svwqySBgslXBmSV5Xk3NXtSy+1pb0JofJQ0EzYgM8e8gN/g+zhYUGWk+
kNsfTaQbpGeeivC0P9EuIMQjI4tCFJwKP30ZMsUbEbC8Igt6E/mBucPUFZlJGcvA86n2PGouzr5/
0emUS0NjcoL88HnN2LillGzNP/kJQCO2gPKRjlDGX9KkIHhaZaW1R6JI3icmgkdKQwU1NGmTl0bc
1VnX9jdknms0KMM1z6tQj9x2Ocv9j4GAqiWTIpyi2GBOjRDSXPZWITfeQViL4NJPuAsdbhrtj/A5
RtUTfbhxW407Xed/jku3kZqYF66RQv9EMbm444ZkzUxobCCCyx3W0Nr1OWmASW5ivglRJghOfna8
2As1+XYutbb2uxq/3l2mSnmEeLkhm4pfqNiuCNh5/VQlg6MCgDQGpCt1fU/tf1uQ99nYuPwhUYme
7PPbKHKzbubOX8GluJ+1nJLgn31Hj7OdGO/XwZLcn2Jw7m61DCloQQAgkA0RoP4PVEjpFaCEr87b
duR3QdD1E9ljeylhU7pV8HE0kxc9jynW7rg5aFNBcVTcdIYCt7O2Wcl6XnAvH2eqlCBwS6XUXolY
INf+y9h6rVq4ysjkk/d/Nuk8SZ9Y8k18z7UcDJ5i4/c6Gqp6d0DaWU8w72gXEhwVjlf53+37fuwT
kY3CR+Skn2j+F/ZWkX9EWFIFm2aTZhhVQe/prtOiKRqI4t5hvLSYUY0ltqrEmAXn9Gq7E2gi+lrg
YvOXuBcLWHlRvKKCL+j/OB/FfDLgh7vNqXcfWphXAW9EUEmHq4Ia7Ot3sVLtKPrH62mLouz88KwU
O/+7j/9l0KPy7hSFKBByohe/3X39ew2vwrB7terReSachOQQtT2MqosIsklTIbRlmvPbuPq2ieCr
V+FaZStLUknBKLJNCwt20d62QU9evp84ZP9t+48x0uLm0qxI74rbxC7MFpZoume2jSxK55TEVAoo
T/uthCoziXA4GywG0pmxtdvMQuSk8V60J+bZmb4RitYEw/Bk5V7zb+UASssh4BGM1tvrjATEyVbL
8LvLBDVz+b1aEOndQI6rVwzb6v6eZfCSdJtYfzSaoahCQivJiT2Jkb7wB4mR5s5EiOiNwn+23v/2
01UMdJWKH4cnGKP8g0b8u8grLUdC4SjW9D54Rm1BBMRGzGt00DyWtB3+pdRLw3p9Afmt4+7Ald5S
YwvqV/yqfUhYVhniYfKuNTR5jNEqMjOYBTmYEkF9OE4aYQTLM6biGl/xuyHsZx0nskaKBg0+Y2Zc
0MCf7qOa8YkgxMr6GB2I8MsFZ2nk0IwZja8OGASFZNRqj036UI/eq0VP19deXDqAxP7yzzQXFmDZ
WGQK3H+i7jS1ZZSleIo0IHL2rFCEm8XoyhgDV3OEZTOR5S4tfAOA0nA6jXrgjlbCFi5OANj6rhFq
s0LfXyW1iI1SCB0bjt8jyFbHaPgG2yVPkI/69TZuVkP/w8z94ruPhBCnyGUw+xfXneGgSCPsIx3q
3Cg89M2x5EIXnP0hMS0W5Q+UO3KADVP2en4lB1sfHE/PIy69fElQHnfRjyiKOK1i3eCNlZ/5IzYv
w0bSMRN38k17VPCfyMpFAbDFXh5p+2LtG84PUsfGESsdORNrpfgC0DJqpQarYeFtfyxU8BfKSIeO
s4gcpw==
`pragma protect end_protected
